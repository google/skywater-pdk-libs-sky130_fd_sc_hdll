* File: sky130_fd_sc_hdll__o221a_2.pxi.spice
* Created: Wed Sep  2 08:44:37 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221A_2%C1 N_C1_c_77_n N_C1_M1007_g N_C1_c_73_n
+ N_C1_M1002_g N_C1_c_74_n N_C1_c_75_n C1 C1 PM_SKY130_FD_SC_HDLL__O221A_2%C1
x_PM_SKY130_FD_SC_HDLL__O221A_2%B1 N_B1_c_106_n N_B1_M1001_g N_B1_c_107_n
+ N_B1_M1000_g B1 B1 PM_SKY130_FD_SC_HDLL__O221A_2%B1
x_PM_SKY130_FD_SC_HDLL__O221A_2%B2 N_B2_c_138_n N_B2_M1003_g N_B2_c_139_n
+ N_B2_M1010_g B2 B2 B2 PM_SKY130_FD_SC_HDLL__O221A_2%B2
x_PM_SKY130_FD_SC_HDLL__O221A_2%A2 N_A2_c_170_n N_A2_M1006_g N_A2_c_171_n
+ N_A2_M1008_g A2 A2 PM_SKY130_FD_SC_HDLL__O221A_2%A2
x_PM_SKY130_FD_SC_HDLL__O221A_2%A1 N_A1_c_201_n N_A1_M1005_g N_A1_c_202_n
+ N_A1_M1004_g A1 A1 PM_SKY130_FD_SC_HDLL__O221A_2%A1
x_PM_SKY130_FD_SC_HDLL__O221A_2%A_38_47# N_A_38_47#_M1002_s N_A_38_47#_M1007_s
+ N_A_38_47#_M1010_d N_A_38_47#_c_233_n N_A_38_47#_M1011_g N_A_38_47#_c_239_n
+ N_A_38_47#_M1009_g N_A_38_47#_c_240_n N_A_38_47#_M1012_g N_A_38_47#_c_234_n
+ N_A_38_47#_M1013_g N_A_38_47#_c_235_n N_A_38_47#_c_249_n N_A_38_47#_c_236_n
+ N_A_38_47#_c_237_n N_A_38_47#_c_242_n N_A_38_47#_c_258_n N_A_38_47#_c_269_n
+ N_A_38_47#_c_279_n N_A_38_47#_c_280_n N_A_38_47#_c_243_n N_A_38_47#_c_244_n
+ N_A_38_47#_c_245_n N_A_38_47#_c_246_n N_A_38_47#_c_275_n N_A_38_47#_c_277_n
+ N_A_38_47#_c_295_n N_A_38_47#_c_238_n PM_SKY130_FD_SC_HDLL__O221A_2%A_38_47#
x_PM_SKY130_FD_SC_HDLL__O221A_2%VPWR N_VPWR_M1007_d N_VPWR_M1005_d
+ N_VPWR_M1012_d N_VPWR_c_367_n N_VPWR_c_368_n N_VPWR_c_369_n N_VPWR_c_370_n
+ N_VPWR_c_371_n N_VPWR_c_372_n N_VPWR_c_373_n N_VPWR_c_374_n VPWR
+ N_VPWR_c_375_n N_VPWR_c_366_n VPWR PM_SKY130_FD_SC_HDLL__O221A_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O221A_2%X N_X_M1011_s N_X_M1009_s N_X_c_449_n
+ N_X_c_450_n N_X_c_454_n N_X_c_455_n N_X_c_443_n N_X_c_444_n X N_X_c_447_n X
+ PM_SKY130_FD_SC_HDLL__O221A_2%X
x_PM_SKY130_FD_SC_HDLL__O221A_2%A_151_47# N_A_151_47#_M1002_d
+ N_A_151_47#_M1003_d N_A_151_47#_c_489_n
+ PM_SKY130_FD_SC_HDLL__O221A_2%A_151_47#
x_PM_SKY130_FD_SC_HDLL__O221A_2%A_245_47# N_A_245_47#_M1001_d
+ N_A_245_47#_M1008_d N_A_245_47#_c_506_n N_A_245_47#_c_507_n
+ N_A_245_47#_c_520_n N_A_245_47#_c_508_n
+ PM_SKY130_FD_SC_HDLL__O221A_2%A_245_47#
x_PM_SKY130_FD_SC_HDLL__O221A_2%VGND N_VGND_M1008_s N_VGND_M1004_d
+ N_VGND_M1013_d N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n N_VGND_c_545_n
+ N_VGND_c_546_n N_VGND_c_547_n N_VGND_c_548_n N_VGND_c_549_n N_VGND_c_550_n
+ N_VGND_c_551_n VGND N_VGND_c_552_n VGND PM_SKY130_FD_SC_HDLL__O221A_2%VGND
cc_1 VNB N_C1_c_73_n 0.0187966f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.975
cc_2 VNB N_C1_c_74_n 0.0360732f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_3 VNB N_C1_c_75_n 0.0118772f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.192
cc_4 VNB C1 0.013421f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_5 VNB N_B1_c_106_n 0.0169369f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.41
cc_6 VNB N_B1_c_107_n 0.0234345f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.975
cc_7 VNB B1 0.00404875f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_8 VNB N_B2_c_138_n 0.0218477f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.41
cc_9 VNB N_B2_c_139_n 0.0283278f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.975
cc_10 VNB B2 0.00222738f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_11 VNB N_A2_c_170_n 0.0312224f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.41
cc_12 VNB N_A2_c_171_n 0.0221572f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.975
cc_13 VNB A2 0.00222688f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_14 VNB N_A1_c_201_n 0.0243241f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.41
cc_15 VNB N_A1_c_202_n 0.0169343f $X=-0.19 $Y=-0.24 $X2=0.68 $Y2=0.975
cc_16 VNB A1 0.00573183f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_17 VNB N_A_38_47#_c_233_n 0.0170601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_38_47#_c_234_n 0.0200861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_38_47#_c_235_n 0.0146062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_38_47#_c_236_n 0.00702036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_38_47#_c_237_n 0.00669912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_38_47#_c_238_n 0.0394644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_366_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_443_n 0.0133842f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.15
cc_25 VNB N_X_c_444_n 0.00414466f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_26 VNB X 0.0220177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_151_47#_c_489_n 0.00268179f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.15
cc_28 VNB N_A_245_47#_c_506_n 0.00429419f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.15
cc_29 VNB N_A_245_47#_c_507_n 0.0264606f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.15
cc_30 VNB N_A_245_47#_c_508_n 0.00253367f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.15
cc_31 VNB N_VGND_c_542_n 0.00469858f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_32 VNB N_VGND_c_543_n 0.00681291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_544_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_545_n 0.0578272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_546_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_547_n 0.020358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_548_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_549_n 0.010578f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_550_n 0.0201421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_551_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_552_n 0.246478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VPB N_C1_c_77_n 0.0197461f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.41
cc_43 VPB N_C1_c_74_n 0.0152679f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.15
cc_44 VPB N_C1_c_75_n 0.00673405f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.192
cc_45 VPB C1 0.00218988f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_46 VPB N_B1_c_107_n 0.0258592f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.975
cc_47 VPB N_B2_c_139_n 0.0318817f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=0.975
cc_48 VPB B2 0.00170303f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.15
cc_49 VPB N_A2_c_170_n 0.033402f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.41
cc_50 VPB A2 0.00166286f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.15
cc_51 VPB N_A1_c_201_n 0.0259222f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.41
cc_52 VPB N_A_38_47#_c_239_n 0.0163537f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_53 VPB N_A_38_47#_c_240_n 0.0180199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_38_47#_c_237_n 0.00575967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_38_47#_c_242_n 0.00808998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_38_47#_c_243_n 0.00463197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_38_47#_c_244_n 0.00142863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_38_47#_c_245_n 0.0011221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_38_47#_c_246_n 0.00158837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_38_47#_c_238_n 0.0216339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_367_n 0.00495553f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_62 VPB N_VPWR_c_368_n 0.00447672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_369_n 0.0140528f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_64 VPB N_VPWR_c_370_n 0.0139511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_371_n 0.024391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_372_n 0.00401341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_373_n 0.0565587f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_374_n 0.00439477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_375_n 0.0156068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_366_n 0.0513124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB X 0.0265406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_447_n 0.00936108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 N_C1_c_73_n N_B1_c_106_n 0.0206764f $X=0.68 $Y=0.975 $X2=-0.19 $Y2=-0.24
cc_74 N_C1_c_77_n N_B1_c_107_n 0.0185566f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C1_c_75_n N_B1_c_107_n 0.0241102f $X=0.655 $Y=1.192 $X2=0 $Y2=0
cc_76 N_C1_c_75_n B1 6.54684e-19 $X=0.655 $Y=1.192 $X2=0 $Y2=0
cc_77 N_C1_c_73_n N_A_38_47#_c_235_n 0.0119732f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_78 N_C1_c_77_n N_A_38_47#_c_249_n 0.010556f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_79 N_C1_c_73_n N_A_38_47#_c_236_n 0.00984489f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_80 N_C1_c_74_n N_A_38_47#_c_236_n 0.0118554f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_81 C1 N_A_38_47#_c_236_n 0.0130074f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_82 N_C1_c_77_n N_A_38_47#_c_237_n 0.00119485f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_83 N_C1_c_73_n N_A_38_47#_c_237_n 0.00611951f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_84 N_C1_c_74_n N_A_38_47#_c_237_n 0.00583306f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_85 N_C1_c_75_n N_A_38_47#_c_237_n 0.0116131f $X=0.655 $Y=1.192 $X2=0 $Y2=0
cc_86 C1 N_A_38_47#_c_237_n 0.0219283f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_87 N_C1_c_77_n N_A_38_47#_c_258_n 5.44998e-19 $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_88 N_C1_c_77_n N_A_38_47#_c_246_n 0.0160601f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_89 N_C1_c_74_n N_A_38_47#_c_246_n 0.0102869f $X=0.555 $Y=1.15 $X2=0 $Y2=0
cc_90 C1 N_A_38_47#_c_246_n 0.00787756f $X=0.23 $Y=1.19 $X2=0 $Y2=0
cc_91 N_C1_c_77_n N_VPWR_c_367_n 0.00284844f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_92 N_C1_c_77_n N_VPWR_c_371_n 0.00681208f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_93 N_C1_c_77_n N_VPWR_c_366_n 0.0132071f $X=0.655 $Y=1.41 $X2=0 $Y2=0
cc_94 N_C1_c_73_n N_A_151_47#_c_489_n 0.0044924f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_95 N_C1_c_73_n N_A_245_47#_c_506_n 2.96875e-19 $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_96 N_C1_c_73_n N_VGND_c_545_n 0.00391671f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_97 N_C1_c_73_n N_VGND_c_552_n 0.00679073f $X=0.68 $Y=0.975 $X2=0 $Y2=0
cc_98 N_B1_c_106_n N_B2_c_138_n 0.0257427f $X=1.15 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_99 N_B1_c_107_n N_B2_c_139_n 0.0871886f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_100 B1 N_B2_c_139_n 0.00122466f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B1_c_107_n B2 0.00164396f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_102 B1 B2 0.0148521f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B1_c_107_n N_A_38_47#_c_249_n 6.28257e-19 $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B1_c_106_n N_A_38_47#_c_237_n 0.00205282f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_c_107_n N_A_38_47#_c_237_n 0.00552626f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_106 B1 N_A_38_47#_c_237_n 0.0162917f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B1_c_107_n N_A_38_47#_c_242_n 0.0177907f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_108 B1 N_A_38_47#_c_242_n 0.0297378f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_109 N_B1_c_107_n N_A_38_47#_c_258_n 0.0056809f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B1_c_107_n N_A_38_47#_c_269_n 0.00674657f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B1_c_107_n N_VPWR_c_367_n 0.0119537f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B1_c_107_n N_VPWR_c_373_n 0.00604528f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_107_n N_VPWR_c_366_n 0.00965599f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B1_c_106_n N_A_151_47#_c_489_n 0.00879018f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B1_c_107_n N_A_151_47#_c_489_n 0.00171606f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_116 B1 N_A_151_47#_c_489_n 0.00437831f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_117 N_B1_c_106_n N_A_245_47#_c_506_n 0.00762262f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_107_n N_A_245_47#_c_506_n 0.00172151f $X=1.185 $Y=1.41 $X2=0 $Y2=0
cc_119 B1 N_A_245_47#_c_506_n 0.0144199f $X=1.09 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B1_c_106_n N_VGND_c_545_n 0.00366111f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_106_n N_VGND_c_552_n 0.00545176f $X=1.15 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B2_c_139_n N_A2_c_170_n 0.0107333f $X=1.61 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_123 B2 N_A2_c_170_n 0.0026414f $X=1.565 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_124 N_B2_c_139_n A2 0.00279124f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_125 B2 A2 0.0331293f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_126 B2 N_A_38_47#_M1010_d 0.00477364f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_127 N_B2_c_139_n N_A_38_47#_c_242_n 0.00138157f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_128 B2 N_A_38_47#_c_242_n 0.0188532f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_129 N_B2_c_139_n N_A_38_47#_c_258_n 0.00363785f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_130 B2 N_A_38_47#_c_258_n 0.00257934f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_131 N_B2_c_139_n N_A_38_47#_c_275_n 0.0112843f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_132 B2 N_A_38_47#_c_275_n 0.0264944f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B2_c_139_n N_A_38_47#_c_277_n 5.16332e-19 $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B2_c_139_n N_VPWR_c_373_n 0.00517074f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B2_c_139_n N_VPWR_c_366_n 0.00810495f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B2_c_138_n N_A_151_47#_c_489_n 0.00830516f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_B2_c_138_n N_A_245_47#_c_507_n 0.00821652f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_B2_c_139_n N_A_245_47#_c_507_n 0.00547992f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B2_c_138_n N_A_245_47#_c_508_n 0.00734899f $X=1.585 $Y=0.995 $X2=0
+ $Y2=0
cc_140 B2 N_A_245_47#_c_508_n 0.0301087f $X=1.565 $Y=1.105 $X2=0 $Y2=0
cc_141 N_B2_c_138_n N_VGND_c_542_n 0.00228706f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_142 N_B2_c_138_n N_VGND_c_545_n 0.00366111f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B2_c_138_n N_VGND_c_552_n 0.00663241f $X=1.585 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A2_c_170_n N_A1_c_201_n 0.094241f $X=2.585 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_145 A2 N_A1_c_201_n 0.00143837f $X=2.25 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_146 N_A2_c_171_n N_A1_c_202_n 0.0103136f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A2_c_170_n A1 0.00147145f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_148 A2 A1 0.0142111f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_149 A2 N_A_38_47#_M1010_d 0.00593972f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A2_c_170_n N_A_38_47#_c_279_n 0.0130879f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A2_c_170_n N_A_38_47#_c_280_n 0.00410101f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_152 A2 N_A_38_47#_c_280_n 0.00567933f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A2_c_170_n N_A_38_47#_c_244_n 0.00115278f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_154 A2 N_A_38_47#_c_244_n 0.013617f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A2_c_170_n N_A_38_47#_c_277_n 7.11161e-19 $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_156 A2 N_A_38_47#_c_277_n 0.0268097f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_157 N_A2_c_170_n N_VPWR_c_373_n 0.00517074f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_170_n N_VPWR_c_366_n 0.00806399f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A2_c_170_n N_A_245_47#_c_507_n 0.00683475f $X=2.585 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A2_c_171_n N_A_245_47#_c_507_n 0.0130702f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_161 A2 N_A_245_47#_c_507_n 0.0298958f $X=2.25 $Y=1.105 $X2=0 $Y2=0
cc_162 N_A2_c_171_n N_A_245_47#_c_520_n 0.0134788f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_171_n N_VGND_c_542_n 0.00534472f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_171_n N_VGND_c_547_n 0.00398883f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_171_n N_VGND_c_552_n 0.0070457f $X=2.61 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_202_n N_A_38_47#_c_233_n 0.012217f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_201_n N_A_38_47#_c_239_n 0.0271337f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A1_c_201_n N_A_38_47#_c_279_n 0.00544624f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A1_c_201_n N_A_38_47#_c_280_n 0.00595691f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_201_n N_A_38_47#_c_243_n 0.0144931f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_171 A1 N_A_38_47#_c_243_n 0.0260955f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_172 N_A1_c_201_n N_A_38_47#_c_244_n 0.00298298f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_173 A1 N_A_38_47#_c_244_n 0.0104746f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A1_c_201_n N_A_38_47#_c_245_n 9.44845e-19 $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_175 A1 N_A_38_47#_c_295_n 0.0173281f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A1_c_201_n N_A_38_47#_c_238_n 0.0262784f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_177 A1 N_A_38_47#_c_238_n 0.0015342f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_178 N_A1_c_201_n N_VPWR_c_368_n 0.0127889f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A1_c_201_n N_VPWR_c_373_n 0.00640609f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A1_c_201_n N_VPWR_c_366_n 0.0106815f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A1_c_201_n N_A_245_47#_c_507_n 0.00265789f $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_c_202_n N_A_245_47#_c_507_n 2.01812e-19 $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_183 A1 N_A_245_47#_c_507_n 0.0124324f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A1_c_201_n N_VGND_c_543_n 2.31083e-19 $X=2.995 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A1_c_202_n N_VGND_c_543_n 0.00283672f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_186 A1 N_VGND_c_543_n 0.0101626f $X=3.15 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A1_c_202_n N_VGND_c_547_n 0.00585385f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_202_n N_VGND_c_552_n 0.0107097f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_38_47#_c_242_n N_VPWR_M1007_d 0.00341819f $X=1.18 $Y=1.557 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_38_47#_c_243_n N_VPWR_M1005_d 0.00242368f $X=3.495 $Y=1.54 $X2=0
+ $Y2=0
cc_191 N_A_38_47#_c_242_n N_VPWR_c_367_n 0.0164467f $X=1.18 $Y=1.557 $X2=0 $Y2=0
cc_192 N_A_38_47#_c_258_n N_VPWR_c_367_n 0.00175043f $X=1.265 $Y=1.875 $X2=0
+ $Y2=0
cc_193 N_A_38_47#_c_269_n N_VPWR_c_367_n 0.0135613f $X=1.35 $Y=1.96 $X2=0 $Y2=0
cc_194 N_A_38_47#_c_239_n N_VPWR_c_368_n 0.00876077f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_38_47#_c_279_n N_VPWR_c_368_n 0.0130546f $X=2.795 $Y=1.96 $X2=0 $Y2=0
cc_196 N_A_38_47#_c_280_n N_VPWR_c_368_n 0.00547057f $X=2.88 $Y=1.875 $X2=0
+ $Y2=0
cc_197 N_A_38_47#_c_243_n N_VPWR_c_368_n 0.0185497f $X=3.495 $Y=1.54 $X2=0 $Y2=0
cc_198 N_A_38_47#_c_239_n N_VPWR_c_370_n 5.08766e-19 $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_38_47#_c_240_n N_VPWR_c_370_n 0.0112193f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_38_47#_c_249_n N_VPWR_c_371_n 0.0210167f $X=0.415 $Y=2.3 $X2=0 $Y2=0
cc_201 N_A_38_47#_c_269_n N_VPWR_c_373_n 0.00236727f $X=1.35 $Y=1.96 $X2=0 $Y2=0
cc_202 N_A_38_47#_c_279_n N_VPWR_c_373_n 0.00695287f $X=2.795 $Y=1.96 $X2=0
+ $Y2=0
cc_203 N_A_38_47#_c_275_n N_VPWR_c_373_n 0.00498588f $X=1.7 $Y=2.17 $X2=0 $Y2=0
cc_204 N_A_38_47#_c_277_n N_VPWR_c_373_n 0.0496909f $X=2.455 $Y=2.17 $X2=0 $Y2=0
cc_205 N_A_38_47#_c_239_n N_VPWR_c_375_n 0.00597712f $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_38_47#_c_240_n N_VPWR_c_375_n 0.00315243f $X=3.995 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_38_47#_M1007_s N_VPWR_c_366_n 0.00343707f $X=0.23 $Y=1.485 $X2=0
+ $Y2=0
cc_208 N_A_38_47#_M1010_d N_VPWR_c_366_n 0.00660656f $X=1.7 $Y=1.485 $X2=0 $Y2=0
cc_209 N_A_38_47#_c_239_n N_VPWR_c_366_n 0.0102395f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_38_47#_c_240_n N_VPWR_c_366_n 0.00378256f $X=3.995 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_38_47#_c_249_n N_VPWR_c_366_n 0.0124902f $X=0.415 $Y=2.3 $X2=0 $Y2=0
cc_212 N_A_38_47#_c_269_n N_VPWR_c_366_n 0.00444983f $X=1.35 $Y=1.96 $X2=0 $Y2=0
cc_213 N_A_38_47#_c_279_n N_VPWR_c_366_n 0.0130047f $X=2.795 $Y=1.96 $X2=0 $Y2=0
cc_214 N_A_38_47#_c_275_n N_VPWR_c_366_n 0.0086825f $X=1.7 $Y=2.17 $X2=0 $Y2=0
cc_215 N_A_38_47#_c_277_n N_VPWR_c_366_n 0.0289141f $X=2.455 $Y=2.17 $X2=0 $Y2=0
cc_216 N_A_38_47#_c_242_n A_255_297# 0.00161167f $X=1.18 $Y=1.557 $X2=-0.19
+ $Y2=-0.24
cc_217 N_A_38_47#_c_258_n A_255_297# 0.00224467f $X=1.265 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_38_47#_c_269_n A_255_297# 3.42807e-19 $X=1.35 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_38_47#_c_275_n A_255_297# 0.00631597f $X=1.7 $Y=2.17 $X2=-0.19
+ $Y2=-0.24
cc_220 N_A_38_47#_c_279_n A_535_297# 0.00450513f $X=2.795 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_38_47#_c_280_n A_535_297# 0.00256872f $X=2.88 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_222 N_A_38_47#_c_244_n A_535_297# 0.00122783f $X=2.965 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_223 N_A_38_47#_c_243_n N_X_M1009_s 0.00242346f $X=3.495 $Y=1.54 $X2=0 $Y2=0
cc_224 N_A_38_47#_c_233_n N_X_c_449_n 0.00514397f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_38_47#_c_239_n N_X_c_450_n 0.00360111f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_38_47#_c_243_n N_X_c_450_n 0.00678757f $X=3.495 $Y=1.54 $X2=0 $Y2=0
cc_227 N_A_38_47#_c_295_n N_X_c_450_n 0.00389232f $X=3.71 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_38_47#_c_238_n N_X_c_450_n 0.0026402f $X=3.995 $Y=1.202 $X2=0 $Y2=0
cc_229 N_A_38_47#_c_239_n N_X_c_454_n 0.00647521f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_38_47#_c_240_n N_X_c_455_n 0.0179209f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_38_47#_c_234_n N_X_c_443_n 0.0166517f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_38_47#_c_233_n N_X_c_444_n 0.00248453f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_38_47#_c_295_n N_X_c_444_n 0.0267239f $X=3.71 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_38_47#_c_238_n N_X_c_444_n 0.00486036f $X=3.995 $Y=1.202 $X2=0 $Y2=0
cc_235 N_A_38_47#_c_240_n X 0.0157642f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_38_47#_c_234_n X 0.0176215f $X=4.02 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_38_47#_c_243_n X 0.00691945f $X=3.495 $Y=1.54 $X2=0 $Y2=0
cc_238 N_A_38_47#_c_245_n X 0.00659725f $X=3.605 $Y=1.455 $X2=0 $Y2=0
cc_239 N_A_38_47#_c_295_n X 0.0107327f $X=3.71 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_38_47#_c_235_n N_A_151_47#_c_489_n 0.0138438f $X=0.335 $Y=0.36 $X2=0
+ $Y2=0
cc_241 N_A_38_47#_c_236_n N_A_151_47#_c_489_n 0.00543362f $X=0.655 $Y=0.805
+ $X2=0 $Y2=0
cc_242 N_A_38_47#_c_237_n N_A_245_47#_c_506_n 0.00263883f $X=0.655 $Y=1.445
+ $X2=0 $Y2=0
cc_243 N_A_38_47#_c_242_n N_A_245_47#_c_506_n 7.70925e-19 $X=1.18 $Y=1.557 $X2=0
+ $Y2=0
cc_244 N_A_38_47#_c_244_n N_A_245_47#_c_507_n 0.00162517f $X=2.965 $Y=1.54 $X2=0
+ $Y2=0
cc_245 N_A_38_47#_c_233_n N_VGND_c_543_n 0.00282267f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_38_47#_c_243_n N_VGND_c_543_n 0.00182844f $X=3.495 $Y=1.54 $X2=0
+ $Y2=0
cc_247 N_A_38_47#_c_234_n N_VGND_c_544_n 0.00438629f $X=4.02 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_A_38_47#_c_235_n N_VGND_c_545_n 0.0221435f $X=0.335 $Y=0.36 $X2=0 $Y2=0
cc_249 N_A_38_47#_c_236_n N_VGND_c_545_n 0.00249731f $X=0.655 $Y=0.805 $X2=0
+ $Y2=0
cc_250 N_A_38_47#_c_233_n N_VGND_c_550_n 0.00541763f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_38_47#_c_234_n N_VGND_c_550_n 0.00439206f $X=4.02 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_38_47#_M1002_s N_VGND_c_552_n 0.00375862f $X=0.19 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_38_47#_c_233_n N_VGND_c_552_n 0.00977145f $X=3.5 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_38_47#_c_234_n N_VGND_c_552_n 0.00719786f $X=4.02 $Y=0.995 $X2=0
+ $Y2=0
cc_255 N_A_38_47#_c_235_n N_VGND_c_552_n 0.0124484f $X=0.335 $Y=0.36 $X2=0 $Y2=0
cc_256 N_A_38_47#_c_236_n N_VGND_c_552_n 0.00470547f $X=0.655 $Y=0.805 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_366_n A_255_297# 0.00300277f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_258 N_VPWR_c_366_n A_535_297# 0.00281834f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_259 N_VPWR_c_366_n N_X_M1009_s 0.0025542f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_260 N_VPWR_c_368_n N_X_c_450_n 0.013649f $X=3.23 $Y=1.96 $X2=0 $Y2=0
cc_261 N_VPWR_c_368_n N_X_c_454_n 0.0314525f $X=3.23 $Y=1.96 $X2=0 $Y2=0
cc_262 N_VPWR_c_370_n N_X_c_454_n 0.0195074f $X=4.23 $Y=2.3 $X2=0 $Y2=0
cc_263 N_VPWR_c_375_n N_X_c_454_n 0.0186169f $X=4.015 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_366_n N_X_c_454_n 0.0110465f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_265 N_VPWR_M1012_d N_X_c_455_n 0.00179278f $X=4.085 $Y=1.485 $X2=0 $Y2=0
cc_266 N_VPWR_c_370_n N_X_c_455_n 0.00784747f $X=4.23 $Y=2.3 $X2=0 $Y2=0
cc_267 N_VPWR_c_375_n N_X_c_455_n 0.00215715f $X=4.015 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_c_366_n N_X_c_455_n 0.00473818f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_M1012_d X 0.00767541f $X=4.085 $Y=1.485 $X2=0 $Y2=0
cc_270 N_VPWR_M1012_d N_X_c_447_n 0.00271208f $X=4.085 $Y=1.485 $X2=0 $Y2=0
cc_271 N_VPWR_c_369_n N_X_c_447_n 0.00158638f $X=4.21 $Y=2.635 $X2=0 $Y2=0
cc_272 N_VPWR_c_370_n N_X_c_447_n 0.0192306f $X=4.23 $Y=2.3 $X2=0 $Y2=0
cc_273 N_VPWR_c_366_n N_X_c_447_n 0.00357059f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_274 N_X_c_443_n N_VGND_M1013_d 0.00320735f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_275 N_X_c_444_n N_VGND_c_543_n 0.00787895f $X=3.925 $Y=0.82 $X2=0 $Y2=0
cc_276 N_X_c_443_n N_VGND_c_544_n 0.013781f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_277 N_X_c_443_n N_VGND_c_549_n 0.00287861f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_278 N_X_c_449_n N_VGND_c_550_n 0.0217742f $X=3.76 $Y=0.39 $X2=0 $Y2=0
cc_279 N_X_c_443_n N_VGND_c_550_n 0.00248202f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_280 N_X_M1011_s N_VGND_c_552_n 0.0030486f $X=3.575 $Y=0.235 $X2=0 $Y2=0
cc_281 N_X_c_449_n N_VGND_c_552_n 0.0142593f $X=3.76 $Y=0.39 $X2=0 $Y2=0
cc_282 N_X_c_443_n N_VGND_c_552_n 0.0105565f $X=4.18 $Y=0.82 $X2=0 $Y2=0
cc_283 N_A_151_47#_c_489_n N_A_245_47#_M1001_d 0.00358294f $X=1.83 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_284 N_A_151_47#_c_489_n N_A_245_47#_c_506_n 0.020948f $X=1.83 $Y=0.38 $X2=0
+ $Y2=0
cc_285 N_A_151_47#_M1003_d N_A_245_47#_c_507_n 0.00397845f $X=1.66 $Y=0.235
+ $X2=0 $Y2=0
cc_286 N_A_151_47#_c_489_n N_A_245_47#_c_507_n 0.0173766f $X=1.83 $Y=0.38 $X2=0
+ $Y2=0
cc_287 N_A_151_47#_c_489_n N_VGND_c_542_n 0.0102968f $X=1.83 $Y=0.38 $X2=0 $Y2=0
cc_288 N_A_151_47#_c_489_n N_VGND_c_545_n 0.0605799f $X=1.83 $Y=0.38 $X2=0 $Y2=0
cc_289 N_A_151_47#_M1002_d N_VGND_c_552_n 0.00257403f $X=0.755 $Y=0.235 $X2=0
+ $Y2=0
cc_290 N_A_151_47#_M1003_d N_VGND_c_552_n 0.00240661f $X=1.66 $Y=0.235 $X2=0
+ $Y2=0
cc_291 N_A_151_47#_c_489_n N_VGND_c_552_n 0.0465191f $X=1.83 $Y=0.38 $X2=0 $Y2=0
cc_292 N_A_245_47#_c_507_n N_VGND_M1008_s 0.00446694f $X=2.605 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_293 N_A_245_47#_c_507_n N_VGND_c_542_n 0.0125492f $X=2.605 $Y=0.82 $X2=0
+ $Y2=0
cc_294 N_A_245_47#_c_520_n N_VGND_c_542_n 0.0212768f $X=2.82 $Y=0.39 $X2=0 $Y2=0
cc_295 N_A_245_47#_c_507_n N_VGND_c_543_n 0.00133683f $X=2.605 $Y=0.82 $X2=0
+ $Y2=0
cc_296 N_A_245_47#_c_507_n N_VGND_c_545_n 0.00384963f $X=2.605 $Y=0.82 $X2=0
+ $Y2=0
cc_297 N_A_245_47#_c_507_n N_VGND_c_547_n 0.00194552f $X=2.605 $Y=0.82 $X2=0
+ $Y2=0
cc_298 N_A_245_47#_c_520_n N_VGND_c_547_n 0.021028f $X=2.82 $Y=0.39 $X2=0 $Y2=0
cc_299 N_A_245_47#_M1001_d N_VGND_c_552_n 0.00231419f $X=1.225 $Y=0.235 $X2=0
+ $Y2=0
cc_300 N_A_245_47#_M1008_d N_VGND_c_552_n 0.00325408f $X=2.685 $Y=0.235 $X2=0
+ $Y2=0
cc_301 N_A_245_47#_c_507_n N_VGND_c_552_n 0.0126587f $X=2.605 $Y=0.82 $X2=0
+ $Y2=0
cc_302 N_A_245_47#_c_520_n N_VGND_c_552_n 0.0139896f $X=2.82 $Y=0.39 $X2=0 $Y2=0
