* File: sky130_fd_sc_hdll__o31ai_1.pex.spice
* Created: Thu Aug 27 19:22:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%A1 1 3 4 6 7 12
c24 7 0 1.7225e-19 $X=0.235 $Y=1.19
r25 12 13 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r26 10 12 31.6932 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.495 $Y2=1.202
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r28 4 13 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r29 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r30 1 12 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r31 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%A2 1 3 4 6 7 8 9 10 17
c33 1 0 1.7225e-19 $X=0.975 $Y=1.41
r34 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r35 9 10 8.13333 $w=4.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.855 $Y=1.87
+ $X2=0.855 $Y2=2.21
r36 8 9 8.13333 $w=4.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.855 $Y=1.53
+ $X2=0.855 $Y2=1.87
r37 7 8 8.13333 $w=4.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.855 $Y=1.19
+ $X2=0.855 $Y2=1.53
r38 7 17 0.717647 $w=4.98e-07 $l=3e-08 $layer=LI1_cond $X=0.855 $Y=1.19
+ $X2=0.855 $Y2=1.16
r39 4 16 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1 $Y=0.995
+ $X2=0.94 $Y2=1.16
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=0.56
r41 1 16 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.94 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%A3 1 3 4 6 9 16 17
r36 16 17 4.37928 $w=2.48e-07 $l=9.5e-08 $layer=LI1_cond $X=1.48 $Y=1.2
+ $X2=1.575 $Y2=1.2
r37 12 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.48
+ $Y=1.16 $X2=1.48 $Y2=1.16
r38 9 17 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=1.61 $Y=1.2 $X2=1.575
+ $Y2=1.2
r39 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.445 $Y=1.41
+ $X2=1.48 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.445 $Y=1.41
+ $X2=1.445 $Y2=1.985
r41 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.42 $Y=0.995
+ $X2=1.48 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.42 $Y=0.995 $X2=1.42
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%B1 1 3 4 6 7 10 17
r28 13 17 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.41 $Y=1.16
+ $X2=2.55 $Y2=1.16
r29 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.16 $X2=2.41 $Y2=1.16
r30 10 12 27.4472 $w=3.6e-07 $l=2.05e-07 $layer=POLY_cond $X=2.205 $Y=1.202
+ $X2=2.41 $Y2=1.202
r31 9 10 19.4139 $w=3.6e-07 $l=1.45e-07 $layer=POLY_cond $X=2.06 $Y=1.202
+ $X2=2.205 $Y2=1.202
r32 7 17 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=2.56 $Y=1.16 $X2=2.55
+ $Y2=1.16
r33 4 10 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.205 $Y=1.41
+ $X2=2.205 $Y2=1.202
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.205 $Y=1.41
+ $X2=2.205 $Y2=1.985
r35 1 9 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.06 $Y=0.995
+ $X2=2.06 $Y2=1.202
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.06 $Y=0.995 $X2=2.06
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%VPWR 1 2 7 9 13 15 19 21 34
r32 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 28 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r35 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 22 30 4.82229 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.42 $Y=2.72
+ $X2=0.202 $Y2=2.72
r39 22 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=0.42 $Y=2.72 $X2=0.69
+ $Y2=2.72
r40 21 33 3.40825 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.557 $Y2=2.72
r41 21 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 19 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 19 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r44 15 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.44 $Y=1.66
+ $X2=2.44 $Y2=2.34
r45 13 33 3.40825 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.44 $Y=2.635
+ $X2=2.557 $Y2=2.72
r46 13 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.44 $Y=2.635
+ $X2=2.44 $Y2=2.34
r47 9 12 23.3929 $w=3.33e-07 $l=6.8e-07 $layer=LI1_cond $X=0.252 $Y=1.66
+ $X2=0.252 $Y2=2.34
r48 7 30 2.98628 $w=3.35e-07 $l=1.07121e-07 $layer=LI1_cond $X=0.252 $Y=2.635
+ $X2=0.202 $Y2=2.72
r49 7 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.252 $Y=2.635
+ $X2=0.252 $Y2=2.34
r50 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.485 $X2=2.44 $Y2=2.34
r51 2 15 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.485 $X2=2.44 $Y2=1.66
r52 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r53 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%Y 1 2 7 8 9 10 11 12 22 36
r26 22 43 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.02 $Y=0.85
+ $X2=2.02 $Y2=0.825
r27 11 12 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=1.87
+ $X2=2.02 $Y2=2.21
r28 11 29 10.0305 $w=2.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.02 $Y=1.87
+ $X2=2.02 $Y2=1.635
r29 10 29 4.48172 $w=2.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.02 $Y=1.53
+ $X2=2.02 $Y2=1.635
r30 9 10 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.02 $Y=1.19 $X2=2.02
+ $Y2=1.53
r31 8 43 4.36048 $w=6.08e-07 $l=3e-08 $layer=LI1_cond $X=2.19 $Y=0.795 $X2=2.19
+ $Y2=0.825
r32 8 41 1.07843 $w=6.08e-07 $l=5.5e-08 $layer=LI1_cond $X=2.19 $Y=0.795
+ $X2=2.19 $Y2=0.74
r33 8 9 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.02 $Y=0.88 $X2=2.02
+ $Y2=1.19
r34 8 22 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=2.02 $Y=0.88 $X2=2.02
+ $Y2=0.85
r35 7 41 4.5098 $w=6.08e-07 $l=2.3e-07 $layer=LI1_cond $X=2.19 $Y=0.51 $X2=2.19
+ $Y2=0.74
r36 7 36 2.15686 $w=6.08e-07 $l=1.1e-07 $layer=LI1_cond $X=2.19 $Y=0.51 $X2=2.19
+ $Y2=0.4
r37 2 29 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.485 $X2=1.97 $Y2=1.635
r38 1 41 182 $w=1.7e-07 $l=5.94559e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.33 $Y2=0.74
r39 1 36 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.33 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%VGND 1 2 7 9 11 15 17 24 25 31
r36 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r37 24 25 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r38 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r39 22 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r40 21 24 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r41 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r42 19 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.21
+ $Y2=0
r43 19 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.295 $Y=0 $X2=1.61
+ $Y2=0
r44 17 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r45 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r46 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0
r47 13 15 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.21 $Y=0.085
+ $X2=1.21 $Y2=0.4
r48 12 28 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r49 11 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.21
+ $Y2=0
r50 11 12 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.345
+ $Y2=0
r51 7 28 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r52 7 9 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r53 2 15 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.075
+ $Y=0.235 $X2=1.21 $Y2=0.4
r54 1 9 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_1%A_119_47# 1 2 9 11 12 15
r33 13 15 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.59 $Y=0.735
+ $X2=1.59 $Y2=0.625
r34 11 13 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.465 $Y=0.82
+ $X2=1.59 $Y2=0.735
r35 11 12 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.465 $Y=0.82
+ $X2=0.895 $Y2=0.82
r36 7 12 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.895 $Y2=0.82
r37 7 9 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.705 $Y2=0.4
r38 2 15 182 $w=1.7e-07 $l=4.52493e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.63 $Y2=0.625
r39 1 9 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

