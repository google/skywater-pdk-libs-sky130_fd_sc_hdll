* File: sky130_fd_sc_hdll__or4_4.pex.spice
* Created: Wed Sep  2 08:49:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4_4%D 1 3 4 6 7 8 14
r31 14 15 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.545 $Y2=1.202
r32 12 14 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.285 $Y=1.202
+ $X2=0.52 $Y2=1.202
r33 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r34 7 8 12.5353 $w=2.83e-07 $l=3.1e-07 $layer=LI1_cond $X=0.227 $Y=0.85
+ $X2=0.227 $Y2=1.16
r35 4 15 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=1.202
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=0.56
r37 1 14 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.202
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41 $X2=0.52
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%C 1 3 4 6 9 12 13 20
r43 18 20 1.44055 $w=3.98e-07 $l=5e-08 $layer=LI1_cond $X=1.13 $Y=1.82 $X2=1.13
+ $Y2=1.87
r44 12 18 0.518599 $w=3.98e-07 $l=1.8e-08 $layer=LI1_cond $X=1.13 $Y=1.802
+ $X2=1.13 $Y2=1.82
r45 12 26 9.1374 $w=3.98e-07 $l=1.82e-07 $layer=LI1_cond $X=1.13 $Y=1.802
+ $X2=1.13 $Y2=1.62
r46 12 13 9.30598 $w=3.98e-07 $l=3.23e-07 $layer=LI1_cond $X=1.13 $Y=1.887
+ $X2=1.13 $Y2=2.21
r47 12 20 0.489788 $w=3.98e-07 $l=1.7e-08 $layer=LI1_cond $X=1.13 $Y=1.887
+ $X2=1.13 $Y2=1.87
r48 9 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=1.015 $Y=1.16
+ $X2=1.015 $Y2=1.62
r49 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.015
+ $Y=1.16 $X2=1.015 $Y2=1.16
r50 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.125 $Y=0.995
+ $X2=1.04 $Y2=1.16
r51 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.125 $Y=0.995
+ $X2=1.125 $Y2=0.56
r52 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.1 $Y=1.41
+ $X2=1.04 $Y2=1.16
r53 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.1 $Y=1.41 $X2=1.1
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%B 1 3 4 6 9 13 14
c38 1 0 5.72837e-20 $X=1.57 $Y=1.41
r39 14 19 7.47531 $w=3.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.685 $Y=2.21
+ $X2=1.685 $Y2=1.97
r40 13 19 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=1.685 $Y=1.87
+ $X2=1.685 $Y2=1.97
r41 12 13 11.8168 $w=3.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.63 $Y=1.45
+ $X2=1.63 $Y2=1.785
r42 9 12 9.95254 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=1.57 $Y=1.16 $X2=1.57
+ $Y2=1.45
r43 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.545
+ $Y=1.16 $X2=1.545 $Y2=1.16
r44 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.57 $Y2=1.16
r45 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.595 $Y=0.995
+ $X2=1.595 $Y2=0.56
r46 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.57 $Y=1.41
+ $X2=1.57 $Y2=1.16
r47 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.57 $Y=1.41 $X2=1.57
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%A 1 3 4 6 7 12 21
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.075
+ $Y=1.16 $X2=2.075 $Y2=1.16
r40 7 21 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.265 $Y=1.53 $X2=2.27
+ $Y2=1.53
r41 7 12 11.0886 $w=2.98e-07 $l=2.85e-07 $layer=LI1_cond $X=2.075 $Y=1.445
+ $X2=2.075 $Y2=1.16
r42 4 11 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.04 $Y=1.41
+ $X2=2.1 $Y2=1.16
r43 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.04 $Y=1.41 $X2=2.04
+ $Y2=1.985
r44 1 11 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.1 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%A_32_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 36 39 42 44 45 48 50 53 54 59 70 79
c137 70 0 5.72837e-20 $X=1.805 $Y=0.74
c138 50 0 1.60701e-19 $X=2.38 $Y=0.74
r139 79 80 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.03 $Y=1.202
+ $X2=4.055 $Y2=1.202
r140 76 77 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.535 $Y=1.202
+ $X2=3.56 $Y2=1.202
r141 75 76 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=3.09 $Y=1.202
+ $X2=3.535 $Y2=1.202
r142 74 75 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.065 $Y=1.202
+ $X2=3.09 $Y2=1.202
r143 71 72 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.595 $Y=1.202
+ $X2=2.62 $Y2=1.202
r144 60 79 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=3.825 $Y=1.202
+ $X2=4.03 $Y2=1.202
r145 60 77 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=3.825 $Y=1.202
+ $X2=3.56 $Y2=1.202
r146 59 60 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.825
+ $Y=1.16 $X2=3.825 $Y2=1.16
r147 57 74 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=2.655 $Y=1.202
+ $X2=3.065 $Y2=1.202
r148 57 72 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=2.655 $Y=1.202
+ $X2=2.62 $Y2=1.202
r149 56 59 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=2.655 $Y=1.16
+ $X2=3.825 $Y2=1.16
r150 56 57 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.655
+ $Y=1.16 $X2=2.655 $Y2=1.16
r151 54 56 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.55 $Y=1.16
+ $X2=2.655 $Y2=1.16
r152 53 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.465 $Y=1.075
+ $X2=2.55 $Y2=1.16
r153 52 53 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.465 $Y=0.825
+ $X2=2.465 $Y2=1.075
r154 51 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.89 $Y=0.74
+ $X2=1.805 $Y2=0.74
r155 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.38 $Y=0.74
+ $X2=2.465 $Y2=0.825
r156 50 51 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.38 $Y=0.74
+ $X2=1.89 $Y2=0.74
r157 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.655
+ $X2=1.805 $Y2=0.74
r158 46 48 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.805 $Y=0.655
+ $X2=1.805 $Y2=0.49
r159 45 69 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.92 $Y=0.74
+ $X2=0.835 $Y2=0.74
r160 44 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.74
+ $X2=1.805 $Y2=0.74
r161 44 45 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.72 $Y=0.74 $X2=0.92
+ $Y2=0.74
r162 40 69 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0.655
+ $X2=0.835 $Y2=0.74
r163 40 42 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.835 $Y=0.655
+ $X2=0.835 $Y2=0.49
r164 38 69 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.65 $Y=0.74
+ $X2=0.835 $Y2=0.74
r165 38 39 35.0971 $w=2.18e-07 $l=6.7e-07 $layer=LI1_cond $X=0.65 $Y=0.825
+ $X2=0.65 $Y2=1.495
r166 34 39 24.0086 $w=1.68e-07 $l=3.68e-07 $layer=LI1_cond $X=0.282 $Y=1.58
+ $X2=0.65 $Y2=1.58
r167 34 36 23.2209 $w=3.33e-07 $l=6.75e-07 $layer=LI1_cond $X=0.282 $Y=1.665
+ $X2=0.282 $Y2=2.34
r168 31 80 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.055 $Y=0.995
+ $X2=4.055 $Y2=1.202
r169 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.055 $Y=0.995
+ $X2=4.055 $Y2=0.56
r170 28 79 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.03 $Y=1.41
+ $X2=4.03 $Y2=1.202
r171 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.03 $Y=1.41
+ $X2=4.03 $Y2=1.985
r172 25 77 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.56 $Y=1.41
+ $X2=3.56 $Y2=1.202
r173 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.56 $Y=1.41
+ $X2=3.56 $Y2=1.985
r174 22 76 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.535 $Y=0.995
+ $X2=3.535 $Y2=1.202
r175 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.535 $Y=0.995
+ $X2=3.535 $Y2=0.56
r176 19 75 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.09 $Y=1.41
+ $X2=3.09 $Y2=1.202
r177 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.09 $Y=1.41
+ $X2=3.09 $Y2=1.985
r178 16 74 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.065 $Y=0.995
+ $X2=3.065 $Y2=1.202
r179 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.065 $Y=0.995
+ $X2=3.065 $Y2=0.56
r180 13 72 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.62 $Y=1.41
+ $X2=2.62 $Y2=1.202
r181 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.62 $Y=1.41
+ $X2=2.62 $Y2=1.985
r182 10 71 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.595 $Y=0.995
+ $X2=2.595 $Y2=1.202
r183 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.595 $Y=0.995
+ $X2=2.595 $Y2=0.56
r184 3 34 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=1.66
r185 3 36 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=2.34
r186 2 48 182 $w=1.7e-07 $l=3.15357e-07 $layer=licon1_NDIFF $count=1 $X=1.67
+ $Y=0.235 $X2=1.805 $Y2=0.49
r187 1 42 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.835 $Y2=0.49
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%VPWR 1 2 3 12 16 18 20 23 24 26 27 28 40 46
+ 50
r55 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r56 43 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r57 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 40 45 3.91173 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.14 $Y=2.72 $X2=4.37
+ $Y2=2.72
r59 40 42 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=4.14 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r62 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 36 50 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 35 36 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 31 35 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 31 50 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 28 50 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 26 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.2 $Y=2.72 $X2=2.99
+ $Y2=2.72
r69 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.2 $Y=2.72
+ $X2=3.325 $Y2=2.72
r70 25 42 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r71 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.325 $Y2=2.72
r72 23 35 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.07 $Y2=2.72
r73 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.205 $Y=2.72
+ $X2=2.33 $Y2=2.72
r74 22 38 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.455 $Y=2.72
+ $X2=2.33 $Y2=2.72
r76 18 45 3.23143 $w=2.5e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.265 $Y=2.635
+ $X2=4.37 $Y2=2.72
r77 18 20 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.265 $Y=2.635
+ $X2=4.265 $Y2=1.96
r78 14 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=2.72
r79 14 16 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.325 $Y=2.635
+ $X2=3.325 $Y2=1.96
r80 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.33 $Y=2.635
+ $X2=2.33 $Y2=2.72
r81 10 12 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.33 $Y=2.635
+ $X2=2.33 $Y2=1.96
r82 3 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.12
+ $Y=1.485 $X2=4.265 $Y2=1.96
r83 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.18
+ $Y=1.485 $X2=3.325 $Y2=1.96
r84 1 12 300 $w=1.7e-07 $l=5.66238e-07 $layer=licon1_PDIFF $count=2 $X=2.13
+ $Y=1.485 $X2=2.33 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%X 1 2 3 4 13 15 19 21 23 24 27 31 33 35 39
+ 41 43 46
r79 43 46 2.85869 $w=2.75e-07 $l=9e-08 $layer=LI1_cond $X=4.347 $Y=0.815
+ $X2=4.347 $Y2=0.905
r80 43 46 0.628605 $w=2.73e-07 $l=1.5e-08 $layer=LI1_cond $X=4.347 $Y=0.92
+ $X2=4.347 $Y2=0.905
r81 42 43 22.4203 $w=2.73e-07 $l=5.35e-07 $layer=LI1_cond $X=4.347 $Y=1.455
+ $X2=4.347 $Y2=0.92
r82 36 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.96 $Y=0.815
+ $X2=3.77 $Y2=0.815
r83 35 43 4.35156 $w=1.8e-07 $l=1.37e-07 $layer=LI1_cond $X=4.21 $Y=0.815
+ $X2=4.347 $Y2=0.815
r84 35 36 15.404 $w=1.78e-07 $l=2.5e-07 $layer=LI1_cond $X=4.21 $Y=0.815
+ $X2=3.96 $Y2=0.815
r85 34 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.92 $Y=1.54
+ $X2=3.795 $Y2=1.54
r86 33 42 7.32204 $w=1.7e-07 $l=1.74396e-07 $layer=LI1_cond $X=4.21 $Y=1.54
+ $X2=4.347 $Y2=1.455
r87 33 34 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=4.21 $Y=1.54
+ $X2=3.92 $Y2=1.54
r88 29 41 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=1.625
+ $X2=3.795 $Y2=1.54
r89 29 31 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.795 $Y=1.625
+ $X2=3.795 $Y2=2.3
r90 25 39 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.77 $Y=0.725 $X2=3.77
+ $Y2=0.815
r91 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.77 $Y=0.725
+ $X2=3.77 $Y2=0.39
r92 23 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.58 $Y=0.815
+ $X2=3.77 $Y2=0.815
r93 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.58 $Y=0.815
+ $X2=3.02 $Y2=0.815
r94 22 38 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.98 $Y=1.54
+ $X2=2.855 $Y2=1.54
r95 21 41 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.67 $Y=1.54
+ $X2=3.795 $Y2=1.54
r96 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.67 $Y=1.54 $X2=2.98
+ $Y2=1.54
r97 17 24 7.0541 $w=1.8e-07 $l=1.63936e-07 $layer=LI1_cond $X=2.895 $Y=0.725
+ $X2=3.02 $Y2=0.815
r98 17 19 11.0635 $w=2.48e-07 $l=2.4e-07 $layer=LI1_cond $X=2.895 $Y=0.725
+ $X2=2.895 $Y2=0.485
r99 13 38 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=1.625
+ $X2=2.855 $Y2=1.54
r100 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.855 $Y=1.625
+ $X2=2.855 $Y2=2.3
r101 4 41 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.485 $X2=3.795 $Y2=1.62
r102 4 31 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.65
+ $Y=1.485 $X2=3.795 $Y2=2.3
r103 3 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.485 $X2=2.855 $Y2=1.62
r104 3 15 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.71
+ $Y=1.485 $X2=2.855 $Y2=2.3
r105 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.61
+ $Y=0.235 $X2=3.795 $Y2=0.39
r106 1 19 182 $w=1.7e-07 $l=3.29773e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.235 $X2=2.855 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_4%VGND 1 2 3 4 5 16 18 20 24 28 32 34 36 39 40
+ 42 43 44 53 61 65 69
c86 42 0 1.60701e-19 $X=3.24 $Y=0
r87 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r88 62 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r89 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r90 58 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r91 56 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r92 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r93 53 64 3.40825 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=4.39
+ $Y2=0
r94 53 55 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.18 $Y=0 $X2=3.91
+ $Y2=0
r95 52 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r96 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r97 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r98 49 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r99 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r100 46 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.5 $Y=0 $X2=1.31
+ $Y2=0
r101 46 48 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.5 $Y=0 $X2=2.07
+ $Y2=0
r102 44 69 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0
+ $X2=0.23 $Y2=0
r103 42 51 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.24 $Y=0 $X2=2.99
+ $Y2=0
r104 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=0 $X2=3.325
+ $Y2=0
r105 41 55 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.91
+ $Y2=0
r106 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.41 $Y=0 $X2=3.325
+ $Y2=0
r107 39 48 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.07
+ $Y2=0
r108 39 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.16 $Y=0 $X2=2.35
+ $Y2=0
r109 38 51 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.99
+ $Y2=0
r110 38 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.54 $Y=0 $X2=2.35
+ $Y2=0
r111 34 64 3.40825 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.265 $Y=0.085
+ $X2=4.39 $Y2=0
r112 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.265 $Y=0.085
+ $X2=4.265 $Y2=0.39
r113 30 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=0.085
+ $X2=3.325 $Y2=0
r114 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.325 $Y=0.085
+ $X2=3.325 $Y2=0.39
r115 26 40 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0
r116 26 28 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0.4
r117 22 61 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0
r118 22 24 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.31 $Y=0.085
+ $X2=1.31 $Y2=0.4
r119 21 58 4.0045 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.37 $Y=0 $X2=0.185
+ $Y2=0
r120 20 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=1.31
+ $Y2=0
r121 20 21 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.12 $Y=0 $X2=0.37
+ $Y2=0
r122 16 58 3.13866 $w=2.5e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.185 $Y2=0
r123 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.245 $Y=0.085
+ $X2=0.245 $Y2=0.42
r124 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.13
+ $Y=0.235 $X2=4.265 $Y2=0.39
r125 4 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.14
+ $Y=0.235 $X2=3.325 $Y2=0.39
r126 3 28 182 $w=1.7e-07 $l=3.5812e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.375 $Y2=0.4
r127 2 24 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.2
+ $Y=0.235 $X2=1.335 $Y2=0.4
r128 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.42
.ends

