* File: sky130_fd_sc_hdll__o21a_4.pxi.spice
* Created: Wed Sep  2 08:43:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21A_4%A_80_21# N_A_80_21#_M1013_s N_A_80_21#_M1001_d
+ N_A_80_21#_M1004_s N_A_80_21#_c_79_n N_A_80_21#_M1005_g N_A_80_21#_c_86_n
+ N_A_80_21#_M1000_g N_A_80_21#_c_80_n N_A_80_21#_M1006_g N_A_80_21#_c_87_n
+ N_A_80_21#_M1002_g N_A_80_21#_c_81_n N_A_80_21#_M1009_g N_A_80_21#_c_88_n
+ N_A_80_21#_M1010_g N_A_80_21#_c_82_n N_A_80_21#_M1018_g N_A_80_21#_c_89_n
+ N_A_80_21#_M1017_g N_A_80_21#_c_90_n N_A_80_21#_c_83_n N_A_80_21#_c_92_n
+ N_A_80_21#_c_84_n N_A_80_21#_c_95_p N_A_80_21#_c_123_p N_A_80_21#_c_135_p
+ N_A_80_21#_c_98_p N_A_80_21#_c_85_n N_A_80_21#_c_106_p N_A_80_21#_c_112_p
+ PM_SKY130_FD_SC_HDLL__O21A_4%A_80_21#
x_PM_SKY130_FD_SC_HDLL__O21A_4%B1 N_B1_c_215_n N_B1_M1001_g N_B1_c_211_n
+ N_B1_M1013_g N_B1_c_216_n N_B1_M1011_g N_B1_c_212_n N_B1_M1015_g B1
+ N_B1_c_213_n N_B1_c_214_n PM_SKY130_FD_SC_HDLL__O21A_4%B1
x_PM_SKY130_FD_SC_HDLL__O21A_4%A1 N_A1_c_262_n N_A1_M1012_g N_A1_c_263_n
+ N_A1_M1014_g N_A1_c_264_n N_A1_M1016_g N_A1_c_265_n N_A1_M1008_g N_A1_c_266_n
+ N_A1_c_276_n N_A1_c_279_n A1 N_A1_c_267_n N_A1_c_272_n
+ PM_SKY130_FD_SC_HDLL__O21A_4%A1
x_PM_SKY130_FD_SC_HDLL__O21A_4%A2 N_A2_c_331_n N_A2_M1003_g N_A2_c_334_n
+ N_A2_M1004_g N_A2_c_332_n N_A2_M1007_g N_A2_c_335_n N_A2_M1019_g A2
+ N_A2_c_333_n N_A2_c_353_n PM_SKY130_FD_SC_HDLL__O21A_4%A2
x_PM_SKY130_FD_SC_HDLL__O21A_4%VPWR N_VPWR_M1000_s N_VPWR_M1002_s N_VPWR_M1017_s
+ N_VPWR_M1011_s N_VPWR_M1008_d N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n
+ N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n VPWR
+ N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_375_n PM_SKY130_FD_SC_HDLL__O21A_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O21A_4%X N_X_M1005_d N_X_M1009_d N_X_M1000_d N_X_M1010_d
+ N_X_c_464_n N_X_c_465_n N_X_c_511_p N_X_c_470_n N_X_c_497_n N_X_c_475_n
+ N_X_c_481_n N_X_c_484_n N_X_c_487_n X N_X_c_462_n X
+ PM_SKY130_FD_SC_HDLL__O21A_4%X
x_PM_SKY130_FD_SC_HDLL__O21A_4%VGND N_VGND_M1005_s N_VGND_M1006_s N_VGND_M1018_s
+ N_VGND_M1012_s N_VGND_M1007_s N_VGND_c_524_n N_VGND_c_525_n N_VGND_c_526_n
+ N_VGND_c_527_n N_VGND_c_528_n N_VGND_c_529_n N_VGND_c_530_n N_VGND_c_531_n
+ N_VGND_c_532_n N_VGND_c_533_n VGND N_VGND_c_534_n N_VGND_c_535_n
+ N_VGND_c_536_n N_VGND_c_537_n N_VGND_c_538_n PM_SKY130_FD_SC_HDLL__O21A_4%VGND
x_PM_SKY130_FD_SC_HDLL__O21A_4%A_525_47# N_A_525_47#_M1013_d N_A_525_47#_M1015_d
+ N_A_525_47#_M1003_d N_A_525_47#_M1016_d N_A_525_47#_c_613_n
+ N_A_525_47#_c_614_n N_A_525_47#_c_618_n PM_SKY130_FD_SC_HDLL__O21A_4%A_525_47#
cc_1 VNB N_A_80_21#_c_79_n 0.0188746f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_80_n 0.017151f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_A_80_21#_c_81_n 0.0169529f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.995
cc_4 VNB N_A_80_21#_c_82_n 0.020128f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.995
cc_5 VNB N_A_80_21#_c_83_n 0.10295f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=1.16
cc_6 VNB N_A_80_21#_c_84_n 0.00364764f $X=-0.19 $Y=-0.24 $X2=3.17 $Y2=0.76
cc_7 VNB N_A_80_21#_c_85_n 0.012317f $X=-0.19 $Y=-0.24 $X2=2.44 $Y2=0.762
cc_8 VNB N_B1_c_211_n 0.0195423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B1_c_212_n 0.0176647f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_10 VNB N_B1_c_213_n 0.00218044f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=1.41
cc_11 VNB N_B1_c_214_n 0.0418269f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=1.985
cc_12 VNB N_A1_c_262_n 0.0179525f $X=-0.19 $Y=-0.24 $X2=3.035 $Y2=0.235
cc_13 VNB N_A1_c_263_n 0.0328439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_264_n 0.0225274f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_265_n 0.0330937f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_16 VNB N_A1_c_266_n 0.00214097f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.985
cc_17 VNB N_A1_c_267_n 0.0174623f $X=-0.19 $Y=-0.24 $X2=1.83 $Y2=1.985
cc_18 VNB N_A2_c_331_n 0.016871f $X=-0.19 $Y=-0.24 $X2=3.035 $Y2=0.235
cc_19 VNB N_A2_c_332_n 0.0171269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A2_c_333_n 0.0422554f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=1.41
cc_21 VNB N_VPWR_c_375_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_462_n 0.00760135f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=1.165
cc_23 VNB X 0.0244575f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=1.16
cc_24 VNB N_VGND_c_524_n 0.0103103f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_25 VNB N_VGND_c_525_n 0.011918f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.56
cc_26 VNB N_VGND_c_526_n 0.00218451f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.995
cc_27 VNB N_VGND_c_527_n 0.016723f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.56
cc_28 VNB N_VGND_c_528_n 0.00774104f $X=-0.19 $Y=-0.24 $X2=1.915 $Y2=0.995
cc_29 VNB N_VGND_c_529_n 4.07777e-19 $X=-0.19 $Y=-0.24 $X2=2.31 $Y2=1.985
cc_30 VNB N_VGND_c_530_n 0.0389992f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.165
cc_31 VNB N_VGND_c_531_n 0.0044932f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_32 VNB N_VGND_c_532_n 0.00546647f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_33 VNB N_VGND_c_533_n 0.0136487f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_534_n 0.0160736f $X=-0.19 $Y=-0.24 $X2=3.17 $Y2=0.76
cc_35 VNB N_VGND_c_535_n 0.0187906f $X=-0.19 $Y=-0.24 $X2=4.685 $Y2=1.99
cc_36 VNB N_VGND_c_536_n 0.300075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_537_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.202
cc_38 VNB N_VGND_c_538_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_39 VNB N_A_525_47#_c_613_n 0.00310297f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.41
cc_40 VNB N_A_525_47#_c_614_n 0.00798832f $X=-0.19 $Y=-0.24 $X2=1.35 $Y2=1.985
cc_41 VPB N_A_80_21#_c_86_n 0.0188287f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.41
cc_42 VPB N_A_80_21#_c_87_n 0.0160052f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.41
cc_43 VPB N_A_80_21#_c_88_n 0.0162781f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.41
cc_44 VPB N_A_80_21#_c_89_n 0.0158373f $X=-0.19 $Y=1.305 $X2=2.31 $Y2=1.41
cc_45 VPB N_A_80_21#_c_90_n 0.012226f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.165
cc_46 VPB N_A_80_21#_c_83_n 0.0610986f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=1.16
cc_47 VPB N_A_80_21#_c_92_n 8.92831e-19 $X=-0.19 $Y=1.305 $X2=2.445 $Y2=1.83
cc_48 VPB N_B1_c_215_n 0.0165873f $X=-0.19 $Y=1.305 $X2=3.035 $Y2=0.235
cc_49 VPB N_B1_c_216_n 0.0175647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_B1_c_213_n 0.00149701f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.41
cc_51 VPB N_B1_c_214_n 0.0228408f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.985
cc_52 VPB N_A1_c_263_n 0.0309823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A1_c_265_n 0.0320398f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_54 VPB N_A1_c_266_n 0.0012417f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.985
cc_55 VPB N_A1_c_267_n 0.00735524f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_56 VPB N_A1_c_272_n 0.0101609f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_57 VPB N_A2_c_334_n 0.01619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A2_c_335_n 0.0165971f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.995
cc_59 VPB N_A2_c_333_n 0.0216759f $X=-0.19 $Y=1.305 $X2=1.35 $Y2=1.41
cc_60 VPB N_VPWR_c_376_n 0.0274705f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=0.56
cc_61 VPB N_VPWR_c_377_n 3.26289e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=0.995
cc_62 VPB N_VPWR_c_378_n 0.00564356f $X=-0.19 $Y=1.305 $X2=1.83 $Y2=1.985
cc_63 VPB N_VPWR_c_379_n 0.0122798f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.995
cc_64 VPB N_VPWR_c_380_n 0.0255024f $X=-0.19 $Y=1.305 $X2=1.915 $Y2=0.56
cc_65 VPB N_VPWR_c_381_n 0.0190198f $X=-0.19 $Y=1.305 $X2=2.31 $Y2=1.985
cc_66 VPB N_VPWR_c_382_n 0.00631318f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=1.165
cc_67 VPB N_VPWR_c_383_n 0.0153494f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_68 VPB N_VPWR_c_384_n 0.0145309f $X=-0.19 $Y=1.305 $X2=2.445 $Y2=1.335
cc_69 VPB N_VPWR_c_385_n 0.0146064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_386_n 0.04369f $X=-0.19 $Y=1.305 $X2=2.44 $Y2=0.762
cc_71 VPB N_VPWR_c_387_n 0.00612933f $X=-0.19 $Y=1.305 $X2=4.685 $Y2=2.02
cc_72 VPB N_VPWR_c_388_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.202
cc_73 VPB N_VPWR_c_389_n 0.00573392f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.202
cc_74 VPB N_VPWR_c_375_n 0.0574779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_X_c_464_n 0.00546147f $X=-0.19 $Y=1.305 $X2=0.87 $Y2=1.985
cc_76 VPB N_X_c_465_n 0.0190662f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=0.995
cc_77 VPB X 0.0128201f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=1.16
cc_78 N_A_80_21#_c_89_n N_B1_c_215_n 0.0311995f $X=2.31 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_80_21#_c_92_n N_B1_c_215_n 0.00627588f $X=2.445 $Y=1.83 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_80_21#_c_95_p N_B1_c_215_n 0.0147918f $X=2.955 $Y=1.957 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_80_21#_c_84_n N_B1_c_211_n 0.0116464f $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_85_n N_B1_c_211_n 0.00454125f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_98_p N_B1_c_216_n 0.0183219f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_84_n N_B1_c_212_n 0.00632215f $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_85 N_A_80_21#_M1001_d N_B1_c_213_n 0.00287485f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_83_n N_B1_c_213_n 3.15696e-19 $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_84_n N_B1_c_213_n 0.0377787f $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_95_p N_B1_c_213_n 0.0104133f $X=2.955 $Y=1.957 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_98_p N_B1_c_213_n 0.00977019f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_85_n N_B1_c_213_n 0.0438518f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_106_p N_B1_c_213_n 0.0174608f $X=3.05 $Y=1.96 $X2=0 $Y2=0
cc_92 N_A_80_21#_c_83_n N_B1_c_214_n 0.016892f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_80_21#_c_84_n N_B1_c_214_n 0.00736715f $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_85_n N_B1_c_214_n 0.00449669f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_106_p N_B1_c_214_n 0.00100311f $X=3.05 $Y=1.96 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_98_p N_A1_c_263_n 0.0185916f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_97 N_A_80_21#_c_112_p N_A1_c_263_n 0.00152341f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_98 N_A_80_21#_c_112_p N_A1_c_265_n 0.00174563f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_99 N_A_80_21#_M1004_s N_A1_c_276_n 0.00355698f $X=4.56 $Y=1.485 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_98_p N_A1_c_276_n 0.0193975f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_112_p N_A1_c_276_n 0.0209957f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_98_p N_A1_c_279_n 0.0238919f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_98_p N_A2_c_334_n 0.010382f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_112_p N_A2_c_334_n 0.0110904f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_112_p N_A2_c_335_n 0.0108362f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_92_n N_VPWR_M1017_s 0.00365721f $X=2.445 $Y=1.83 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_95_p N_VPWR_M1017_s 0.00489156f $X=2.955 $Y=1.957 $X2=0
+ $Y2=0
cc_108 N_A_80_21#_c_123_p N_VPWR_M1017_s 0.00113906f $X=2.565 $Y=1.957 $X2=0
+ $Y2=0
cc_109 N_A_80_21#_c_98_p N_VPWR_M1011_s 0.0177523f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_86_n N_VPWR_c_376_n 0.0250826f $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_87_n N_VPWR_c_376_n 6.00901e-19 $X=1.35 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_80_21#_c_86_n N_VPWR_c_377_n 6.36327e-19 $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_80_21#_c_87_n N_VPWR_c_377_n 0.0145038f $X=1.35 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_88_n N_VPWR_c_377_n 0.0109673f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_89_n N_VPWR_c_377_n 6.00901e-19 $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_98_p N_VPWR_c_378_n 0.0253598f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_112_p N_VPWR_c_378_n 0.00459043f $X=4.685 $Y=1.99 $X2=0
+ $Y2=0
cc_118 N_A_80_21#_c_112_p N_VPWR_c_380_n 0.0142916f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_119 N_A_80_21#_c_95_p N_VPWR_c_381_n 0.00330094f $X=2.955 $Y=1.957 $X2=0
+ $Y2=0
cc_120 N_A_80_21#_c_135_p N_VPWR_c_381_n 0.0165836f $X=3.05 $Y=2.3 $X2=0 $Y2=0
cc_121 N_A_80_21#_c_98_p N_VPWR_c_381_n 0.00481355f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_122 N_A_80_21#_c_86_n N_VPWR_c_384_n 0.00642146f $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_80_21#_c_87_n N_VPWR_c_384_n 0.00447018f $X=1.35 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_80_21#_c_88_n N_VPWR_c_385_n 0.00642146f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_80_21#_c_89_n N_VPWR_c_385_n 0.00438099f $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_80_21#_c_98_p N_VPWR_c_386_n 0.010345f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_127 N_A_80_21#_c_112_p N_VPWR_c_386_n 0.0196466f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_128 N_A_80_21#_c_88_n N_VPWR_c_389_n 5.34966e-19 $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_80_21#_c_89_n N_VPWR_c_389_n 0.00933723f $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_80_21#_c_95_p N_VPWR_c_389_n 0.00863002f $X=2.955 $Y=1.957 $X2=0
+ $Y2=0
cc_131 N_A_80_21#_c_123_p N_VPWR_c_389_n 0.0140817f $X=2.565 $Y=1.957 $X2=0
+ $Y2=0
cc_132 N_A_80_21#_M1001_d N_VPWR_c_375_n 0.00316828f $X=2.9 $Y=1.485 $X2=0 $Y2=0
cc_133 N_A_80_21#_M1004_s N_VPWR_c_375_n 0.00240217f $X=4.56 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_A_80_21#_c_86_n N_VPWR_c_375_n 0.0107337f $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_80_21#_c_87_n N_VPWR_c_375_n 0.00766229f $X=1.35 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_80_21#_c_88_n N_VPWR_c_375_n 0.0107337f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_80_21#_c_89_n N_VPWR_c_375_n 0.00730029f $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_80_21#_c_95_p N_VPWR_c_375_n 0.00625016f $X=2.955 $Y=1.957 $X2=0
+ $Y2=0
cc_139 N_A_80_21#_c_123_p N_VPWR_c_375_n 0.00140781f $X=2.565 $Y=1.957 $X2=0
+ $Y2=0
cc_140 N_A_80_21#_c_135_p N_VPWR_c_375_n 0.00913903f $X=3.05 $Y=2.3 $X2=0 $Y2=0
cc_141 N_A_80_21#_c_98_p N_VPWR_c_375_n 0.0274858f $X=4.495 $Y=1.99 $X2=0 $Y2=0
cc_142 N_A_80_21#_c_112_p N_VPWR_c_375_n 0.0138432f $X=4.685 $Y=1.99 $X2=0 $Y2=0
cc_143 N_A_80_21#_c_86_n N_X_c_464_n 0.0184107f $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_80_21#_c_90_n N_X_c_464_n 0.0300828f $X=2.315 $Y=1.165 $X2=0 $Y2=0
cc_145 N_A_80_21#_c_83_n N_X_c_464_n 0.00634591f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_80_21#_c_80_n N_X_c_470_n 0.0106979f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_80_21#_c_81_n N_X_c_470_n 0.0104591f $X=1.435 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_80_21#_c_82_n N_X_c_470_n 0.00536307f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_80_21#_c_83_n N_X_c_470_n 0.0067559f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_80_21#_c_85_n N_X_c_470_n 0.00587745f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_151 N_A_80_21#_c_87_n N_X_c_475_n 0.0149729f $X=1.35 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_80_21#_c_88_n N_X_c_475_n 0.0162133f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_80_21#_c_89_n N_X_c_475_n 0.00116864f $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_80_21#_c_90_n N_X_c_475_n 0.0586661f $X=2.315 $Y=1.165 $X2=0 $Y2=0
cc_155 N_A_80_21#_c_83_n N_X_c_475_n 0.00299718f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_80_21#_c_92_n N_X_c_475_n 0.0137331f $X=2.445 $Y=1.83 $X2=0 $Y2=0
cc_157 N_A_80_21#_c_89_n N_X_c_481_n 0.00533329f $X=2.31 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_80_21#_c_92_n N_X_c_481_n 0.00933464f $X=2.445 $Y=1.83 $X2=0 $Y2=0
cc_159 N_A_80_21#_c_123_p N_X_c_481_n 0.0201226f $X=2.565 $Y=1.957 $X2=0 $Y2=0
cc_160 N_A_80_21#_c_79_n N_X_c_484_n 0.0143761f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_80_21#_c_90_n N_X_c_484_n 0.0793739f $X=2.315 $Y=1.165 $X2=0 $Y2=0
cc_162 N_A_80_21#_c_83_n N_X_c_484_n 0.00337291f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_80_21#_c_90_n N_X_c_487_n 0.0147777f $X=2.315 $Y=1.165 $X2=0 $Y2=0
cc_164 N_A_80_21#_c_83_n N_X_c_487_n 0.00142106f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_80_21#_c_79_n X 0.016142f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_80_21#_c_86_n X 0.00332236f $X=0.87 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_80_21#_c_90_n X 0.0278999f $X=2.315 $Y=1.165 $X2=0 $Y2=0
cc_168 N_A_80_21#_c_83_n X 0.0022064f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_80_21#_c_98_p A_826_297# 0.0038039f $X=4.495 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_80_21#_c_79_n N_VGND_c_525_n 0.00966928f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_80_21#_c_80_n N_VGND_c_525_n 0.00118056f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_80_21#_c_80_n N_VGND_c_526_n 0.0016992f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_80_21#_c_81_n N_VGND_c_526_n 0.00817928f $X=1.435 $Y=0.995 $X2=0
+ $Y2=0
cc_174 N_A_80_21#_c_82_n N_VGND_c_526_n 0.00108517f $X=1.915 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_80_21#_c_81_n N_VGND_c_527_n 0.00351072f $X=1.435 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_80_21#_c_82_n N_VGND_c_527_n 0.00558173f $X=1.915 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_80_21#_c_82_n N_VGND_c_528_n 0.00336831f $X=1.915 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_80_21#_c_90_n N_VGND_c_528_n 0.00946301f $X=2.315 $Y=1.165 $X2=0
+ $Y2=0
cc_179 N_A_80_21#_c_83_n N_VGND_c_528_n 0.00567011f $X=2.195 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_80_21#_c_85_n N_VGND_c_528_n 0.00224089f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_181 N_A_80_21#_c_84_n N_VGND_c_530_n 3.56478e-19 $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_182 N_A_80_21#_c_85_n N_VGND_c_530_n 0.00425926f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_183 N_A_80_21#_c_79_n N_VGND_c_534_n 0.00353537f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_80_21#_c_80_n N_VGND_c_534_n 0.00422112f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_80_21#_M1013_s N_VGND_c_536_n 0.00216833f $X=3.035 $Y=0.235 $X2=0
+ $Y2=0
cc_186 N_A_80_21#_c_79_n N_VGND_c_536_n 0.00428642f $X=0.475 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_80_21#_c_80_n N_VGND_c_536_n 0.0059085f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_80_21#_c_81_n N_VGND_c_536_n 0.00424612f $X=1.435 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_80_21#_c_82_n N_VGND_c_536_n 0.0112026f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_80_21#_c_84_n N_VGND_c_536_n 0.00204802f $X=3.17 $Y=0.76 $X2=0 $Y2=0
cc_191 N_A_80_21#_c_85_n N_VGND_c_536_n 0.00668324f $X=2.44 $Y=0.762 $X2=0 $Y2=0
cc_192 N_A_80_21#_c_84_n N_A_525_47#_M1013_d 0.00750608f $X=3.17 $Y=0.76
+ $X2=-0.19 $Y2=-0.24
cc_193 N_A_80_21#_M1013_s N_A_525_47#_c_613_n 0.00305179f $X=3.035 $Y=0.235
+ $X2=0 $Y2=0
cc_194 N_A_80_21#_c_84_n N_A_525_47#_c_613_n 0.0442241f $X=3.17 $Y=0.76 $X2=0
+ $Y2=0
cc_195 N_A_80_21#_c_84_n N_A_525_47#_c_618_n 0.01063f $X=3.17 $Y=0.76 $X2=0
+ $Y2=0
cc_196 N_B1_c_212_n N_A1_c_262_n 0.0142332f $X=3.38 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_197 N_B1_c_216_n N_A1_c_263_n 0.0255321f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_213_n N_A1_c_263_n 0.00257386f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_c_214_n N_A1_c_263_n 0.0186263f $X=3.34 $Y=1.202 $X2=0 $Y2=0
cc_200 N_B1_c_216_n N_A1_c_266_n 3.30378e-19 $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B1_c_213_n N_A1_c_266_n 0.0251297f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_202 N_B1_c_214_n N_A1_c_266_n 0.00116539f $X=3.34 $Y=1.202 $X2=0 $Y2=0
cc_203 N_B1_c_216_n N_A1_c_279_n 0.00276964f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B1_c_216_n N_VPWR_c_378_n 0.00587295f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B1_c_215_n N_VPWR_c_381_n 0.00467604f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B1_c_216_n N_VPWR_c_381_n 0.00506535f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B1_c_215_n N_VPWR_c_389_n 0.00769171f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B1_c_216_n N_VPWR_c_389_n 0.00101916f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_215_n N_VPWR_c_375_n 0.00542545f $X=2.81 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B1_c_216_n N_VPWR_c_375_n 0.00739241f $X=3.34 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B1_c_211_n N_VGND_c_528_n 0.00217307f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B1_c_212_n N_VGND_c_529_n 8.57813e-19 $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B1_c_211_n N_VGND_c_530_n 0.00357877f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_212_n N_VGND_c_530_n 0.00357877f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B1_c_211_n N_VGND_c_536_n 0.00655123f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B1_c_212_n N_VGND_c_536_n 0.00569584f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B1_c_211_n N_A_525_47#_c_613_n 0.00912735f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B1_c_212_n N_A_525_47#_c_613_n 0.0123547f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_213_n N_A_525_47#_c_613_n 0.00245524f $X=3.32 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B1_c_212_n N_A_525_47#_c_618_n 0.0063644f $X=3.38 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A1_c_262_n N_A2_c_331_n 0.0239928f $X=3.985 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_222 N_A1_c_263_n N_A2_c_334_n 0.0639383f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A1_c_266_n N_A2_c_334_n 5.26034e-19 $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A1_c_276_n N_A2_c_334_n 0.0145798f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_225 N_A1_c_264_n N_A2_c_332_n 0.0226992f $X=5.405 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A1_c_265_n N_A2_c_335_n 0.0508339f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A1_c_276_n N_A2_c_335_n 0.018939f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_228 N_A1_c_267_n N_A2_c_335_n 4.53944e-19 $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A1_c_263_n N_A2_c_333_n 0.024642f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A1_c_265_n N_A2_c_333_n 0.0261251f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A1_c_266_n N_A2_c_333_n 0.00191128f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A1_c_276_n N_A2_c_333_n 0.00843868f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_233 N_A1_c_267_n N_A2_c_333_n 0.0016748f $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A1_c_263_n N_A2_c_353_n 0.0011681f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A1_c_265_n N_A2_c_353_n 0.00114226f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_266_n N_A2_c_353_n 0.0163973f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A1_c_276_n N_A2_c_353_n 0.0425646f $X=5.41 $Y=1.6 $X2=0 $Y2=0
cc_238 N_A1_c_267_n N_A2_c_353_n 0.0153249f $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A1_c_279_n N_VPWR_M1011_s 0.00429182f $X=4.115 $Y=1.6 $X2=0 $Y2=0
cc_240 N_A1_c_272_n N_VPWR_M1008_d 0.00424303f $X=5.645 $Y=1.495 $X2=0 $Y2=0
cc_241 N_A1_c_263_n N_VPWR_c_378_n 0.00666331f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A1_c_265_n N_VPWR_c_380_n 0.0208268f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A1_c_272_n N_VPWR_c_380_n 0.0251255f $X=5.645 $Y=1.495 $X2=0 $Y2=0
cc_244 N_A1_c_263_n N_VPWR_c_386_n 0.00506535f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A1_c_265_n N_VPWR_c_386_n 0.00447018f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A1_c_263_n N_VPWR_c_375_n 0.00719994f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A1_c_265_n N_VPWR_c_375_n 0.00776557f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A1_c_276_n A_826_297# 0.00678231f $X=5.41 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_249 N_A1_c_276_n A_1008_297# 0.013935f $X=5.41 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_250 N_A1_c_262_n N_VGND_c_529_n 0.00632487f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A1_c_262_n N_VGND_c_530_n 0.00407353f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A1_c_264_n N_VGND_c_532_n 0.0144186f $X=5.405 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A1_c_264_n N_VGND_c_535_n 0.0035176f $X=5.405 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A1_c_262_n N_VGND_c_536_n 0.00502672f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A1_c_264_n N_VGND_c_536_n 0.00517023f $X=5.405 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A1_c_262_n N_A_525_47#_c_614_n 0.00988092f $X=3.985 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A1_c_263_n N_A_525_47#_c_614_n 9.56499e-19 $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_c_264_n N_A_525_47#_c_614_n 0.0122857f $X=5.405 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A1_c_265_n N_A_525_47#_c_614_n 0.00140671f $X=5.43 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_266_n N_A_525_47#_c_614_n 0.0130949f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A1_c_267_n N_A_525_47#_c_614_n 0.0270518f $X=5.495 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A1_c_263_n N_A_525_47#_c_618_n 0.00270105f $X=4.04 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_266_n N_A_525_47#_c_618_n 0.00855765f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A2_c_335_n N_VPWR_c_380_n 0.00284923f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A2_c_334_n N_VPWR_c_386_n 0.00481901f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A2_c_335_n N_VPWR_c_386_n 0.00681596f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A2_c_334_n N_VPWR_c_375_n 0.00643974f $X=4.47 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A2_c_335_n N_VPWR_c_375_n 0.0122809f $X=4.95 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A2_c_331_n N_VGND_c_529_n 0.00806659f $X=4.445 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A2_c_332_n N_VGND_c_529_n 0.00105862f $X=4.925 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A2_c_331_n N_VGND_c_532_n 0.00106058f $X=4.445 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A2_c_332_n N_VGND_c_532_n 0.00814859f $X=4.925 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A2_c_331_n N_VGND_c_533_n 0.00351072f $X=4.445 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A2_c_332_n N_VGND_c_533_n 0.0035176f $X=4.925 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A2_c_331_n N_VGND_c_536_n 0.00424612f $X=4.445 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A2_c_332_n N_VGND_c_536_n 0.00424616f $X=4.925 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A2_c_331_n N_A_525_47#_c_614_n 0.0112845f $X=4.445 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A2_c_332_n N_A_525_47#_c_614_n 0.00996055f $X=4.925 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A2_c_333_n N_A_525_47#_c_614_n 0.00662408f $X=4.935 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A2_c_353_n N_A_525_47#_c_614_n 0.0348066f $X=4.935 $Y=1.16 $X2=0 $Y2=0
cc_281 N_VPWR_c_375_n N_X_M1000_d 0.00621163f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_375_n N_X_M1010_d 0.00655879f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_M1000_s N_X_c_464_n 0.00678317f $X=0.455 $Y=1.485 $X2=0 $Y2=0
cc_284 N_VPWR_c_376_n N_X_c_464_n 0.0261645f $X=0.58 $Y=1.955 $X2=0 $Y2=0
cc_285 N_VPWR_c_384_n N_X_c_497_n 0.0131506f $X=1.375 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_375_n N_X_c_497_n 0.00722976f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_M1002_s N_X_c_475_n 0.00363854f $X=1.44 $Y=1.485 $X2=0 $Y2=0
cc_288 N_VPWR_c_377_n N_X_c_475_n 0.0209901f $X=1.59 $Y=1.955 $X2=0 $Y2=0
cc_289 N_VPWR_c_385_n N_X_c_481_n 0.0124822f $X=2.335 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_c_389_n N_X_c_481_n 0.015123f $X=2.57 $Y=2.34 $X2=0 $Y2=0
cc_291 N_VPWR_c_375_n N_X_c_481_n 0.00684987f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_292 N_VPWR_c_375_n A_826_297# 0.00284794f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_293 N_VPWR_c_375_n A_1008_297# 0.0128237f $X=5.75 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_294 N_X_c_462_n N_VGND_M1005_s 0.00301407f $X=0.22 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_295 X N_VGND_M1005_s 3.71677e-19 $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_296 N_X_c_470_n N_VGND_M1006_s 0.00427121f $X=1.7 $Y=0.71 $X2=0 $Y2=0
cc_297 N_X_c_484_n N_VGND_c_525_n 0.00167305f $X=0.645 $Y=0.71 $X2=0 $Y2=0
cc_298 N_X_c_462_n N_VGND_c_525_n 0.0209438f $X=0.22 $Y=0.805 $X2=0 $Y2=0
cc_299 N_X_c_470_n N_VGND_c_526_n 0.0181676f $X=1.7 $Y=0.71 $X2=0 $Y2=0
cc_300 N_X_c_470_n N_VGND_c_527_n 0.00772466f $X=1.7 $Y=0.71 $X2=0 $Y2=0
cc_301 N_X_c_511_p N_VGND_c_534_n 0.00669276f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_302 N_X_c_484_n N_VGND_c_534_n 0.00324423f $X=0.645 $Y=0.71 $X2=0 $Y2=0
cc_303 N_X_M1005_d N_VGND_c_536_n 0.00378648f $X=0.55 $Y=0.235 $X2=0 $Y2=0
cc_304 N_X_M1009_d N_VGND_c_536_n 0.00375928f $X=1.51 $Y=0.235 $X2=0 $Y2=0
cc_305 N_X_c_511_p N_VGND_c_536_n 0.011034f $X=0.74 $Y=0.72 $X2=0 $Y2=0
cc_306 N_X_c_470_n N_VGND_c_536_n 0.0146499f $X=1.7 $Y=0.71 $X2=0 $Y2=0
cc_307 N_X_c_484_n N_VGND_c_536_n 0.0059446f $X=0.645 $Y=0.71 $X2=0 $Y2=0
cc_308 N_X_c_462_n N_VGND_c_536_n 0.00147807f $X=0.22 $Y=0.805 $X2=0 $Y2=0
cc_309 N_VGND_c_536_n N_A_525_47#_M1013_d 0.00209344f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_310 N_VGND_c_536_n N_A_525_47#_M1015_d 0.00372626f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_311 N_VGND_c_536_n N_A_525_47#_M1003_d 0.00375928f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_536_n N_A_525_47#_M1016_d 0.0036111f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_313 N_VGND_c_528_n N_A_525_47#_c_613_n 0.0145167f $X=2.18 $Y=0.38 $X2=0 $Y2=0
cc_314 N_VGND_c_530_n N_A_525_47#_c_613_n 0.0554826f $X=4.055 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_536_n N_A_525_47#_c_613_n 0.0349279f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_M1012_s N_A_525_47#_c_614_n 0.00887205f $X=4.06 $Y=0.235 $X2=0
+ $Y2=0
cc_317 N_VGND_M1007_s N_A_525_47#_c_614_n 0.00875471f $X=5 $Y=0.235 $X2=0 $Y2=0
cc_318 N_VGND_c_529_n N_A_525_47#_c_614_n 0.0167638f $X=4.22 $Y=0.36 $X2=0 $Y2=0
cc_319 N_VGND_c_530_n N_A_525_47#_c_614_n 0.00272761f $X=4.055 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_532_n N_A_525_47#_c_614_n 0.0196989f $X=5.165 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_533_n N_A_525_47#_c_614_n 0.00939327f $X=4.975 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_535_n N_A_525_47#_c_614_n 0.00821053f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_536_n N_A_525_47#_c_614_n 0.0361194f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_324 N_VGND_c_530_n N_A_525_47#_c_618_n 0.0216097f $X=4.055 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_536_n N_A_525_47#_c_618_n 0.0125507f $X=5.75 $Y=0 $X2=0 $Y2=0
