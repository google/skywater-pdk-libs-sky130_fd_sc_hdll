* File: sky130_fd_sc_hdll__muxb16to1_4.pex.spice
* Created: Thu Aug 27 19:11:38 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VNB 9 10 11
r1126 9 11 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=25.99 $Y=4.8
+ $X2=25.99 $Y2=4.93
r1127 9 10 5.16612 $w=2.88e-07 $l=1.3e-07 $layer=LI1_cond $X=25.99 $Y=0.64
+ $X2=25.99 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPB 7 8 9 10 11 26
c742 7 0 0.00193304f $X=51.665 $Y=2.635
r743 10 11 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=25.99 $Y=3.23
+ $X2=25.99 $Y2=3.57
r744 8 9 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=25.99 $Y=1.87
+ $X2=25.99 $Y2=2.21
r745 8 26 5.56352 $w=2.88e-07 $l=1.4e-07 $layer=LI1_cond $X=25.99 $Y=1.87
+ $X2=25.99 $Y2=1.73
r746 7 10 91 $w=1.7e-07 $l=2.89396e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=25.905 $Y=3.04 $X2=25.99 $Y2=3.29
r747 7 26 91 $w=1.7e-07 $l=2.43824e-07 $layer=licon1_NTAP_notbjt $count=2
+ $X=25.905 $Y=1.525 $X2=25.99 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[0] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r90 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.905 $Y2=1.16
r91 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=1.62 $Y=1.16
+ $X2=1.88 $Y2=1.16
r92 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r93 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.46 $Y=1.16
+ $X2=1.62 $Y2=1.16
r94 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.16
+ $X2=1.46 $Y2=1.16
r95 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.965 $Y2=1.16
r96 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r97 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=1.16 $X2=0.94
+ $Y2=1.16
r98 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r99 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=1.19
+ $X2=1.62 $Y2=1.19
r100 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=1.19
+ $X2=0.94 $Y2=1.19
r101 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.16 $X2=1.28 $Y2=1.16
r102 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=0.965 $Y2=1.16
r103 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=1.28 $Y2=1.16
r104 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.435 $Y2=1.16
r105 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.28 $Y2=1.16
r106 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=0.94 $Y2=1.19
r107 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.905 $Y=1.295
+ $X2=1.905 $Y2=1.16
r108 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.905 $Y=1.295
+ $X2=1.905 $Y2=1.985
r109 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.16
r110 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r111 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.16
r112 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r113 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.16
r114 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.985
r115 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r116 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.985
r117 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.16
r118 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r119 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.16
r120 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r121 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.16
r122 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[8] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r86 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=4.28
+ $X2=1.905 $Y2=4.28
r87 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=1.62 $Y=4.28
+ $X2=1.88 $Y2=4.28
r88 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=4.28 $X2=1.62 $Y2=4.28
r89 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.46 $Y=4.28
+ $X2=1.62 $Y2=4.28
r90 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=4.28
+ $X2=1.46 $Y2=4.28
r91 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=4.28
+ $X2=0.965 $Y2=4.28
r92 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94
+ $Y=4.28 $X2=0.94 $Y2=4.28
r93 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=4.28 $X2=0.94
+ $Y2=4.28
r94 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=4.28
+ $X2=0.52 $Y2=4.28
r95 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=4.25
+ $X2=1.62 $Y2=4.25
r96 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=4.25
+ $X2=0.94 $Y2=4.25
r97 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=4.28 $X2=1.28 $Y2=4.28
r98 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=4.28
+ $X2=0.965 $Y2=4.28
r99 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=1.055 $Y=4.28
+ $X2=1.28 $Y2=4.28
r100 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.345 $Y=4.28
+ $X2=1.435 $Y2=4.28
r101 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=1.345 $Y=4.28
+ $X2=1.28 $Y2=4.28
r102 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=4.25
+ $X2=0.94 $Y2=4.25
r103 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.905 $Y=4.145
+ $X2=1.905 $Y2=4.28
r104 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.905 $Y=4.145
+ $X2=1.905 $Y2=3.455
r105 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.88 $Y=4.415
+ $X2=1.88 $Y2=4.28
r106 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=4.415
+ $X2=1.88 $Y2=4.88
r107 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.46 $Y=4.415
+ $X2=1.46 $Y2=4.28
r108 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=4.415
+ $X2=1.46 $Y2=4.88
r109 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=4.145
+ $X2=1.435 $Y2=4.28
r110 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.435 $Y=4.145
+ $X2=1.435 $Y2=3.455
r111 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=4.145
+ $X2=0.965 $Y2=4.28
r112 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=4.145
+ $X2=0.965 $Y2=3.455
r113 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=4.415
+ $X2=0.94 $Y2=4.28
r114 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=4.415
+ $X2=0.94 $Y2=4.88
r115 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=4.415
+ $X2=0.52 $Y2=4.28
r116 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=4.415
+ $X2=0.52 $Y2=4.88
r117 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=4.145
+ $X2=0.495 $Y2=4.28
r118 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=4.145
+ $X2=0.495 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c118 22 0 9.37986e-20 $X=4.305 $Y=1.475
c119 20 0 1.10627e-19 $X=4.215 $Y=1.4
c120 17 0 9.37986e-20 $X=3.835 $Y=1.475
c121 12 0 9.37986e-20 $X=3.365 $Y=1.475
c122 7 0 9.37986e-20 $X=2.895 $Y=1.475
r123 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=1.77
+ $X2=5.585 $Y2=1.605
r124 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=1.395
+ $X2=5.505 $Y2=1.23
r125 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.505 $Y=1.395
+ $X2=5.505 $Y2=1.605
r126 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=1.065
+ $X2=5.505 $Y2=1.23
r127 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.505 $Y=1.065
+ $X2=5.505 $Y2=0.825
r128 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=0.7
+ $X2=5.545 $Y2=0.825
r129 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=0.7
+ $X2=5.545 $Y2=0.445
r130 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=4.875 $Y=1.23
+ $X2=4.625 $Y2=1.23
r131 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.23 $X2=4.875 $Y2=1.23
r132 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=4.535 $Y=1.285
+ $X2=4.625 $Y2=1.23
r133 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.535 $Y=1.23
+ $X2=4.875 $Y2=1.23
r134 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.23 $X2=4.535 $Y2=1.23
r135 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=1.23
+ $X2=5.505 $Y2=1.23
r136 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=5.42 $Y=1.23
+ $X2=4.875 $Y2=1.23
r137 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.535 $Y2=1.285
r138 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.305 $Y2=1.965
r139 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.925 $Y=1.4
+ $X2=3.835 $Y2=1.4
r140 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.215 $Y=1.4
+ $X2=4.305 $Y2=1.475
r141 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.215 $Y=1.4
+ $X2=3.925 $Y2=1.4
r142 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=1.475
+ $X2=3.835 $Y2=1.4
r143 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.835 $Y=1.475
+ $X2=3.835 $Y2=1.965
r144 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=1.4
+ $X2=3.365 $Y2=1.4
r145 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.745 $Y=1.4
+ $X2=3.835 $Y2=1.4
r146 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.745 $Y=1.4
+ $X2=3.455 $Y2=1.4
r147 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.475
+ $X2=3.365 $Y2=1.4
r148 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.365 $Y=1.475
+ $X2=3.365 $Y2=1.965
r149 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.275 $Y=1.4
+ $X2=3.365 $Y2=1.4
r150 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.275 $Y=1.4
+ $X2=2.985 $Y2=1.4
r151 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.895 $Y=1.475
+ $X2=2.985 $Y2=1.4
r152 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.895 $Y=1.475
+ $X2=2.895 $Y2=1.965
r153 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.625 $X2=5.585 $Y2=1.77
r154 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.45
+ $Y=0.235 $X2=5.585 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c124 22 0 9.37986e-20 $X=4.305 $Y=3.965
c125 20 0 1.10627e-19 $X=4.215 $Y=4.04
c126 17 0 9.37986e-20 $X=3.835 $Y=3.965
c127 12 0 9.37986e-20 $X=3.365 $Y=3.965
c128 7 0 9.37986e-20 $X=2.895 $Y=3.965
r129 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=4.74
+ $X2=5.545 $Y2=4.615
r130 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=4.74
+ $X2=5.545 $Y2=4.995
r131 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=4.375
+ $X2=5.505 $Y2=4.21
r132 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.505 $Y=4.375
+ $X2=5.505 $Y2=4.615
r133 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=4.045
+ $X2=5.505 $Y2=4.21
r134 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.505 $Y=4.045
+ $X2=5.505 $Y2=3.835
r135 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=3.67
+ $X2=5.585 $Y2=3.835
r136 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=5.585 $Y=3.67
+ $X2=5.585 $Y2=3.14
r137 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=4.875 $Y=4.21
+ $X2=4.625 $Y2=4.21
r138 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=4.21 $X2=4.875 $Y2=4.21
r139 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=4.535 $Y=4.155
+ $X2=4.625 $Y2=4.21
r140 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.535 $Y=4.21
+ $X2=4.875 $Y2=4.21
r141 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=4.21 $X2=4.535 $Y2=4.21
r142 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=4.21
+ $X2=5.505 $Y2=4.21
r143 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=5.42 $Y=4.21
+ $X2=4.875 $Y2=4.21
r144 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=4.305 $Y=3.965
+ $X2=4.535 $Y2=4.155
r145 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=4.305 $Y=3.965
+ $X2=4.305 $Y2=3.475
r146 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.925 $Y=4.04
+ $X2=3.835 $Y2=4.04
r147 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.215 $Y=4.04
+ $X2=4.305 $Y2=3.965
r148 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.215 $Y=4.04
+ $X2=3.925 $Y2=4.04
r149 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=3.965
+ $X2=3.835 $Y2=4.04
r150 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.835 $Y=3.965
+ $X2=3.835 $Y2=3.475
r151 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=4.04
+ $X2=3.365 $Y2=4.04
r152 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.745 $Y=4.04
+ $X2=3.835 $Y2=4.04
r153 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.745 $Y=4.04
+ $X2=3.455 $Y2=4.04
r154 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=3.965
+ $X2=3.365 $Y2=4.04
r155 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.365 $Y=3.965
+ $X2=3.365 $Y2=3.475
r156 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.275 $Y=4.04
+ $X2=3.365 $Y2=4.04
r157 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.275 $Y=4.04
+ $X2=2.985 $Y2=4.04
r158 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.895 $Y=3.965
+ $X2=2.985 $Y2=4.04
r159 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.895 $Y=3.965
+ $X2=2.895 $Y2=3.475
r160 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=2.995 $X2=5.585 $Y2=3.14
r161 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.45
+ $Y=4.785 $X2=5.585 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[0] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c117 11 0 1.3204e-19 $X=3.66 $Y=0.255
r118 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.2
+ $Y=1.16 $X2=6.2 $Y2=1.16
r119 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=5.82 $Y=1.55
+ $X2=6.027 $Y2=1.16
r120 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.82 $Y=1.55
+ $X2=5.82 $Y2=2.035
r121 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.795 $Y=0.735
+ $X2=5.795 $Y2=0.445
r122 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.45 $Y=0.81 $X2=5.35
+ $Y2=0.81
r123 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=6.027 $Y2=1.16
r124 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=5.795 $Y2=0.735
r125 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=5.45 $Y2=0.81
r126 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=5.375 $Y=0.735
+ $X2=5.35 $Y2=0.81
r127 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.375 $Y=0.735
+ $X2=5.375 $Y2=0.445
r128 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.35 $Y=1.55
+ $X2=5.35 $Y2=2.035
r129 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.35 $Y=1.45 $X2=5.35
+ $Y2=1.55
r130 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.35 $Y=0.885
+ $X2=5.35 $Y2=0.81
r131 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=5.35 $Y=0.885
+ $X2=5.35 $Y2=1.45
r132 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.25 $Y=0.81 $X2=5.35
+ $Y2=0.81
r133 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.25 $Y=0.81
+ $X2=4.915 $Y2=0.81
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=0.735
+ $X2=4.915 $Y2=0.81
r135 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.84 $Y2=0.735
r136 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=0.18
+ $X2=4.08 $Y2=0.18
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=0.18
+ $X2=4.84 $Y2=0.255
r138 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.765 $Y=0.18
+ $X2=4.155 $Y2=0.18
r139 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.08 $Y=0.255
+ $X2=4.08 $Y2=0.18
r140 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.08 $Y=0.255
+ $X2=4.08 $Y2=0.59
r141 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=0.18
+ $X2=3.66 $Y2=0.18
r142 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.005 $Y=0.18
+ $X2=4.08 $Y2=0.18
r143 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.005 $Y=0.18
+ $X2=3.735 $Y2=0.18
r144 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.18
r145 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.59
r146 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.315 $Y=0.18
+ $X2=3.24 $Y2=0.18
r147 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.66 $Y2=0.18
r148 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.315 $Y2=0.18
r149 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.24 $Y=0.255
+ $X2=3.24 $Y2=0.18
r150 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.24 $Y=0.255
+ $X2=3.24 $Y2=0.59
r151 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=0.18
+ $X2=3.24 $Y2=0.18
r152 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.165 $Y=0.18
+ $X2=2.895 $Y2=0.18
r153 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.82 $Y=0.255
+ $X2=2.895 $Y2=0.18
r154 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.82 $Y=0.255
+ $X2=2.82 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[8] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c125 11 0 1.3204e-19 $X=3.66 $Y=5.185
r126 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.2
+ $Y=4.28 $X2=6.2 $Y2=4.28
r127 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=5.82 $Y=3.89
+ $X2=6.027 $Y2=4.28
r128 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.82 $Y=3.89
+ $X2=5.82 $Y2=3.405
r129 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.795 $Y=4.705
+ $X2=5.795 $Y2=4.995
r130 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.45 $Y=4.63 $X2=5.35
+ $Y2=4.63
r131 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.72 $Y=4.63
+ $X2=5.795 $Y2=4.705
r132 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=5.72 $Y=4.63
+ $X2=6.027 $Y2=4.28
r133 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.72 $Y=4.63
+ $X2=5.45 $Y2=4.63
r134 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=5.375 $Y=4.705
+ $X2=5.35 $Y2=4.63
r135 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.375 $Y=4.705
+ $X2=5.375 $Y2=4.995
r136 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.35 $Y=3.89
+ $X2=5.35 $Y2=3.405
r137 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.35 $Y=4.555
+ $X2=5.35 $Y2=4.63
r138 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.35 $Y=3.99 $X2=5.35
+ $Y2=3.89
r139 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=5.35 $Y=3.99
+ $X2=5.35 $Y2=4.555
r140 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.25 $Y=4.63 $X2=5.35
+ $Y2=4.63
r141 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.25 $Y=4.63
+ $X2=4.915 $Y2=4.63
r142 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=4.705
+ $X2=4.915 $Y2=4.63
r143 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.84 $Y=4.705
+ $X2=4.84 $Y2=5.185
r144 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=5.26
+ $X2=4.08 $Y2=5.26
r145 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=5.26
+ $X2=4.84 $Y2=5.185
r146 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.765 $Y=5.26
+ $X2=4.155 $Y2=5.26
r147 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.08 $Y=5.185
+ $X2=4.08 $Y2=5.26
r148 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.08 $Y=5.185
+ $X2=4.08 $Y2=4.85
r149 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=5.26
+ $X2=3.66 $Y2=5.26
r150 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.005 $Y=5.26
+ $X2=4.08 $Y2=5.26
r151 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.005 $Y=5.26
+ $X2=3.735 $Y2=5.26
r152 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=5.185
+ $X2=3.66 $Y2=5.26
r153 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.66 $Y=5.185
+ $X2=3.66 $Y2=4.85
r154 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.315 $Y=5.26
+ $X2=3.24 $Y2=5.26
r155 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=5.26
+ $X2=3.66 $Y2=5.26
r156 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.585 $Y=5.26
+ $X2=3.315 $Y2=5.26
r157 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.24 $Y=5.185
+ $X2=3.24 $Y2=5.26
r158 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.24 $Y=5.185
+ $X2=3.24 $Y2=4.85
r159 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=5.26
+ $X2=3.24 $Y2=5.26
r160 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.165 $Y=5.26
+ $X2=2.895 $Y2=5.26
r161 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.82 $Y=5.185
+ $X2=2.895 $Y2=5.26
r162 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.82 $Y=5.185
+ $X2=2.82 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[1] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c120 30 0 1.3204e-19 $X=9.22 $Y=0.255
r121 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=7.02 $Y2=1.16
r122 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.06 $Y=0.255
+ $X2=10.06 $Y2=0.59
r123 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.715 $Y=0.18
+ $X2=9.64 $Y2=0.18
r124 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=10.06 $Y2=0.255
r125 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=9.715 $Y2=0.18
r126 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.18
r127 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.59
r128 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.295 $Y=0.18
+ $X2=9.22 $Y2=0.18
r129 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.64 $Y2=0.18
r130 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.295 $Y2=0.18
r131 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.18
r132 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.59
r133 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.875 $Y=0.18
+ $X2=8.8 $Y2=0.18
r134 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=9.22 $Y2=0.18
r135 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=8.875 $Y2=0.18
r136 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.8 $Y=0.255
+ $X2=8.8 $Y2=0.18
r137 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.8 $Y=0.255
+ $X2=8.8 $Y2=0.59
r138 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.725 $Y=0.18
+ $X2=8.8 $Y2=0.18
r139 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.725 $Y=0.18
+ $X2=8.115 $Y2=0.18
r140 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.04 $Y=0.255
+ $X2=8.115 $Y2=0.18
r141 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.04 $Y=0.255
+ $X2=8.04 $Y2=0.735
r142 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.63 $Y=0.81 $X2=7.53
+ $Y2=0.81
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.965 $Y=0.81
+ $X2=8.04 $Y2=0.735
r144 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.965 $Y=0.81
+ $X2=7.63 $Y2=0.81
r145 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.53 $Y=1.55
+ $X2=7.53 $Y2=2.035
r146 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.53 $Y=1.45 $X2=7.53
+ $Y2=1.55
r147 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=7.53 $Y=0.885
+ $X2=7.53 $Y2=0.81
r148 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=7.53 $Y=0.885
+ $X2=7.53 $Y2=1.45
r149 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.505 $Y=0.735
+ $X2=7.53 $Y2=0.81
r150 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.505 $Y=0.735
+ $X2=7.505 $Y2=0.445
r151 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.16 $Y=0.81 $X2=7.06
+ $Y2=0.81
r152 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.43 $Y=0.81 $X2=7.53
+ $Y2=0.81
r153 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.43 $Y=0.81
+ $X2=7.16 $Y2=0.81
r154 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.085 $Y=0.735
+ $X2=7.06 $Y2=0.81
r155 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.085 $Y=0.735
+ $X2=7.085 $Y2=0.445
r156 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.06 $Y=1.55
+ $X2=7.06 $Y2=2.035
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=7.06 $Y=1.16
+ $X2=7.06 $Y2=1.55
r158 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.02
+ $Y=1.16 $X2=7.02 $Y2=1.16
r159 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=7.06 $Y=1.16
+ $X2=7.06 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[9] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c128 30 0 1.3204e-19 $X=9.22 $Y=5.185
r129 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.67 $Y=4.28
+ $X2=7.02 $Y2=4.28
r130 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.06 $Y=5.185
+ $X2=10.06 $Y2=4.85
r131 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.715 $Y=5.26
+ $X2=9.64 $Y2=5.26
r132 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.985 $Y=5.26
+ $X2=10.06 $Y2=5.185
r133 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.985 $Y=5.26
+ $X2=9.715 $Y2=5.26
r134 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.64 $Y=5.185
+ $X2=9.64 $Y2=5.26
r135 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.64 $Y=5.185
+ $X2=9.64 $Y2=4.85
r136 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.295 $Y=5.26
+ $X2=9.22 $Y2=5.26
r137 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.565 $Y=5.26
+ $X2=9.64 $Y2=5.26
r138 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.565 $Y=5.26
+ $X2=9.295 $Y2=5.26
r139 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=5.185
+ $X2=9.22 $Y2=5.26
r140 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.22 $Y=5.185
+ $X2=9.22 $Y2=4.85
r141 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.875 $Y=5.26
+ $X2=8.8 $Y2=5.26
r142 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=5.26
+ $X2=9.22 $Y2=5.26
r143 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.145 $Y=5.26
+ $X2=8.875 $Y2=5.26
r144 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.8 $Y=5.185
+ $X2=8.8 $Y2=5.26
r145 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.8 $Y=5.185
+ $X2=8.8 $Y2=4.85
r146 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.725 $Y=5.26
+ $X2=8.8 $Y2=5.26
r147 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.725 $Y=5.26
+ $X2=8.115 $Y2=5.26
r148 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.04 $Y=5.185
+ $X2=8.115 $Y2=5.26
r149 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.04 $Y=4.705
+ $X2=8.04 $Y2=5.185
r150 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.63 $Y=4.63 $X2=7.53
+ $Y2=4.63
r151 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.965 $Y=4.63
+ $X2=8.04 $Y2=4.705
r152 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.965 $Y=4.63
+ $X2=7.63 $Y2=4.63
r153 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.53 $Y=3.89
+ $X2=7.53 $Y2=3.405
r154 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.505 $Y=4.705
+ $X2=7.53 $Y2=4.63
r155 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.505 $Y=4.705
+ $X2=7.505 $Y2=4.995
r156 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=7.53 $Y=4.555
+ $X2=7.53 $Y2=4.63
r157 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.53 $Y=3.99 $X2=7.53
+ $Y2=3.89
r158 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=7.53 $Y=3.99
+ $X2=7.53 $Y2=4.555
r159 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.16 $Y=4.63 $X2=7.06
+ $Y2=4.63
r160 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.43 $Y=4.63 $X2=7.53
+ $Y2=4.63
r161 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.43 $Y=4.63
+ $X2=7.16 $Y2=4.63
r162 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.085 $Y=4.705
+ $X2=7.06 $Y2=4.63
r163 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.085 $Y=4.705
+ $X2=7.085 $Y2=4.995
r164 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.06 $Y=3.89
+ $X2=7.06 $Y2=3.405
r165 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=7.06 $Y=4.28
+ $X2=7.06 $Y2=4.63
r166 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.02
+ $Y=4.28 $X2=7.02 $Y2=4.28
r167 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=7.06 $Y=4.28
+ $X2=7.06 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c116 22 0 9.37986e-20 $X=9.985 $Y=1.475
c117 20 0 1.74242e-19 $X=9.895 $Y=1.4
c118 17 0 9.37986e-20 $X=9.515 $Y=1.475
c119 12 0 9.37986e-20 $X=9.045 $Y=1.475
c120 7 0 9.37986e-20 $X=8.575 $Y=1.475
r121 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=8.345 $Y=1.285
+ $X2=8.255 $Y2=1.23
r122 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.345
+ $Y=1.23 $X2=8.345 $Y2=1.23
r123 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=8.005 $Y=1.23
+ $X2=8.255 $Y2=1.23
r124 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.005 $Y=1.23
+ $X2=8.345 $Y2=1.23
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.005
+ $Y=1.23 $X2=8.005 $Y2=1.23
r126 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=1.23
+ $X2=7.375 $Y2=1.23
r127 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=7.46 $Y=1.23
+ $X2=8.005 $Y2=1.23
r128 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=1.395
+ $X2=7.375 $Y2=1.23
r129 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.375 $Y=1.395
+ $X2=7.375 $Y2=1.605
r130 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=1.065
+ $X2=7.375 $Y2=1.23
r131 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.375 $Y=1.065
+ $X2=7.375 $Y2=0.825
r132 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=0.7
+ $X2=7.335 $Y2=0.825
r133 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=0.7
+ $X2=7.335 $Y2=0.445
r134 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=1.77
+ $X2=7.295 $Y2=1.605
r135 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.985 $Y=1.475
+ $X2=9.985 $Y2=1.965
r136 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.605 $Y=1.4
+ $X2=9.515 $Y2=1.4
r137 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.895 $Y=1.4
+ $X2=9.985 $Y2=1.475
r138 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.895 $Y=1.4
+ $X2=9.605 $Y2=1.4
r139 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.515 $Y=1.475
+ $X2=9.515 $Y2=1.4
r140 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.515 $Y=1.475
+ $X2=9.515 $Y2=1.965
r141 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.135 $Y=1.4
+ $X2=9.045 $Y2=1.4
r142 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.425 $Y=1.4
+ $X2=9.515 $Y2=1.4
r143 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.425 $Y=1.4
+ $X2=9.135 $Y2=1.4
r144 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.045 $Y=1.475
+ $X2=9.045 $Y2=1.4
r145 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.045 $Y=1.475
+ $X2=9.045 $Y2=1.965
r146 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.955 $Y=1.4
+ $X2=9.045 $Y2=1.4
r147 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.955 $Y=1.4
+ $X2=8.665 $Y2=1.4
r148 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.665 $Y2=1.4
r149 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.345 $Y2=1.285
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.575 $Y2=1.965
r151 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.15
+ $Y=1.625 $X2=7.295 $Y2=1.77
r152 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.235 $X2=7.295 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_599# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c122 22 0 9.37986e-20 $X=9.985 $Y=3.965
c123 20 0 1.74242e-19 $X=9.895 $Y=4.04
c124 17 0 9.37986e-20 $X=9.515 $Y=3.965
c125 12 0 9.37986e-20 $X=9.045 $Y=3.965
c126 7 0 9.37986e-20 $X=8.575 $Y=3.965
r127 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=8.345 $Y=4.155
+ $X2=8.255 $Y2=4.21
r128 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.345
+ $Y=4.21 $X2=8.345 $Y2=4.21
r129 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=8.005 $Y=4.21
+ $X2=8.255 $Y2=4.21
r130 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.005 $Y=4.21
+ $X2=8.345 $Y2=4.21
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.005
+ $Y=4.21 $X2=8.005 $Y2=4.21
r132 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=4.21
+ $X2=7.375 $Y2=4.21
r133 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=7.46 $Y=4.21
+ $X2=8.005 $Y2=4.21
r134 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=4.375
+ $X2=7.375 $Y2=4.21
r135 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.375 $Y=4.375
+ $X2=7.375 $Y2=4.615
r136 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=4.045
+ $X2=7.375 $Y2=4.21
r137 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.375 $Y=4.045
+ $X2=7.375 $Y2=3.835
r138 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=4.74
+ $X2=7.335 $Y2=4.615
r139 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=4.74
+ $X2=7.335 $Y2=4.995
r140 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=3.67
+ $X2=7.295 $Y2=3.835
r141 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=7.295 $Y=3.67
+ $X2=7.295 $Y2=3.14
r142 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.985 $Y=3.965
+ $X2=9.985 $Y2=3.475
r143 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.605 $Y=4.04
+ $X2=9.515 $Y2=4.04
r144 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.895 $Y=4.04
+ $X2=9.985 $Y2=3.965
r145 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.895 $Y=4.04
+ $X2=9.605 $Y2=4.04
r146 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.515 $Y=3.965
+ $X2=9.515 $Y2=4.04
r147 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.515 $Y=3.965
+ $X2=9.515 $Y2=3.475
r148 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.135 $Y=4.04
+ $X2=9.045 $Y2=4.04
r149 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.425 $Y=4.04
+ $X2=9.515 $Y2=4.04
r150 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.425 $Y=4.04
+ $X2=9.135 $Y2=4.04
r151 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.045 $Y=3.965
+ $X2=9.045 $Y2=4.04
r152 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.045 $Y=3.965
+ $X2=9.045 $Y2=3.475
r153 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.955 $Y=4.04
+ $X2=9.045 $Y2=4.04
r154 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.955 $Y=4.04
+ $X2=8.665 $Y2=4.04
r155 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.575 $Y=3.965
+ $X2=8.665 $Y2=4.04
r156 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=8.575 $Y=3.965
+ $X2=8.345 $Y2=4.155
r157 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=8.575 $Y=3.965
+ $X2=8.575 $Y2=3.475
r158 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.15
+ $Y=2.995 $X2=7.295 $Y2=3.14
r159 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=4.785 $X2=7.295 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[1] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r93 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=1.16
+ $X2=12.385 $Y2=1.16
r94 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=12.28 $Y=1.16
+ $X2=12.36 $Y2=1.16
r95 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.28
+ $Y=1.16 $X2=12.28 $Y2=1.16
r96 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=11.94 $Y=1.16
+ $X2=12.28 $Y2=1.16
r97 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=1.16
+ $X2=11.94 $Y2=1.16
r98 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.42 $Y=1.16
+ $X2=11.445 $Y2=1.16
r99 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=11.26 $Y=1.16
+ $X2=11.42 $Y2=1.16
r100 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=1.16 $X2=11.26 $Y2=1.16
r101 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=11 $Y=1.16
+ $X2=11.26 $Y2=1.16
r102 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.975 $Y=1.16
+ $X2=11 $Y2=1.16
r103 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.6 $Y=1.19
+ $X2=11.26 $Y2=1.19
r104 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.6
+ $Y=1.16 $X2=11.6 $Y2=1.16
r105 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.535 $Y=1.16
+ $X2=11.445 $Y2=1.16
r106 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=11.535 $Y=1.16
+ $X2=11.6 $Y2=1.16
r107 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.825 $Y=1.16
+ $X2=11.915 $Y2=1.16
r108 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=11.825 $Y=1.16
+ $X2=11.6 $Y2=1.16
r109 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=12.19 $Y=1.19
+ $X2=12.28 $Y2=1.19
r110 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.19 $Y=1.19
+ $X2=11.6 $Y2=1.19
r111 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.16
r112 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.985
r113 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=1.16
r114 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=0.56
r115 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=1.16
r116 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=0.56
r117 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.16
r118 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.985
r119 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.445 $Y=1.295
+ $X2=11.445 $Y2=1.16
r120 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.445 $Y=1.295
+ $X2=11.445 $Y2=1.985
r121 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.42 $Y=1.025
+ $X2=11.42 $Y2=1.16
r122 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.42 $Y=1.025
+ $X2=11.42 $Y2=0.56
r123 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11 $Y=1.025 $X2=11
+ $Y2=1.16
r124 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11 $Y=1.025 $X2=11
+ $Y2=0.56
r125 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.975 $Y=1.295
+ $X2=10.975 $Y2=1.16
r126 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=10.975 $Y=1.295
+ $X2=10.975 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[9] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r91 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=4.28
+ $X2=12.385 $Y2=4.28
r92 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=12.28 $Y=4.28
+ $X2=12.36 $Y2=4.28
r93 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.28
+ $Y=4.28 $X2=12.28 $Y2=4.28
r94 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=11.94 $Y=4.28
+ $X2=12.28 $Y2=4.28
r95 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=4.28
+ $X2=11.94 $Y2=4.28
r96 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.42 $Y=4.28
+ $X2=11.445 $Y2=4.28
r97 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=11.26 $Y=4.28
+ $X2=11.42 $Y2=4.28
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=4.28 $X2=11.26 $Y2=4.28
r99 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=11 $Y=4.28 $X2=11.26
+ $Y2=4.28
r100 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.975 $Y=4.28
+ $X2=11 $Y2=4.28
r101 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.6 $Y=4.25
+ $X2=11.26 $Y2=4.25
r102 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.6
+ $Y=4.28 $X2=11.6 $Y2=4.28
r103 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.535 $Y=4.28
+ $X2=11.445 $Y2=4.28
r104 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=11.535 $Y=4.28
+ $X2=11.6 $Y2=4.28
r105 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.825 $Y=4.28
+ $X2=11.915 $Y2=4.28
r106 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=11.825 $Y=4.28
+ $X2=11.6 $Y2=4.28
r107 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=12.19 $Y=4.25
+ $X2=12.28 $Y2=4.25
r108 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.19 $Y=4.25
+ $X2=11.6 $Y2=4.25
r109 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=4.145
+ $X2=12.385 $Y2=4.28
r110 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=4.145
+ $X2=12.385 $Y2=3.455
r111 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=4.415
+ $X2=12.36 $Y2=4.28
r112 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=4.415
+ $X2=12.36 $Y2=4.88
r113 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=4.415
+ $X2=11.94 $Y2=4.28
r114 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=4.415
+ $X2=11.94 $Y2=4.88
r115 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=4.145
+ $X2=11.915 $Y2=4.28
r116 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=4.145
+ $X2=11.915 $Y2=3.455
r117 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.445 $Y=4.145
+ $X2=11.445 $Y2=4.28
r118 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.445 $Y=4.145
+ $X2=11.445 $Y2=3.455
r119 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.42 $Y=4.415
+ $X2=11.42 $Y2=4.28
r120 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.42 $Y=4.415
+ $X2=11.42 $Y2=4.88
r121 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11 $Y=4.415 $X2=11
+ $Y2=4.28
r122 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11 $Y=4.415 $X2=11
+ $Y2=4.88
r123 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.975 $Y=4.145
+ $X2=10.975 $Y2=4.28
r124 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=10.975 $Y=4.145
+ $X2=10.975 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[2] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r95 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.76 $Y=1.16
+ $X2=14.785 $Y2=1.16
r96 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=14.5 $Y=1.16
+ $X2=14.76 $Y2=1.16
r97 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.5
+ $Y=1.16 $X2=14.5 $Y2=1.16
r98 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=14.34 $Y=1.16
+ $X2=14.5 $Y2=1.16
r99 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.315 $Y=1.16
+ $X2=14.34 $Y2=1.16
r100 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=1.16
+ $X2=13.845 $Y2=1.16
r101 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.82
+ $Y=1.16 $X2=13.82 $Y2=1.16
r102 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=13.4 $Y=1.16
+ $X2=13.82 $Y2=1.16
r103 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=1.16
+ $X2=13.4 $Y2=1.16
r104 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=1.19
+ $X2=14.5 $Y2=1.19
r105 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=1.19
+ $X2=13.82 $Y2=1.19
r106 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.16
+ $Y=1.16 $X2=14.16 $Y2=1.16
r107 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=13.935 $Y=1.16
+ $X2=13.845 $Y2=1.16
r108 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=13.935 $Y=1.16
+ $X2=14.16 $Y2=1.16
r109 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=14.225 $Y=1.16
+ $X2=14.315 $Y2=1.16
r110 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=14.225 $Y=1.16
+ $X2=14.16 $Y2=1.16
r111 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.57 $Y=1.19
+ $X2=13.82 $Y2=1.19
r112 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.785 $Y=1.295
+ $X2=14.785 $Y2=1.16
r113 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.785 $Y=1.295
+ $X2=14.785 $Y2=1.985
r114 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.76 $Y=1.025
+ $X2=14.76 $Y2=1.16
r115 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.76 $Y=1.025
+ $X2=14.76 $Y2=0.56
r116 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.34 $Y=1.025
+ $X2=14.34 $Y2=1.16
r117 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.34 $Y=1.025
+ $X2=14.34 $Y2=0.56
r118 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.315 $Y=1.295
+ $X2=14.315 $Y2=1.16
r119 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.315 $Y=1.295
+ $X2=14.315 $Y2=1.985
r120 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.16
r121 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.985
r122 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=1.16
r123 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=0.56
r124 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=1.16
r125 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=0.56
r126 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.16
r127 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[10] 3 7 11 15 19 23 27 31 33 35 36
+ 51 53
r91 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.76 $Y=4.28
+ $X2=14.785 $Y2=4.28
r92 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=14.5 $Y=4.28
+ $X2=14.76 $Y2=4.28
r93 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.5
+ $Y=4.28 $X2=14.5 $Y2=4.28
r94 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=14.34 $Y=4.28
+ $X2=14.5 $Y2=4.28
r95 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.315 $Y=4.28
+ $X2=14.34 $Y2=4.28
r96 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=4.28
+ $X2=13.845 $Y2=4.28
r97 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.82
+ $Y=4.28 $X2=13.82 $Y2=4.28
r98 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=13.4 $Y=4.28
+ $X2=13.82 $Y2=4.28
r99 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=4.28
+ $X2=13.4 $Y2=4.28
r100 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=4.25
+ $X2=14.5 $Y2=4.25
r101 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=4.25
+ $X2=13.82 $Y2=4.25
r102 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.16
+ $Y=4.28 $X2=14.16 $Y2=4.28
r103 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=13.935 $Y=4.28
+ $X2=13.845 $Y2=4.28
r104 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=13.935 $Y=4.28
+ $X2=14.16 $Y2=4.28
r105 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=14.225 $Y=4.28
+ $X2=14.315 $Y2=4.28
r106 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=14.225 $Y=4.28
+ $X2=14.16 $Y2=4.28
r107 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.57 $Y=4.25
+ $X2=13.82 $Y2=4.25
r108 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.785 $Y=4.145
+ $X2=14.785 $Y2=4.28
r109 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.785 $Y=4.145
+ $X2=14.785 $Y2=3.455
r110 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.76 $Y=4.415
+ $X2=14.76 $Y2=4.28
r111 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.76 $Y=4.415
+ $X2=14.76 $Y2=4.88
r112 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.34 $Y=4.415
+ $X2=14.34 $Y2=4.28
r113 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.34 $Y=4.415
+ $X2=14.34 $Y2=4.88
r114 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.315 $Y=4.145
+ $X2=14.315 $Y2=4.28
r115 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.315 $Y=4.145
+ $X2=14.315 $Y2=3.455
r116 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=4.145
+ $X2=13.845 $Y2=4.28
r117 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=4.145
+ $X2=13.845 $Y2=3.455
r118 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=4.415
+ $X2=13.82 $Y2=4.28
r119 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=4.415
+ $X2=13.82 $Y2=4.88
r120 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=4.415
+ $X2=13.4 $Y2=4.28
r121 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=4.415
+ $X2=13.4 $Y2=4.88
r122 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=4.145
+ $X2=13.375 $Y2=4.28
r123 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=4.145
+ $X2=13.375 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c119 22 0 9.37986e-20 $X=17.185 $Y=1.475
c120 20 0 1.10627e-19 $X=17.095 $Y=1.4
c121 17 0 9.37986e-20 $X=16.715 $Y=1.475
c122 12 0 9.37986e-20 $X=16.245 $Y=1.475
c123 11 0 1.74242e-19 $X=15.865 $Y=1.4
c124 7 0 9.37986e-20 $X=15.775 $Y=1.475
r125 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=1.77
+ $X2=18.465 $Y2=1.605
r126 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=1.395
+ $X2=18.385 $Y2=1.23
r127 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=18.385 $Y=1.395
+ $X2=18.385 $Y2=1.605
r128 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=1.065
+ $X2=18.385 $Y2=1.23
r129 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=18.385 $Y=1.065
+ $X2=18.385 $Y2=0.825
r130 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=18.425 $Y=0.7
+ $X2=18.425 $Y2=0.825
r131 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=18.425 $Y=0.7
+ $X2=18.425 $Y2=0.445
r132 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=17.755 $Y=1.23
+ $X2=17.505 $Y2=1.23
r133 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.755
+ $Y=1.23 $X2=17.755 $Y2=1.23
r134 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=17.415
+ $Y=1.285 $X2=17.505 $Y2=1.23
r135 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=17.415 $Y=1.23
+ $X2=17.755 $Y2=1.23
r136 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.415
+ $Y=1.23 $X2=17.415 $Y2=1.23
r137 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.3 $Y=1.23
+ $X2=18.385 $Y2=1.23
r138 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=18.3 $Y=1.23
+ $X2=17.755 $Y2=1.23
r139 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=17.185
+ $Y=1.475 $X2=17.415 $Y2=1.285
r140 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=17.185 $Y=1.475
+ $X2=17.185 $Y2=1.965
r141 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.805 $Y=1.4
+ $X2=16.715 $Y2=1.4
r142 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.095 $Y=1.4
+ $X2=17.185 $Y2=1.475
r143 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.095 $Y=1.4
+ $X2=16.805 $Y2=1.4
r144 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.715 $Y=1.475
+ $X2=16.715 $Y2=1.4
r145 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.715 $Y=1.475
+ $X2=16.715 $Y2=1.965
r146 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.335 $Y=1.4
+ $X2=16.245 $Y2=1.4
r147 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.625 $Y=1.4
+ $X2=16.715 $Y2=1.4
r148 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.625 $Y=1.4
+ $X2=16.335 $Y2=1.4
r149 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.245 $Y=1.475
+ $X2=16.245 $Y2=1.4
r150 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.245 $Y=1.475
+ $X2=16.245 $Y2=1.965
r151 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.155 $Y=1.4
+ $X2=16.245 $Y2=1.4
r152 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.155 $Y=1.4
+ $X2=15.865 $Y2=1.4
r153 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=15.775 $Y=1.475
+ $X2=15.865 $Y2=1.4
r154 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.775 $Y=1.475
+ $X2=15.775 $Y2=1.965
r155 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.32
+ $Y=1.625 $X2=18.465 $Y2=1.77
r156 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.33
+ $Y=0.235 $X2=18.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c125 22 0 9.37986e-20 $X=17.185 $Y=3.965
c126 20 0 1.10627e-19 $X=17.095 $Y=4.04
c127 17 0 9.37986e-20 $X=16.715 $Y=3.965
c128 12 0 9.37986e-20 $X=16.245 $Y=3.965
c129 11 0 1.74242e-19 $X=15.865 $Y=4.04
c130 7 0 9.37986e-20 $X=15.775 $Y=3.965
r131 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=18.425 $Y=4.74
+ $X2=18.425 $Y2=4.615
r132 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=18.425 $Y=4.74
+ $X2=18.425 $Y2=4.995
r133 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=4.375
+ $X2=18.385 $Y2=4.21
r134 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=18.385 $Y=4.375
+ $X2=18.385 $Y2=4.615
r135 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=4.045
+ $X2=18.385 $Y2=4.21
r136 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=18.385 $Y=4.045
+ $X2=18.385 $Y2=3.835
r137 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=3.67
+ $X2=18.465 $Y2=3.835
r138 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=18.465 $Y=3.67
+ $X2=18.465 $Y2=3.14
r139 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=17.755 $Y=4.21
+ $X2=17.505 $Y2=4.21
r140 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.755
+ $Y=4.21 $X2=17.755 $Y2=4.21
r141 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=17.415
+ $Y=4.155 $X2=17.505 $Y2=4.21
r142 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=17.415 $Y=4.21
+ $X2=17.755 $Y2=4.21
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.415
+ $Y=4.21 $X2=17.415 $Y2=4.21
r144 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.3 $Y=4.21
+ $X2=18.385 $Y2=4.21
r145 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=18.3 $Y=4.21
+ $X2=17.755 $Y2=4.21
r146 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=17.185
+ $Y=3.965 $X2=17.415 $Y2=4.155
r147 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=17.185 $Y=3.965
+ $X2=17.185 $Y2=3.475
r148 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.805 $Y=4.04
+ $X2=16.715 $Y2=4.04
r149 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.095 $Y=4.04
+ $X2=17.185 $Y2=3.965
r150 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.095 $Y=4.04
+ $X2=16.805 $Y2=4.04
r151 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.715 $Y=3.965
+ $X2=16.715 $Y2=4.04
r152 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.715 $Y=3.965
+ $X2=16.715 $Y2=3.475
r153 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.335 $Y=4.04
+ $X2=16.245 $Y2=4.04
r154 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.625 $Y=4.04
+ $X2=16.715 $Y2=4.04
r155 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.625 $Y=4.04
+ $X2=16.335 $Y2=4.04
r156 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.245 $Y=3.965
+ $X2=16.245 $Y2=4.04
r157 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.245 $Y=3.965
+ $X2=16.245 $Y2=3.475
r158 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.155 $Y=4.04
+ $X2=16.245 $Y2=4.04
r159 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.155 $Y=4.04
+ $X2=15.865 $Y2=4.04
r160 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=15.775 $Y=3.965
+ $X2=15.865 $Y2=4.04
r161 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.775 $Y=3.965
+ $X2=15.775 $Y2=3.475
r162 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.32
+ $Y=2.995 $X2=18.465 $Y2=3.14
r163 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.33
+ $Y=4.785 $X2=18.465 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[2] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c117 11 0 1.3204e-19 $X=16.54 $Y=0.255
r118 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.08
+ $Y=1.16 $X2=19.08 $Y2=1.16
r119 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=18.7 $Y=1.55
+ $X2=18.907 $Y2=1.16
r120 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.7 $Y=1.55
+ $X2=18.7 $Y2=2.035
r121 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.675 $Y=0.735
+ $X2=18.675 $Y2=0.445
r122 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.33 $Y=0.81
+ $X2=18.23 $Y2=0.81
r123 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.907 $Y2=1.16
r124 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.675 $Y2=0.735
r125 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.33 $Y2=0.81
r126 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=18.255 $Y=0.735
+ $X2=18.23 $Y2=0.81
r127 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.255 $Y=0.735
+ $X2=18.255 $Y2=0.445
r128 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.23 $Y=1.55
+ $X2=18.23 $Y2=2.035
r129 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=18.23 $Y=1.45 $X2=18.23
+ $Y2=1.55
r130 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=18.23 $Y=0.885
+ $X2=18.23 $Y2=0.81
r131 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=18.23 $Y=0.885
+ $X2=18.23 $Y2=1.45
r132 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.13 $Y=0.81
+ $X2=18.23 $Y2=0.81
r133 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=18.13 $Y=0.81
+ $X2=17.795 $Y2=0.81
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.72 $Y=0.735
+ $X2=17.795 $Y2=0.81
r135 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.72 $Y=0.255
+ $X2=17.72 $Y2=0.735
r136 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.035 $Y=0.18
+ $X2=16.96 $Y2=0.18
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.645 $Y=0.18
+ $X2=17.72 $Y2=0.255
r138 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=17.645 $Y=0.18
+ $X2=17.035 $Y2=0.18
r139 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.96 $Y=0.255
+ $X2=16.96 $Y2=0.18
r140 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.96 $Y=0.255
+ $X2=16.96 $Y2=0.59
r141 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.615 $Y=0.18
+ $X2=16.54 $Y2=0.18
r142 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.885 $Y=0.18
+ $X2=16.96 $Y2=0.18
r143 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.885 $Y=0.18
+ $X2=16.615 $Y2=0.18
r144 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.54 $Y=0.255
+ $X2=16.54 $Y2=0.18
r145 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.54 $Y=0.255
+ $X2=16.54 $Y2=0.59
r146 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.195 $Y=0.18
+ $X2=16.12 $Y2=0.18
r147 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.465 $Y=0.18
+ $X2=16.54 $Y2=0.18
r148 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.465 $Y=0.18
+ $X2=16.195 $Y2=0.18
r149 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.12 $Y=0.255
+ $X2=16.12 $Y2=0.18
r150 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.12 $Y=0.255
+ $X2=16.12 $Y2=0.59
r151 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.045 $Y=0.18
+ $X2=16.12 $Y2=0.18
r152 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.045 $Y=0.18
+ $X2=15.775 $Y2=0.18
r153 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.7 $Y=0.255
+ $X2=15.775 $Y2=0.18
r154 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.7 $Y=0.255
+ $X2=15.7 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[10] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c125 11 0 1.3204e-19 $X=16.54 $Y=5.185
r126 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.08
+ $Y=4.28 $X2=19.08 $Y2=4.28
r127 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=18.7 $Y=3.89
+ $X2=18.907 $Y2=4.28
r128 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.7 $Y=3.89
+ $X2=18.7 $Y2=3.405
r129 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.675 $Y=4.705
+ $X2=18.675 $Y2=4.995
r130 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.33 $Y=4.63
+ $X2=18.23 $Y2=4.63
r131 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=18.6 $Y=4.63
+ $X2=18.675 $Y2=4.705
r132 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=18.6 $Y=4.63
+ $X2=18.907 $Y2=4.28
r133 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=18.6 $Y=4.63
+ $X2=18.33 $Y2=4.63
r134 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=18.255 $Y=4.705
+ $X2=18.23 $Y2=4.63
r135 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.255 $Y=4.705
+ $X2=18.255 $Y2=4.995
r136 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.23 $Y=3.89
+ $X2=18.23 $Y2=3.405
r137 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=18.23 $Y=4.555
+ $X2=18.23 $Y2=4.63
r138 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=18.23 $Y=3.99 $X2=18.23
+ $Y2=3.89
r139 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=18.23 $Y=3.99
+ $X2=18.23 $Y2=4.555
r140 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.13 $Y=4.63
+ $X2=18.23 $Y2=4.63
r141 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=18.13 $Y=4.63
+ $X2=17.795 $Y2=4.63
r142 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.72 $Y=4.705
+ $X2=17.795 $Y2=4.63
r143 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.72 $Y=4.705
+ $X2=17.72 $Y2=5.185
r144 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.035 $Y=5.26
+ $X2=16.96 $Y2=5.26
r145 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.645 $Y=5.26
+ $X2=17.72 $Y2=5.185
r146 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=17.645 $Y=5.26
+ $X2=17.035 $Y2=5.26
r147 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.96 $Y=5.185
+ $X2=16.96 $Y2=5.26
r148 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.96 $Y=5.185
+ $X2=16.96 $Y2=4.85
r149 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.615 $Y=5.26
+ $X2=16.54 $Y2=5.26
r150 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.885 $Y=5.26
+ $X2=16.96 $Y2=5.26
r151 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.885 $Y=5.26
+ $X2=16.615 $Y2=5.26
r152 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.54 $Y=5.185
+ $X2=16.54 $Y2=5.26
r153 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.54 $Y=5.185
+ $X2=16.54 $Y2=4.85
r154 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.195 $Y=5.26
+ $X2=16.12 $Y2=5.26
r155 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.465 $Y=5.26
+ $X2=16.54 $Y2=5.26
r156 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.465 $Y=5.26
+ $X2=16.195 $Y2=5.26
r157 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.12 $Y=5.185
+ $X2=16.12 $Y2=5.26
r158 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.12 $Y=5.185
+ $X2=16.12 $Y2=4.85
r159 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.045 $Y=5.26
+ $X2=16.12 $Y2=5.26
r160 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.045 $Y=5.26
+ $X2=15.775 $Y2=5.26
r161 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.7 $Y=5.185
+ $X2=15.775 $Y2=5.26
r162 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.7 $Y=5.185
+ $X2=15.7 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[3] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c120 30 0 1.3204e-19 $X=22.1 $Y=0.255
r121 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=19.55 $Y=1.16
+ $X2=19.9 $Y2=1.16
r122 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.94 $Y=0.255
+ $X2=22.94 $Y2=0.59
r123 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.595 $Y=0.18
+ $X2=22.52 $Y2=0.18
r124 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=22.865 $Y=0.18
+ $X2=22.94 $Y2=0.255
r125 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.865 $Y=0.18
+ $X2=22.595 $Y2=0.18
r126 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.52 $Y=0.255
+ $X2=22.52 $Y2=0.18
r127 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.52 $Y=0.255
+ $X2=22.52 $Y2=0.59
r128 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.175 $Y=0.18
+ $X2=22.1 $Y2=0.18
r129 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.445 $Y=0.18
+ $X2=22.52 $Y2=0.18
r130 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.445 $Y=0.18
+ $X2=22.175 $Y2=0.18
r131 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.1 $Y=0.255
+ $X2=22.1 $Y2=0.18
r132 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.1 $Y=0.255
+ $X2=22.1 $Y2=0.59
r133 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.755 $Y=0.18
+ $X2=21.68 $Y2=0.18
r134 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.025 $Y=0.18
+ $X2=22.1 $Y2=0.18
r135 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.025 $Y=0.18
+ $X2=21.755 $Y2=0.18
r136 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.68 $Y=0.255
+ $X2=21.68 $Y2=0.18
r137 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.68 $Y=0.255
+ $X2=21.68 $Y2=0.59
r138 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.605 $Y=0.18
+ $X2=21.68 $Y2=0.18
r139 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=21.605 $Y=0.18
+ $X2=20.995 $Y2=0.18
r140 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.92 $Y=0.255
+ $X2=20.995 $Y2=0.18
r141 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=20.92 $Y=0.255
+ $X2=20.92 $Y2=0.735
r142 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.51 $Y=0.81
+ $X2=20.41 $Y2=0.81
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.845 $Y=0.81
+ $X2=20.92 $Y2=0.735
r144 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=20.845 $Y=0.81
+ $X2=20.51 $Y2=0.81
r145 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=20.41 $Y=1.55
+ $X2=20.41 $Y2=2.035
r146 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=20.41 $Y=1.45 $X2=20.41
+ $Y2=1.55
r147 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=20.41 $Y=0.885
+ $X2=20.41 $Y2=0.81
r148 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=20.41 $Y=0.885
+ $X2=20.41 $Y2=1.45
r149 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=20.385 $Y=0.735
+ $X2=20.41 $Y2=0.81
r150 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=20.385 $Y=0.735
+ $X2=20.385 $Y2=0.445
r151 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.04 $Y=0.81
+ $X2=19.94 $Y2=0.81
r152 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.31 $Y=0.81
+ $X2=20.41 $Y2=0.81
r153 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=20.31 $Y=0.81
+ $X2=20.04 $Y2=0.81
r154 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=19.965 $Y=0.735
+ $X2=19.94 $Y2=0.81
r155 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=19.965 $Y=0.735
+ $X2=19.965 $Y2=0.445
r156 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=19.94 $Y=1.55
+ $X2=19.94 $Y2=2.035
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=19.94 $Y=1.16
+ $X2=19.94 $Y2=1.55
r158 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.9
+ $Y=1.16 $X2=19.9 $Y2=1.16
r159 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=19.94 $Y=1.16
+ $X2=19.94 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[11] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c128 30 0 1.3204e-19 $X=22.1 $Y=5.185
r129 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=19.55 $Y=4.28
+ $X2=19.9 $Y2=4.28
r130 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.94 $Y=5.185
+ $X2=22.94 $Y2=4.85
r131 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.595 $Y=5.26
+ $X2=22.52 $Y2=5.26
r132 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=22.865 $Y=5.26
+ $X2=22.94 $Y2=5.185
r133 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.865 $Y=5.26
+ $X2=22.595 $Y2=5.26
r134 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.52 $Y=5.185
+ $X2=22.52 $Y2=5.26
r135 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.52 $Y=5.185
+ $X2=22.52 $Y2=4.85
r136 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.175 $Y=5.26
+ $X2=22.1 $Y2=5.26
r137 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.445 $Y=5.26
+ $X2=22.52 $Y2=5.26
r138 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.445 $Y=5.26
+ $X2=22.175 $Y2=5.26
r139 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.1 $Y=5.185
+ $X2=22.1 $Y2=5.26
r140 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.1 $Y=5.185
+ $X2=22.1 $Y2=4.85
r141 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.755 $Y=5.26
+ $X2=21.68 $Y2=5.26
r142 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.025 $Y=5.26
+ $X2=22.1 $Y2=5.26
r143 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.025 $Y=5.26
+ $X2=21.755 $Y2=5.26
r144 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.68 $Y=5.185
+ $X2=21.68 $Y2=5.26
r145 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.68 $Y=5.185
+ $X2=21.68 $Y2=4.85
r146 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.605 $Y=5.26
+ $X2=21.68 $Y2=5.26
r147 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=21.605 $Y=5.26
+ $X2=20.995 $Y2=5.26
r148 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.92 $Y=5.185
+ $X2=20.995 $Y2=5.26
r149 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=20.92 $Y=4.705
+ $X2=20.92 $Y2=5.185
r150 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.51 $Y=4.63
+ $X2=20.41 $Y2=4.63
r151 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.845 $Y=4.63
+ $X2=20.92 $Y2=4.705
r152 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=20.845 $Y=4.63
+ $X2=20.51 $Y2=4.63
r153 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=20.41 $Y=3.89
+ $X2=20.41 $Y2=3.405
r154 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=20.385 $Y=4.705
+ $X2=20.41 $Y2=4.63
r155 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=20.385 $Y=4.705
+ $X2=20.385 $Y2=4.995
r156 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=20.41 $Y=4.555
+ $X2=20.41 $Y2=4.63
r157 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=20.41 $Y=3.99 $X2=20.41
+ $Y2=3.89
r158 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=20.41 $Y=3.99
+ $X2=20.41 $Y2=4.555
r159 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.04 $Y=4.63
+ $X2=19.94 $Y2=4.63
r160 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.31 $Y=4.63
+ $X2=20.41 $Y2=4.63
r161 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=20.31 $Y=4.63
+ $X2=20.04 $Y2=4.63
r162 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=19.965 $Y=4.705
+ $X2=19.94 $Y2=4.63
r163 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=19.965 $Y=4.705
+ $X2=19.965 $Y2=4.995
r164 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=19.94 $Y=3.89
+ $X2=19.94 $Y2=3.405
r165 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=19.94 $Y=4.28
+ $X2=19.94 $Y2=4.63
r166 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.9
+ $Y=4.28 $X2=19.9 $Y2=4.28
r167 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=19.94 $Y=4.28
+ $X2=19.94 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c116 22 0 9.37986e-20 $X=22.865 $Y=1.475
c117 20 0 1.74242e-19 $X=22.775 $Y=1.4
c118 17 0 9.37986e-20 $X=22.395 $Y=1.475
c119 12 0 9.37986e-20 $X=21.925 $Y=1.475
c120 7 0 9.37986e-20 $X=21.455 $Y=1.475
r121 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=21.225
+ $Y=1.285 $X2=21.135 $Y2=1.23
r122 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.225
+ $Y=1.23 $X2=21.225 $Y2=1.23
r123 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=20.885 $Y=1.23
+ $X2=21.135 $Y2=1.23
r124 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=20.885 $Y=1.23
+ $X2=21.225 $Y2=1.23
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.885
+ $Y=1.23 $X2=20.885 $Y2=1.23
r126 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.34 $Y=1.23
+ $X2=20.255 $Y2=1.23
r127 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=20.34 $Y=1.23
+ $X2=20.885 $Y2=1.23
r128 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=1.395
+ $X2=20.255 $Y2=1.23
r129 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=20.255 $Y=1.395
+ $X2=20.255 $Y2=1.605
r130 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=1.065
+ $X2=20.255 $Y2=1.23
r131 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=20.255 $Y=1.065
+ $X2=20.255 $Y2=0.825
r132 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=20.215 $Y=0.7
+ $X2=20.215 $Y2=0.825
r133 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=20.215 $Y=0.7
+ $X2=20.215 $Y2=0.445
r134 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.175 $Y=1.77
+ $X2=20.175 $Y2=1.605
r135 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.865 $Y=1.475
+ $X2=22.865 $Y2=1.965
r136 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.485 $Y=1.4
+ $X2=22.395 $Y2=1.4
r137 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=22.775 $Y=1.4
+ $X2=22.865 $Y2=1.475
r138 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.775 $Y=1.4
+ $X2=22.485 $Y2=1.4
r139 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=22.395 $Y=1.475
+ $X2=22.395 $Y2=1.4
r140 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.395 $Y=1.475
+ $X2=22.395 $Y2=1.965
r141 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.015 $Y=1.4
+ $X2=21.925 $Y2=1.4
r142 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.305 $Y=1.4
+ $X2=22.395 $Y2=1.4
r143 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.305 $Y=1.4
+ $X2=22.015 $Y2=1.4
r144 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=21.925 $Y=1.475
+ $X2=21.925 $Y2=1.4
r145 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.925 $Y=1.475
+ $X2=21.925 $Y2=1.965
r146 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.835 $Y=1.4
+ $X2=21.925 $Y2=1.4
r147 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.835 $Y=1.4
+ $X2=21.545 $Y2=1.4
r148 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.545 $Y2=1.4
r149 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.225 $Y2=1.285
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.455 $Y2=1.965
r151 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.03
+ $Y=1.625 $X2=20.175 $Y2=1.77
r152 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.04
+ $Y=0.235 $X2=20.175 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_599# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c122 22 0 9.37986e-20 $X=22.865 $Y=3.965
c123 20 0 1.74242e-19 $X=22.775 $Y=4.04
c124 17 0 9.37986e-20 $X=22.395 $Y=3.965
c125 12 0 9.37986e-20 $X=21.925 $Y=3.965
c126 7 0 9.37986e-20 $X=21.455 $Y=3.965
r127 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=21.225
+ $Y=4.155 $X2=21.135 $Y2=4.21
r128 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.225
+ $Y=4.21 $X2=21.225 $Y2=4.21
r129 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=20.885 $Y=4.21
+ $X2=21.135 $Y2=4.21
r130 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=20.885 $Y=4.21
+ $X2=21.225 $Y2=4.21
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.885
+ $Y=4.21 $X2=20.885 $Y2=4.21
r132 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.34 $Y=4.21
+ $X2=20.255 $Y2=4.21
r133 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=20.34 $Y=4.21
+ $X2=20.885 $Y2=4.21
r134 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=4.375
+ $X2=20.255 $Y2=4.21
r135 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=20.255 $Y=4.375
+ $X2=20.255 $Y2=4.615
r136 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=4.045
+ $X2=20.255 $Y2=4.21
r137 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=20.255 $Y=4.045
+ $X2=20.255 $Y2=3.835
r138 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=20.215 $Y=4.74
+ $X2=20.215 $Y2=4.615
r139 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=20.215 $Y=4.74
+ $X2=20.215 $Y2=4.995
r140 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.175 $Y=3.67
+ $X2=20.175 $Y2=3.835
r141 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=20.175 $Y=3.67
+ $X2=20.175 $Y2=3.14
r142 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.865 $Y=3.965
+ $X2=22.865 $Y2=3.475
r143 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.485 $Y=4.04
+ $X2=22.395 $Y2=4.04
r144 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=22.775 $Y=4.04
+ $X2=22.865 $Y2=3.965
r145 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.775 $Y=4.04
+ $X2=22.485 $Y2=4.04
r146 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=22.395 $Y=3.965
+ $X2=22.395 $Y2=4.04
r147 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.395 $Y=3.965
+ $X2=22.395 $Y2=3.475
r148 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.015 $Y=4.04
+ $X2=21.925 $Y2=4.04
r149 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.305 $Y=4.04
+ $X2=22.395 $Y2=4.04
r150 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.305 $Y=4.04
+ $X2=22.015 $Y2=4.04
r151 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=21.925 $Y=3.965
+ $X2=21.925 $Y2=4.04
r152 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.925 $Y=3.965
+ $X2=21.925 $Y2=3.475
r153 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.835 $Y=4.04
+ $X2=21.925 $Y2=4.04
r154 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.835 $Y=4.04
+ $X2=21.545 $Y2=4.04
r155 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=21.455 $Y=3.965
+ $X2=21.545 $Y2=4.04
r156 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=21.455 $Y=3.965
+ $X2=21.225 $Y2=4.155
r157 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.455 $Y=3.965
+ $X2=21.455 $Y2=3.475
r158 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.03
+ $Y=2.995 $X2=20.175 $Y2=3.14
r159 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.04
+ $Y=4.785 $X2=20.175 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[3] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r94 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=1.16
+ $X2=25.265 $Y2=1.16
r95 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=25.16 $Y=1.16
+ $X2=25.24 $Y2=1.16
r96 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=25.16
+ $Y=1.16 $X2=25.16 $Y2=1.16
r97 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=24.82 $Y=1.16
+ $X2=25.16 $Y2=1.16
r98 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=1.16
+ $X2=24.82 $Y2=1.16
r99 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.3 $Y=1.16
+ $X2=24.325 $Y2=1.16
r100 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=24.14 $Y=1.16
+ $X2=24.3 $Y2=1.16
r101 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.14
+ $Y=1.16 $X2=24.14 $Y2=1.16
r102 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=23.88 $Y=1.16
+ $X2=24.14 $Y2=1.16
r103 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=23.855 $Y=1.16
+ $X2=23.88 $Y2=1.16
r104 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=24.48 $Y=1.19
+ $X2=24.14 $Y2=1.19
r105 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.48
+ $Y=1.16 $X2=24.48 $Y2=1.16
r106 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.415 $Y=1.16
+ $X2=24.325 $Y2=1.16
r107 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=24.415 $Y=1.16
+ $X2=24.48 $Y2=1.16
r108 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.705 $Y=1.16
+ $X2=24.795 $Y2=1.16
r109 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=24.705 $Y=1.16
+ $X2=24.48 $Y2=1.16
r110 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=25.07 $Y=1.19
+ $X2=25.16 $Y2=1.19
r111 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=25.07 $Y=1.19
+ $X2=24.48 $Y2=1.19
r112 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.16
r113 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.985
r114 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=1.16
r115 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=0.56
r116 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=1.16
r117 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=0.56
r118 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.16
r119 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.985
r120 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.325 $Y=1.295
+ $X2=24.325 $Y2=1.16
r121 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.325 $Y=1.295
+ $X2=24.325 $Y2=1.985
r122 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.3 $Y=1.025
+ $X2=24.3 $Y2=1.16
r123 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.3 $Y=1.025
+ $X2=24.3 $Y2=0.56
r124 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=23.88 $Y=1.025
+ $X2=23.88 $Y2=1.16
r125 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=23.88 $Y=1.025
+ $X2=23.88 $Y2=0.56
r126 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.855 $Y=1.295
+ $X2=23.855 $Y2=1.16
r127 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=23.855 $Y=1.295
+ $X2=23.855 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[11] 3 7 11 15 19 23 27 31 33 35 36
+ 52 54
r92 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=4.28
+ $X2=25.265 $Y2=4.28
r93 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=25.16 $Y=4.28
+ $X2=25.24 $Y2=4.28
r94 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=25.16
+ $Y=4.28 $X2=25.16 $Y2=4.28
r95 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=24.82 $Y=4.28
+ $X2=25.16 $Y2=4.28
r96 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=4.28
+ $X2=24.82 $Y2=4.28
r97 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.3 $Y=4.28
+ $X2=24.325 $Y2=4.28
r98 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=24.14 $Y=4.28
+ $X2=24.3 $Y2=4.28
r99 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.14
+ $Y=4.28 $X2=24.14 $Y2=4.28
r100 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=23.88 $Y=4.28
+ $X2=24.14 $Y2=4.28
r101 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=23.855 $Y=4.28
+ $X2=23.88 $Y2=4.28
r102 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=24.48 $Y=4.25
+ $X2=24.14 $Y2=4.25
r103 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.48
+ $Y=4.28 $X2=24.48 $Y2=4.28
r104 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.415 $Y=4.28
+ $X2=24.325 $Y2=4.28
r105 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=24.415 $Y=4.28
+ $X2=24.48 $Y2=4.28
r106 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.705 $Y=4.28
+ $X2=24.795 $Y2=4.28
r107 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=24.705 $Y=4.28
+ $X2=24.48 $Y2=4.28
r108 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=25.07 $Y=4.25
+ $X2=25.16 $Y2=4.25
r109 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=25.07 $Y=4.25
+ $X2=24.48 $Y2=4.25
r110 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=4.145
+ $X2=25.265 $Y2=4.28
r111 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=4.145
+ $X2=25.265 $Y2=3.455
r112 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=4.415
+ $X2=25.24 $Y2=4.28
r113 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=4.415
+ $X2=25.24 $Y2=4.88
r114 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=4.415
+ $X2=24.82 $Y2=4.28
r115 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=4.415
+ $X2=24.82 $Y2=4.88
r116 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=4.145
+ $X2=24.795 $Y2=4.28
r117 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=4.145
+ $X2=24.795 $Y2=3.455
r118 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.325 $Y=4.145
+ $X2=24.325 $Y2=4.28
r119 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.325 $Y=4.145
+ $X2=24.325 $Y2=3.455
r120 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.3 $Y=4.415
+ $X2=24.3 $Y2=4.28
r121 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.3 $Y=4.415
+ $X2=24.3 $Y2=4.88
r122 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=23.88 $Y=4.415
+ $X2=23.88 $Y2=4.28
r123 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=23.88 $Y=4.415
+ $X2=23.88 $Y2=4.88
r124 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.855 $Y=4.145
+ $X2=23.855 $Y2=4.28
r125 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=23.855 $Y=4.145
+ $X2=23.855 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[4] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r96 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=28.1 $Y=1.16
+ $X2=28.125 $Y2=1.16
r97 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=27.84 $Y=1.16
+ $X2=28.1 $Y2=1.16
r98 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=27.84
+ $Y=1.16 $X2=27.84 $Y2=1.16
r99 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=27.68 $Y=1.16
+ $X2=27.84 $Y2=1.16
r100 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=27.655 $Y=1.16
+ $X2=27.68 $Y2=1.16
r101 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=27.16 $Y=1.16
+ $X2=27.185 $Y2=1.16
r102 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=27.16
+ $Y=1.16 $X2=27.16 $Y2=1.16
r103 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=26.74 $Y=1.16
+ $X2=27.16 $Y2=1.16
r104 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=26.715 $Y=1.16
+ $X2=26.74 $Y2=1.16
r105 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=27.5 $Y=1.19
+ $X2=27.84 $Y2=1.19
r106 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=27.5 $Y=1.19
+ $X2=27.16 $Y2=1.19
r107 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=27.5
+ $Y=1.16 $X2=27.5 $Y2=1.16
r108 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=27.275 $Y=1.16
+ $X2=27.185 $Y2=1.16
r109 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=27.275 $Y=1.16
+ $X2=27.5 $Y2=1.16
r110 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=27.565 $Y=1.16
+ $X2=27.655 $Y2=1.16
r111 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=27.565 $Y=1.16
+ $X2=27.5 $Y2=1.16
r112 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=26.91 $Y=1.19
+ $X2=27.16 $Y2=1.19
r113 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=28.125 $Y=1.295
+ $X2=28.125 $Y2=1.16
r114 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=28.125 $Y=1.295
+ $X2=28.125 $Y2=1.985
r115 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=28.1 $Y=1.025
+ $X2=28.1 $Y2=1.16
r116 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=28.1 $Y=1.025
+ $X2=28.1 $Y2=0.56
r117 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=27.68 $Y=1.025
+ $X2=27.68 $Y2=1.16
r118 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=27.68 $Y=1.025
+ $X2=27.68 $Y2=0.56
r119 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=27.655 $Y=1.295
+ $X2=27.655 $Y2=1.16
r120 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=27.655 $Y=1.295
+ $X2=27.655 $Y2=1.985
r121 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=27.185 $Y=1.295
+ $X2=27.185 $Y2=1.16
r122 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=27.185 $Y=1.295
+ $X2=27.185 $Y2=1.985
r123 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=27.16 $Y=1.025
+ $X2=27.16 $Y2=1.16
r124 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=27.16 $Y=1.025
+ $X2=27.16 $Y2=0.56
r125 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=26.74 $Y=1.025
+ $X2=26.74 $Y2=1.16
r126 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=26.74 $Y=1.025
+ $X2=26.74 $Y2=0.56
r127 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=26.715 $Y=1.295
+ $X2=26.715 $Y2=1.16
r128 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=26.715 $Y=1.295
+ $X2=26.715 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[12] 3 7 11 15 19 23 27 31 33 35 36
+ 51 53
r92 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=28.1 $Y=4.28
+ $X2=28.125 $Y2=4.28
r93 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=27.84 $Y=4.28
+ $X2=28.1 $Y2=4.28
r94 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=27.84
+ $Y=4.28 $X2=27.84 $Y2=4.28
r95 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=27.68 $Y=4.28
+ $X2=27.84 $Y2=4.28
r96 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=27.655 $Y=4.28
+ $X2=27.68 $Y2=4.28
r97 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=27.16 $Y=4.28
+ $X2=27.185 $Y2=4.28
r98 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=27.16
+ $Y=4.28 $X2=27.16 $Y2=4.28
r99 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=26.74 $Y=4.28
+ $X2=27.16 $Y2=4.28
r100 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=26.715 $Y=4.28
+ $X2=26.74 $Y2=4.28
r101 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=27.5 $Y=4.25
+ $X2=27.84 $Y2=4.25
r102 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=27.5 $Y=4.25
+ $X2=27.16 $Y2=4.25
r103 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=27.5
+ $Y=4.28 $X2=27.5 $Y2=4.28
r104 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=27.275 $Y=4.28
+ $X2=27.185 $Y2=4.28
r105 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=27.275 $Y=4.28
+ $X2=27.5 $Y2=4.28
r106 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=27.565 $Y=4.28
+ $X2=27.655 $Y2=4.28
r107 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=27.565 $Y=4.28
+ $X2=27.5 $Y2=4.28
r108 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=26.91 $Y=4.25
+ $X2=27.16 $Y2=4.25
r109 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=28.125 $Y=4.145
+ $X2=28.125 $Y2=4.28
r110 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=28.125 $Y=4.145
+ $X2=28.125 $Y2=3.455
r111 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=28.1 $Y=4.415
+ $X2=28.1 $Y2=4.28
r112 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=28.1 $Y=4.415
+ $X2=28.1 $Y2=4.88
r113 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=27.68 $Y=4.415
+ $X2=27.68 $Y2=4.28
r114 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=27.68 $Y=4.415
+ $X2=27.68 $Y2=4.88
r115 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=27.655 $Y=4.145
+ $X2=27.655 $Y2=4.28
r116 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=27.655 $Y=4.145
+ $X2=27.655 $Y2=3.455
r117 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=27.185 $Y=4.145
+ $X2=27.185 $Y2=4.28
r118 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=27.185 $Y=4.145
+ $X2=27.185 $Y2=3.455
r119 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=27.16 $Y=4.415
+ $X2=27.16 $Y2=4.28
r120 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=27.16 $Y=4.415
+ $X2=27.16 $Y2=4.88
r121 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=26.74 $Y=4.415
+ $X2=26.74 $Y2=4.28
r122 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=26.74 $Y=4.415
+ $X2=26.74 $Y2=4.88
r123 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=26.715 $Y=4.145
+ $X2=26.715 $Y2=4.28
r124 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=26.715 $Y=4.145
+ $X2=26.715 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c119 22 0 9.37986e-20 $X=30.525 $Y=1.475
c120 20 0 1.10627e-19 $X=30.435 $Y=1.4
c121 17 0 9.37986e-20 $X=30.055 $Y=1.475
c122 12 0 9.37986e-20 $X=29.585 $Y=1.475
c123 11 0 1.74242e-19 $X=29.205 $Y=1.4
c124 7 0 9.37986e-20 $X=29.115 $Y=1.475
r125 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=31.805 $Y=1.77
+ $X2=31.805 $Y2=1.605
r126 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=31.725 $Y=1.395
+ $X2=31.725 $Y2=1.23
r127 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=31.725 $Y=1.395
+ $X2=31.725 $Y2=1.605
r128 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=31.725 $Y=1.065
+ $X2=31.725 $Y2=1.23
r129 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=31.725 $Y=1.065
+ $X2=31.725 $Y2=0.825
r130 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=31.765 $Y=0.7
+ $X2=31.765 $Y2=0.825
r131 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=31.765 $Y=0.7
+ $X2=31.765 $Y2=0.445
r132 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=31.095 $Y=1.23
+ $X2=30.845 $Y2=1.23
r133 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=31.095
+ $Y=1.23 $X2=31.095 $Y2=1.23
r134 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=30.755
+ $Y=1.285 $X2=30.845 $Y2=1.23
r135 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=30.755 $Y=1.23
+ $X2=31.095 $Y2=1.23
r136 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=30.755
+ $Y=1.23 $X2=30.755 $Y2=1.23
r137 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=31.64 $Y=1.23
+ $X2=31.725 $Y2=1.23
r138 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=31.64 $Y=1.23
+ $X2=31.095 $Y2=1.23
r139 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=30.525
+ $Y=1.475 $X2=30.755 $Y2=1.285
r140 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=30.525 $Y=1.475
+ $X2=30.525 $Y2=1.965
r141 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=30.145 $Y=1.4
+ $X2=30.055 $Y2=1.4
r142 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=30.435 $Y=1.4
+ $X2=30.525 $Y2=1.475
r143 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=30.435 $Y=1.4
+ $X2=30.145 $Y2=1.4
r144 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=30.055 $Y=1.475
+ $X2=30.055 $Y2=1.4
r145 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=30.055 $Y=1.475
+ $X2=30.055 $Y2=1.965
r146 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.675 $Y=1.4
+ $X2=29.585 $Y2=1.4
r147 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.965 $Y=1.4
+ $X2=30.055 $Y2=1.4
r148 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=29.965 $Y=1.4
+ $X2=29.675 $Y2=1.4
r149 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=29.585 $Y=1.475
+ $X2=29.585 $Y2=1.4
r150 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=29.585 $Y=1.475
+ $X2=29.585 $Y2=1.965
r151 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.495 $Y=1.4
+ $X2=29.585 $Y2=1.4
r152 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=29.495 $Y=1.4
+ $X2=29.205 $Y2=1.4
r153 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=29.115 $Y=1.475
+ $X2=29.205 $Y2=1.4
r154 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=29.115 $Y=1.475
+ $X2=29.115 $Y2=1.965
r155 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=31.66
+ $Y=1.625 $X2=31.805 $Y2=1.77
r156 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=31.67
+ $Y=0.235 $X2=31.805 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c125 22 0 9.37986e-20 $X=30.525 $Y=3.965
c126 20 0 1.10627e-19 $X=30.435 $Y=4.04
c127 17 0 9.37986e-20 $X=30.055 $Y=3.965
c128 12 0 9.37986e-20 $X=29.585 $Y=3.965
c129 11 0 1.74242e-19 $X=29.205 $Y=4.04
c130 7 0 9.37986e-20 $X=29.115 $Y=3.965
r131 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=31.765 $Y=4.74
+ $X2=31.765 $Y2=4.615
r132 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=31.765 $Y=4.74
+ $X2=31.765 $Y2=4.995
r133 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=31.725 $Y=4.375
+ $X2=31.725 $Y2=4.21
r134 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=31.725 $Y=4.375
+ $X2=31.725 $Y2=4.615
r135 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=31.725 $Y=4.045
+ $X2=31.725 $Y2=4.21
r136 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=31.725 $Y=4.045
+ $X2=31.725 $Y2=3.835
r137 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=31.805 $Y=3.67
+ $X2=31.805 $Y2=3.835
r138 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=31.805 $Y=3.67
+ $X2=31.805 $Y2=3.14
r139 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=31.095 $Y=4.21
+ $X2=30.845 $Y2=4.21
r140 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=31.095
+ $Y=4.21 $X2=31.095 $Y2=4.21
r141 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=30.755
+ $Y=4.155 $X2=30.845 $Y2=4.21
r142 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=30.755 $Y=4.21
+ $X2=31.095 $Y2=4.21
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=30.755
+ $Y=4.21 $X2=30.755 $Y2=4.21
r144 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=31.64 $Y=4.21
+ $X2=31.725 $Y2=4.21
r145 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=31.64 $Y=4.21
+ $X2=31.095 $Y2=4.21
r146 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=30.525
+ $Y=3.965 $X2=30.755 $Y2=4.155
r147 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=30.525 $Y=3.965
+ $X2=30.525 $Y2=3.475
r148 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=30.145 $Y=4.04
+ $X2=30.055 $Y2=4.04
r149 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=30.435 $Y=4.04
+ $X2=30.525 $Y2=3.965
r150 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=30.435 $Y=4.04
+ $X2=30.145 $Y2=4.04
r151 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=30.055 $Y=3.965
+ $X2=30.055 $Y2=4.04
r152 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=30.055 $Y=3.965
+ $X2=30.055 $Y2=3.475
r153 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.675 $Y=4.04
+ $X2=29.585 $Y2=4.04
r154 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.965 $Y=4.04
+ $X2=30.055 $Y2=4.04
r155 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=29.965 $Y=4.04
+ $X2=29.675 $Y2=4.04
r156 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=29.585 $Y=3.965
+ $X2=29.585 $Y2=4.04
r157 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=29.585 $Y=3.965
+ $X2=29.585 $Y2=3.475
r158 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=29.495 $Y=4.04
+ $X2=29.585 $Y2=4.04
r159 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=29.495 $Y=4.04
+ $X2=29.205 $Y2=4.04
r160 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=29.115 $Y=3.965
+ $X2=29.205 $Y2=4.04
r161 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=29.115 $Y=3.965
+ $X2=29.115 $Y2=3.475
r162 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=31.66
+ $Y=2.995 $X2=31.805 $Y2=3.14
r163 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=31.67
+ $Y=4.785 $X2=31.805 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[4] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c117 11 0 1.3204e-19 $X=29.88 $Y=0.255
r118 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=32.42
+ $Y=1.16 $X2=32.42 $Y2=1.16
r119 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=32.04 $Y=1.55
+ $X2=32.247 $Y2=1.16
r120 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=32.04 $Y=1.55
+ $X2=32.04 $Y2=2.035
r121 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=32.015 $Y=0.735
+ $X2=32.015 $Y2=0.445
r122 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=31.67 $Y=0.81
+ $X2=31.57 $Y2=0.81
r123 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=31.94 $Y=0.81
+ $X2=32.247 $Y2=1.16
r124 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=31.94 $Y=0.81
+ $X2=32.015 $Y2=0.735
r125 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=31.94 $Y=0.81
+ $X2=31.67 $Y2=0.81
r126 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=31.595 $Y=0.735
+ $X2=31.57 $Y2=0.81
r127 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=31.595 $Y=0.735
+ $X2=31.595 $Y2=0.445
r128 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=31.57 $Y=1.55
+ $X2=31.57 $Y2=2.035
r129 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=31.57 $Y=1.45 $X2=31.57
+ $Y2=1.55
r130 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=31.57 $Y=0.885
+ $X2=31.57 $Y2=0.81
r131 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=31.57 $Y=0.885
+ $X2=31.57 $Y2=1.45
r132 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=31.47 $Y=0.81
+ $X2=31.57 $Y2=0.81
r133 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=31.47 $Y=0.81
+ $X2=31.135 $Y2=0.81
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=31.06 $Y=0.735
+ $X2=31.135 $Y2=0.81
r135 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=31.06 $Y=0.255
+ $X2=31.06 $Y2=0.735
r136 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.375 $Y=0.18
+ $X2=30.3 $Y2=0.18
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=30.985 $Y=0.18
+ $X2=31.06 $Y2=0.255
r138 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=30.985 $Y=0.18
+ $X2=30.375 $Y2=0.18
r139 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.3 $Y=0.255
+ $X2=30.3 $Y2=0.18
r140 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=30.3 $Y=0.255
+ $X2=30.3 $Y2=0.59
r141 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.955 $Y=0.18
+ $X2=29.88 $Y2=0.18
r142 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.225 $Y=0.18
+ $X2=30.3 $Y2=0.18
r143 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=30.225 $Y=0.18
+ $X2=29.955 $Y2=0.18
r144 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.88 $Y=0.255
+ $X2=29.88 $Y2=0.18
r145 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.88 $Y=0.255
+ $X2=29.88 $Y2=0.59
r146 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.535 $Y=0.18
+ $X2=29.46 $Y2=0.18
r147 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.805 $Y=0.18
+ $X2=29.88 $Y2=0.18
r148 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=29.805 $Y=0.18
+ $X2=29.535 $Y2=0.18
r149 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.46 $Y=0.255
+ $X2=29.46 $Y2=0.18
r150 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.46 $Y=0.255
+ $X2=29.46 $Y2=0.59
r151 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.385 $Y=0.18
+ $X2=29.46 $Y2=0.18
r152 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=29.385 $Y=0.18
+ $X2=29.115 $Y2=0.18
r153 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=29.04 $Y=0.255
+ $X2=29.115 $Y2=0.18
r154 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.04 $Y=0.255
+ $X2=29.04 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[12] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c125 11 0 1.3204e-19 $X=29.88 $Y=5.185
r126 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=32.42
+ $Y=4.28 $X2=32.42 $Y2=4.28
r127 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=32.04 $Y=3.89
+ $X2=32.247 $Y2=4.28
r128 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=32.04 $Y=3.89
+ $X2=32.04 $Y2=3.405
r129 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=32.015 $Y=4.705
+ $X2=32.015 $Y2=4.995
r130 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=31.67 $Y=4.63
+ $X2=31.57 $Y2=4.63
r131 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=31.94 $Y=4.63
+ $X2=32.015 $Y2=4.705
r132 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=31.94 $Y=4.63
+ $X2=32.247 $Y2=4.28
r133 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=31.94 $Y=4.63
+ $X2=31.67 $Y2=4.63
r134 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=31.595 $Y=4.705
+ $X2=31.57 $Y2=4.63
r135 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=31.595 $Y=4.705
+ $X2=31.595 $Y2=4.995
r136 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=31.57 $Y=3.89
+ $X2=31.57 $Y2=3.405
r137 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=31.57 $Y=4.555
+ $X2=31.57 $Y2=4.63
r138 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=31.57 $Y=3.99 $X2=31.57
+ $Y2=3.89
r139 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=31.57 $Y=3.99
+ $X2=31.57 $Y2=4.555
r140 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=31.47 $Y=4.63
+ $X2=31.57 $Y2=4.63
r141 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=31.47 $Y=4.63
+ $X2=31.135 $Y2=4.63
r142 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=31.06 $Y=4.705
+ $X2=31.135 $Y2=4.63
r143 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=31.06 $Y=4.705
+ $X2=31.06 $Y2=5.185
r144 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.375 $Y=5.26
+ $X2=30.3 $Y2=5.26
r145 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=30.985 $Y=5.26
+ $X2=31.06 $Y2=5.185
r146 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=30.985 $Y=5.26
+ $X2=30.375 $Y2=5.26
r147 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.3 $Y=5.185
+ $X2=30.3 $Y2=5.26
r148 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=30.3 $Y=5.185
+ $X2=30.3 $Y2=4.85
r149 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.955 $Y=5.26
+ $X2=29.88 $Y2=5.26
r150 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=30.225 $Y=5.26
+ $X2=30.3 $Y2=5.26
r151 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=30.225 $Y=5.26
+ $X2=29.955 $Y2=5.26
r152 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.88 $Y=5.185
+ $X2=29.88 $Y2=5.26
r153 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.88 $Y=5.185
+ $X2=29.88 $Y2=4.85
r154 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.535 $Y=5.26
+ $X2=29.46 $Y2=5.26
r155 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.805 $Y=5.26
+ $X2=29.88 $Y2=5.26
r156 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=29.805 $Y=5.26
+ $X2=29.535 $Y2=5.26
r157 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.46 $Y=5.185
+ $X2=29.46 $Y2=5.26
r158 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.46 $Y=5.185
+ $X2=29.46 $Y2=4.85
r159 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=29.385 $Y=5.26
+ $X2=29.46 $Y2=5.26
r160 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=29.385 $Y=5.26
+ $X2=29.115 $Y2=5.26
r161 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=29.04 $Y=5.185
+ $X2=29.115 $Y2=5.26
r162 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=29.04 $Y=5.185
+ $X2=29.04 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[5] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c120 30 0 1.3204e-19 $X=35.44 $Y=0.255
r121 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=32.89 $Y=1.16
+ $X2=33.24 $Y2=1.16
r122 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=36.28 $Y=0.255
+ $X2=36.28 $Y2=0.59
r123 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.935 $Y=0.18
+ $X2=35.86 $Y2=0.18
r124 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=36.205 $Y=0.18
+ $X2=36.28 $Y2=0.255
r125 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=36.205 $Y=0.18
+ $X2=35.935 $Y2=0.18
r126 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.86 $Y=0.255
+ $X2=35.86 $Y2=0.18
r127 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.86 $Y=0.255
+ $X2=35.86 $Y2=0.59
r128 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.515 $Y=0.18
+ $X2=35.44 $Y2=0.18
r129 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.785 $Y=0.18
+ $X2=35.86 $Y2=0.18
r130 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=35.785 $Y=0.18
+ $X2=35.515 $Y2=0.18
r131 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.44 $Y=0.255
+ $X2=35.44 $Y2=0.18
r132 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.44 $Y=0.255
+ $X2=35.44 $Y2=0.59
r133 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.095 $Y=0.18
+ $X2=35.02 $Y2=0.18
r134 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.365 $Y=0.18
+ $X2=35.44 $Y2=0.18
r135 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=35.365 $Y=0.18
+ $X2=35.095 $Y2=0.18
r136 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.02 $Y=0.255
+ $X2=35.02 $Y2=0.18
r137 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.02 $Y=0.255
+ $X2=35.02 $Y2=0.59
r138 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=34.945 $Y=0.18
+ $X2=35.02 $Y2=0.18
r139 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=34.945 $Y=0.18
+ $X2=34.335 $Y2=0.18
r140 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=34.26 $Y=0.255
+ $X2=34.335 $Y2=0.18
r141 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=34.26 $Y=0.255
+ $X2=34.26 $Y2=0.735
r142 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.85 $Y=0.81
+ $X2=33.75 $Y2=0.81
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=34.185 $Y=0.81
+ $X2=34.26 $Y2=0.735
r144 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=34.185 $Y=0.81
+ $X2=33.85 $Y2=0.81
r145 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=33.75 $Y=1.55
+ $X2=33.75 $Y2=2.035
r146 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=33.75 $Y=1.45 $X2=33.75
+ $Y2=1.55
r147 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=33.75 $Y=0.885
+ $X2=33.75 $Y2=0.81
r148 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=33.75 $Y=0.885
+ $X2=33.75 $Y2=1.45
r149 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=33.725 $Y=0.735
+ $X2=33.75 $Y2=0.81
r150 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=33.725 $Y=0.735
+ $X2=33.725 $Y2=0.445
r151 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.38 $Y=0.81
+ $X2=33.28 $Y2=0.81
r152 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.65 $Y=0.81
+ $X2=33.75 $Y2=0.81
r153 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=33.65 $Y=0.81
+ $X2=33.38 $Y2=0.81
r154 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=33.305 $Y=0.735
+ $X2=33.28 $Y2=0.81
r155 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=33.305 $Y=0.735
+ $X2=33.305 $Y2=0.445
r156 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=33.28 $Y=1.55
+ $X2=33.28 $Y2=2.035
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=33.28 $Y=1.16
+ $X2=33.28 $Y2=1.55
r158 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=33.24
+ $Y=1.16 $X2=33.24 $Y2=1.16
r159 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=33.28 $Y=1.16
+ $X2=33.28 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[13] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c128 30 0 1.3204e-19 $X=35.44 $Y=5.185
r129 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=32.89 $Y=4.28
+ $X2=33.24 $Y2=4.28
r130 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=36.28 $Y=5.185
+ $X2=36.28 $Y2=4.85
r131 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.935 $Y=5.26
+ $X2=35.86 $Y2=5.26
r132 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=36.205 $Y=5.26
+ $X2=36.28 $Y2=5.185
r133 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=36.205 $Y=5.26
+ $X2=35.935 $Y2=5.26
r134 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.86 $Y=5.185
+ $X2=35.86 $Y2=5.26
r135 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.86 $Y=5.185
+ $X2=35.86 $Y2=4.85
r136 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.515 $Y=5.26
+ $X2=35.44 $Y2=5.26
r137 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.785 $Y=5.26
+ $X2=35.86 $Y2=5.26
r138 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=35.785 $Y=5.26
+ $X2=35.515 $Y2=5.26
r139 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.44 $Y=5.185
+ $X2=35.44 $Y2=5.26
r140 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.44 $Y=5.185
+ $X2=35.44 $Y2=4.85
r141 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.095 $Y=5.26
+ $X2=35.02 $Y2=5.26
r142 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.365 $Y=5.26
+ $X2=35.44 $Y2=5.26
r143 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=35.365 $Y=5.26
+ $X2=35.095 $Y2=5.26
r144 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=35.02 $Y=5.185
+ $X2=35.02 $Y2=5.26
r145 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=35.02 $Y=5.185
+ $X2=35.02 $Y2=4.85
r146 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=34.945 $Y=5.26
+ $X2=35.02 $Y2=5.26
r147 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=34.945 $Y=5.26
+ $X2=34.335 $Y2=5.26
r148 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=34.26 $Y=5.185
+ $X2=34.335 $Y2=5.26
r149 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=34.26 $Y=4.705
+ $X2=34.26 $Y2=5.185
r150 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.85 $Y=4.63
+ $X2=33.75 $Y2=4.63
r151 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=34.185 $Y=4.63
+ $X2=34.26 $Y2=4.705
r152 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=34.185 $Y=4.63
+ $X2=33.85 $Y2=4.63
r153 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=33.75 $Y=3.89
+ $X2=33.75 $Y2=3.405
r154 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=33.725 $Y=4.705
+ $X2=33.75 $Y2=4.63
r155 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=33.725 $Y=4.705
+ $X2=33.725 $Y2=4.995
r156 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=33.75 $Y=4.555
+ $X2=33.75 $Y2=4.63
r157 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=33.75 $Y=3.99 $X2=33.75
+ $Y2=3.89
r158 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=33.75 $Y=3.99
+ $X2=33.75 $Y2=4.555
r159 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.38 $Y=4.63
+ $X2=33.28 $Y2=4.63
r160 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=33.65 $Y=4.63
+ $X2=33.75 $Y2=4.63
r161 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=33.65 $Y=4.63
+ $X2=33.38 $Y2=4.63
r162 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=33.305 $Y=4.705
+ $X2=33.28 $Y2=4.63
r163 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=33.305 $Y=4.705
+ $X2=33.305 $Y2=4.995
r164 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=33.28 $Y=3.89
+ $X2=33.28 $Y2=3.405
r165 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=33.28 $Y=4.28
+ $X2=33.28 $Y2=4.63
r166 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=33.24
+ $Y=4.28 $X2=33.24 $Y2=4.28
r167 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=33.28 $Y=4.28
+ $X2=33.28 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c116 22 0 9.37986e-20 $X=36.205 $Y=1.475
c117 20 0 1.74242e-19 $X=36.115 $Y=1.4
c118 17 0 9.37986e-20 $X=35.735 $Y=1.475
c119 12 0 9.37986e-20 $X=35.265 $Y=1.475
c120 7 0 9.37986e-20 $X=34.795 $Y=1.475
r121 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=34.565
+ $Y=1.285 $X2=34.475 $Y2=1.23
r122 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=34.565
+ $Y=1.23 $X2=34.565 $Y2=1.23
r123 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=34.225 $Y=1.23
+ $X2=34.475 $Y2=1.23
r124 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=34.225 $Y=1.23
+ $X2=34.565 $Y2=1.23
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=34.225
+ $Y=1.23 $X2=34.225 $Y2=1.23
r126 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=33.68 $Y=1.23
+ $X2=33.595 $Y2=1.23
r127 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=33.68 $Y=1.23
+ $X2=34.225 $Y2=1.23
r128 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=33.595 $Y=1.395
+ $X2=33.595 $Y2=1.23
r129 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=33.595 $Y=1.395
+ $X2=33.595 $Y2=1.605
r130 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=33.595 $Y=1.065
+ $X2=33.595 $Y2=1.23
r131 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=33.595 $Y=1.065
+ $X2=33.595 $Y2=0.825
r132 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=33.555 $Y=0.7
+ $X2=33.555 $Y2=0.825
r133 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=33.555 $Y=0.7
+ $X2=33.555 $Y2=0.445
r134 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=33.515 $Y=1.77
+ $X2=33.515 $Y2=1.605
r135 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=36.205 $Y=1.475
+ $X2=36.205 $Y2=1.965
r136 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.825 $Y=1.4
+ $X2=35.735 $Y2=1.4
r137 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=36.115 $Y=1.4
+ $X2=36.205 $Y2=1.475
r138 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=36.115 $Y=1.4
+ $X2=35.825 $Y2=1.4
r139 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=35.735 $Y=1.475
+ $X2=35.735 $Y2=1.4
r140 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=35.735 $Y=1.475
+ $X2=35.735 $Y2=1.965
r141 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.355 $Y=1.4
+ $X2=35.265 $Y2=1.4
r142 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.645 $Y=1.4
+ $X2=35.735 $Y2=1.4
r143 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=35.645 $Y=1.4
+ $X2=35.355 $Y2=1.4
r144 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=35.265 $Y=1.475
+ $X2=35.265 $Y2=1.4
r145 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=35.265 $Y=1.475
+ $X2=35.265 $Y2=1.965
r146 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.175 $Y=1.4
+ $X2=35.265 $Y2=1.4
r147 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=35.175 $Y=1.4
+ $X2=34.885 $Y2=1.4
r148 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=34.795 $Y=1.475
+ $X2=34.885 $Y2=1.4
r149 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=34.795 $Y=1.475
+ $X2=34.565 $Y2=1.285
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=34.795 $Y=1.475
+ $X2=34.795 $Y2=1.965
r151 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=33.37
+ $Y=1.625 $X2=33.515 $Y2=1.77
r152 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=33.38
+ $Y=0.235 $X2=33.515 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_599# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c122 22 0 9.37986e-20 $X=36.205 $Y=3.965
c123 20 0 1.74242e-19 $X=36.115 $Y=4.04
c124 17 0 9.37986e-20 $X=35.735 $Y=3.965
c125 12 0 9.37986e-20 $X=35.265 $Y=3.965
c126 7 0 9.37986e-20 $X=34.795 $Y=3.965
r127 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=34.565
+ $Y=4.155 $X2=34.475 $Y2=4.21
r128 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=34.565
+ $Y=4.21 $X2=34.565 $Y2=4.21
r129 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=34.225 $Y=4.21
+ $X2=34.475 $Y2=4.21
r130 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=34.225 $Y=4.21
+ $X2=34.565 $Y2=4.21
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=34.225
+ $Y=4.21 $X2=34.225 $Y2=4.21
r132 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=33.68 $Y=4.21
+ $X2=33.595 $Y2=4.21
r133 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=33.68 $Y=4.21
+ $X2=34.225 $Y2=4.21
r134 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=33.595 $Y=4.375
+ $X2=33.595 $Y2=4.21
r135 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=33.595 $Y=4.375
+ $X2=33.595 $Y2=4.615
r136 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=33.595 $Y=4.045
+ $X2=33.595 $Y2=4.21
r137 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=33.595 $Y=4.045
+ $X2=33.595 $Y2=3.835
r138 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=33.555 $Y=4.74
+ $X2=33.555 $Y2=4.615
r139 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=33.555 $Y=4.74
+ $X2=33.555 $Y2=4.995
r140 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=33.515 $Y=3.67
+ $X2=33.515 $Y2=3.835
r141 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=33.515 $Y=3.67
+ $X2=33.515 $Y2=3.14
r142 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=36.205 $Y=3.965
+ $X2=36.205 $Y2=3.475
r143 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.825 $Y=4.04
+ $X2=35.735 $Y2=4.04
r144 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=36.115 $Y=4.04
+ $X2=36.205 $Y2=3.965
r145 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=36.115 $Y=4.04
+ $X2=35.825 $Y2=4.04
r146 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=35.735 $Y=3.965
+ $X2=35.735 $Y2=4.04
r147 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=35.735 $Y=3.965
+ $X2=35.735 $Y2=3.475
r148 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.355 $Y=4.04
+ $X2=35.265 $Y2=4.04
r149 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.645 $Y=4.04
+ $X2=35.735 $Y2=4.04
r150 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=35.645 $Y=4.04
+ $X2=35.355 $Y2=4.04
r151 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=35.265 $Y=3.965
+ $X2=35.265 $Y2=4.04
r152 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=35.265 $Y=3.965
+ $X2=35.265 $Y2=3.475
r153 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=35.175 $Y=4.04
+ $X2=35.265 $Y2=4.04
r154 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=35.175 $Y=4.04
+ $X2=34.885 $Y2=4.04
r155 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=34.795 $Y=3.965
+ $X2=34.885 $Y2=4.04
r156 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=34.795 $Y=3.965
+ $X2=34.565 $Y2=4.155
r157 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=34.795 $Y=3.965
+ $X2=34.795 $Y2=3.475
r158 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=33.37
+ $Y=2.995 $X2=33.515 $Y2=3.14
r159 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=33.38
+ $Y=4.785 $X2=33.515 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[5] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r93 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=38.58 $Y=1.16
+ $X2=38.605 $Y2=1.16
r94 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=38.5 $Y=1.16 $X2=38.58
+ $Y2=1.16
r95 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=38.5
+ $Y=1.16 $X2=38.5 $Y2=1.16
r96 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=38.16 $Y=1.16
+ $X2=38.5 $Y2=1.16
r97 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=38.135 $Y=1.16
+ $X2=38.16 $Y2=1.16
r98 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=37.64 $Y=1.16
+ $X2=37.665 $Y2=1.16
r99 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=37.48 $Y=1.16
+ $X2=37.64 $Y2=1.16
r100 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=37.48
+ $Y=1.16 $X2=37.48 $Y2=1.16
r101 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=37.22 $Y=1.16
+ $X2=37.48 $Y2=1.16
r102 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=37.195 $Y=1.16
+ $X2=37.22 $Y2=1.16
r103 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=37.82 $Y=1.19
+ $X2=37.48 $Y2=1.19
r104 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=37.82
+ $Y=1.16 $X2=37.82 $Y2=1.16
r105 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=37.755 $Y=1.16
+ $X2=37.665 $Y2=1.16
r106 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=37.755 $Y=1.16
+ $X2=37.82 $Y2=1.16
r107 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=38.045 $Y=1.16
+ $X2=38.135 $Y2=1.16
r108 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=38.045 $Y=1.16
+ $X2=37.82 $Y2=1.16
r109 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=38.41 $Y=1.19
+ $X2=38.5 $Y2=1.19
r110 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=38.41 $Y=1.19
+ $X2=37.82 $Y2=1.19
r111 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=38.605 $Y=1.295
+ $X2=38.605 $Y2=1.16
r112 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=38.605 $Y=1.295
+ $X2=38.605 $Y2=1.985
r113 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=38.58 $Y=1.025
+ $X2=38.58 $Y2=1.16
r114 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=38.58 $Y=1.025
+ $X2=38.58 $Y2=0.56
r115 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=38.16 $Y=1.025
+ $X2=38.16 $Y2=1.16
r116 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=38.16 $Y=1.025
+ $X2=38.16 $Y2=0.56
r117 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=38.135 $Y=1.295
+ $X2=38.135 $Y2=1.16
r118 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=38.135 $Y=1.295
+ $X2=38.135 $Y2=1.985
r119 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=37.665 $Y=1.295
+ $X2=37.665 $Y2=1.16
r120 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=37.665 $Y=1.295
+ $X2=37.665 $Y2=1.985
r121 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=37.64 $Y=1.025
+ $X2=37.64 $Y2=1.16
r122 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=37.64 $Y=1.025
+ $X2=37.64 $Y2=0.56
r123 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=37.22 $Y=1.025
+ $X2=37.22 $Y2=1.16
r124 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=37.22 $Y=1.025
+ $X2=37.22 $Y2=0.56
r125 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=37.195 $Y=1.295
+ $X2=37.195 $Y2=1.16
r126 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=37.195 $Y=1.295
+ $X2=37.195 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[13] 3 7 11 15 19 23 27 31 33 35 36
+ 52 54
r91 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=38.58 $Y=4.28
+ $X2=38.605 $Y2=4.28
r92 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=38.5 $Y=4.28 $X2=38.58
+ $Y2=4.28
r93 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=38.5
+ $Y=4.28 $X2=38.5 $Y2=4.28
r94 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=38.16 $Y=4.28
+ $X2=38.5 $Y2=4.28
r95 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=38.135 $Y=4.28
+ $X2=38.16 $Y2=4.28
r96 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=37.64 $Y=4.28
+ $X2=37.665 $Y2=4.28
r97 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=37.48 $Y=4.28
+ $X2=37.64 $Y2=4.28
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=37.48
+ $Y=4.28 $X2=37.48 $Y2=4.28
r99 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=37.22 $Y=4.28
+ $X2=37.48 $Y2=4.28
r100 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=37.195 $Y=4.28
+ $X2=37.22 $Y2=4.28
r101 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=37.82 $Y=4.25
+ $X2=37.48 $Y2=4.25
r102 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=37.82
+ $Y=4.28 $X2=37.82 $Y2=4.28
r103 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=37.755 $Y=4.28
+ $X2=37.665 $Y2=4.28
r104 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=37.755 $Y=4.28
+ $X2=37.82 $Y2=4.28
r105 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=38.045 $Y=4.28
+ $X2=38.135 $Y2=4.28
r106 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=38.045 $Y=4.28
+ $X2=37.82 $Y2=4.28
r107 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=38.41 $Y=4.25
+ $X2=38.5 $Y2=4.25
r108 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=38.41 $Y=4.25
+ $X2=37.82 $Y2=4.25
r109 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=38.605 $Y=4.145
+ $X2=38.605 $Y2=4.28
r110 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=38.605 $Y=4.145
+ $X2=38.605 $Y2=3.455
r111 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=38.58 $Y=4.415
+ $X2=38.58 $Y2=4.28
r112 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=38.58 $Y=4.415
+ $X2=38.58 $Y2=4.88
r113 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=38.16 $Y=4.415
+ $X2=38.16 $Y2=4.28
r114 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=38.16 $Y=4.415
+ $X2=38.16 $Y2=4.88
r115 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=38.135 $Y=4.145
+ $X2=38.135 $Y2=4.28
r116 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=38.135 $Y=4.145
+ $X2=38.135 $Y2=3.455
r117 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=37.665 $Y=4.145
+ $X2=37.665 $Y2=4.28
r118 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=37.665 $Y=4.145
+ $X2=37.665 $Y2=3.455
r119 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=37.64 $Y=4.415
+ $X2=37.64 $Y2=4.28
r120 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=37.64 $Y=4.415
+ $X2=37.64 $Y2=4.88
r121 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=37.22 $Y=4.415
+ $X2=37.22 $Y2=4.28
r122 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=37.22 $Y=4.415
+ $X2=37.22 $Y2=4.88
r123 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=37.195 $Y=4.145
+ $X2=37.195 $Y2=4.28
r124 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=37.195 $Y=4.145
+ $X2=37.195 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[6] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r95 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.98 $Y=1.16
+ $X2=41.005 $Y2=1.16
r96 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=40.72 $Y=1.16
+ $X2=40.98 $Y2=1.16
r97 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=40.72
+ $Y=1.16 $X2=40.72 $Y2=1.16
r98 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=40.56 $Y=1.16
+ $X2=40.72 $Y2=1.16
r99 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.535 $Y=1.16
+ $X2=40.56 $Y2=1.16
r100 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.04 $Y=1.16
+ $X2=40.065 $Y2=1.16
r101 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=40.04
+ $Y=1.16 $X2=40.04 $Y2=1.16
r102 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=39.62 $Y=1.16
+ $X2=40.04 $Y2=1.16
r103 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=39.595 $Y=1.16
+ $X2=39.62 $Y2=1.16
r104 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=40.38 $Y=1.19
+ $X2=40.72 $Y2=1.19
r105 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=40.38 $Y=1.19
+ $X2=40.04 $Y2=1.19
r106 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=40.38
+ $Y=1.16 $X2=40.38 $Y2=1.16
r107 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=40.155 $Y=1.16
+ $X2=40.065 $Y2=1.16
r108 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=40.155 $Y=1.16
+ $X2=40.38 $Y2=1.16
r109 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=40.445 $Y=1.16
+ $X2=40.535 $Y2=1.16
r110 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=40.445 $Y=1.16
+ $X2=40.38 $Y2=1.16
r111 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=39.79 $Y=1.19
+ $X2=40.04 $Y2=1.19
r112 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=41.005 $Y=1.295
+ $X2=41.005 $Y2=1.16
r113 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=41.005 $Y=1.295
+ $X2=41.005 $Y2=1.985
r114 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.98 $Y=1.025
+ $X2=40.98 $Y2=1.16
r115 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.98 $Y=1.025
+ $X2=40.98 $Y2=0.56
r116 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.56 $Y=1.025
+ $X2=40.56 $Y2=1.16
r117 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.56 $Y=1.025
+ $X2=40.56 $Y2=0.56
r118 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=40.535 $Y=1.295
+ $X2=40.535 $Y2=1.16
r119 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=40.535 $Y=1.295
+ $X2=40.535 $Y2=1.985
r120 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=40.065 $Y=1.295
+ $X2=40.065 $Y2=1.16
r121 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=40.065 $Y=1.295
+ $X2=40.065 $Y2=1.985
r122 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.04 $Y=1.025
+ $X2=40.04 $Y2=1.16
r123 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.04 $Y=1.025
+ $X2=40.04 $Y2=0.56
r124 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=39.62 $Y=1.025
+ $X2=39.62 $Y2=1.16
r125 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=39.62 $Y=1.025
+ $X2=39.62 $Y2=0.56
r126 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=39.595 $Y=1.295
+ $X2=39.595 $Y2=1.16
r127 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=39.595 $Y=1.295
+ $X2=39.595 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[14] 3 7 11 15 19 23 27 31 33 35 36
+ 51 53
r91 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.98 $Y=4.28
+ $X2=41.005 $Y2=4.28
r92 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=40.72 $Y=4.28
+ $X2=40.98 $Y2=4.28
r93 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=40.72
+ $Y=4.28 $X2=40.72 $Y2=4.28
r94 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=40.56 $Y=4.28
+ $X2=40.72 $Y2=4.28
r95 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.535 $Y=4.28
+ $X2=40.56 $Y2=4.28
r96 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=40.04 $Y=4.28
+ $X2=40.065 $Y2=4.28
r97 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=40.04
+ $Y=4.28 $X2=40.04 $Y2=4.28
r98 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=39.62 $Y=4.28
+ $X2=40.04 $Y2=4.28
r99 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=39.595 $Y=4.28
+ $X2=39.62 $Y2=4.28
r100 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=40.38 $Y=4.25
+ $X2=40.72 $Y2=4.25
r101 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=40.38 $Y=4.25
+ $X2=40.04 $Y2=4.25
r102 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=40.38
+ $Y=4.28 $X2=40.38 $Y2=4.28
r103 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=40.155 $Y=4.28
+ $X2=40.065 $Y2=4.28
r104 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=40.155 $Y=4.28
+ $X2=40.38 $Y2=4.28
r105 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=40.445 $Y=4.28
+ $X2=40.535 $Y2=4.28
r106 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=40.445 $Y=4.28
+ $X2=40.38 $Y2=4.28
r107 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=39.79 $Y=4.25
+ $X2=40.04 $Y2=4.25
r108 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=41.005 $Y=4.145
+ $X2=41.005 $Y2=4.28
r109 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=41.005 $Y=4.145
+ $X2=41.005 $Y2=3.455
r110 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.98 $Y=4.415
+ $X2=40.98 $Y2=4.28
r111 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.98 $Y=4.415
+ $X2=40.98 $Y2=4.88
r112 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.56 $Y=4.415
+ $X2=40.56 $Y2=4.28
r113 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.56 $Y=4.415
+ $X2=40.56 $Y2=4.88
r114 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=40.535 $Y=4.145
+ $X2=40.535 $Y2=4.28
r115 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=40.535 $Y=4.145
+ $X2=40.535 $Y2=3.455
r116 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=40.065 $Y=4.145
+ $X2=40.065 $Y2=4.28
r117 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=40.065 $Y=4.145
+ $X2=40.065 $Y2=3.455
r118 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=40.04 $Y=4.415
+ $X2=40.04 $Y2=4.28
r119 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=40.04 $Y=4.415
+ $X2=40.04 $Y2=4.88
r120 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=39.62 $Y=4.415
+ $X2=39.62 $Y2=4.28
r121 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=39.62 $Y=4.415
+ $X2=39.62 $Y2=4.88
r122 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=39.595 $Y=4.145
+ $X2=39.595 $Y2=4.28
r123 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=39.595 $Y=4.145
+ $X2=39.595 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c119 22 0 9.37986e-20 $X=43.405 $Y=1.475
c120 20 0 1.10627e-19 $X=43.315 $Y=1.4
c121 17 0 9.37986e-20 $X=42.935 $Y=1.475
c122 12 0 9.37986e-20 $X=42.465 $Y=1.475
c123 11 0 1.74242e-19 $X=42.085 $Y=1.4
c124 7 0 9.37986e-20 $X=41.995 $Y=1.475
r125 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=44.685 $Y=1.77
+ $X2=44.685 $Y2=1.605
r126 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=44.605 $Y=1.395
+ $X2=44.605 $Y2=1.23
r127 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=44.605 $Y=1.395
+ $X2=44.605 $Y2=1.605
r128 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=44.605 $Y=1.065
+ $X2=44.605 $Y2=1.23
r129 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=44.605 $Y=1.065
+ $X2=44.605 $Y2=0.825
r130 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=44.645 $Y=0.7
+ $X2=44.645 $Y2=0.825
r131 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=44.645 $Y=0.7
+ $X2=44.645 $Y2=0.445
r132 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=43.975 $Y=1.23
+ $X2=43.725 $Y2=1.23
r133 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=43.975
+ $Y=1.23 $X2=43.975 $Y2=1.23
r134 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=43.635
+ $Y=1.285 $X2=43.725 $Y2=1.23
r135 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=43.635 $Y=1.23
+ $X2=43.975 $Y2=1.23
r136 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=43.635
+ $Y=1.23 $X2=43.635 $Y2=1.23
r137 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=44.52 $Y=1.23
+ $X2=44.605 $Y2=1.23
r138 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=44.52 $Y=1.23
+ $X2=43.975 $Y2=1.23
r139 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=43.405
+ $Y=1.475 $X2=43.635 $Y2=1.285
r140 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=43.405 $Y=1.475
+ $X2=43.405 $Y2=1.965
r141 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=43.025 $Y=1.4
+ $X2=42.935 $Y2=1.4
r142 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=43.315 $Y=1.4
+ $X2=43.405 $Y2=1.475
r143 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=43.315 $Y=1.4
+ $X2=43.025 $Y2=1.4
r144 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=42.935 $Y=1.475
+ $X2=42.935 $Y2=1.4
r145 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=42.935 $Y=1.475
+ $X2=42.935 $Y2=1.965
r146 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.555 $Y=1.4
+ $X2=42.465 $Y2=1.4
r147 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.845 $Y=1.4
+ $X2=42.935 $Y2=1.4
r148 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=42.845 $Y=1.4
+ $X2=42.555 $Y2=1.4
r149 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=42.465 $Y=1.475
+ $X2=42.465 $Y2=1.4
r150 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=42.465 $Y=1.475
+ $X2=42.465 $Y2=1.965
r151 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.375 $Y=1.4
+ $X2=42.465 $Y2=1.4
r152 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=42.375 $Y=1.4
+ $X2=42.085 $Y2=1.4
r153 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=41.995 $Y=1.475
+ $X2=42.085 $Y2=1.4
r154 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=41.995 $Y=1.475
+ $X2=41.995 $Y2=1.965
r155 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=44.54
+ $Y=1.625 $X2=44.685 $Y2=1.77
r156 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=44.55
+ $Y=0.235 $X2=44.685 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c125 22 0 9.37986e-20 $X=43.405 $Y=3.965
c126 20 0 1.10627e-19 $X=43.315 $Y=4.04
c127 17 0 9.37986e-20 $X=42.935 $Y=3.965
c128 12 0 9.37986e-20 $X=42.465 $Y=3.965
c129 11 0 1.74242e-19 $X=42.085 $Y=4.04
c130 7 0 9.37986e-20 $X=41.995 $Y=3.965
r131 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=44.645 $Y=4.74
+ $X2=44.645 $Y2=4.615
r132 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=44.645 $Y=4.74
+ $X2=44.645 $Y2=4.995
r133 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=44.605 $Y=4.375
+ $X2=44.605 $Y2=4.21
r134 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=44.605 $Y=4.375
+ $X2=44.605 $Y2=4.615
r135 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=44.605 $Y=4.045
+ $X2=44.605 $Y2=4.21
r136 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=44.605 $Y=4.045
+ $X2=44.605 $Y2=3.835
r137 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=44.685 $Y=3.67
+ $X2=44.685 $Y2=3.835
r138 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=44.685 $Y=3.67
+ $X2=44.685 $Y2=3.14
r139 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=43.975 $Y=4.21
+ $X2=43.725 $Y2=4.21
r140 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=43.975
+ $Y=4.21 $X2=43.975 $Y2=4.21
r141 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=43.635
+ $Y=4.155 $X2=43.725 $Y2=4.21
r142 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=43.635 $Y=4.21
+ $X2=43.975 $Y2=4.21
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=43.635
+ $Y=4.21 $X2=43.635 $Y2=4.21
r144 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=44.52 $Y=4.21
+ $X2=44.605 $Y2=4.21
r145 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=44.52 $Y=4.21
+ $X2=43.975 $Y2=4.21
r146 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=43.405
+ $Y=3.965 $X2=43.635 $Y2=4.155
r147 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=43.405 $Y=3.965
+ $X2=43.405 $Y2=3.475
r148 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=43.025 $Y=4.04
+ $X2=42.935 $Y2=4.04
r149 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=43.315 $Y=4.04
+ $X2=43.405 $Y2=3.965
r150 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=43.315 $Y=4.04
+ $X2=43.025 $Y2=4.04
r151 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=42.935 $Y=3.965
+ $X2=42.935 $Y2=4.04
r152 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=42.935 $Y=3.965
+ $X2=42.935 $Y2=3.475
r153 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.555 $Y=4.04
+ $X2=42.465 $Y2=4.04
r154 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.845 $Y=4.04
+ $X2=42.935 $Y2=4.04
r155 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=42.845 $Y=4.04
+ $X2=42.555 $Y2=4.04
r156 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=42.465 $Y=3.965
+ $X2=42.465 $Y2=4.04
r157 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=42.465 $Y=3.965
+ $X2=42.465 $Y2=3.475
r158 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=42.375 $Y=4.04
+ $X2=42.465 $Y2=4.04
r159 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=42.375 $Y=4.04
+ $X2=42.085 $Y2=4.04
r160 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=41.995 $Y=3.965
+ $X2=42.085 $Y2=4.04
r161 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=41.995 $Y=3.965
+ $X2=41.995 $Y2=3.475
r162 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=44.54
+ $Y=2.995 $X2=44.685 $Y2=3.14
r163 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=44.55
+ $Y=4.785 $X2=44.685 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[6] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c117 11 0 1.3204e-19 $X=42.76 $Y=0.255
r118 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=45.3
+ $Y=1.16 $X2=45.3 $Y2=1.16
r119 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=44.92 $Y=1.55
+ $X2=45.127 $Y2=1.16
r120 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=44.92 $Y=1.55
+ $X2=44.92 $Y2=2.035
r121 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=44.895 $Y=0.735
+ $X2=44.895 $Y2=0.445
r122 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=44.55 $Y=0.81
+ $X2=44.45 $Y2=0.81
r123 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=44.82 $Y=0.81
+ $X2=45.127 $Y2=1.16
r124 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=44.82 $Y=0.81
+ $X2=44.895 $Y2=0.735
r125 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=44.82 $Y=0.81
+ $X2=44.55 $Y2=0.81
r126 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=44.475 $Y=0.735
+ $X2=44.45 $Y2=0.81
r127 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=44.475 $Y=0.735
+ $X2=44.475 $Y2=0.445
r128 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=44.45 $Y=1.55
+ $X2=44.45 $Y2=2.035
r129 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=44.45 $Y=1.45 $X2=44.45
+ $Y2=1.55
r130 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=44.45 $Y=0.885
+ $X2=44.45 $Y2=0.81
r131 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=44.45 $Y=0.885
+ $X2=44.45 $Y2=1.45
r132 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=44.35 $Y=0.81
+ $X2=44.45 $Y2=0.81
r133 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=44.35 $Y=0.81
+ $X2=44.015 $Y2=0.81
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=43.94 $Y=0.735
+ $X2=44.015 $Y2=0.81
r135 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=43.94 $Y=0.255
+ $X2=43.94 $Y2=0.735
r136 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.255 $Y=0.18
+ $X2=43.18 $Y2=0.18
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=43.865 $Y=0.18
+ $X2=43.94 $Y2=0.255
r138 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=43.865 $Y=0.18
+ $X2=43.255 $Y2=0.18
r139 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.18 $Y=0.255
+ $X2=43.18 $Y2=0.18
r140 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=43.18 $Y=0.255
+ $X2=43.18 $Y2=0.59
r141 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.835 $Y=0.18
+ $X2=42.76 $Y2=0.18
r142 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.105 $Y=0.18
+ $X2=43.18 $Y2=0.18
r143 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=43.105 $Y=0.18
+ $X2=42.835 $Y2=0.18
r144 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.76 $Y=0.255
+ $X2=42.76 $Y2=0.18
r145 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=42.76 $Y=0.255
+ $X2=42.76 $Y2=0.59
r146 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.415 $Y=0.18
+ $X2=42.34 $Y2=0.18
r147 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.685 $Y=0.18
+ $X2=42.76 $Y2=0.18
r148 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=42.685 $Y=0.18
+ $X2=42.415 $Y2=0.18
r149 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.34 $Y=0.255
+ $X2=42.34 $Y2=0.18
r150 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=42.34 $Y=0.255
+ $X2=42.34 $Y2=0.59
r151 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.265 $Y=0.18
+ $X2=42.34 $Y2=0.18
r152 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=42.265 $Y=0.18
+ $X2=41.995 $Y2=0.18
r153 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=41.92 $Y=0.255
+ $X2=41.995 $Y2=0.18
r154 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=41.92 $Y=0.255
+ $X2=41.92 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[14] 1 3 4 5 6 8 9 11 13 14 16 18 19
+ 22 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c125 11 0 1.3204e-19 $X=42.76 $Y=5.185
r126 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=45.3
+ $Y=4.28 $X2=45.3 $Y2=4.28
r127 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=44.92 $Y=3.89
+ $X2=45.127 $Y2=4.28
r128 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=44.92 $Y=3.89
+ $X2=44.92 $Y2=3.405
r129 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=44.895 $Y=4.705
+ $X2=44.895 $Y2=4.995
r130 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=44.55 $Y=4.63
+ $X2=44.45 $Y2=4.63
r131 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=44.82 $Y=4.63
+ $X2=44.895 $Y2=4.705
r132 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=44.82 $Y=4.63
+ $X2=45.127 $Y2=4.28
r133 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=44.82 $Y=4.63
+ $X2=44.55 $Y2=4.63
r134 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=44.475 $Y=4.705
+ $X2=44.45 $Y2=4.63
r135 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=44.475 $Y=4.705
+ $X2=44.475 $Y2=4.995
r136 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=44.45 $Y=3.89
+ $X2=44.45 $Y2=3.405
r137 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=44.45 $Y=4.555
+ $X2=44.45 $Y2=4.63
r138 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=44.45 $Y=3.99 $X2=44.45
+ $Y2=3.89
r139 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=44.45 $Y=3.99
+ $X2=44.45 $Y2=4.555
r140 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=44.35 $Y=4.63
+ $X2=44.45 $Y2=4.63
r141 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=44.35 $Y=4.63
+ $X2=44.015 $Y2=4.63
r142 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=43.94 $Y=4.705
+ $X2=44.015 $Y2=4.63
r143 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=43.94 $Y=4.705
+ $X2=43.94 $Y2=5.185
r144 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.255 $Y=5.26
+ $X2=43.18 $Y2=5.26
r145 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=43.865 $Y=5.26
+ $X2=43.94 $Y2=5.185
r146 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=43.865 $Y=5.26
+ $X2=43.255 $Y2=5.26
r147 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.18 $Y=5.185
+ $X2=43.18 $Y2=5.26
r148 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=43.18 $Y=5.185
+ $X2=43.18 $Y2=4.85
r149 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.835 $Y=5.26
+ $X2=42.76 $Y2=5.26
r150 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=43.105 $Y=5.26
+ $X2=43.18 $Y2=5.26
r151 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=43.105 $Y=5.26
+ $X2=42.835 $Y2=5.26
r152 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.76 $Y=5.185
+ $X2=42.76 $Y2=5.26
r153 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=42.76 $Y=5.185
+ $X2=42.76 $Y2=4.85
r154 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.415 $Y=5.26
+ $X2=42.34 $Y2=5.26
r155 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.685 $Y=5.26
+ $X2=42.76 $Y2=5.26
r156 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=42.685 $Y=5.26
+ $X2=42.415 $Y2=5.26
r157 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.34 $Y=5.185
+ $X2=42.34 $Y2=5.26
r158 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=42.34 $Y=5.185
+ $X2=42.34 $Y2=4.85
r159 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=42.265 $Y=5.26
+ $X2=42.34 $Y2=5.26
r160 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=42.265 $Y=5.26
+ $X2=41.995 $Y2=5.26
r161 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=41.92 $Y=5.185
+ $X2=41.995 $Y2=5.26
r162 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=41.92 $Y=5.185
+ $X2=41.92 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[7] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c120 30 0 1.3204e-19 $X=48.32 $Y=0.255
r121 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=45.77 $Y=1.16
+ $X2=46.12 $Y2=1.16
r122 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=49.16 $Y=0.255
+ $X2=49.16 $Y2=0.59
r123 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.815 $Y=0.18
+ $X2=48.74 $Y2=0.18
r124 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=49.085 $Y=0.18
+ $X2=49.16 $Y2=0.255
r125 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=49.085 $Y=0.18
+ $X2=48.815 $Y2=0.18
r126 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.74 $Y=0.255
+ $X2=48.74 $Y2=0.18
r127 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=48.74 $Y=0.255
+ $X2=48.74 $Y2=0.59
r128 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.395 $Y=0.18
+ $X2=48.32 $Y2=0.18
r129 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.665 $Y=0.18
+ $X2=48.74 $Y2=0.18
r130 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=48.665 $Y=0.18
+ $X2=48.395 $Y2=0.18
r131 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.32 $Y=0.255
+ $X2=48.32 $Y2=0.18
r132 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=48.32 $Y=0.255
+ $X2=48.32 $Y2=0.59
r133 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.975 $Y=0.18
+ $X2=47.9 $Y2=0.18
r134 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.245 $Y=0.18
+ $X2=48.32 $Y2=0.18
r135 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=48.245 $Y=0.18
+ $X2=47.975 $Y2=0.18
r136 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.9 $Y=0.255
+ $X2=47.9 $Y2=0.18
r137 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=47.9 $Y=0.255
+ $X2=47.9 $Y2=0.59
r138 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.825 $Y=0.18
+ $X2=47.9 $Y2=0.18
r139 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=47.825 $Y=0.18
+ $X2=47.215 $Y2=0.18
r140 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=47.14 $Y=0.255
+ $X2=47.215 $Y2=0.18
r141 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=47.14 $Y=0.255
+ $X2=47.14 $Y2=0.735
r142 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.73 $Y=0.81
+ $X2=46.63 $Y2=0.81
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=47.065 $Y=0.81
+ $X2=47.14 $Y2=0.735
r144 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=47.065 $Y=0.81
+ $X2=46.73 $Y2=0.81
r145 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=46.63 $Y=1.55
+ $X2=46.63 $Y2=2.035
r146 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=46.63 $Y=1.45 $X2=46.63
+ $Y2=1.55
r147 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=46.63 $Y=0.885
+ $X2=46.63 $Y2=0.81
r148 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=46.63 $Y=0.885
+ $X2=46.63 $Y2=1.45
r149 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=46.605 $Y=0.735
+ $X2=46.63 $Y2=0.81
r150 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=46.605 $Y=0.735
+ $X2=46.605 $Y2=0.445
r151 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.26 $Y=0.81
+ $X2=46.16 $Y2=0.81
r152 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.53 $Y=0.81
+ $X2=46.63 $Y2=0.81
r153 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=46.53 $Y=0.81
+ $X2=46.26 $Y2=0.81
r154 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=46.185 $Y=0.735
+ $X2=46.16 $Y2=0.81
r155 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=46.185 $Y=0.735
+ $X2=46.185 $Y2=0.445
r156 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=46.16 $Y=1.55
+ $X2=46.16 $Y2=2.035
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=46.16 $Y=1.16
+ $X2=46.16 $Y2=1.55
r158 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=46.12
+ $Y=1.16 $X2=46.12 $Y2=1.16
r159 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=46.16 $Y=1.16
+ $X2=46.16 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[15] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c128 30 0 1.3204e-19 $X=48.32 $Y=5.185
r129 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=45.77 $Y=4.28
+ $X2=46.12 $Y2=4.28
r130 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=49.16 $Y=5.185
+ $X2=49.16 $Y2=4.85
r131 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.815 $Y=5.26
+ $X2=48.74 $Y2=5.26
r132 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=49.085 $Y=5.26
+ $X2=49.16 $Y2=5.185
r133 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=49.085 $Y=5.26
+ $X2=48.815 $Y2=5.26
r134 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.74 $Y=5.185
+ $X2=48.74 $Y2=5.26
r135 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=48.74 $Y=5.185
+ $X2=48.74 $Y2=4.85
r136 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.395 $Y=5.26
+ $X2=48.32 $Y2=5.26
r137 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.665 $Y=5.26
+ $X2=48.74 $Y2=5.26
r138 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=48.665 $Y=5.26
+ $X2=48.395 $Y2=5.26
r139 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.32 $Y=5.185
+ $X2=48.32 $Y2=5.26
r140 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=48.32 $Y=5.185
+ $X2=48.32 $Y2=4.85
r141 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.975 $Y=5.26
+ $X2=47.9 $Y2=5.26
r142 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=48.245 $Y=5.26
+ $X2=48.32 $Y2=5.26
r143 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=48.245 $Y=5.26
+ $X2=47.975 $Y2=5.26
r144 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.9 $Y=5.185
+ $X2=47.9 $Y2=5.26
r145 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=47.9 $Y=5.185
+ $X2=47.9 $Y2=4.85
r146 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=47.825 $Y=5.26
+ $X2=47.9 $Y2=5.26
r147 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=47.825 $Y=5.26
+ $X2=47.215 $Y2=5.26
r148 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=47.14 $Y=5.185
+ $X2=47.215 $Y2=5.26
r149 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=47.14 $Y=4.705
+ $X2=47.14 $Y2=5.185
r150 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.73 $Y=4.63
+ $X2=46.63 $Y2=4.63
r151 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=47.065 $Y=4.63
+ $X2=47.14 $Y2=4.705
r152 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=47.065 $Y=4.63
+ $X2=46.73 $Y2=4.63
r153 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=46.63 $Y=3.89
+ $X2=46.63 $Y2=3.405
r154 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=46.605 $Y=4.705
+ $X2=46.63 $Y2=4.63
r155 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=46.605 $Y=4.705
+ $X2=46.605 $Y2=4.995
r156 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=46.63 $Y=4.555
+ $X2=46.63 $Y2=4.63
r157 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=46.63 $Y=3.99 $X2=46.63
+ $Y2=3.89
r158 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=46.63 $Y=3.99
+ $X2=46.63 $Y2=4.555
r159 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.26 $Y=4.63
+ $X2=46.16 $Y2=4.63
r160 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=46.53 $Y=4.63
+ $X2=46.63 $Y2=4.63
r161 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=46.53 $Y=4.63
+ $X2=46.26 $Y2=4.63
r162 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=46.185 $Y=4.705
+ $X2=46.16 $Y2=4.63
r163 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=46.185 $Y=4.705
+ $X2=46.185 $Y2=4.995
r164 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=46.16 $Y=3.89
+ $X2=46.16 $Y2=3.405
r165 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=46.16 $Y=4.28
+ $X2=46.16 $Y2=4.63
r166 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=46.12
+ $Y=4.28 $X2=46.12 $Y2=4.28
r167 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=46.16 $Y=4.28
+ $X2=46.16 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c115 22 0 9.37986e-20 $X=49.085 $Y=1.475
c116 17 0 9.37986e-20 $X=48.615 $Y=1.475
c117 12 0 9.37986e-20 $X=48.145 $Y=1.475
c118 7 0 9.37986e-20 $X=47.675 $Y=1.475
r119 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=47.445
+ $Y=1.285 $X2=47.355 $Y2=1.23
r120 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=47.445
+ $Y=1.23 $X2=47.445 $Y2=1.23
r121 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=47.105 $Y=1.23
+ $X2=47.355 $Y2=1.23
r122 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=47.105 $Y=1.23
+ $X2=47.445 $Y2=1.23
r123 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=47.105
+ $Y=1.23 $X2=47.105 $Y2=1.23
r124 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=46.56 $Y=1.23
+ $X2=46.475 $Y2=1.23
r125 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=46.56 $Y=1.23
+ $X2=47.105 $Y2=1.23
r126 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=46.475 $Y=1.395
+ $X2=46.475 $Y2=1.23
r127 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=46.475 $Y=1.395
+ $X2=46.475 $Y2=1.605
r128 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=46.475 $Y=1.065
+ $X2=46.475 $Y2=1.23
r129 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=46.475 $Y=1.065
+ $X2=46.475 $Y2=0.825
r130 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=46.435 $Y=0.7
+ $X2=46.435 $Y2=0.825
r131 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=46.435 $Y=0.7
+ $X2=46.435 $Y2=0.445
r132 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=46.395 $Y=1.77
+ $X2=46.395 $Y2=1.605
r133 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=49.085 $Y=1.475
+ $X2=49.085 $Y2=1.965
r134 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.705 $Y=1.4
+ $X2=48.615 $Y2=1.4
r135 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=48.995 $Y=1.4
+ $X2=49.085 $Y2=1.475
r136 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.995 $Y=1.4
+ $X2=48.705 $Y2=1.4
r137 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=48.615 $Y=1.475
+ $X2=48.615 $Y2=1.4
r138 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=48.615 $Y=1.475
+ $X2=48.615 $Y2=1.965
r139 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.235 $Y=1.4
+ $X2=48.145 $Y2=1.4
r140 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.525 $Y=1.4
+ $X2=48.615 $Y2=1.4
r141 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.525 $Y=1.4
+ $X2=48.235 $Y2=1.4
r142 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=48.145 $Y=1.475
+ $X2=48.145 $Y2=1.4
r143 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=48.145 $Y=1.475
+ $X2=48.145 $Y2=1.965
r144 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.055 $Y=1.4
+ $X2=48.145 $Y2=1.4
r145 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.055 $Y=1.4
+ $X2=47.765 $Y2=1.4
r146 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=47.675 $Y=1.475
+ $X2=47.765 $Y2=1.4
r147 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=47.675 $Y=1.475
+ $X2=47.445 $Y2=1.285
r148 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=47.675 $Y=1.475
+ $X2=47.675 $Y2=1.965
r149 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=46.25
+ $Y=1.625 $X2=46.395 $Y2=1.77
r150 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=46.26
+ $Y=0.235 $X2=46.395 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_599# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c121 22 0 9.37986e-20 $X=49.085 $Y=3.965
c122 17 0 9.37986e-20 $X=48.615 $Y=3.965
c123 12 0 9.37986e-20 $X=48.145 $Y=3.965
c124 7 0 9.37986e-20 $X=47.675 $Y=3.965
r125 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=47.445
+ $Y=4.155 $X2=47.355 $Y2=4.21
r126 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=47.445
+ $Y=4.21 $X2=47.445 $Y2=4.21
r127 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=47.105 $Y=4.21
+ $X2=47.355 $Y2=4.21
r128 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=47.105 $Y=4.21
+ $X2=47.445 $Y2=4.21
r129 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=47.105
+ $Y=4.21 $X2=47.105 $Y2=4.21
r130 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=46.56 $Y=4.21
+ $X2=46.475 $Y2=4.21
r131 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=46.56 $Y=4.21
+ $X2=47.105 $Y2=4.21
r132 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=46.475 $Y=4.375
+ $X2=46.475 $Y2=4.21
r133 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=46.475 $Y=4.375
+ $X2=46.475 $Y2=4.615
r134 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=46.475 $Y=4.045
+ $X2=46.475 $Y2=4.21
r135 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=46.475 $Y=4.045
+ $X2=46.475 $Y2=3.835
r136 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=46.435 $Y=4.74
+ $X2=46.435 $Y2=4.615
r137 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=46.435 $Y=4.74
+ $X2=46.435 $Y2=4.995
r138 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=46.395 $Y=3.67
+ $X2=46.395 $Y2=3.835
r139 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=46.395 $Y=3.67
+ $X2=46.395 $Y2=3.14
r140 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=49.085 $Y=3.965
+ $X2=49.085 $Y2=3.475
r141 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.705 $Y=4.04
+ $X2=48.615 $Y2=4.04
r142 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=48.995 $Y=4.04
+ $X2=49.085 $Y2=3.965
r143 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.995 $Y=4.04
+ $X2=48.705 $Y2=4.04
r144 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=48.615 $Y=3.965
+ $X2=48.615 $Y2=4.04
r145 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=48.615 $Y=3.965
+ $X2=48.615 $Y2=3.475
r146 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.235 $Y=4.04
+ $X2=48.145 $Y2=4.04
r147 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.525 $Y=4.04
+ $X2=48.615 $Y2=4.04
r148 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.525 $Y=4.04
+ $X2=48.235 $Y2=4.04
r149 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=48.145 $Y=3.965
+ $X2=48.145 $Y2=4.04
r150 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=48.145 $Y=3.965
+ $X2=48.145 $Y2=3.475
r151 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=48.055 $Y=4.04
+ $X2=48.145 $Y2=4.04
r152 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=48.055 $Y=4.04
+ $X2=47.765 $Y2=4.04
r153 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=47.675 $Y=3.965
+ $X2=47.765 $Y2=4.04
r154 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=47.675 $Y=3.965
+ $X2=47.445 $Y2=4.155
r155 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=47.675 $Y=3.965
+ $X2=47.675 $Y2=3.475
r156 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=46.25
+ $Y=2.995 $X2=46.395 $Y2=3.14
r157 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=46.26
+ $Y=4.785 $X2=46.395 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[7] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r88 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=51.46 $Y=1.16
+ $X2=51.485 $Y2=1.16
r89 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=51.38 $Y=1.16
+ $X2=51.46 $Y2=1.16
r90 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=51.38
+ $Y=1.16 $X2=51.38 $Y2=1.16
r91 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=51.04 $Y=1.16
+ $X2=51.38 $Y2=1.16
r92 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=51.015 $Y=1.16
+ $X2=51.04 $Y2=1.16
r93 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=50.52 $Y=1.16
+ $X2=50.545 $Y2=1.16
r94 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=50.36 $Y=1.16
+ $X2=50.52 $Y2=1.16
r95 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=50.36
+ $Y=1.16 $X2=50.36 $Y2=1.16
r96 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=50.1 $Y=1.16
+ $X2=50.36 $Y2=1.16
r97 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=50.075 $Y=1.16
+ $X2=50.1 $Y2=1.16
r98 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=50.7 $Y=1.19
+ $X2=50.36 $Y2=1.19
r99 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=50.7
+ $Y=1.16 $X2=50.7 $Y2=1.16
r100 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=50.635 $Y=1.16
+ $X2=50.545 $Y2=1.16
r101 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=50.635 $Y=1.16
+ $X2=50.7 $Y2=1.16
r102 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=50.925 $Y=1.16
+ $X2=51.015 $Y2=1.16
r103 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=50.925 $Y=1.16
+ $X2=50.7 $Y2=1.16
r104 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=51.29 $Y=1.19
+ $X2=51.38 $Y2=1.19
r105 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=51.29 $Y=1.19
+ $X2=50.7 $Y2=1.19
r106 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=51.485 $Y=1.295
+ $X2=51.485 $Y2=1.16
r107 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=51.485 $Y=1.295
+ $X2=51.485 $Y2=1.985
r108 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=51.46 $Y=1.025
+ $X2=51.46 $Y2=1.16
r109 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=51.46 $Y=1.025
+ $X2=51.46 $Y2=0.56
r110 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=51.04 $Y=1.025
+ $X2=51.04 $Y2=1.16
r111 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=51.04 $Y=1.025
+ $X2=51.04 $Y2=0.56
r112 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=51.015 $Y=1.295
+ $X2=51.015 $Y2=1.16
r113 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=51.015 $Y=1.295
+ $X2=51.015 $Y2=1.985
r114 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=50.545 $Y=1.295
+ $X2=50.545 $Y2=1.16
r115 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=50.545 $Y=1.295
+ $X2=50.545 $Y2=1.985
r116 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=50.52 $Y=1.025
+ $X2=50.52 $Y2=1.16
r117 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=50.52 $Y=1.025
+ $X2=50.52 $Y2=0.56
r118 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=50.1 $Y=1.025
+ $X2=50.1 $Y2=1.16
r119 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=50.1 $Y=1.025
+ $X2=50.1 $Y2=0.56
r120 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=50.075 $Y=1.295
+ $X2=50.075 $Y2=1.16
r121 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=50.075 $Y=1.295
+ $X2=50.075 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[15] 3 7 11 15 19 23 27 31 33 35 36
+ 52 54
r86 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=51.46 $Y=4.28
+ $X2=51.485 $Y2=4.28
r87 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=51.38 $Y=4.28
+ $X2=51.46 $Y2=4.28
r88 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=51.38
+ $Y=4.28 $X2=51.38 $Y2=4.28
r89 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=51.04 $Y=4.28
+ $X2=51.38 $Y2=4.28
r90 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=51.015 $Y=4.28
+ $X2=51.04 $Y2=4.28
r91 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=50.52 $Y=4.28
+ $X2=50.545 $Y2=4.28
r92 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=50.36 $Y=4.28
+ $X2=50.52 $Y2=4.28
r93 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=50.36
+ $Y=4.28 $X2=50.36 $Y2=4.28
r94 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=50.1 $Y=4.28
+ $X2=50.36 $Y2=4.28
r95 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=50.075 $Y=4.28
+ $X2=50.1 $Y2=4.28
r96 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=50.7 $Y=4.25
+ $X2=50.36 $Y2=4.25
r97 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=50.7
+ $Y=4.28 $X2=50.7 $Y2=4.28
r98 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=50.635 $Y=4.28
+ $X2=50.545 $Y2=4.28
r99 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=50.635 $Y=4.28
+ $X2=50.7 $Y2=4.28
r100 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=50.925 $Y=4.28
+ $X2=51.015 $Y2=4.28
r101 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=50.925 $Y=4.28
+ $X2=50.7 $Y2=4.28
r102 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=51.29 $Y=4.25
+ $X2=51.38 $Y2=4.25
r103 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=51.29 $Y=4.25
+ $X2=50.7 $Y2=4.25
r104 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=51.485 $Y=4.145
+ $X2=51.485 $Y2=4.28
r105 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=51.485 $Y=4.145
+ $X2=51.485 $Y2=3.455
r106 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=51.46 $Y=4.415
+ $X2=51.46 $Y2=4.28
r107 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=51.46 $Y=4.415
+ $X2=51.46 $Y2=4.88
r108 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=51.04 $Y=4.415
+ $X2=51.04 $Y2=4.28
r109 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=51.04 $Y=4.415
+ $X2=51.04 $Y2=4.88
r110 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=51.015 $Y=4.145
+ $X2=51.015 $Y2=4.28
r111 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=51.015 $Y=4.145
+ $X2=51.015 $Y2=3.455
r112 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=50.545 $Y=4.145
+ $X2=50.545 $Y2=4.28
r113 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=50.545 $Y=4.145
+ $X2=50.545 $Y2=3.455
r114 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=50.52 $Y=4.415
+ $X2=50.52 $Y2=4.28
r115 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=50.52 $Y=4.415
+ $X2=50.52 $Y2=4.88
r116 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=50.1 $Y=4.415
+ $X2=50.1 $Y2=4.28
r117 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=50.1 $Y=4.415
+ $X2=50.1 $Y2=4.88
r118 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=50.075 $Y=4.145
+ $X2=50.075 $Y2=4.28
r119 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=50.075 $Y=4.145
+ $X2=50.075 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 243 249 255 259 261 265 269 273 277
+ 281 285 287 291 295 299 303 307 311 315 319 323 329 333 337 343 349 353 355
+ 359 363 367 371 375 379 381 385 389 393 397 401 405 409 413 417 423 429 435
+ 441 445 447 451 455 459 463 467 471 473 477 481 485 489 493 497 501 505 509
+ 515 519 523 529 535 539 541 545 549 553 557 561 565 567 571 575 579 583 587
+ 591 595 599 603 609 614 615 616 617 618 619 620 622 623 625 626 627 628 629
+ 630 631 633 634 636 637 638 639 640 641 642 644 645 647 648 649 650 651 652
+ 653 655 656 657 658 659 660 661 662 663 664 665 675 682 702 706 711 718 738
+ 742 747 752 759 779 783 788 795 815 819 825 828 831 834 837 840 843 846 849
+ 852 855 858 861 864 867 870 873 876 879 882 885 888 891 894
c1554 819 0 3.95698e-19 $X=51.585 $Y=2.72
c1555 815 0 3.95698e-19 $X=50.645 $Y=2.72
c1556 795 0 3.94334e-19 $X=41.63 $Y=2.72
c1557 788 0 3.95698e-19 $X=40.165 $Y=2.72
c1558 783 0 3.95698e-19 $X=38.705 $Y=2.72
c1559 779 0 3.95698e-19 $X=37.765 $Y=2.72
c1560 759 0 3.94334e-19 $X=28.75 $Y=2.72
c1561 752 0 3.95698e-19 $X=27.285 $Y=2.72
c1562 742 0 3.95698e-19 $X=25.365 $Y=2.72
c1563 738 0 3.95698e-19 $X=24.425 $Y=2.72
c1564 718 0 3.94334e-19 $X=15.41 $Y=2.72
c1565 711 0 3.95698e-19 $X=13.945 $Y=2.72
c1566 706 0 3.95698e-19 $X=12.485 $Y=2.72
c1567 702 0 3.95698e-19 $X=11.545 $Y=2.72
c1568 682 0 3.94334e-19 $X=2.53 $Y=2.72
c1569 675 0 3.95698e-19 $X=1.065 $Y=2.72
c1570 655 0 3.94334e-19 $X=49.705 $Y=2.72
c1571 651 0 3.94334e-19 $X=47.03 $Y=2.72
c1572 647 0 3.94334e-19 $X=44.05 $Y=2.72
c1573 644 0 3.94334e-19 $X=36.825 $Y=2.72
c1574 640 0 3.94334e-19 $X=34.15 $Y=2.72
c1575 636 0 3.94334e-19 $X=31.17 $Y=2.72
c1576 633 0 3.94334e-19 $X=23.485 $Y=2.72
c1577 629 0 3.94334e-19 $X=20.81 $Y=2.72
c1578 625 0 3.94334e-19 $X=17.83 $Y=2.72
c1579 622 0 3.94334e-19 $X=10.605 $Y=2.72
c1580 618 0 3.94334e-19 $X=7.93 $Y=2.72
c1581 614 0 3.94334e-19 $X=4.95 $Y=2.72
c1582 541 0 3.95698e-19 $X=41.105 $Y=2.72
c1583 447 0 3.95698e-19 $X=28.225 $Y=2.72
c1584 355 0 3.95698e-19 $X=14.885 $Y=2.72
c1585 261 0 3.95698e-19 $X=2.005 $Y=2.72
c1586 76 0 1.36925e-19 $X=49.715 $Y=2.955
c1587 75 0 1.36925e-19 $X=49.715 $Y=1.485
c1588 66 0 9.57576e-20 $X=41.095 $Y=2.955
c1589 65 0 9.57576e-20 $X=41.095 $Y=1.485
c1590 64 0 1.91515e-19 $X=40.155 $Y=2.955
c1591 63 0 1.91515e-19 $X=40.155 $Y=1.485
c1592 58 0 1.91515e-19 $X=37.755 $Y=2.955
c1593 57 0 1.91515e-19 $X=37.755 $Y=1.485
c1594 56 0 9.57576e-20 $X=36.835 $Y=2.955
c1595 55 0 9.57576e-20 $X=36.835 $Y=1.485
c1596 46 0 9.57576e-20 $X=28.215 $Y=2.955
c1597 45 0 9.57576e-20 $X=28.215 $Y=1.485
c1598 44 0 1.91515e-19 $X=27.275 $Y=2.955
c1599 43 0 1.91515e-19 $X=27.275 $Y=1.485
c1600 38 0 1.91515e-19 $X=24.415 $Y=2.955
c1601 37 0 1.91515e-19 $X=24.415 $Y=1.485
c1602 36 0 9.57576e-20 $X=23.495 $Y=2.955
c1603 35 0 9.57576e-20 $X=23.495 $Y=1.485
c1604 26 0 9.57576e-20 $X=14.875 $Y=2.955
c1605 25 0 9.57576e-20 $X=14.875 $Y=1.485
c1606 24 0 1.91515e-19 $X=13.935 $Y=2.955
c1607 23 0 1.91515e-19 $X=13.935 $Y=1.485
c1608 18 0 1.91515e-19 $X=11.535 $Y=2.955
c1609 17 0 1.91515e-19 $X=11.535 $Y=1.485
c1610 16 0 9.57576e-20 $X=10.615 $Y=2.955
c1611 15 0 9.57576e-20 $X=10.615 $Y=1.485
c1612 6 0 1.36925e-19 $X=1.995 $Y=2.955
c1613 5 0 1.36925e-19 $X=1.995 $Y=1.485
r1614 891 892 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=50.83 $Y=2.72
+ $X2=50.83 $Y2=2.72
r1615 888 889 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=45.77 $Y=2.72
+ $X2=45.77 $Y2=2.72
r1616 885 886 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=41.17 $Y=2.72
+ $X2=41.17 $Y2=2.72
r1617 883 886 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=40.25 $Y=2.72
+ $X2=41.17 $Y2=2.72
r1618 882 883 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=40.25 $Y=2.72
+ $X2=40.25 $Y2=2.72
r1619 873 874 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=37.95 $Y=2.72
+ $X2=37.95 $Y2=2.72
r1620 870 871 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=32.89 $Y=2.72
+ $X2=32.89 $Y2=2.72
r1621 867 868 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=28.29 $Y=2.72
+ $X2=28.29 $Y2=2.72
r1622 865 868 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=27.37 $Y=2.72
+ $X2=28.29 $Y2=2.72
r1623 864 865 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.37 $Y=2.72
+ $X2=27.37 $Y2=2.72
r1624 855 856 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1625 852 853 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1626 849 850 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r1627 847 850 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.95 $Y2=2.72
r1628 846 847 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r1629 837 838 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1630 834 835 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1631 831 832 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r1632 829 832 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r1633 828 829 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r1634 823 892 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.29 $Y=2.72
+ $X2=50.83 $Y2=2.72
r1635 822 823 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.29 $Y=2.72
+ $X2=51.29 $Y2=2.72
r1636 820 891 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.915 $Y=2.72
+ $X2=50.78 $Y2=2.72
r1637 820 822 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=50.915 $Y=2.72
+ $X2=51.29 $Y2=2.72
r1638 819 894 3.05049 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=51.585 $Y=2.72
+ $X2=51.782 $Y2=2.72
r1639 819 822 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=51.585 $Y=2.72
+ $X2=51.29 $Y2=2.72
r1640 818 892 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=50.37 $Y=2.72
+ $X2=50.83 $Y2=2.72
r1641 817 818 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=50.37 $Y=2.72
+ $X2=50.37 $Y2=2.72
r1642 815 891 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.645 $Y=2.72
+ $X2=50.78 $Y2=2.72
r1643 815 817 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=50.645 $Y=2.72
+ $X2=50.37 $Y2=2.72
r1644 813 818 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=49.45 $Y=2.72
+ $X2=50.37 $Y2=2.72
r1645 812 813 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=49.45 $Y=2.72
+ $X2=49.45 $Y2=2.72
r1646 810 813 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=47.15 $Y=2.72
+ $X2=49.45 $Y2=2.72
r1647 809 810 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=47.15 $Y=2.72
+ $X2=47.15 $Y2=2.72
r1648 807 810 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=46.69 $Y=2.72
+ $X2=47.15 $Y2=2.72
r1649 807 889 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=46.69 $Y=2.72
+ $X2=45.77 $Y2=2.72
r1650 806 807 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=46.69 $Y=2.72
+ $X2=46.69 $Y2=2.72
r1651 804 888 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=46.06 $Y=2.72
+ $X2=45.91 $Y2=2.72
r1652 804 806 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=46.06 $Y=2.72
+ $X2=46.69 $Y2=2.72
r1653 803 889 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=44.85 $Y=2.72
+ $X2=45.77 $Y2=2.72
r1654 802 803 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=44.85 $Y=2.72
+ $X2=44.85 $Y2=2.72
r1655 800 803 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=43.93 $Y=2.72
+ $X2=44.85 $Y2=2.72
r1656 799 800 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=43.93 $Y=2.72
+ $X2=43.93 $Y2=2.72
r1657 796 800 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=41.63 $Y=2.72
+ $X2=43.93 $Y2=2.72
r1658 796 886 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=41.63 $Y=2.72
+ $X2=41.17 $Y2=2.72
r1659 795 796 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=41.63 $Y=2.72
+ $X2=41.63 $Y2=2.72
r1660 793 885 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=41.375 $Y=2.72
+ $X2=41.24 $Y2=2.72
r1661 793 795 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=41.375 $Y=2.72
+ $X2=41.63 $Y2=2.72
r1662 792 883 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.79 $Y=2.72
+ $X2=40.25 $Y2=2.72
r1663 791 792 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.79 $Y=2.72
+ $X2=39.79 $Y2=2.72
r1664 789 879 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=39.495 $Y=2.72
+ $X2=39.36 $Y2=2.72
r1665 789 791 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=39.495 $Y=2.72
+ $X2=39.79 $Y2=2.72
r1666 788 882 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.165 $Y=2.72
+ $X2=40.3 $Y2=2.72
r1667 788 791 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=40.165 $Y=2.72
+ $X2=39.79 $Y2=2.72
r1668 787 874 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.41 $Y=2.72
+ $X2=37.95 $Y2=2.72
r1669 786 787 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.41 $Y=2.72
+ $X2=38.41 $Y2=2.72
r1670 784 873 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=38.035 $Y=2.72
+ $X2=37.9 $Y2=2.72
r1671 784 786 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=38.035 $Y=2.72
+ $X2=38.41 $Y2=2.72
r1672 783 876 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=38.705 $Y=2.72
+ $X2=38.84 $Y2=2.72
r1673 783 786 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=38.705 $Y=2.72
+ $X2=38.41 $Y2=2.72
r1674 782 874 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=37.49 $Y=2.72
+ $X2=37.95 $Y2=2.72
r1675 781 782 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=37.49 $Y=2.72
+ $X2=37.49 $Y2=2.72
r1676 779 873 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=37.765 $Y=2.72
+ $X2=37.9 $Y2=2.72
r1677 779 781 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=37.765 $Y=2.72
+ $X2=37.49 $Y2=2.72
r1678 777 782 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=36.57 $Y=2.72
+ $X2=37.49 $Y2=2.72
r1679 776 777 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=36.57 $Y=2.72
+ $X2=36.57 $Y2=2.72
r1680 774 777 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=34.27 $Y=2.72
+ $X2=36.57 $Y2=2.72
r1681 773 774 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=34.27 $Y=2.72
+ $X2=34.27 $Y2=2.72
r1682 771 774 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=33.81 $Y=2.72
+ $X2=34.27 $Y2=2.72
r1683 771 871 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=33.81 $Y=2.72
+ $X2=32.89 $Y2=2.72
r1684 770 771 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=33.81 $Y=2.72
+ $X2=33.81 $Y2=2.72
r1685 768 870 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=33.18 $Y=2.72
+ $X2=33.03 $Y2=2.72
r1686 768 770 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=33.18 $Y=2.72
+ $X2=33.81 $Y2=2.72
r1687 767 871 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.97 $Y=2.72
+ $X2=32.89 $Y2=2.72
r1688 766 767 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=31.97 $Y=2.72
+ $X2=31.97 $Y2=2.72
r1689 764 767 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.05 $Y=2.72
+ $X2=31.97 $Y2=2.72
r1690 763 764 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=31.05 $Y=2.72
+ $X2=31.05 $Y2=2.72
r1691 760 764 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=28.75 $Y=2.72
+ $X2=31.05 $Y2=2.72
r1692 760 868 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=28.75 $Y=2.72
+ $X2=28.29 $Y2=2.72
r1693 759 760 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=28.75 $Y=2.72
+ $X2=28.75 $Y2=2.72
r1694 757 867 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=28.495 $Y=2.72
+ $X2=28.36 $Y2=2.72
r1695 757 759 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=28.495 $Y=2.72
+ $X2=28.75 $Y2=2.72
r1696 756 865 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.91 $Y=2.72
+ $X2=27.37 $Y2=2.72
r1697 755 756 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.91 $Y=2.72
+ $X2=26.91 $Y2=2.72
r1698 753 861 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=26.615 $Y=2.72
+ $X2=26.48 $Y2=2.72
r1699 753 755 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=26.615 $Y=2.72
+ $X2=26.91 $Y2=2.72
r1700 752 864 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.285 $Y=2.72
+ $X2=27.42 $Y2=2.72
r1701 752 755 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=27.285 $Y=2.72
+ $X2=26.91 $Y2=2.72
r1702 748 858 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=25.635 $Y=2.72
+ $X2=25.5 $Y2=2.72
r1703 748 750 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=25.635 $Y=2.72
+ $X2=25.99 $Y2=2.72
r1704 747 861 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=26.345 $Y=2.72
+ $X2=26.48 $Y2=2.72
r1705 747 750 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=26.345 $Y=2.72
+ $X2=25.99 $Y2=2.72
r1706 746 856 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.07 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1707 745 746 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1708 743 855 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.695 $Y=2.72
+ $X2=24.56 $Y2=2.72
r1709 743 745 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=24.695 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1710 742 858 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=25.365 $Y=2.72
+ $X2=25.5 $Y2=2.72
r1711 742 745 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.365 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1712 741 856 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=2.72
+ $X2=24.61 $Y2=2.72
r1713 740 741 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=2.72
+ $X2=24.15 $Y2=2.72
r1714 738 855 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.425 $Y=2.72
+ $X2=24.56 $Y2=2.72
r1715 738 740 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=24.425 $Y=2.72
+ $X2=24.15 $Y2=2.72
r1716 736 741 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=2.72
+ $X2=24.15 $Y2=2.72
r1717 735 736 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.23 $Y=2.72
+ $X2=23.23 $Y2=2.72
r1718 733 736 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=2.72
+ $X2=23.23 $Y2=2.72
r1719 732 733 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.93 $Y=2.72
+ $X2=20.93 $Y2=2.72
r1720 730 733 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=20.93 $Y2=2.72
r1721 730 853 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1722 729 730 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=2.72
+ $X2=20.47 $Y2=2.72
r1723 727 852 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.84 $Y=2.72
+ $X2=19.69 $Y2=2.72
r1724 727 729 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=19.84 $Y=2.72
+ $X2=20.47 $Y2=2.72
r1725 726 853 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=18.63 $Y=2.72
+ $X2=19.55 $Y2=2.72
r1726 725 726 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1727 723 726 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.71 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1728 722 723 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=2.72
+ $X2=17.71 $Y2=2.72
r1729 719 723 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=17.71 $Y2=2.72
r1730 719 850 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=14.95 $Y2=2.72
r1731 718 719 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r1732 716 849 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.155 $Y=2.72
+ $X2=15.02 $Y2=2.72
r1733 716 718 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=15.155 $Y=2.72
+ $X2=15.41 $Y2=2.72
r1734 715 847 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r1735 714 715 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1736 712 843 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.275 $Y=2.72
+ $X2=13.14 $Y2=2.72
r1737 712 714 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.275 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1738 711 846 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.945 $Y=2.72
+ $X2=14.08 $Y2=2.72
r1739 711 714 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.945 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1740 710 838 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1741 709 710 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1742 707 837 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=11.68 $Y2=2.72
r1743 707 709 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1744 706 840 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.485 $Y=2.72
+ $X2=12.62 $Y2=2.72
r1745 706 709 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.485 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1746 705 838 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r1747 704 705 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r1748 702 837 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.545 $Y=2.72
+ $X2=11.68 $Y2=2.72
r1749 702 704 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.545 $Y=2.72
+ $X2=11.27 $Y2=2.72
r1750 700 705 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r1751 699 700 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r1752 697 700 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r1753 696 697 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r1754 694 697 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r1755 694 835 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1756 693 694 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r1757 691 834 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=6.81 $Y2=2.72
r1758 691 693 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=7.59 $Y2=2.72
r1759 690 835 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r1760 689 690 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1761 687 690 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1762 686 687 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r1763 683 687 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r1764 683 832 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r1765 682 683 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r1766 680 831 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r1767 680 682 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.53 $Y2=2.72
r1768 679 829 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r1769 678 679 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1770 676 825 3.05049 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r1771 676 678 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1772 675 828 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r1773 675 678 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1774 665 823 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.75 $Y=2.72
+ $X2=51.29 $Y2=2.72
r1775 665 894 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.75 $Y=2.72
+ $X2=51.75 $Y2=2.72
r1776 664 792 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.33 $Y=2.72
+ $X2=39.79 $Y2=2.72
r1777 664 879 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.33 $Y=2.72
+ $X2=39.33 $Y2=2.72
r1778 663 664 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=2.72
+ $X2=39.33 $Y2=2.72
r1779 663 787 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=2.72
+ $X2=38.41 $Y2=2.72
r1780 663 876 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.87 $Y=2.72
+ $X2=38.87 $Y2=2.72
r1781 662 756 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.45 $Y=2.72
+ $X2=26.91 $Y2=2.72
r1782 662 861 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.45 $Y=2.72
+ $X2=26.45 $Y2=2.72
r1783 661 662 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.99 $Y=2.72
+ $X2=26.45 $Y2=2.72
r1784 661 750 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.99 $Y=2.72
+ $X2=25.99 $Y2=2.72
r1785 660 661 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=2.72
+ $X2=25.99 $Y2=2.72
r1786 660 746 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=2.72
+ $X2=25.07 $Y2=2.72
r1787 660 858 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=2.72
+ $X2=25.53 $Y2=2.72
r1788 659 715 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r1789 659 843 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1790 658 659 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r1791 658 710 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r1792 658 840 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r1793 657 679 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r1794 657 825 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r1795 655 812 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=49.705 $Y=2.72
+ $X2=49.45 $Y2=2.72
r1796 655 656 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=49.705 $Y=2.72
+ $X2=49.84 $Y2=2.72
r1797 654 817 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=49.975 $Y=2.72
+ $X2=50.37 $Y2=2.72
r1798 654 656 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=49.975 $Y=2.72
+ $X2=49.84 $Y2=2.72
r1799 652 806 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=46.755 $Y=2.72
+ $X2=46.69 $Y2=2.72
r1800 652 653 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=46.755 $Y=2.72
+ $X2=46.892 $Y2=2.72
r1801 651 809 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=47.03 $Y=2.72
+ $X2=47.15 $Y2=2.72
r1802 651 653 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=47.03 $Y=2.72
+ $X2=46.892 $Y2=2.72
r1803 649 802 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=45.02 $Y=2.72
+ $X2=44.85 $Y2=2.72
r1804 649 650 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=45.02 $Y=2.72
+ $X2=45.17 $Y2=2.72
r1805 647 799 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=44.05 $Y=2.72
+ $X2=43.93 $Y2=2.72
r1806 647 648 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=44.05 $Y=2.72
+ $X2=44.187 $Y2=2.72
r1807 646 802 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=44.325 $Y=2.72
+ $X2=44.85 $Y2=2.72
r1808 646 648 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=44.325 $Y=2.72
+ $X2=44.187 $Y2=2.72
r1809 644 776 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=36.825 $Y=2.72
+ $X2=36.57 $Y2=2.72
r1810 644 645 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=36.825 $Y=2.72
+ $X2=36.96 $Y2=2.72
r1811 643 781 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=37.095 $Y=2.72
+ $X2=37.49 $Y2=2.72
r1812 643 645 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=37.095 $Y=2.72
+ $X2=36.96 $Y2=2.72
r1813 641 770 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=33.875 $Y=2.72
+ $X2=33.81 $Y2=2.72
r1814 641 642 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=33.875 $Y=2.72
+ $X2=34.012 $Y2=2.72
r1815 640 773 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=34.15 $Y=2.72
+ $X2=34.27 $Y2=2.72
r1816 640 642 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=34.15 $Y=2.72
+ $X2=34.012 $Y2=2.72
r1817 638 766 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=32.14 $Y=2.72
+ $X2=31.97 $Y2=2.72
r1818 638 639 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=32.14 $Y=2.72
+ $X2=32.29 $Y2=2.72
r1819 636 763 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=31.17 $Y=2.72
+ $X2=31.05 $Y2=2.72
r1820 636 637 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=31.17 $Y=2.72
+ $X2=31.307 $Y2=2.72
r1821 635 766 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=31.445 $Y=2.72
+ $X2=31.97 $Y2=2.72
r1822 635 637 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=31.445 $Y=2.72
+ $X2=31.307 $Y2=2.72
r1823 633 735 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=23.485 $Y=2.72
+ $X2=23.23 $Y2=2.72
r1824 633 634 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=23.485 $Y=2.72
+ $X2=23.62 $Y2=2.72
r1825 632 740 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=23.755 $Y=2.72
+ $X2=24.15 $Y2=2.72
r1826 632 634 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=23.755 $Y=2.72
+ $X2=23.62 $Y2=2.72
r1827 630 729 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=20.535 $Y=2.72
+ $X2=20.47 $Y2=2.72
r1828 630 631 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=20.535 $Y=2.72
+ $X2=20.672 $Y2=2.72
r1829 629 732 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=20.81 $Y=2.72
+ $X2=20.93 $Y2=2.72
r1830 629 631 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=20.81 $Y=2.72
+ $X2=20.672 $Y2=2.72
r1831 627 725 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=18.8 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1832 627 628 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.8 $Y=2.72
+ $X2=18.95 $Y2=2.72
r1833 625 722 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=17.83 $Y=2.72
+ $X2=17.71 $Y2=2.72
r1834 625 626 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=17.83 $Y=2.72
+ $X2=17.967 $Y2=2.72
r1835 624 725 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=18.105 $Y=2.72
+ $X2=18.63 $Y2=2.72
r1836 624 626 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=18.105 $Y=2.72
+ $X2=17.967 $Y2=2.72
r1837 622 699 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.605 $Y=2.72
+ $X2=10.35 $Y2=2.72
r1838 622 623 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.605 $Y=2.72
+ $X2=10.74 $Y2=2.72
r1839 621 704 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=11.27 $Y2=2.72
r1840 621 623 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=10.74 $Y2=2.72
r1841 619 693 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.655 $Y=2.72
+ $X2=7.59 $Y2=2.72
r1842 619 620 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.655 $Y=2.72
+ $X2=7.792 $Y2=2.72
r1843 618 696 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.93 $Y=2.72
+ $X2=8.05 $Y2=2.72
r1844 618 620 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=7.93 $Y=2.72
+ $X2=7.792 $Y2=2.72
r1845 616 689 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1846 616 617 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.07 $Y2=2.72
r1847 614 686 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=4.83 $Y2=2.72
r1848 614 615 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=5.087 $Y2=2.72
r1849 613 689 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.75 $Y2=2.72
r1850 613 615 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.087 $Y2=2.72
r1851 609 611 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=51.72 $Y=3.1
+ $X2=51.72 $Y2=3.78
r1852 607 894 3.46198 $w=2.7e-07 $l=1.11781e-07 $layer=LI1_cond $X=51.72
+ $Y=2.805 $X2=51.782 $Y2=2.72
r1853 607 609 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=51.72 $Y=2.805
+ $X2=51.72 $Y2=3.1
r1854 603 606 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=51.72 $Y=1.66
+ $X2=51.72 $Y2=2.34
r1855 601 894 3.46198 $w=2.7e-07 $l=1.11781e-07 $layer=LI1_cond $X=51.72
+ $Y=2.635 $X2=51.782 $Y2=2.72
r1856 601 606 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=51.72 $Y=2.635
+ $X2=51.72 $Y2=2.34
r1857 597 891 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=50.78 $Y=2.805
+ $X2=50.78 $Y2=2.72
r1858 597 599 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=50.78 $Y=2.805
+ $X2=50.78 $Y2=3.1
r1859 593 891 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=50.78 $Y=2.635
+ $X2=50.78 $Y2=2.72
r1860 593 595 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=50.78 $Y=2.635
+ $X2=50.78 $Y2=2
r1861 589 656 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=49.84 $Y=2.805
+ $X2=49.84 $Y2=2.72
r1862 589 591 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=49.84 $Y=2.805
+ $X2=49.84 $Y2=3.1
r1863 585 656 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=49.84 $Y=2.635
+ $X2=49.84 $Y2=2.72
r1864 585 587 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=49.84 $Y=2.635
+ $X2=49.84 $Y2=2
r1865 581 653 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=46.892 $Y=2.805
+ $X2=46.892 $Y2=2.72
r1866 581 583 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=46.892 $Y=2.805
+ $X2=46.892 $Y2=3.14
r1867 577 653 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=46.892 $Y=2.635
+ $X2=46.892 $Y2=2.72
r1868 577 579 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=46.892 $Y=2.635
+ $X2=46.892 $Y2=1.77
r1869 573 888 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=45.91 $Y=2.805
+ $X2=45.91 $Y2=2.72
r1870 573 575 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=45.91 $Y=2.805
+ $X2=45.91 $Y2=3.14
r1871 569 888 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=45.91 $Y=2.635
+ $X2=45.91 $Y2=2.72
r1872 569 571 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=45.91 $Y=2.635
+ $X2=45.91 $Y2=1.77
r1873 568 650 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=45.32 $Y=2.72
+ $X2=45.17 $Y2=2.72
r1874 567 888 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=45.76 $Y=2.72
+ $X2=45.91 $Y2=2.72
r1875 567 568 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=45.76 $Y=2.72
+ $X2=45.32 $Y2=2.72
r1876 563 650 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=45.17 $Y=2.805
+ $X2=45.17 $Y2=2.72
r1877 563 565 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=45.17 $Y=2.805
+ $X2=45.17 $Y2=3.14
r1878 559 650 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=45.17 $Y=2.635
+ $X2=45.17 $Y2=2.72
r1879 559 561 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=45.17 $Y=2.635
+ $X2=45.17 $Y2=1.77
r1880 555 648 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=44.187 $Y=2.805
+ $X2=44.187 $Y2=2.72
r1881 555 557 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=44.187 $Y=2.805
+ $X2=44.187 $Y2=3.14
r1882 551 648 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=44.187 $Y=2.635
+ $X2=44.187 $Y2=2.72
r1883 551 553 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=44.187 $Y=2.635
+ $X2=44.187 $Y2=1.77
r1884 547 885 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=41.24 $Y=2.805
+ $X2=41.24 $Y2=2.72
r1885 547 549 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=41.24 $Y=2.805
+ $X2=41.24 $Y2=3.1
r1886 543 885 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=41.24 $Y=2.635
+ $X2=41.24 $Y2=2.72
r1887 543 545 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=41.24 $Y=2.635
+ $X2=41.24 $Y2=2
r1888 542 882 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.435 $Y=2.72
+ $X2=40.3 $Y2=2.72
r1889 541 885 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=41.105 $Y=2.72
+ $X2=41.24 $Y2=2.72
r1890 541 542 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=41.105 $Y=2.72
+ $X2=40.435 $Y2=2.72
r1891 537 882 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=40.3 $Y=2.805
+ $X2=40.3 $Y2=2.72
r1892 537 539 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=40.3 $Y=2.805
+ $X2=40.3 $Y2=3.1
r1893 533 882 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=40.3 $Y=2.635
+ $X2=40.3 $Y2=2.72
r1894 533 535 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=40.3 $Y=2.635
+ $X2=40.3 $Y2=2
r1895 529 531 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=39.36 $Y=3.1
+ $X2=39.36 $Y2=3.78
r1896 527 879 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=39.36 $Y=2.805
+ $X2=39.36 $Y2=2.72
r1897 527 529 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=39.36 $Y=2.805
+ $X2=39.36 $Y2=3.1
r1898 523 526 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=39.36 $Y=1.66
+ $X2=39.36 $Y2=2.34
r1899 521 879 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=39.36 $Y=2.635
+ $X2=39.36 $Y2=2.72
r1900 521 526 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=39.36 $Y=2.635
+ $X2=39.36 $Y2=2.34
r1901 520 876 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=38.975 $Y=2.72
+ $X2=38.84 $Y2=2.72
r1902 519 879 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=39.225 $Y=2.72
+ $X2=39.36 $Y2=2.72
r1903 519 520 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=39.225 $Y=2.72
+ $X2=38.975 $Y2=2.72
r1904 515 517 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=38.84 $Y=3.1
+ $X2=38.84 $Y2=3.78
r1905 513 876 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=38.84 $Y=2.805
+ $X2=38.84 $Y2=2.72
r1906 513 515 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=38.84 $Y=2.805
+ $X2=38.84 $Y2=3.1
r1907 509 512 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=38.84 $Y=1.66
+ $X2=38.84 $Y2=2.34
r1908 507 876 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=38.84 $Y=2.635
+ $X2=38.84 $Y2=2.72
r1909 507 512 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=38.84 $Y=2.635
+ $X2=38.84 $Y2=2.34
r1910 503 873 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=37.9 $Y=2.805
+ $X2=37.9 $Y2=2.72
r1911 503 505 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=37.9 $Y=2.805
+ $X2=37.9 $Y2=3.1
r1912 499 873 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=37.9 $Y=2.635
+ $X2=37.9 $Y2=2.72
r1913 499 501 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=37.9 $Y=2.635
+ $X2=37.9 $Y2=2
r1914 495 645 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=36.96 $Y=2.805
+ $X2=36.96 $Y2=2.72
r1915 495 497 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=36.96 $Y=2.805
+ $X2=36.96 $Y2=3.1
r1916 491 645 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=36.96 $Y=2.635
+ $X2=36.96 $Y2=2.72
r1917 491 493 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=36.96 $Y=2.635
+ $X2=36.96 $Y2=2
r1918 487 642 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=34.012 $Y=2.805
+ $X2=34.012 $Y2=2.72
r1919 487 489 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=34.012 $Y=2.805
+ $X2=34.012 $Y2=3.14
r1920 483 642 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=34.012 $Y=2.635
+ $X2=34.012 $Y2=2.72
r1921 483 485 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=34.012 $Y=2.635
+ $X2=34.012 $Y2=1.77
r1922 479 870 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=33.03 $Y=2.805
+ $X2=33.03 $Y2=2.72
r1923 479 481 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=33.03 $Y=2.805
+ $X2=33.03 $Y2=3.14
r1924 475 870 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=33.03 $Y=2.635
+ $X2=33.03 $Y2=2.72
r1925 475 477 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=33.03 $Y=2.635
+ $X2=33.03 $Y2=1.77
r1926 474 639 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=32.44 $Y=2.72
+ $X2=32.29 $Y2=2.72
r1927 473 870 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=32.88 $Y=2.72
+ $X2=33.03 $Y2=2.72
r1928 473 474 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=32.88 $Y=2.72
+ $X2=32.44 $Y2=2.72
r1929 469 639 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=32.29 $Y=2.805
+ $X2=32.29 $Y2=2.72
r1930 469 471 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=32.29 $Y=2.805
+ $X2=32.29 $Y2=3.14
r1931 465 639 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=32.29 $Y=2.635
+ $X2=32.29 $Y2=2.72
r1932 465 467 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=32.29 $Y=2.635
+ $X2=32.29 $Y2=1.77
r1933 461 637 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=31.307 $Y=2.805
+ $X2=31.307 $Y2=2.72
r1934 461 463 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=31.307 $Y=2.805
+ $X2=31.307 $Y2=3.14
r1935 457 637 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=31.307 $Y=2.635
+ $X2=31.307 $Y2=2.72
r1936 457 459 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=31.307 $Y=2.635
+ $X2=31.307 $Y2=1.77
r1937 453 867 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=28.36 $Y=2.805
+ $X2=28.36 $Y2=2.72
r1938 453 455 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=28.36 $Y=2.805
+ $X2=28.36 $Y2=3.1
r1939 449 867 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=28.36 $Y=2.635
+ $X2=28.36 $Y2=2.72
r1940 449 451 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=28.36 $Y=2.635
+ $X2=28.36 $Y2=2
r1941 448 864 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.555 $Y=2.72
+ $X2=27.42 $Y2=2.72
r1942 447 867 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=28.225 $Y=2.72
+ $X2=28.36 $Y2=2.72
r1943 447 448 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=28.225 $Y=2.72
+ $X2=27.555 $Y2=2.72
r1944 443 864 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=27.42 $Y=2.805
+ $X2=27.42 $Y2=2.72
r1945 443 445 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=27.42 $Y=2.805
+ $X2=27.42 $Y2=3.1
r1946 439 864 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=27.42 $Y=2.635
+ $X2=27.42 $Y2=2.72
r1947 439 441 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=27.42 $Y=2.635
+ $X2=27.42 $Y2=2
r1948 435 437 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=26.48 $Y=3.1
+ $X2=26.48 $Y2=3.78
r1949 433 861 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=26.48 $Y=2.805
+ $X2=26.48 $Y2=2.72
r1950 433 435 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=26.48 $Y=2.805
+ $X2=26.48 $Y2=3.1
r1951 429 432 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=26.48 $Y=1.66
+ $X2=26.48 $Y2=2.34
r1952 427 861 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=26.48 $Y=2.635
+ $X2=26.48 $Y2=2.72
r1953 427 432 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=26.48 $Y=2.635
+ $X2=26.48 $Y2=2.34
r1954 423 425 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=25.5 $Y=3.1
+ $X2=25.5 $Y2=3.78
r1955 421 858 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=25.5 $Y=2.805
+ $X2=25.5 $Y2=2.72
r1956 421 423 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.5 $Y=2.805
+ $X2=25.5 $Y2=3.1
r1957 417 420 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=25.5 $Y=1.66
+ $X2=25.5 $Y2=2.34
r1958 415 858 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=25.5 $Y=2.635
+ $X2=25.5 $Y2=2.72
r1959 415 420 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.5 $Y=2.635
+ $X2=25.5 $Y2=2.34
r1960 411 855 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=2.805
+ $X2=24.56 $Y2=2.72
r1961 411 413 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=24.56 $Y=2.805
+ $X2=24.56 $Y2=3.1
r1962 407 855 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=2.635
+ $X2=24.56 $Y2=2.72
r1963 407 409 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=24.56 $Y=2.635
+ $X2=24.56 $Y2=2
r1964 403 634 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.62 $Y=2.805
+ $X2=23.62 $Y2=2.72
r1965 403 405 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=23.62 $Y=2.805
+ $X2=23.62 $Y2=3.1
r1966 399 634 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.62 $Y=2.635
+ $X2=23.62 $Y2=2.72
r1967 399 401 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=23.62 $Y=2.635
+ $X2=23.62 $Y2=2
r1968 395 631 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=20.672 $Y=2.805
+ $X2=20.672 $Y2=2.72
r1969 395 397 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=20.672 $Y=2.805
+ $X2=20.672 $Y2=3.14
r1970 391 631 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=20.672 $Y=2.635
+ $X2=20.672 $Y2=2.72
r1971 391 393 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=20.672 $Y=2.635
+ $X2=20.672 $Y2=1.77
r1972 387 852 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.69 $Y=2.805
+ $X2=19.69 $Y2=2.72
r1973 387 389 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=19.69 $Y=2.805
+ $X2=19.69 $Y2=3.14
r1974 383 852 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.69 $Y=2.635
+ $X2=19.69 $Y2=2.72
r1975 383 385 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=19.69 $Y=2.635
+ $X2=19.69 $Y2=1.77
r1976 382 628 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.1 $Y=2.72
+ $X2=18.95 $Y2=2.72
r1977 381 852 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.54 $Y=2.72
+ $X2=19.69 $Y2=2.72
r1978 381 382 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=19.54 $Y=2.72
+ $X2=19.1 $Y2=2.72
r1979 377 628 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.95 $Y=2.805
+ $X2=18.95 $Y2=2.72
r1980 377 379 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=18.95 $Y=2.805
+ $X2=18.95 $Y2=3.14
r1981 373 628 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.95 $Y=2.635
+ $X2=18.95 $Y2=2.72
r1982 373 375 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=18.95 $Y=2.635
+ $X2=18.95 $Y2=1.77
r1983 369 626 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=17.967 $Y=2.805
+ $X2=17.967 $Y2=2.72
r1984 369 371 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=17.967 $Y=2.805
+ $X2=17.967 $Y2=3.14
r1985 365 626 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=17.967 $Y=2.635
+ $X2=17.967 $Y2=2.72
r1986 365 367 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=17.967 $Y=2.635
+ $X2=17.967 $Y2=1.77
r1987 361 849 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.02 $Y=2.805
+ $X2=15.02 $Y2=2.72
r1988 361 363 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.02 $Y=2.805
+ $X2=15.02 $Y2=3.1
r1989 357 849 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.02 $Y=2.635
+ $X2=15.02 $Y2=2.72
r1990 357 359 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=15.02 $Y=2.635
+ $X2=15.02 $Y2=2
r1991 356 846 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.215 $Y=2.72
+ $X2=14.08 $Y2=2.72
r1992 355 849 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=15.02 $Y2=2.72
r1993 355 356 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=14.215 $Y2=2.72
r1994 351 846 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=2.805
+ $X2=14.08 $Y2=2.72
r1995 351 353 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.08 $Y=2.805
+ $X2=14.08 $Y2=3.1
r1996 347 846 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=2.635
+ $X2=14.08 $Y2=2.72
r1997 347 349 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.08 $Y=2.635
+ $X2=14.08 $Y2=2
r1998 343 345 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.14 $Y=3.1
+ $X2=13.14 $Y2=3.78
r1999 341 843 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=2.805
+ $X2=13.14 $Y2=2.72
r2000 341 343 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.14 $Y=2.805
+ $X2=13.14 $Y2=3.1
r2001 337 340 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.14 $Y=1.66
+ $X2=13.14 $Y2=2.34
r2002 335 843 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=2.635
+ $X2=13.14 $Y2=2.72
r2003 335 340 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.14 $Y=2.635
+ $X2=13.14 $Y2=2.34
r2004 334 840 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.755 $Y=2.72
+ $X2=12.62 $Y2=2.72
r2005 333 843 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.005 $Y=2.72
+ $X2=13.14 $Y2=2.72
r2006 333 334 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.005 $Y=2.72
+ $X2=12.755 $Y2=2.72
r2007 329 331 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.62 $Y=3.1
+ $X2=12.62 $Y2=3.78
r2008 327 840 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.62 $Y=2.805
+ $X2=12.62 $Y2=2.72
r2009 327 329 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.62 $Y=2.805
+ $X2=12.62 $Y2=3.1
r2010 323 326 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.62 $Y=1.66
+ $X2=12.62 $Y2=2.34
r2011 321 840 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.62 $Y=2.635
+ $X2=12.62 $Y2=2.72
r2012 321 326 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.62 $Y=2.635
+ $X2=12.62 $Y2=2.34
r2013 317 837 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=2.805
+ $X2=11.68 $Y2=2.72
r2014 317 319 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.68 $Y=2.805
+ $X2=11.68 $Y2=3.1
r2015 313 837 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=2.635
+ $X2=11.68 $Y2=2.72
r2016 313 315 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.68 $Y=2.635
+ $X2=11.68 $Y2=2
r2017 309 623 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=2.805
+ $X2=10.74 $Y2=2.72
r2018 309 311 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.74 $Y=2.805
+ $X2=10.74 $Y2=3.1
r2019 305 623 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=2.635
+ $X2=10.74 $Y2=2.72
r2020 305 307 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.74 $Y=2.635
+ $X2=10.74 $Y2=2
r2021 301 620 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.792 $Y=2.805
+ $X2=7.792 $Y2=2.72
r2022 301 303 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=7.792 $Y=2.805
+ $X2=7.792 $Y2=3.14
r2023 297 620 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.792 $Y=2.635
+ $X2=7.792 $Y2=2.72
r2024 297 299 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=7.792 $Y=2.635
+ $X2=7.792 $Y2=1.77
r2025 293 834 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=2.805
+ $X2=6.81 $Y2=2.72
r2026 293 295 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.81 $Y=2.805
+ $X2=6.81 $Y2=3.14
r2027 289 834 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=2.635
+ $X2=6.81 $Y2=2.72
r2028 289 291 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=6.81 $Y=2.635
+ $X2=6.81 $Y2=1.77
r2029 288 617 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.22 $Y=2.72
+ $X2=6.07 $Y2=2.72
r2030 287 834 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.66 $Y=2.72
+ $X2=6.81 $Y2=2.72
r2031 287 288 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.66 $Y=2.72
+ $X2=6.22 $Y2=2.72
r2032 283 617 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.805
+ $X2=6.07 $Y2=2.72
r2033 283 285 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=6.07 $Y=2.805
+ $X2=6.07 $Y2=3.14
r2034 279 617 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.635
+ $X2=6.07 $Y2=2.72
r2035 279 281 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=6.07 $Y=2.635
+ $X2=6.07 $Y2=1.77
r2036 275 615 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.087 $Y=2.805
+ $X2=5.087 $Y2=2.72
r2037 275 277 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=5.087 $Y=2.805
+ $X2=5.087 $Y2=3.14
r2038 271 615 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=2.72
r2039 271 273 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=1.77
r2040 267 831 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.805
+ $X2=2.14 $Y2=2.72
r2041 267 269 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.14 $Y=2.805
+ $X2=2.14 $Y2=3.1
r2042 263 831 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r2043 263 265 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r2044 262 828 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r2045 261 831 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r2046 261 262 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r2047 257 828 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.805
+ $X2=1.2 $Y2=2.72
r2048 257 259 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.805
+ $X2=1.2 $Y2=3.1
r2049 253 828 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r2050 253 255 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r2051 249 251 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=3.1
+ $X2=0.26 $Y2=3.78
r2052 247 825 3.46198 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.805
+ $X2=0.197 $Y2=2.72
r2053 247 249 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.805
+ $X2=0.26 $Y2=3.1
r2054 243 246 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r2055 241 825 3.46198 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.197 $Y2=2.72
r2056 241 246 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r2057 80 611 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1
+ $X=51.575 $Y=2.955 $X2=51.72 $Y2=3.78
r2058 80 609 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=51.575 $Y=2.955 $X2=51.72 $Y2=3.1
r2059 79 606 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=51.575 $Y=1.485 $X2=51.72 $Y2=2.34
r2060 79 603 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1
+ $X=51.575 $Y=1.485 $X2=51.72 $Y2=1.66
r2061 78 599 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=50.635 $Y=2.955 $X2=50.78 $Y2=3.1
r2062 77 595 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=50.635 $Y=1.485 $X2=50.78 $Y2=2
r2063 76 591 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2
+ $X=49.715 $Y=2.955 $X2=49.84 $Y2=3.1
r2064 75 587 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2
+ $X=49.715 $Y=1.485 $X2=49.84 $Y2=2
r2065 74 583 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=46.72
+ $Y=2.995 $X2=46.865 $Y2=3.14
r2066 73 579 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=46.72
+ $Y=1.625 $X2=46.865 $Y2=1.77
r2067 72 575 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=45.8
+ $Y=2.995 $X2=45.925 $Y2=3.14
r2068 71 571 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=45.8
+ $Y=1.625 $X2=45.925 $Y2=1.77
r2069 70 565 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=45.01
+ $Y=2.995 $X2=45.155 $Y2=3.14
r2070 69 561 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=45.01
+ $Y=1.625 $X2=45.155 $Y2=1.77
r2071 68 557 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=44.09
+ $Y=2.995 $X2=44.215 $Y2=3.14
r2072 67 553 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=44.09
+ $Y=1.625 $X2=44.215 $Y2=1.77
r2073 66 549 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=41.095 $Y=2.955 $X2=41.24 $Y2=3.1
r2074 65 545 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=41.095 $Y=1.485 $X2=41.24 $Y2=2
r2075 64 539 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=40.155 $Y=2.955 $X2=40.3 $Y2=3.1
r2076 63 535 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=40.155 $Y=1.485 $X2=40.3 $Y2=2
r2077 62 531 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1
+ $X=39.235 $Y=2.955 $X2=39.36 $Y2=3.78
r2078 62 529 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1
+ $X=39.235 $Y=2.955 $X2=39.36 $Y2=3.1
r2079 61 526 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1
+ $X=39.235 $Y=1.485 $X2=39.36 $Y2=2.34
r2080 61 523 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1
+ $X=39.235 $Y=1.485 $X2=39.36 $Y2=1.66
r2081 60 517 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1
+ $X=38.695 $Y=2.955 $X2=38.84 $Y2=3.78
r2082 60 515 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=38.695 $Y=2.955 $X2=38.84 $Y2=3.1
r2083 59 512 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=38.695 $Y=1.485 $X2=38.84 $Y2=2.34
r2084 59 509 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1
+ $X=38.695 $Y=1.485 $X2=38.84 $Y2=1.66
r2085 58 505 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=37.755 $Y=2.955 $X2=37.9 $Y2=3.1
r2086 57 501 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=37.755 $Y=1.485 $X2=37.9 $Y2=2
r2087 56 497 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2
+ $X=36.835 $Y=2.955 $X2=36.96 $Y2=3.1
r2088 55 493 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2
+ $X=36.835 $Y=1.485 $X2=36.96 $Y2=2
r2089 54 489 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=33.84
+ $Y=2.995 $X2=33.985 $Y2=3.14
r2090 53 485 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=33.84
+ $Y=1.625 $X2=33.985 $Y2=1.77
r2091 52 481 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=32.92
+ $Y=2.995 $X2=33.045 $Y2=3.14
r2092 51 477 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=32.92
+ $Y=1.625 $X2=33.045 $Y2=1.77
r2093 50 471 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=32.13
+ $Y=2.995 $X2=32.275 $Y2=3.14
r2094 49 467 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=32.13
+ $Y=1.625 $X2=32.275 $Y2=1.77
r2095 48 463 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=31.21
+ $Y=2.995 $X2=31.335 $Y2=3.14
r2096 47 459 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=31.21
+ $Y=1.625 $X2=31.335 $Y2=1.77
r2097 46 455 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=28.215 $Y=2.955 $X2=28.36 $Y2=3.1
r2098 45 451 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=28.215 $Y=1.485 $X2=28.36 $Y2=2
r2099 44 445 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=27.275 $Y=2.955 $X2=27.42 $Y2=3.1
r2100 43 441 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=27.275 $Y=1.485 $X2=27.42 $Y2=2
r2101 42 437 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1
+ $X=26.355 $Y=2.955 $X2=26.48 $Y2=3.78
r2102 42 435 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1
+ $X=26.355 $Y=2.955 $X2=26.48 $Y2=3.1
r2103 41 432 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1
+ $X=26.355 $Y=1.485 $X2=26.48 $Y2=2.34
r2104 41 429 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1
+ $X=26.355 $Y=1.485 $X2=26.48 $Y2=1.66
r2105 40 425 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1
+ $X=25.355 $Y=2.955 $X2=25.5 $Y2=3.78
r2106 40 423 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=25.355 $Y=2.955 $X2=25.5 $Y2=3.1
r2107 39 420 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=25.355 $Y=1.485 $X2=25.5 $Y2=2.34
r2108 39 417 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1
+ $X=25.355 $Y=1.485 $X2=25.5 $Y2=1.66
r2109 38 413 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=24.415 $Y=2.955 $X2=24.56 $Y2=3.1
r2110 37 409 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=24.415 $Y=1.485 $X2=24.56 $Y2=2
r2111 36 405 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2
+ $X=23.495 $Y=2.955 $X2=23.62 $Y2=3.1
r2112 35 401 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2
+ $X=23.495 $Y=1.485 $X2=23.62 $Y2=2
r2113 34 397 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.5
+ $Y=2.995 $X2=20.645 $Y2=3.14
r2114 33 393 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.5
+ $Y=1.625 $X2=20.645 $Y2=1.77
r2115 32 389 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=19.58
+ $Y=2.995 $X2=19.705 $Y2=3.14
r2116 31 385 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=19.58
+ $Y=1.625 $X2=19.705 $Y2=1.77
r2117 30 379 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.79
+ $Y=2.995 $X2=18.935 $Y2=3.14
r2118 29 375 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.79
+ $Y=1.625 $X2=18.935 $Y2=1.77
r2119 28 371 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=17.87
+ $Y=2.995 $X2=17.995 $Y2=3.14
r2120 27 367 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=17.87
+ $Y=1.625 $X2=17.995 $Y2=1.77
r2121 26 363 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=14.875 $Y=2.955 $X2=15.02 $Y2=3.1
r2122 25 359 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=14.875 $Y=1.485 $X2=15.02 $Y2=2
r2123 24 353 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=13.935 $Y=2.955 $X2=14.08 $Y2=3.1
r2124 23 349 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=13.935 $Y=1.485 $X2=14.08 $Y2=2
r2125 22 345 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1
+ $X=13.015 $Y=2.955 $X2=13.14 $Y2=3.78
r2126 22 343 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1
+ $X=13.015 $Y=2.955 $X2=13.14 $Y2=3.1
r2127 21 340 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1
+ $X=13.015 $Y=1.485 $X2=13.14 $Y2=2.34
r2128 21 337 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1
+ $X=13.015 $Y=1.485 $X2=13.14 $Y2=1.66
r2129 20 331 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1
+ $X=12.475 $Y=2.955 $X2=12.62 $Y2=3.78
r2130 20 329 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1
+ $X=12.475 $Y=2.955 $X2=12.62 $Y2=3.1
r2131 19 326 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1
+ $X=12.475 $Y=1.485 $X2=12.62 $Y2=2.34
r2132 19 323 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1
+ $X=12.475 $Y=1.485 $X2=12.62 $Y2=1.66
r2133 18 319 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=11.535 $Y=2.955 $X2=11.68 $Y2=3.1
r2134 17 315 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2
+ $X=11.535 $Y=1.485 $X2=11.68 $Y2=2
r2135 16 311 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2
+ $X=10.615 $Y=2.955 $X2=10.74 $Y2=3.1
r2136 15 307 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2
+ $X=10.615 $Y=1.485 $X2=10.74 $Y2=2
r2137 14 303 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.62
+ $Y=2.995 $X2=7.765 $Y2=3.14
r2138 13 299 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.62
+ $Y=1.625 $X2=7.765 $Y2=1.77
r2139 12 295 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.7
+ $Y=2.995 $X2=6.825 $Y2=3.14
r2140 11 291 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.7
+ $Y=1.625 $X2=6.825 $Y2=1.77
r2141 10 285 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=2.995 $X2=6.055 $Y2=3.14
r2142 9 281 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.625 $X2=6.055 $Y2=1.77
r2143 8 277 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=2.995 $X2=5.115 $Y2=3.14
r2144 7 273 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=1.625 $X2=5.115 $Y2=1.77
r2145 6 269 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=2.955 $X2=2.14 $Y2=3.1
r2146 5 265 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r2147 4 259 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=2.955 $X2=1.2 $Y2=3.1
r2148 3 255 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r2149 2 251 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.78
r2150 2 249 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.955 $X2=0.26 $Y2=3.1
r2151 1 246 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r2152 1 243 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_297# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 37 41 49 59 63 68
c116 63 0 1.3204e-19 $X=3.6 $Y=1.7
c117 49 0 1.97167e-19 $X=4.55 $Y=2.225
c118 33 0 1.87597e-19 $X=4.405 $Y=2.225
c119 32 0 1.97167e-19 $X=2.795 $Y=2.225
c120 31 0 1.87597e-19 $X=3.455 $Y=2.225
c121 30 0 1.97849e-19 $X=1.815 $Y=2.225
c122 29 0 1.36925e-19 $X=2.505 $Y=2.225
c123 28 0 1.97849e-19 $X=0.875 $Y=2.225
r124 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=4.555 $Y=2.225
+ $X2=4.555 $Y2=1.73
r125 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=2.225
+ $X2=4.55 $Y2=2.225
r126 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=3.6 $Y=2.225
+ $X2=3.6 $Y2=1.7
r127 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=2.225
+ $X2=3.6 $Y2=2.225
r128 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=2.645 $Y=2.225
+ $X2=2.645 $Y2=1.7
r129 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.65 $Y=2.225
+ $X2=2.65 $Y2=2.225
r130 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.67 $Y=2.225
+ $X2=1.67 $Y2=2.225
r131 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=2.225
+ $X2=0.73 $Y2=2.225
r132 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=2.225
+ $X2=3.6 $Y2=2.225
r133 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.405 $Y=2.225
+ $X2=4.55 $Y2=2.225
r134 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=4.405 $Y=2.225
+ $X2=3.745 $Y2=2.225
r135 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.795 $Y=2.225
+ $X2=2.65 $Y2=2.225
r136 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=2.225
+ $X2=3.6 $Y2=2.225
r137 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=3.455 $Y=2.225
+ $X2=2.795 $Y2=2.225
r138 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.815 $Y=2.225
+ $X2=1.67 $Y2=2.225
r139 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.505 $Y=2.225
+ $X2=2.65 $Y2=2.225
r140 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=2.505 $Y=2.225
+ $X2=1.815 $Y2=2.225
r141 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=2.225
+ $X2=0.73 $Y2=2.225
r142 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.525 $Y=2.225
+ $X2=1.67 $Y2=2.225
r143 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.525 $Y=2.225
+ $X2=0.875 $Y2=2.225
r144 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=1.7
r145 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.225
r146 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r147 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.225
r148 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r149 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r150 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=2.645 $Y2=1.665
r151 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=1.835 $Y2=1.58
r152 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r153 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r154 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r155 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.555 $X2=4.54 $Y2=1.73
r156 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.555 $X2=3.6 $Y2=1.7
r157 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.555 $X2=2.66 $Y2=1.7
r158 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r159 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r160 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r161 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_591# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 49 53 56 59 62 66
c116 62 0 1.3204e-19 $X=3.6 $Y=3.21
c117 49 0 1.97167e-19 $X=4.55 $Y=3.215
c118 33 0 1.87597e-19 $X=4.405 $Y=3.215
c119 32 0 1.97167e-19 $X=2.795 $Y=3.215
c120 31 0 1.87597e-19 $X=3.455 $Y=3.215
c121 30 0 1.97849e-19 $X=1.815 $Y=3.215
c122 29 0 1.36925e-19 $X=2.505 $Y=3.215
c123 28 0 1.97849e-19 $X=0.875 $Y=3.215
r124 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.55 $Y=3.215
+ $X2=4.55 $Y2=3.215
r125 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.6 $Y=3.215
+ $X2=3.6 $Y2=3.215
r126 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.65 $Y=3.215
+ $X2=2.65 $Y2=3.215
r127 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.67 $Y=3.215
+ $X2=1.67 $Y2=3.215
r128 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=3.215
+ $X2=0.73 $Y2=3.215
r129 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.745 $Y=3.215
+ $X2=3.6 $Y2=3.215
r130 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.405 $Y=3.215
+ $X2=4.55 $Y2=3.215
r131 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=4.405 $Y=3.215
+ $X2=3.745 $Y2=3.215
r132 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.795 $Y=3.215
+ $X2=2.65 $Y2=3.215
r133 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=3.215
+ $X2=3.6 $Y2=3.215
r134 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=3.455 $Y=3.215
+ $X2=2.795 $Y2=3.215
r135 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.815 $Y=3.215
+ $X2=1.67 $Y2=3.215
r136 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.505 $Y=3.215
+ $X2=2.65 $Y2=3.215
r137 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=2.505 $Y=3.215
+ $X2=1.815 $Y2=3.215
r138 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=3.215
+ $X2=0.73 $Y2=3.215
r139 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.525 $Y=3.215
+ $X2=1.67 $Y2=3.215
r140 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.525 $Y=3.215
+ $X2=0.875 $Y2=3.215
r141 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=2.645 $Y=3.775
+ $X2=2.645 $Y2=3.21
r142 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=3.775
+ $X2=1.67 $Y2=3.1
r143 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=3.775
+ $X2=1.67 $Y2=3.86
r144 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=3.775
+ $X2=0.73 $Y2=3.1
r145 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=3.775
+ $X2=0.73 $Y2=3.86
r146 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=3.86
+ $X2=1.67 $Y2=3.86
r147 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.495 $Y=3.86
+ $X2=2.645 $Y2=3.775
r148 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.495 $Y=3.86
+ $X2=1.835 $Y2=3.86
r149 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=3.86
+ $X2=0.73 $Y2=3.86
r150 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=3.86
+ $X2=1.67 $Y2=3.86
r151 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=3.86
+ $X2=0.895 $Y2=3.86
r152 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=3.065 $X2=4.54 $Y2=3.21
r153 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=3.065 $X2=3.6 $Y2=3.21
r154 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=3.065 $X2=2.66 $Y2=3.21
r155 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=2.955 $X2=1.67 $Y2=3.1
r156 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=2.955 $X2=1.67 $Y2=3.78
r157 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.955 $X2=0.73 $Y2=3.1
r158 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.955 $X2=0.73 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 194 197
+ 199 203 207 211 215 217 219 222 226 229 231 235 239 243 247 249 251 254 258
+ 261 263 267 271 275 279 281 283 286 290 293 295 299 303 307 311 313 315 318
+ 322 326 327 330 332 334 336 338 340 342 344 346 350 351 354 358 359 362 364
+ 366 368 370 372 374 376 378 382 383 386 390 391 394 396 398 400 402 404 406
+ 408 410 414 415 418 422 423 426 428 430 432 434 436 438 440 442 446 447 449
+ 450 451 452 453 454 455 456 457 458 459 460 461 462 463 464 465 466 467 468
+ 469 470 471 472 473 474 475 476 477 481 485 489 493 497 501 505 509 513 517
+ 521 525 527 530 532 535 536 537 538 539 540 541 542 543 544 545 546 547 548
+ 549 550 551 552 588 597 606 615 620 625 634 643 648 653 662 671 676 681 690
+ 699 704 706
c1894 471 0 3.48484e-19 $X=42.085 $Y=3.57
c1895 469 0 3.48484e-19 $X=42.085 $Y=1.87
c1896 463 0 3.48484e-19 $X=29.205 $Y=3.57
c1897 461 0 3.48484e-19 $X=29.205 $Y=1.87
c1898 455 0 3.48484e-19 $X=15.865 $Y=3.57
c1899 453 0 3.48484e-19 $X=15.865 $Y=1.87
c1900 436 0 1.20815e-19 $X=48.01 $Y=4.225
c1901 434 0 1.20815e-19 $X=48.01 $Y=1.215
c1902 432 0 1.20815e-19 $X=43.07 $Y=4.225
c1903 430 0 1.20815e-19 $X=43.07 $Y=1.215
c1904 404 0 1.20815e-19 $X=35.13 $Y=4.225
c1905 402 0 1.20815e-19 $X=35.13 $Y=1.215
c1906 400 0 1.20815e-19 $X=30.19 $Y=4.225
c1907 398 0 1.20815e-19 $X=30.19 $Y=1.215
c1908 372 0 1.20815e-19 $X=21.79 $Y=4.225
c1909 370 0 1.20815e-19 $X=21.79 $Y=1.215
c1910 368 0 1.20815e-19 $X=16.85 $Y=4.225
c1911 366 0 1.20815e-19 $X=16.85 $Y=1.215
c1912 340 0 1.20815e-19 $X=8.91 $Y=4.225
c1913 338 0 1.20815e-19 $X=8.91 $Y=1.215
c1914 336 0 1.20815e-19 $X=3.97 $Y=4.225
c1915 334 0 1.20815e-19 $X=3.97 $Y=1.215
r1916 699 701 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=48.85 $Y=1.7
+ $X2=48.85 $Y2=3.21
r1917 694 696 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=47.91 $Y=3.21
+ $X2=47.91 $Y2=3.57
r1918 690 694 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=47.91 $Y=1.7
+ $X2=47.91 $Y2=3.21
r1919 685 687 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=43.17 $Y=3.21
+ $X2=43.17 $Y2=3.57
r1920 681 685 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=43.17 $Y=1.7
+ $X2=43.17 $Y2=3.21
r1921 676 678 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=42.23 $Y=1.7
+ $X2=42.23 $Y2=3.21
r1922 671 673 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=35.97 $Y=1.7
+ $X2=35.97 $Y2=3.21
r1923 666 668 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=35.03 $Y=3.21
+ $X2=35.03 $Y2=3.57
r1924 662 666 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=35.03 $Y=1.7
+ $X2=35.03 $Y2=3.21
r1925 657 659 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=30.29 $Y=3.21
+ $X2=30.29 $Y2=3.57
r1926 653 657 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=30.29 $Y=1.7
+ $X2=30.29 $Y2=3.21
r1927 648 650 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=29.35 $Y=1.7
+ $X2=29.35 $Y2=3.21
r1928 643 645 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=22.63 $Y=1.7
+ $X2=22.63 $Y2=3.21
r1929 638 640 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=21.69 $Y=3.21
+ $X2=21.69 $Y2=3.57
r1930 634 638 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=21.69 $Y=1.7
+ $X2=21.69 $Y2=3.21
r1931 629 631 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=16.95 $Y=3.21
+ $X2=16.95 $Y2=3.57
r1932 625 629 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=16.95 $Y=1.7
+ $X2=16.95 $Y2=3.21
r1933 620 622 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=16.01 $Y=1.7
+ $X2=16.01 $Y2=3.21
r1934 615 617 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=9.75 $Y=1.7
+ $X2=9.75 $Y2=3.21
r1935 610 612 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=8.81 $Y=3.21
+ $X2=8.81 $Y2=3.57
r1936 606 610 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=8.81 $Y=1.7
+ $X2=8.81 $Y2=3.21
r1937 601 603 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.07 $Y=3.21
+ $X2=4.07 $Y2=3.57
r1938 597 601 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=4.07 $Y=1.7
+ $X2=4.07 $Y2=3.21
r1939 592 594 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.13 $Y=3.21
+ $X2=3.13 $Y2=3.57
r1940 588 592 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=3.13 $Y=1.7
+ $X2=3.13 $Y2=3.21
r1941 552 696 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=47.91 $Y=3.57
+ $X2=47.91 $Y2=3.57
r1942 551 690 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=47.91 $Y=1.87
+ $X2=47.91 $Y2=1.87
r1943 550 687 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=43.17 $Y=3.57
+ $X2=43.17 $Y2=3.57
r1944 549 681 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=43.17 $Y=1.87
+ $X2=43.17 $Y2=1.87
r1945 548 668 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.03 $Y=3.57
+ $X2=35.03 $Y2=3.57
r1946 547 662 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.03 $Y=1.87
+ $X2=35.03 $Y2=1.87
r1947 546 659 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=30.29 $Y=3.57
+ $X2=30.29 $Y2=3.57
r1948 545 653 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=30.29 $Y=1.87
+ $X2=30.29 $Y2=1.87
r1949 544 640 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.69 $Y=3.57
+ $X2=21.69 $Y2=3.57
r1950 543 634 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.69 $Y=1.87
+ $X2=21.69 $Y2=1.87
r1951 542 631 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.95 $Y=3.57
+ $X2=16.95 $Y2=3.57
r1952 541 625 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.95 $Y=1.87
+ $X2=16.95 $Y2=1.87
r1953 540 612 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.81 $Y=3.57
+ $X2=8.81 $Y2=3.57
r1954 539 606 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.81 $Y=1.87
+ $X2=8.81 $Y2=1.87
r1955 538 706 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=3.925 $Y=3.57
+ $X2=3.275 $Y2=3.57
r1956 538 603 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=3.57
+ $X2=4.07 $Y2=3.57
r1957 537 704 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=3.925 $Y=1.87
+ $X2=3.275 $Y2=1.87
r1958 537 597 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=1.87
+ $X2=4.07 $Y2=1.87
r1959 536 706 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.13 $Y=3.57
+ $X2=3.275 $Y2=3.57
r1960 536 594 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.13 $Y=3.57
+ $X2=3.13 $Y2=3.57
r1961 535 704 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.13 $Y=1.87
+ $X2=3.275 $Y2=1.87
r1962 535 588 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.13 $Y=1.87
+ $X2=3.13 $Y2=1.87
r1963 533 701 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=48.85 $Y=3.57
+ $X2=48.85 $Y2=3.21
r1964 532 533 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=48.85 $Y=3.57
+ $X2=48.85 $Y2=3.57
r1965 530 552 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=48.705 $Y=3.57
+ $X2=48.055 $Y2=3.57
r1966 530 532 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.705 $Y=3.57
+ $X2=48.85 $Y2=3.57
r1967 527 699 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=48.85 $Y=1.87
+ $X2=48.85 $Y2=1.87
r1968 525 551 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=48.705 $Y=1.87
+ $X2=48.055 $Y2=1.87
r1969 525 527 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.705 $Y=1.87
+ $X2=48.85 $Y2=1.87
r1970 524 678 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=42.23 $Y=3.57
+ $X2=42.23 $Y2=3.21
r1971 523 524 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=42.23 $Y=3.57
+ $X2=42.23 $Y2=3.57
r1972 521 550 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=42.375 $Y=3.57
+ $X2=43.025 $Y2=3.57
r1973 521 523 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.375 $Y=3.57
+ $X2=42.23 $Y2=3.57
r1974 519 676 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=42.23 $Y=1.87
+ $X2=42.23 $Y2=1.87
r1975 517 549 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=42.375 $Y=1.87
+ $X2=43.025 $Y2=1.87
r1976 517 519 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.375 $Y=1.87
+ $X2=42.23 $Y2=1.87
r1977 516 673 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=35.97 $Y=3.57
+ $X2=35.97 $Y2=3.21
r1978 515 516 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.97 $Y=3.57
+ $X2=35.97 $Y2=3.57
r1979 513 548 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=35.825 $Y=3.57
+ $X2=35.175 $Y2=3.57
r1980 513 515 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.825 $Y=3.57
+ $X2=35.97 $Y2=3.57
r1981 511 671 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.97 $Y=1.87
+ $X2=35.97 $Y2=1.87
r1982 509 547 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=35.825 $Y=1.87
+ $X2=35.175 $Y2=1.87
r1983 509 511 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.825 $Y=1.87
+ $X2=35.97 $Y2=1.87
r1984 508 650 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=29.35 $Y=3.57
+ $X2=29.35 $Y2=3.21
r1985 507 508 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=29.35 $Y=3.57
+ $X2=29.35 $Y2=3.57
r1986 505 546 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=29.495 $Y=3.57
+ $X2=30.145 $Y2=3.57
r1987 505 507 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.495 $Y=3.57
+ $X2=29.35 $Y2=3.57
r1988 503 648 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=29.35 $Y=1.87
+ $X2=29.35 $Y2=1.87
r1989 501 545 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=29.495 $Y=1.87
+ $X2=30.145 $Y2=1.87
r1990 501 503 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.495 $Y=1.87
+ $X2=29.35 $Y2=1.87
r1991 500 645 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=22.63 $Y=3.57
+ $X2=22.63 $Y2=3.21
r1992 499 500 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.63 $Y=3.57
+ $X2=22.63 $Y2=3.57
r1993 497 544 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=22.485 $Y=3.57
+ $X2=21.835 $Y2=3.57
r1994 497 499 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.485 $Y=3.57
+ $X2=22.63 $Y2=3.57
r1995 495 643 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.63 $Y=1.87
+ $X2=22.63 $Y2=1.87
r1996 493 543 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=22.485 $Y=1.87
+ $X2=21.835 $Y2=1.87
r1997 493 495 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.485 $Y=1.87
+ $X2=22.63 $Y2=1.87
r1998 492 622 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=16.01 $Y=3.57
+ $X2=16.01 $Y2=3.21
r1999 491 492 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.01 $Y=3.57
+ $X2=16.01 $Y2=3.57
r2000 489 542 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=16.155 $Y=3.57
+ $X2=16.805 $Y2=3.57
r2001 489 491 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.155 $Y=3.57
+ $X2=16.01 $Y2=3.57
r2002 487 620 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.01 $Y=1.87
+ $X2=16.01 $Y2=1.87
r2003 485 541 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=16.155 $Y=1.87
+ $X2=16.805 $Y2=1.87
r2004 485 487 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.155 $Y=1.87
+ $X2=16.01 $Y2=1.87
r2005 484 617 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.75 $Y=3.57
+ $X2=9.75 $Y2=3.21
r2006 483 484 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.75 $Y=3.57
+ $X2=9.75 $Y2=3.57
r2007 481 540 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=9.605 $Y=3.57
+ $X2=8.955 $Y2=3.57
r2008 481 483 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.605 $Y=3.57
+ $X2=9.75 $Y2=3.57
r2009 479 615 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.75 $Y=1.87
+ $X2=9.75 $Y2=1.87
r2010 477 539 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=9.605 $Y=1.87
+ $X2=8.955 $Y2=1.87
r2011 477 479 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.605 $Y=1.87
+ $X2=9.75 $Y2=1.87
r2012 476 550 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=43.315 $Y=3.57
+ $X2=43.11 $Y2=3.57
r2013 475 552 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=47.765 $Y=3.57
+ $X2=47.91 $Y2=3.57
r2014 475 476 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=47.765 $Y=3.57
+ $X2=43.315 $Y2=3.57
r2015 474 549 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=43.315 $Y=1.87
+ $X2=43.11 $Y2=1.87
r2016 473 551 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=47.765 $Y=1.87
+ $X2=47.91 $Y2=1.87
r2017 473 474 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=47.765 $Y=1.87
+ $X2=43.315 $Y2=1.87
r2018 472 515 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.115 $Y=3.57
+ $X2=35.97 $Y2=3.57
r2019 471 523 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.085 $Y=3.57
+ $X2=42.23 $Y2=3.57
r2020 471 472 7.3886 $w=1.4e-07 $l=5.97e-06 $layer=MET1_cond $X=42.085 $Y=3.57
+ $X2=36.115 $Y2=3.57
r2021 470 511 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.115 $Y=1.87
+ $X2=35.97 $Y2=1.87
r2022 469 519 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.085 $Y=1.87
+ $X2=42.23 $Y2=1.87
r2023 469 470 7.3886 $w=1.4e-07 $l=5.97e-06 $layer=MET1_cond $X=42.085 $Y=1.87
+ $X2=36.115 $Y2=1.87
r2024 468 546 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=30.435 $Y=3.57
+ $X2=30.23 $Y2=3.57
r2025 467 548 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=34.885 $Y=3.57
+ $X2=35.03 $Y2=3.57
r2026 467 468 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=34.885 $Y=3.57
+ $X2=30.435 $Y2=3.57
r2027 466 545 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=30.435 $Y=1.87
+ $X2=30.23 $Y2=1.87
r2028 465 547 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=34.885 $Y=1.87
+ $X2=35.03 $Y2=1.87
r2029 465 466 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=34.885 $Y=1.87
+ $X2=30.435 $Y2=1.87
r2030 464 499 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.775 $Y=3.57
+ $X2=22.63 $Y2=3.57
r2031 463 507 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.205 $Y=3.57
+ $X2=29.35 $Y2=3.57
r2032 463 464 7.95791 $w=1.4e-07 $l=6.43e-06 $layer=MET1_cond $X=29.205 $Y=3.57
+ $X2=22.775 $Y2=3.57
r2033 462 495 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.775 $Y=1.87
+ $X2=22.63 $Y2=1.87
r2034 461 503 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.205 $Y=1.87
+ $X2=29.35 $Y2=1.87
r2035 461 462 7.95791 $w=1.4e-07 $l=6.43e-06 $layer=MET1_cond $X=29.205 $Y=1.87
+ $X2=22.775 $Y2=1.87
r2036 460 542 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=17.095 $Y=3.57
+ $X2=16.89 $Y2=3.57
r2037 459 544 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.545 $Y=3.57
+ $X2=21.69 $Y2=3.57
r2038 459 460 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=21.545 $Y=3.57
+ $X2=17.095 $Y2=3.57
r2039 458 541 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=17.095 $Y=1.87
+ $X2=16.89 $Y2=1.87
r2040 457 543 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.545 $Y=1.87
+ $X2=21.69 $Y2=1.87
r2041 457 458 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=21.545 $Y=1.87
+ $X2=17.095 $Y2=1.87
r2042 456 483 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.895 $Y=3.57
+ $X2=9.75 $Y2=3.57
r2043 455 491 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.865 $Y=3.57
+ $X2=16.01 $Y2=3.57
r2044 455 456 7.3886 $w=1.4e-07 $l=5.97e-06 $layer=MET1_cond $X=15.865 $Y=3.57
+ $X2=9.895 $Y2=3.57
r2045 454 479 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.895 $Y=1.87
+ $X2=9.75 $Y2=1.87
r2046 453 487 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.865 $Y=1.87
+ $X2=16.01 $Y2=1.87
r2047 453 454 7.3886 $w=1.4e-07 $l=5.97e-06 $layer=MET1_cond $X=15.865 $Y=1.87
+ $X2=9.895 $Y2=1.87
r2048 452 538 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=4.215 $Y=3.57
+ $X2=4.01 $Y2=3.57
r2049 451 540 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.665 $Y=3.57
+ $X2=8.81 $Y2=3.57
r2050 451 452 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=8.665 $Y=3.57
+ $X2=4.215 $Y2=3.57
r2051 450 537 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=4.215 $Y=1.87
+ $X2=4.01 $Y2=1.87
r2052 449 539 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.665 $Y=1.87
+ $X2=8.81 $Y2=1.87
r2053 449 450 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=8.665 $Y=1.87
+ $X2=4.215 $Y2=1.87
r2054 446 447 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=48.95 $Y=4.76
+ $X2=48.95 $Y2=4.555
r2055 442 444 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=48.95 $Y=0.68
+ $X2=48.95 $Y2=0.885
r2056 439 533 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=48.85 $Y=4.075
+ $X2=48.85 $Y2=3.57
r2057 439 440 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=48.85 $Y=4.075
+ $X2=48.85 $Y2=4.225
r2058 437 699 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=48.85 $Y=1.365
+ $X2=48.85 $Y2=1.7
r2059 437 438 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=48.85 $Y=1.365
+ $X2=48.85 $Y2=1.215
r2060 435 696 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=47.91 $Y=4.075
+ $X2=47.91 $Y2=3.57
r2061 435 436 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=47.91
+ $Y=4.075 $X2=48.01 $Y2=4.225
r2062 433 690 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=47.91 $Y=1.365
+ $X2=47.91 $Y2=1.7
r2063 433 434 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=47.91
+ $Y=1.365 $X2=48.01 $Y2=1.215
r2064 431 687 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=43.17 $Y=4.075
+ $X2=43.17 $Y2=3.57
r2065 431 432 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=43.17
+ $Y=4.075 $X2=43.07 $Y2=4.225
r2066 429 681 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=43.17 $Y=1.365
+ $X2=43.17 $Y2=1.7
r2067 429 430 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=43.17
+ $Y=1.365 $X2=43.07 $Y2=1.215
r2068 427 524 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=42.23 $Y=4.075
+ $X2=42.23 $Y2=3.57
r2069 427 428 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=42.23 $Y=4.075
+ $X2=42.23 $Y2=4.225
r2070 425 676 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=42.23 $Y=1.365
+ $X2=42.23 $Y2=1.7
r2071 425 426 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=42.23 $Y=1.365
+ $X2=42.23 $Y2=1.215
r2072 422 423 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=42.13 $Y=4.76
+ $X2=42.13 $Y2=4.555
r2073 418 420 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=42.13 $Y=0.68
+ $X2=42.13 $Y2=0.885
r2074 414 415 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=36.07 $Y=4.76
+ $X2=36.07 $Y2=4.555
r2075 410 412 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=36.07 $Y=0.68
+ $X2=36.07 $Y2=0.885
r2076 407 516 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=35.97 $Y=4.075
+ $X2=35.97 $Y2=3.57
r2077 407 408 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=35.97 $Y=4.075
+ $X2=35.97 $Y2=4.225
r2078 405 671 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=35.97 $Y=1.365
+ $X2=35.97 $Y2=1.7
r2079 405 406 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=35.97 $Y=1.365
+ $X2=35.97 $Y2=1.215
r2080 403 668 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=35.03 $Y=4.075
+ $X2=35.03 $Y2=3.57
r2081 403 404 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=35.03
+ $Y=4.075 $X2=35.13 $Y2=4.225
r2082 401 662 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=35.03 $Y=1.365
+ $X2=35.03 $Y2=1.7
r2083 401 402 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=35.03
+ $Y=1.365 $X2=35.13 $Y2=1.215
r2084 399 659 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=30.29 $Y=4.075
+ $X2=30.29 $Y2=3.57
r2085 399 400 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=30.29
+ $Y=4.075 $X2=30.19 $Y2=4.225
r2086 397 653 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=30.29 $Y=1.365
+ $X2=30.29 $Y2=1.7
r2087 397 398 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=30.29
+ $Y=1.365 $X2=30.19 $Y2=1.215
r2088 395 508 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=29.35 $Y=4.075
+ $X2=29.35 $Y2=3.57
r2089 395 396 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=29.35 $Y=4.075
+ $X2=29.35 $Y2=4.225
r2090 393 648 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=29.35 $Y=1.365
+ $X2=29.35 $Y2=1.7
r2091 393 394 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=29.35 $Y=1.365
+ $X2=29.35 $Y2=1.215
r2092 390 391 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=29.25 $Y=4.76
+ $X2=29.25 $Y2=4.555
r2093 386 388 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=29.25 $Y=0.68
+ $X2=29.25 $Y2=0.885
r2094 382 383 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=22.73 $Y=4.76
+ $X2=22.73 $Y2=4.555
r2095 378 380 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=22.73 $Y=0.68
+ $X2=22.73 $Y2=0.885
r2096 375 500 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=22.63 $Y=4.075
+ $X2=22.63 $Y2=3.57
r2097 375 376 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=22.63 $Y=4.075
+ $X2=22.63 $Y2=4.225
r2098 373 643 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=22.63 $Y=1.365
+ $X2=22.63 $Y2=1.7
r2099 373 374 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=22.63 $Y=1.365
+ $X2=22.63 $Y2=1.215
r2100 371 640 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=21.69 $Y=4.075
+ $X2=21.69 $Y2=3.57
r2101 371 372 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.69
+ $Y=4.075 $X2=21.79 $Y2=4.225
r2102 369 634 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=21.69 $Y=1.365
+ $X2=21.69 $Y2=1.7
r2103 369 370 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.69
+ $Y=1.365 $X2=21.79 $Y2=1.215
r2104 367 631 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=16.95 $Y=4.075
+ $X2=16.95 $Y2=3.57
r2105 367 368 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.95
+ $Y=4.075 $X2=16.85 $Y2=4.225
r2106 365 625 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=16.95 $Y=1.365
+ $X2=16.95 $Y2=1.7
r2107 365 366 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.95
+ $Y=1.365 $X2=16.85 $Y2=1.215
r2108 363 492 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=16.01 $Y=4.075
+ $X2=16.01 $Y2=3.57
r2109 363 364 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=16.01 $Y=4.075
+ $X2=16.01 $Y2=4.225
r2110 361 620 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=16.01 $Y=1.365
+ $X2=16.01 $Y2=1.7
r2111 361 362 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=16.01 $Y=1.365
+ $X2=16.01 $Y2=1.215
r2112 358 359 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.91 $Y=4.76
+ $X2=15.91 $Y2=4.555
r2113 354 356 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.91 $Y=0.68
+ $X2=15.91 $Y2=0.885
r2114 350 351 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.85 $Y=4.76
+ $X2=9.85 $Y2=4.555
r2115 346 348 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.85 $Y=0.68
+ $X2=9.85 $Y2=0.885
r2116 343 484 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.75 $Y=4.075
+ $X2=9.75 $Y2=3.57
r2117 343 344 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=9.75 $Y=4.075
+ $X2=9.75 $Y2=4.225
r2118 341 615 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.75 $Y=1.365
+ $X2=9.75 $Y2=1.7
r2119 341 342 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=9.75 $Y=1.365
+ $X2=9.75 $Y2=1.215
r2120 339 612 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=8.81 $Y=4.075
+ $X2=8.81 $Y2=3.57
r2121 339 340 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=8.81 $Y=4.075
+ $X2=8.91 $Y2=4.225
r2122 337 606 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.81 $Y=1.365
+ $X2=8.81 $Y2=1.7
r2123 337 338 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=8.81 $Y=1.365
+ $X2=8.91 $Y2=1.215
r2124 335 603 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=4.07 $Y=4.075
+ $X2=4.07 $Y2=3.57
r2125 335 336 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=4.07 $Y=4.075
+ $X2=3.97 $Y2=4.225
r2126 333 597 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=1.365
+ $X2=4.07 $Y2=1.7
r2127 333 334 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=4.07 $Y=1.365
+ $X2=3.97 $Y2=1.215
r2128 331 594 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=3.13 $Y=4.075
+ $X2=3.13 $Y2=3.57
r2129 331 332 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=4.075
+ $X2=3.13 $Y2=4.225
r2130 329 588 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.13 $Y=1.365
+ $X2=3.13 $Y2=1.7
r2131 329 330 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=1.365
+ $X2=3.13 $Y2=1.215
r2132 326 327 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.03 $Y=4.76
+ $X2=3.03 $Y2=4.555
r2133 322 324 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.03 $Y=0.68
+ $X2=3.03 $Y2=0.885
r2134 319 440 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=48.9 $Y=4.375
+ $X2=48.85 $Y2=4.225
r2135 319 447 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=48.9 $Y=4.375
+ $X2=48.9 $Y2=4.555
r2136 318 438 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=48.9 $Y=1.065
+ $X2=48.85 $Y2=1.215
r2137 318 444 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=48.9 $Y=1.065
+ $X2=48.9 $Y2=0.885
r2138 316 436 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=48.275 $Y=4.225
+ $X2=48.01 $Y2=4.225
r2139 315 440 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=48.685 $Y=4.225
+ $X2=48.85 $Y2=4.225
r2140 315 316 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=48.685 $Y=4.225
+ $X2=48.275 $Y2=4.225
r2141 314 434 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=48.275 $Y=1.215
+ $X2=48.01 $Y2=1.215
r2142 313 438 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=48.685 $Y=1.215
+ $X2=48.85 $Y2=1.215
r2143 313 314 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=48.685 $Y=1.215
+ $X2=48.275 $Y2=1.215
r2144 309 436 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=48.11
+ $Y=4.375 $X2=48.01 $Y2=4.225
r2145 309 311 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=48.11 $Y=4.375
+ $X2=48.11 $Y2=4.76
r2146 305 434 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=48.11
+ $Y=1.065 $X2=48.01 $Y2=1.215
r2147 305 307 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=48.11 $Y=1.065
+ $X2=48.11 $Y2=0.68
r2148 301 432 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=42.97
+ $Y=4.375 $X2=43.07 $Y2=4.225
r2149 301 303 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=42.97 $Y=4.375
+ $X2=42.97 $Y2=4.76
r2150 297 430 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=42.97
+ $Y=1.065 $X2=43.07 $Y2=1.215
r2151 297 299 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=42.97 $Y=1.065
+ $X2=42.97 $Y2=0.68
r2152 296 428 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=42.395 $Y=4.225
+ $X2=42.23 $Y2=4.225
r2153 295 432 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=42.805 $Y=4.225
+ $X2=43.07 $Y2=4.225
r2154 295 296 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=42.805 $Y=4.225
+ $X2=42.395 $Y2=4.225
r2155 294 426 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=42.395 $Y=1.215
+ $X2=42.23 $Y2=1.215
r2156 293 430 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=42.805 $Y=1.215
+ $X2=43.07 $Y2=1.215
r2157 293 294 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=42.805 $Y=1.215
+ $X2=42.395 $Y2=1.215
r2158 291 428 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=42.18
+ $Y=4.375 $X2=42.23 $Y2=4.225
r2159 291 423 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=42.18 $Y=4.375
+ $X2=42.18 $Y2=4.555
r2160 290 426 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=42.18
+ $Y=1.065 $X2=42.23 $Y2=1.215
r2161 290 420 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=42.18 $Y=1.065
+ $X2=42.18 $Y2=0.885
r2162 287 408 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=36.02
+ $Y=4.375 $X2=35.97 $Y2=4.225
r2163 287 415 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=36.02 $Y=4.375
+ $X2=36.02 $Y2=4.555
r2164 286 406 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=36.02
+ $Y=1.065 $X2=35.97 $Y2=1.215
r2165 286 412 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=36.02 $Y=1.065
+ $X2=36.02 $Y2=0.885
r2166 284 404 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=35.395 $Y=4.225
+ $X2=35.13 $Y2=4.225
r2167 283 408 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=35.805 $Y=4.225
+ $X2=35.97 $Y2=4.225
r2168 283 284 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=35.805 $Y=4.225
+ $X2=35.395 $Y2=4.225
r2169 282 402 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=35.395 $Y=1.215
+ $X2=35.13 $Y2=1.215
r2170 281 406 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=35.805 $Y=1.215
+ $X2=35.97 $Y2=1.215
r2171 281 282 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=35.805 $Y=1.215
+ $X2=35.395 $Y2=1.215
r2172 277 404 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=35.23
+ $Y=4.375 $X2=35.13 $Y2=4.225
r2173 277 279 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=35.23 $Y=4.375
+ $X2=35.23 $Y2=4.76
r2174 273 402 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=35.23
+ $Y=1.065 $X2=35.13 $Y2=1.215
r2175 273 275 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=35.23 $Y=1.065
+ $X2=35.23 $Y2=0.68
r2176 269 400 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=30.09
+ $Y=4.375 $X2=30.19 $Y2=4.225
r2177 269 271 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=30.09 $Y=4.375
+ $X2=30.09 $Y2=4.76
r2178 265 398 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=30.09
+ $Y=1.065 $X2=30.19 $Y2=1.215
r2179 265 267 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=30.09 $Y=1.065
+ $X2=30.09 $Y2=0.68
r2180 264 396 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=29.515 $Y=4.225
+ $X2=29.35 $Y2=4.225
r2181 263 400 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=29.925 $Y=4.225
+ $X2=30.19 $Y2=4.225
r2182 263 264 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=29.925 $Y=4.225
+ $X2=29.515 $Y2=4.225
r2183 262 394 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=29.515 $Y=1.215
+ $X2=29.35 $Y2=1.215
r2184 261 398 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=29.925 $Y=1.215
+ $X2=30.19 $Y2=1.215
r2185 261 262 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=29.925 $Y=1.215
+ $X2=29.515 $Y2=1.215
r2186 259 396 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=29.3 $Y=4.375
+ $X2=29.35 $Y2=4.225
r2187 259 391 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=29.3 $Y=4.375
+ $X2=29.3 $Y2=4.555
r2188 258 394 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=29.3 $Y=1.065
+ $X2=29.35 $Y2=1.215
r2189 258 388 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=29.3 $Y=1.065
+ $X2=29.3 $Y2=0.885
r2190 255 376 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=22.68
+ $Y=4.375 $X2=22.63 $Y2=4.225
r2191 255 383 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=22.68 $Y=4.375
+ $X2=22.68 $Y2=4.555
r2192 254 374 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=22.68
+ $Y=1.065 $X2=22.63 $Y2=1.215
r2193 254 380 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=22.68 $Y=1.065
+ $X2=22.68 $Y2=0.885
r2194 252 372 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=22.055 $Y=4.225
+ $X2=21.79 $Y2=4.225
r2195 251 376 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=22.465 $Y=4.225
+ $X2=22.63 $Y2=4.225
r2196 251 252 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=22.465 $Y=4.225
+ $X2=22.055 $Y2=4.225
r2197 250 370 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=22.055 $Y=1.215
+ $X2=21.79 $Y2=1.215
r2198 249 374 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=22.465 $Y=1.215
+ $X2=22.63 $Y2=1.215
r2199 249 250 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=22.465 $Y=1.215
+ $X2=22.055 $Y2=1.215
r2200 245 372 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.89
+ $Y=4.375 $X2=21.79 $Y2=4.225
r2201 245 247 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=21.89 $Y=4.375
+ $X2=21.89 $Y2=4.76
r2202 241 370 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.89
+ $Y=1.065 $X2=21.79 $Y2=1.215
r2203 241 243 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=21.89 $Y=1.065
+ $X2=21.89 $Y2=0.68
r2204 237 368 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.75
+ $Y=4.375 $X2=16.85 $Y2=4.225
r2205 237 239 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=16.75 $Y=4.375
+ $X2=16.75 $Y2=4.76
r2206 233 366 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.75
+ $Y=1.065 $X2=16.85 $Y2=1.215
r2207 233 235 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=16.75 $Y=1.065
+ $X2=16.75 $Y2=0.68
r2208 232 364 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.175 $Y=4.225
+ $X2=16.01 $Y2=4.225
r2209 231 368 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=16.585 $Y=4.225
+ $X2=16.85 $Y2=4.225
r2210 231 232 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=16.585 $Y=4.225
+ $X2=16.175 $Y2=4.225
r2211 230 362 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.175 $Y=1.215
+ $X2=16.01 $Y2=1.215
r2212 229 366 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=16.585 $Y=1.215
+ $X2=16.85 $Y2=1.215
r2213 229 230 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=16.585 $Y=1.215
+ $X2=16.175 $Y2=1.215
r2214 227 364 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=15.96
+ $Y=4.375 $X2=16.01 $Y2=4.225
r2215 227 359 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=15.96 $Y=4.375
+ $X2=15.96 $Y2=4.555
r2216 226 362 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=15.96
+ $Y=1.065 $X2=16.01 $Y2=1.215
r2217 226 356 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=15.96 $Y=1.065
+ $X2=15.96 $Y2=0.885
r2218 223 344 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=9.8 $Y=4.375
+ $X2=9.75 $Y2=4.225
r2219 223 351 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.8 $Y=4.375
+ $X2=9.8 $Y2=4.555
r2220 222 342 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=9.8 $Y=1.065
+ $X2=9.75 $Y2=1.215
r2221 222 348 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.8 $Y=1.065
+ $X2=9.8 $Y2=0.885
r2222 220 340 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=9.175 $Y=4.225
+ $X2=8.91 $Y2=4.225
r2223 219 344 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=4.225
+ $X2=9.75 $Y2=4.225
r2224 219 220 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=9.585 $Y=4.225
+ $X2=9.175 $Y2=4.225
r2225 218 338 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=9.175 $Y=1.215
+ $X2=8.91 $Y2=1.215
r2226 217 342 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=1.215
+ $X2=9.75 $Y2=1.215
r2227 217 218 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=9.585 $Y=1.215
+ $X2=9.175 $Y2=1.215
r2228 213 340 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.01 $Y=4.375
+ $X2=8.91 $Y2=4.225
r2229 213 215 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.01 $Y=4.375
+ $X2=9.01 $Y2=4.76
r2230 209 338 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.01 $Y=1.065
+ $X2=8.91 $Y2=1.215
r2231 209 211 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.01 $Y=1.065
+ $X2=9.01 $Y2=0.68
r2232 205 336 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=3.87 $Y=4.375
+ $X2=3.97 $Y2=4.225
r2233 205 207 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.87 $Y=4.375
+ $X2=3.87 $Y2=4.76
r2234 201 334 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.97 $Y2=1.215
r2235 201 203 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.87 $Y2=0.68
r2236 200 332 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=4.225
+ $X2=3.13 $Y2=4.225
r2237 199 336 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=3.705 $Y=4.225
+ $X2=3.97 $Y2=4.225
r2238 199 200 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.705 $Y=4.225
+ $X2=3.295 $Y2=4.225
r2239 198 330 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.215
+ $X2=3.13 $Y2=1.215
r2240 197 334 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=3.705 $Y=1.215
+ $X2=3.97 $Y2=1.215
r2241 197 198 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.705 $Y=1.215
+ $X2=3.295 $Y2=1.215
r2242 195 332 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.08 $Y=4.375
+ $X2=3.13 $Y2=4.225
r2243 195 327 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.08 $Y=4.375
+ $X2=3.08 $Y2=4.555
r2244 194 330 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.08 $Y=1.065
+ $X2=3.13 $Y2=1.215
r2245 194 324 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.08 $Y=1.065
+ $X2=3.08 $Y2=0.885
r2246 64 701 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=48.705 $Y=3.065 $X2=48.85 $Y2=3.21
r2247 63 699 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=48.705 $Y=1.555 $X2=48.85 $Y2=1.7
r2248 62 694 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=47.765 $Y=3.065 $X2=47.91 $Y2=3.21
r2249 61 690 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=47.765 $Y=1.555 $X2=47.91 $Y2=1.7
r2250 60 685 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=43.025 $Y=3.065 $X2=43.17 $Y2=3.21
r2251 59 681 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=43.025 $Y=1.555 $X2=43.17 $Y2=1.7
r2252 58 678 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=42.085 $Y=3.065 $X2=42.23 $Y2=3.21
r2253 57 676 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=42.085 $Y=1.555 $X2=42.23 $Y2=1.7
r2254 56 673 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=35.825 $Y=3.065 $X2=35.97 $Y2=3.21
r2255 55 671 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=35.825 $Y=1.555 $X2=35.97 $Y2=1.7
r2256 54 666 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=34.885 $Y=3.065 $X2=35.03 $Y2=3.21
r2257 53 662 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=34.885 $Y=1.555 $X2=35.03 $Y2=1.7
r2258 52 657 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=30.145 $Y=3.065 $X2=30.29 $Y2=3.21
r2259 51 653 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=30.145 $Y=1.555 $X2=30.29 $Y2=1.7
r2260 50 650 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=29.205 $Y=3.065 $X2=29.35 $Y2=3.21
r2261 49 648 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=29.205 $Y=1.555 $X2=29.35 $Y2=1.7
r2262 48 645 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=22.485 $Y=3.065 $X2=22.63 $Y2=3.21
r2263 47 643 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=22.485 $Y=1.555 $X2=22.63 $Y2=1.7
r2264 46 638 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=21.545 $Y=3.065 $X2=21.69 $Y2=3.21
r2265 45 634 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=21.545 $Y=1.555 $X2=21.69 $Y2=1.7
r2266 44 629 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=16.805 $Y=3.065 $X2=16.95 $Y2=3.21
r2267 43 625 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=16.805 $Y=1.555 $X2=16.95 $Y2=1.7
r2268 42 622 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=15.865 $Y=3.065 $X2=16.01 $Y2=3.21
r2269 41 620 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=15.865 $Y=1.555 $X2=16.01 $Y2=1.7
r2270 40 617 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=3.065 $X2=9.75 $Y2=3.21
r2271 39 615 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=1.555 $X2=9.75 $Y2=1.7
r2272 38 610 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.665
+ $Y=3.065 $X2=8.81 $Y2=3.21
r2273 37 606 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.665
+ $Y=1.555 $X2=8.81 $Y2=1.7
r2274 36 601 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=3.065 $X2=4.07 $Y2=3.21
r2275 35 597 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.555 $X2=4.07 $Y2=1.7
r2276 34 592 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=3.065 $X2=3.13 $Y2=3.21
r2277 33 588 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.555 $X2=3.13 $Y2=1.7
r2278 32 446 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=48.815 $Y=4.59 $X2=48.95 $Y2=4.76
r2279 31 442 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=48.815 $Y=0.33 $X2=48.95 $Y2=0.68
r2280 30 311 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=47.975 $Y=4.59 $X2=48.11 $Y2=4.76
r2281 29 307 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=47.975 $Y=0.33 $X2=48.11 $Y2=0.68
r2282 28 303 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=42.835 $Y=4.59 $X2=42.97 $Y2=4.76
r2283 27 299 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=42.835 $Y=0.33 $X2=42.97 $Y2=0.68
r2284 26 422 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=41.995 $Y=4.59 $X2=42.13 $Y2=4.76
r2285 25 418 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=41.995 $Y=0.33 $X2=42.13 $Y2=0.68
r2286 24 414 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=35.935 $Y=4.59 $X2=36.07 $Y2=4.76
r2287 23 410 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=35.935 $Y=0.33 $X2=36.07 $Y2=0.68
r2288 22 279 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=35.095 $Y=4.59 $X2=35.23 $Y2=4.76
r2289 21 275 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=35.095 $Y=0.33 $X2=35.23 $Y2=0.68
r2290 20 271 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=29.955 $Y=4.59 $X2=30.09 $Y2=4.76
r2291 19 267 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=29.955 $Y=0.33 $X2=30.09 $Y2=0.68
r2292 18 390 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=29.115 $Y=4.59 $X2=29.25 $Y2=4.76
r2293 17 386 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=29.115 $Y=0.33 $X2=29.25 $Y2=0.68
r2294 16 382 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=22.595 $Y=4.59 $X2=22.73 $Y2=4.76
r2295 15 378 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=22.595 $Y=0.33 $X2=22.73 $Y2=0.68
r2296 14 247 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=21.755 $Y=4.59 $X2=21.89 $Y2=4.76
r2297 13 243 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=21.755 $Y=0.33 $X2=21.89 $Y2=0.68
r2298 12 239 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=16.615 $Y=4.59 $X2=16.75 $Y2=4.76
r2299 11 235 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=16.615 $Y=0.33 $X2=16.75 $Y2=0.68
r2300 10 358 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=15.775 $Y=4.59 $X2=15.91 $Y2=4.76
r2301 9 354 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=15.775
+ $Y=0.33 $X2=15.91 $Y2=0.68
r2302 8 350 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=4.59 $X2=9.85 $Y2=4.76
r2303 7 346 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=0.33 $X2=9.85 $Y2=0.68
r2304 6 215 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=4.59 $X2=9.01 $Y2=4.76
r2305 5 211 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=0.33 $X2=9.01 $Y2=0.68
r2306 4 207 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=4.59 $X2=3.87 $Y2=4.76
r2307 3 203 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.33 $X2=3.87 $Y2=0.68
r2308 2 326 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=4.59 $X2=3.03 $Y2=4.76
r2309 1 322 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.33 $X2=3.03 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_311# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 47 49 50 53 58 63
c131 58 0 1.3204e-19 $X=9.28 $Y=1.7
c132 49 0 1.97849e-19 $X=12.15 $Y=2.225
c133 34 0 1.97849e-19 $X=11.355 $Y=2.225
c134 33 0 1.91515e-19 $X=12.005 $Y=2.225
c135 32 0 1.97167e-19 $X=10.375 $Y=2.225
c136 31 0 9.57576e-20 $X=11.065 $Y=2.225
c137 29 0 1.87597e-19 $X=10.085 $Y=2.225
c138 28 0 1.97167e-19 $X=8.475 $Y=2.225
c139 27 0 1.87597e-19 $X=9.135 $Y=2.225
r140 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.15 $Y=2.225
+ $X2=12.15 $Y2=2.225
r141 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.21 $Y=2.225
+ $X2=11.21 $Y2=2.225
r142 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=10.235 $Y=2.225
+ $X2=10.235 $Y2=1.7
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.23 $Y=2.225
+ $X2=10.23 $Y2=2.225
r144 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.28 $Y=2.225
+ $X2=9.28 $Y2=1.7
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=2.225
+ $X2=9.28 $Y2=2.225
r146 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=8.325 $Y=2.225
+ $X2=8.325 $Y2=1.73
r147 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.33 $Y=2.225
+ $X2=8.33 $Y2=2.225
r148 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.355 $Y=2.225
+ $X2=11.21 $Y2=2.225
r149 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.005 $Y=2.225
+ $X2=12.15 $Y2=2.225
r150 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=12.005 $Y=2.225
+ $X2=11.355 $Y2=2.225
r151 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.375 $Y=2.225
+ $X2=10.23 $Y2=2.225
r152 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.065 $Y=2.225
+ $X2=11.21 $Y2=2.225
r153 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=11.065 $Y=2.225
+ $X2=10.375 $Y2=2.225
r154 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.425 $Y=2.225
+ $X2=9.28 $Y2=2.225
r155 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.085 $Y=2.225
+ $X2=10.23 $Y2=2.225
r156 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=10.085 $Y=2.225
+ $X2=9.425 $Y2=2.225
r157 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.475 $Y=2.225
+ $X2=8.33 $Y2=2.225
r158 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.135 $Y=2.225
+ $X2=9.28 $Y2=2.225
r159 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=9.135 $Y=2.225
+ $X2=8.475 $Y2=2.225
r160 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=12.15 $Y=1.665
+ $X2=12.15 $Y2=2.225
r161 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.15 $Y=1.665
+ $X2=12.15 $Y2=1.58
r162 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=11.21 $Y=1.665
+ $X2=11.21 $Y2=2.225
r163 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=1.665
+ $X2=11.21 $Y2=1.58
r164 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=10.235 $Y=1.665
+ $X2=10.235 $Y2=1.7
r165 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=1.58
+ $X2=11.21 $Y2=1.58
r166 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=1.58
+ $X2=12.15 $Y2=1.58
r167 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=1.58
+ $X2=11.375 $Y2=1.58
r168 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.385 $Y=1.58
+ $X2=10.235 $Y2=1.665
r169 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=1.58
+ $X2=11.21 $Y2=1.58
r170 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.045 $Y=1.58
+ $X2=10.385 $Y2=1.58
r171 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=2.34
r172 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=1.66
r173 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.485 $X2=11.21 $Y2=2.34
r174 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.485 $X2=11.21 $Y2=1.66
r175 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.075
+ $Y=1.555 $X2=10.22 $Y2=1.7
r176 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.135
+ $Y=1.555 $X2=9.28 $Y2=1.7
r177 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=8.215
+ $Y=1.555 $X2=8.34 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_613# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 49 53 57 61 64 67
c131 57 0 1.3204e-19 $X=9.28 $Y=3.21
c132 49 0 1.97849e-19 $X=12.15 $Y=3.215
c133 34 0 1.97849e-19 $X=11.355 $Y=3.215
c134 33 0 1.91515e-19 $X=12.005 $Y=3.215
c135 32 0 1.97167e-19 $X=10.375 $Y=3.215
c136 31 0 9.57576e-20 $X=11.065 $Y=3.215
c137 29 0 1.87597e-19 $X=10.085 $Y=3.215
c138 28 0 1.97167e-19 $X=8.475 $Y=3.215
c139 27 0 1.87597e-19 $X=9.135 $Y=3.215
r140 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.15 $Y=3.215
+ $X2=12.15 $Y2=3.215
r141 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.21 $Y=3.215
+ $X2=11.21 $Y2=3.215
r142 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.23 $Y=3.215
+ $X2=10.23 $Y2=3.215
r143 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.28 $Y=3.215
+ $X2=9.28 $Y2=3.215
r144 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.33 $Y=3.215
+ $X2=8.33 $Y2=3.215
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.355 $Y=3.215
+ $X2=11.21 $Y2=3.215
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=12.005 $Y=3.215
+ $X2=12.15 $Y2=3.215
r147 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=12.005 $Y=3.215
+ $X2=11.355 $Y2=3.215
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.375 $Y=3.215
+ $X2=10.23 $Y2=3.215
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.065 $Y=3.215
+ $X2=11.21 $Y2=3.215
r150 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=11.065 $Y=3.215
+ $X2=10.375 $Y2=3.215
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.425 $Y=3.215
+ $X2=9.28 $Y2=3.215
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.085 $Y=3.215
+ $X2=10.23 $Y2=3.215
r153 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=10.085 $Y=3.215
+ $X2=9.425 $Y2=3.215
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.475 $Y=3.215
+ $X2=8.33 $Y2=3.215
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.135 $Y=3.215
+ $X2=9.28 $Y2=3.215
r156 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=9.135 $Y=3.215
+ $X2=8.475 $Y2=3.215
r157 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.15 $Y=3.775
+ $X2=12.15 $Y2=3.1
r158 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.15 $Y=3.775
+ $X2=12.15 $Y2=3.86
r159 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.21 $Y=3.775
+ $X2=11.21 $Y2=3.1
r160 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=3.775
+ $X2=11.21 $Y2=3.86
r161 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=10.235 $Y=3.775
+ $X2=10.235 $Y2=3.21
r162 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=3.86
+ $X2=11.21 $Y2=3.86
r163 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=3.86
+ $X2=12.15 $Y2=3.86
r164 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=3.86
+ $X2=11.375 $Y2=3.86
r165 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.385 $Y=3.86
+ $X2=10.235 $Y2=3.775
r166 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=3.86
+ $X2=11.21 $Y2=3.86
r167 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.045 $Y=3.86
+ $X2=10.385 $Y2=3.86
r168 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=2.955 $X2=12.15 $Y2=3.1
r169 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=2.955 $X2=12.15 $Y2=3.78
r170 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=2.955 $X2=11.21 $Y2=3.1
r171 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=2.955 $X2=11.21 $Y2=3.78
r172 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.075
+ $Y=3.065 $X2=10.22 $Y2=3.21
r173 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.135
+ $Y=3.065 $X2=9.28 $Y2=3.21
r174 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.215
+ $Y=3.065 $X2=8.34 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_297# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 37 41 49 59 63 68
c128 63 0 1.3204e-19 $X=16.48 $Y=1.7
c129 49 0 1.97167e-19 $X=17.43 $Y=2.225
c130 33 0 1.87597e-19 $X=17.285 $Y=2.225
c131 32 0 1.97167e-19 $X=15.675 $Y=2.225
c132 31 0 1.87597e-19 $X=16.335 $Y=2.225
c133 30 0 1.97849e-19 $X=14.695 $Y=2.225
c134 29 0 9.57576e-20 $X=15.385 $Y=2.225
c135 28 0 1.97849e-19 $X=13.755 $Y=2.225
c136 27 0 1.91515e-19 $X=14.405 $Y=2.225
r137 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=17.435 $Y=2.225
+ $X2=17.435 $Y2=1.73
r138 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.43 $Y=2.225
+ $X2=17.43 $Y2=2.225
r139 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=16.48 $Y=2.225
+ $X2=16.48 $Y2=1.7
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.48 $Y=2.225
+ $X2=16.48 $Y2=2.225
r141 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=15.525 $Y=2.225
+ $X2=15.525 $Y2=1.7
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.53 $Y=2.225
+ $X2=15.53 $Y2=2.225
r143 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.55 $Y=2.225
+ $X2=14.55 $Y2=2.225
r144 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.61 $Y=2.225
+ $X2=13.61 $Y2=2.225
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.625 $Y=2.225
+ $X2=16.48 $Y2=2.225
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.285 $Y=2.225
+ $X2=17.43 $Y2=2.225
r147 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=17.285 $Y=2.225
+ $X2=16.625 $Y2=2.225
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.675 $Y=2.225
+ $X2=15.53 $Y2=2.225
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.335 $Y=2.225
+ $X2=16.48 $Y2=2.225
r150 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=16.335 $Y=2.225
+ $X2=15.675 $Y2=2.225
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.695 $Y=2.225
+ $X2=14.55 $Y2=2.225
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.385 $Y=2.225
+ $X2=15.53 $Y2=2.225
r153 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=15.385 $Y=2.225
+ $X2=14.695 $Y2=2.225
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.755 $Y=2.225
+ $X2=13.61 $Y2=2.225
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.405 $Y=2.225
+ $X2=14.55 $Y2=2.225
r156 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=14.405 $Y=2.225
+ $X2=13.755 $Y2=2.225
r157 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=15.525 $Y=1.665
+ $X2=15.525 $Y2=1.7
r158 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=14.55 $Y=1.665
+ $X2=14.55 $Y2=2.225
r159 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.55 $Y=1.665
+ $X2=14.55 $Y2=1.58
r160 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=13.61 $Y=1.665
+ $X2=13.61 $Y2=2.225
r161 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.61 $Y=1.665
+ $X2=13.61 $Y2=1.58
r162 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=1.58
+ $X2=14.55 $Y2=1.58
r163 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=15.375 $Y=1.58
+ $X2=15.525 $Y2=1.665
r164 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=15.375 $Y=1.58
+ $X2=14.715 $Y2=1.58
r165 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.775 $Y=1.58
+ $X2=13.61 $Y2=1.58
r166 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=1.58
+ $X2=14.55 $Y2=1.58
r167 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=1.58
+ $X2=13.775 $Y2=1.58
r168 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=17.275
+ $Y=1.555 $X2=17.42 $Y2=1.73
r169 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.335
+ $Y=1.555 $X2=16.48 $Y2=1.7
r170 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=15.415
+ $Y=1.555 $X2=15.54 $Y2=1.7
r171 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=1.485 $X2=14.55 $Y2=2.34
r172 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=1.485 $X2=14.55 $Y2=1.66
r173 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=2.34
r174 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_591# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 49 53 56 59 62 66
c128 62 0 1.3204e-19 $X=16.48 $Y=3.21
c129 49 0 1.97167e-19 $X=17.43 $Y=3.215
c130 33 0 1.87597e-19 $X=17.285 $Y=3.215
c131 32 0 1.97167e-19 $X=15.675 $Y=3.215
c132 31 0 1.87597e-19 $X=16.335 $Y=3.215
c133 30 0 1.97849e-19 $X=14.695 $Y=3.215
c134 29 0 9.57576e-20 $X=15.385 $Y=3.215
c135 28 0 1.97849e-19 $X=13.755 $Y=3.215
c136 27 0 1.91515e-19 $X=14.405 $Y=3.215
r137 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.43 $Y=3.215
+ $X2=17.43 $Y2=3.215
r138 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.48 $Y=3.215
+ $X2=16.48 $Y2=3.215
r139 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.53 $Y=3.215
+ $X2=15.53 $Y2=3.215
r140 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.55 $Y=3.215
+ $X2=14.55 $Y2=3.215
r141 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.61 $Y=3.215
+ $X2=13.61 $Y2=3.215
r142 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.625 $Y=3.215
+ $X2=16.48 $Y2=3.215
r143 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.285 $Y=3.215
+ $X2=17.43 $Y2=3.215
r144 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=17.285 $Y=3.215
+ $X2=16.625 $Y2=3.215
r145 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.675 $Y=3.215
+ $X2=15.53 $Y2=3.215
r146 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.335 $Y=3.215
+ $X2=16.48 $Y2=3.215
r147 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=16.335 $Y=3.215
+ $X2=15.675 $Y2=3.215
r148 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.695 $Y=3.215
+ $X2=14.55 $Y2=3.215
r149 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.385 $Y=3.215
+ $X2=15.53 $Y2=3.215
r150 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=15.385 $Y=3.215
+ $X2=14.695 $Y2=3.215
r151 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.755 $Y=3.215
+ $X2=13.61 $Y2=3.215
r152 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.405 $Y=3.215
+ $X2=14.55 $Y2=3.215
r153 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=14.405 $Y=3.215
+ $X2=13.755 $Y2=3.215
r154 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=15.525 $Y=3.775
+ $X2=15.525 $Y2=3.21
r155 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.55 $Y=3.775
+ $X2=14.55 $Y2=3.1
r156 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.55 $Y=3.775
+ $X2=14.55 $Y2=3.86
r157 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.61 $Y=3.775
+ $X2=13.61 $Y2=3.1
r158 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.61 $Y=3.775
+ $X2=13.61 $Y2=3.86
r159 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=3.86
+ $X2=14.55 $Y2=3.86
r160 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=15.375 $Y=3.86
+ $X2=15.525 $Y2=3.775
r161 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=15.375 $Y=3.86
+ $X2=14.715 $Y2=3.86
r162 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.775 $Y=3.86
+ $X2=13.61 $Y2=3.86
r163 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=3.86
+ $X2=14.55 $Y2=3.86
r164 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=3.86
+ $X2=13.775 $Y2=3.86
r165 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=17.275
+ $Y=3.065 $X2=17.42 $Y2=3.21
r166 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.335
+ $Y=3.065 $X2=16.48 $Y2=3.21
r167 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=15.415
+ $Y=3.065 $X2=15.54 $Y2=3.21
r168 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=2.955 $X2=14.55 $Y2=3.1
r169 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=2.955 $X2=14.55 $Y2=3.78
r170 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=2.955 $X2=13.61 $Y2=3.1
r171 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=2.955 $X2=13.61 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_311# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 47 49 50 53 58 63
c131 58 0 1.3204e-19 $X=22.16 $Y=1.7
c132 49 0 1.97849e-19 $X=25.03 $Y=2.225
c133 34 0 1.97849e-19 $X=24.235 $Y=2.225
c134 33 0 1.91515e-19 $X=24.885 $Y=2.225
c135 32 0 1.97167e-19 $X=23.255 $Y=2.225
c136 31 0 9.57576e-20 $X=23.945 $Y=2.225
c137 29 0 1.87597e-19 $X=22.965 $Y=2.225
c138 28 0 1.97167e-19 $X=21.355 $Y=2.225
c139 27 0 1.87597e-19 $X=22.015 $Y=2.225
r140 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.03 $Y=2.225
+ $X2=25.03 $Y2=2.225
r141 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.09 $Y=2.225
+ $X2=24.09 $Y2=2.225
r142 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=23.115 $Y=2.225
+ $X2=23.115 $Y2=1.7
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.11 $Y=2.225
+ $X2=23.11 $Y2=2.225
r144 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=22.16 $Y=2.225
+ $X2=22.16 $Y2=1.7
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.16 $Y=2.225
+ $X2=22.16 $Y2=2.225
r146 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=21.205 $Y=2.225
+ $X2=21.205 $Y2=1.73
r147 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.21 $Y=2.225
+ $X2=21.21 $Y2=2.225
r148 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.235 $Y=2.225
+ $X2=24.09 $Y2=2.225
r149 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.885 $Y=2.225
+ $X2=25.03 $Y2=2.225
r150 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=24.885 $Y=2.225
+ $X2=24.235 $Y2=2.225
r151 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.255 $Y=2.225
+ $X2=23.11 $Y2=2.225
r152 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.945 $Y=2.225
+ $X2=24.09 $Y2=2.225
r153 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=23.945 $Y=2.225
+ $X2=23.255 $Y2=2.225
r154 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.305 $Y=2.225
+ $X2=22.16 $Y2=2.225
r155 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.965 $Y=2.225
+ $X2=23.11 $Y2=2.225
r156 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.965 $Y=2.225
+ $X2=22.305 $Y2=2.225
r157 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.355 $Y=2.225
+ $X2=21.21 $Y2=2.225
r158 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.015 $Y=2.225
+ $X2=22.16 $Y2=2.225
r159 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.015 $Y=2.225
+ $X2=21.355 $Y2=2.225
r160 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=25.03 $Y=1.665
+ $X2=25.03 $Y2=2.225
r161 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.03 $Y=1.665
+ $X2=25.03 $Y2=1.58
r162 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=24.09 $Y=1.665
+ $X2=24.09 $Y2=2.225
r163 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=24.09 $Y=1.665
+ $X2=24.09 $Y2=1.58
r164 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=23.115 $Y=1.665
+ $X2=23.115 $Y2=1.7
r165 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=1.58
+ $X2=24.09 $Y2=1.58
r166 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.865 $Y=1.58
+ $X2=25.03 $Y2=1.58
r167 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=1.58
+ $X2=24.255 $Y2=1.58
r168 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=23.265 $Y=1.58
+ $X2=23.115 $Y2=1.665
r169 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=1.58
+ $X2=24.09 $Y2=1.58
r170 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=23.925 $Y=1.58
+ $X2=23.265 $Y2=1.58
r171 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=2.34
r172 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=1.66
r173 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=1.485 $X2=24.09 $Y2=2.34
r174 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=1.485 $X2=24.09 $Y2=1.66
r175 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.955
+ $Y=1.555 $X2=23.1 $Y2=1.7
r176 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.015
+ $Y=1.555 $X2=22.16 $Y2=1.7
r177 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=21.095
+ $Y=1.555 $X2=21.22 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_613# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 49 53 57 61 64 67
c131 57 0 1.3204e-19 $X=22.16 $Y=3.21
c132 49 0 1.97849e-19 $X=25.03 $Y=3.215
c133 34 0 1.97849e-19 $X=24.235 $Y=3.215
c134 33 0 1.91515e-19 $X=24.885 $Y=3.215
c135 32 0 1.97167e-19 $X=23.255 $Y=3.215
c136 31 0 9.57576e-20 $X=23.945 $Y=3.215
c137 29 0 1.87597e-19 $X=22.965 $Y=3.215
c138 28 0 1.97167e-19 $X=21.355 $Y=3.215
c139 27 0 1.87597e-19 $X=22.015 $Y=3.215
r140 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.03 $Y=3.215
+ $X2=25.03 $Y2=3.215
r141 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.09 $Y=3.215
+ $X2=24.09 $Y2=3.215
r142 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.11 $Y=3.215
+ $X2=23.11 $Y2=3.215
r143 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.16 $Y=3.215
+ $X2=22.16 $Y2=3.215
r144 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.21 $Y=3.215
+ $X2=21.21 $Y2=3.215
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.235 $Y=3.215
+ $X2=24.09 $Y2=3.215
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.885 $Y=3.215
+ $X2=25.03 $Y2=3.215
r147 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=24.885 $Y=3.215
+ $X2=24.235 $Y2=3.215
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.255 $Y=3.215
+ $X2=23.11 $Y2=3.215
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=23.945 $Y=3.215
+ $X2=24.09 $Y2=3.215
r150 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=23.945 $Y=3.215
+ $X2=23.255 $Y2=3.215
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.305 $Y=3.215
+ $X2=22.16 $Y2=3.215
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.965 $Y=3.215
+ $X2=23.11 $Y2=3.215
r153 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.965 $Y=3.215
+ $X2=22.305 $Y2=3.215
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.355 $Y=3.215
+ $X2=21.21 $Y2=3.215
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.015 $Y=3.215
+ $X2=22.16 $Y2=3.215
r156 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.015 $Y=3.215
+ $X2=21.355 $Y2=3.215
r157 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=25.03 $Y=3.775
+ $X2=25.03 $Y2=3.1
r158 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.03 $Y=3.775
+ $X2=25.03 $Y2=3.86
r159 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=24.09 $Y=3.775
+ $X2=24.09 $Y2=3.1
r160 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=24.09 $Y=3.775
+ $X2=24.09 $Y2=3.86
r161 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=23.115 $Y=3.775
+ $X2=23.115 $Y2=3.21
r162 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=3.86
+ $X2=24.09 $Y2=3.86
r163 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.865 $Y=3.86
+ $X2=25.03 $Y2=3.86
r164 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=3.86
+ $X2=24.255 $Y2=3.86
r165 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=23.265 $Y=3.86
+ $X2=23.115 $Y2=3.775
r166 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=3.86
+ $X2=24.09 $Y2=3.86
r167 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=23.925 $Y=3.86
+ $X2=23.265 $Y2=3.86
r168 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=2.955 $X2=25.03 $Y2=3.1
r169 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=2.955 $X2=25.03 $Y2=3.78
r170 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=2.955 $X2=24.09 $Y2=3.1
r171 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=2.955 $X2=24.09 $Y2=3.78
r172 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.955
+ $Y=3.065 $X2=23.1 $Y2=3.21
r173 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.015
+ $Y=3.065 $X2=22.16 $Y2=3.21
r174 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=21.095
+ $Y=3.065 $X2=21.22 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_297# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 37 41 49 59 63 68
c128 63 0 1.3204e-19 $X=29.82 $Y=1.7
c129 49 0 1.97167e-19 $X=30.77 $Y=2.225
c130 33 0 1.87597e-19 $X=30.625 $Y=2.225
c131 32 0 1.97167e-19 $X=29.015 $Y=2.225
c132 31 0 1.87597e-19 $X=29.675 $Y=2.225
c133 30 0 1.97849e-19 $X=28.035 $Y=2.225
c134 29 0 9.57576e-20 $X=28.725 $Y=2.225
c135 28 0 1.97849e-19 $X=27.095 $Y=2.225
c136 27 0 1.91515e-19 $X=27.745 $Y=2.225
r137 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=30.775 $Y=2.225
+ $X2=30.775 $Y2=1.73
r138 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=30.77 $Y=2.225
+ $X2=30.77 $Y2=2.225
r139 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=29.82 $Y=2.225
+ $X2=29.82 $Y2=1.7
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=29.82 $Y=2.225
+ $X2=29.82 $Y2=2.225
r141 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=28.865 $Y=2.225
+ $X2=28.865 $Y2=1.7
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=28.87 $Y=2.225
+ $X2=28.87 $Y2=2.225
r143 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.89 $Y=2.225
+ $X2=27.89 $Y2=2.225
r144 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.95 $Y=2.225
+ $X2=26.95 $Y2=2.225
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.965 $Y=2.225
+ $X2=29.82 $Y2=2.225
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=30.625 $Y=2.225
+ $X2=30.77 $Y2=2.225
r147 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=30.625 $Y=2.225
+ $X2=29.965 $Y2=2.225
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.015 $Y=2.225
+ $X2=28.87 $Y2=2.225
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.675 $Y=2.225
+ $X2=29.82 $Y2=2.225
r150 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=29.675 $Y=2.225
+ $X2=29.015 $Y2=2.225
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=28.035 $Y=2.225
+ $X2=27.89 $Y2=2.225
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=28.725 $Y=2.225
+ $X2=28.87 $Y2=2.225
r153 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=28.725 $Y=2.225
+ $X2=28.035 $Y2=2.225
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=27.095 $Y=2.225
+ $X2=26.95 $Y2=2.225
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=27.745 $Y=2.225
+ $X2=27.89 $Y2=2.225
r156 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=27.745 $Y=2.225
+ $X2=27.095 $Y2=2.225
r157 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=28.865 $Y=1.665
+ $X2=28.865 $Y2=1.7
r158 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=27.89 $Y=1.665
+ $X2=27.89 $Y2=2.225
r159 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=27.89 $Y=1.665
+ $X2=27.89 $Y2=1.58
r160 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=26.95 $Y=1.665
+ $X2=26.95 $Y2=2.225
r161 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=26.95 $Y=1.665
+ $X2=26.95 $Y2=1.58
r162 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=28.055 $Y=1.58
+ $X2=27.89 $Y2=1.58
r163 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=28.715 $Y=1.58
+ $X2=28.865 $Y2=1.665
r164 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=28.715 $Y=1.58
+ $X2=28.055 $Y2=1.58
r165 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.115 $Y=1.58
+ $X2=26.95 $Y2=1.58
r166 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.725 $Y=1.58
+ $X2=27.89 $Y2=1.58
r167 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=27.725 $Y=1.58
+ $X2=27.115 $Y2=1.58
r168 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=30.615
+ $Y=1.555 $X2=30.76 $Y2=1.73
r169 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=29.675
+ $Y=1.555 $X2=29.82 $Y2=1.7
r170 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=28.755
+ $Y=1.555 $X2=28.88 $Y2=1.7
r171 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=27.745
+ $Y=1.485 $X2=27.89 $Y2=2.34
r172 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=27.745
+ $Y=1.485 $X2=27.89 $Y2=1.66
r173 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=26.805
+ $Y=1.485 $X2=26.95 $Y2=2.34
r174 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=26.805
+ $Y=1.485 $X2=26.95 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_591# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 49 53 56 59 62 66
c128 62 0 1.3204e-19 $X=29.82 $Y=3.21
c129 49 0 1.97167e-19 $X=30.77 $Y=3.215
c130 33 0 1.87597e-19 $X=30.625 $Y=3.215
c131 32 0 1.97167e-19 $X=29.015 $Y=3.215
c132 31 0 1.87597e-19 $X=29.675 $Y=3.215
c133 30 0 1.97849e-19 $X=28.035 $Y=3.215
c134 29 0 9.57576e-20 $X=28.725 $Y=3.215
c135 28 0 1.97849e-19 $X=27.095 $Y=3.215
c136 27 0 1.91515e-19 $X=27.745 $Y=3.215
r137 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=30.77 $Y=3.215
+ $X2=30.77 $Y2=3.215
r138 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=29.82 $Y=3.215
+ $X2=29.82 $Y2=3.215
r139 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=28.87 $Y=3.215
+ $X2=28.87 $Y2=3.215
r140 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.89 $Y=3.215
+ $X2=27.89 $Y2=3.215
r141 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.95 $Y=3.215
+ $X2=26.95 $Y2=3.215
r142 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.965 $Y=3.215
+ $X2=29.82 $Y2=3.215
r143 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=30.625 $Y=3.215
+ $X2=30.77 $Y2=3.215
r144 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=30.625 $Y=3.215
+ $X2=29.965 $Y2=3.215
r145 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.015 $Y=3.215
+ $X2=28.87 $Y2=3.215
r146 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=29.675 $Y=3.215
+ $X2=29.82 $Y2=3.215
r147 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=29.675 $Y=3.215
+ $X2=29.015 $Y2=3.215
r148 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=28.035 $Y=3.215
+ $X2=27.89 $Y2=3.215
r149 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=28.725 $Y=3.215
+ $X2=28.87 $Y2=3.215
r150 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=28.725 $Y=3.215
+ $X2=28.035 $Y2=3.215
r151 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=27.095 $Y=3.215
+ $X2=26.95 $Y2=3.215
r152 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=27.745 $Y=3.215
+ $X2=27.89 $Y2=3.215
r153 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=27.745 $Y=3.215
+ $X2=27.095 $Y2=3.215
r154 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=28.865 $Y=3.775
+ $X2=28.865 $Y2=3.21
r155 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=27.89 $Y=3.775
+ $X2=27.89 $Y2=3.1
r156 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=27.89 $Y=3.775
+ $X2=27.89 $Y2=3.86
r157 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=26.95 $Y=3.775
+ $X2=26.95 $Y2=3.1
r158 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=26.95 $Y=3.775
+ $X2=26.95 $Y2=3.86
r159 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=28.055 $Y=3.86
+ $X2=27.89 $Y2=3.86
r160 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=28.715 $Y=3.86
+ $X2=28.865 $Y2=3.775
r161 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=28.715 $Y=3.86
+ $X2=28.055 $Y2=3.86
r162 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.115 $Y=3.86
+ $X2=26.95 $Y2=3.86
r163 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.725 $Y=3.86
+ $X2=27.89 $Y2=3.86
r164 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=27.725 $Y=3.86
+ $X2=27.115 $Y2=3.86
r165 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=30.615
+ $Y=3.065 $X2=30.76 $Y2=3.21
r166 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=29.675
+ $Y=3.065 $X2=29.82 $Y2=3.21
r167 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=28.755
+ $Y=3.065 $X2=28.88 $Y2=3.21
r168 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=27.745
+ $Y=2.955 $X2=27.89 $Y2=3.1
r169 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=27.745
+ $Y=2.955 $X2=27.89 $Y2=3.78
r170 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=26.805
+ $Y=2.955 $X2=26.95 $Y2=3.1
r171 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=26.805
+ $Y=2.955 $X2=26.95 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_311# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 47 49 50 53 58 63
c131 58 0 1.3204e-19 $X=35.5 $Y=1.7
c132 49 0 1.97849e-19 $X=38.37 $Y=2.225
c133 34 0 1.97849e-19 $X=37.575 $Y=2.225
c134 33 0 1.91515e-19 $X=38.225 $Y=2.225
c135 32 0 1.97167e-19 $X=36.595 $Y=2.225
c136 31 0 9.57576e-20 $X=37.285 $Y=2.225
c137 29 0 1.87597e-19 $X=36.305 $Y=2.225
c138 28 0 1.97167e-19 $X=34.695 $Y=2.225
c139 27 0 1.87597e-19 $X=35.355 $Y=2.225
r140 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.37 $Y=2.225
+ $X2=38.37 $Y2=2.225
r141 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=37.43 $Y=2.225
+ $X2=37.43 $Y2=2.225
r142 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=36.455 $Y=2.225
+ $X2=36.455 $Y2=1.7
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=36.45 $Y=2.225
+ $X2=36.45 $Y2=2.225
r144 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=35.5 $Y=2.225
+ $X2=35.5 $Y2=1.7
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.5 $Y=2.225
+ $X2=35.5 $Y2=2.225
r146 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=34.545 $Y=2.225
+ $X2=34.545 $Y2=1.73
r147 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=34.55 $Y=2.225
+ $X2=34.55 $Y2=2.225
r148 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=37.575 $Y=2.225
+ $X2=37.43 $Y2=2.225
r149 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=38.225 $Y=2.225
+ $X2=38.37 $Y2=2.225
r150 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=38.225 $Y=2.225
+ $X2=37.575 $Y2=2.225
r151 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.595 $Y=2.225
+ $X2=36.45 $Y2=2.225
r152 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=37.285 $Y=2.225
+ $X2=37.43 $Y2=2.225
r153 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=37.285 $Y=2.225
+ $X2=36.595 $Y2=2.225
r154 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.645 $Y=2.225
+ $X2=35.5 $Y2=2.225
r155 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.305 $Y=2.225
+ $X2=36.45 $Y2=2.225
r156 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=36.305 $Y=2.225
+ $X2=35.645 $Y2=2.225
r157 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=34.695 $Y=2.225
+ $X2=34.55 $Y2=2.225
r158 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.355 $Y=2.225
+ $X2=35.5 $Y2=2.225
r159 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=35.355 $Y=2.225
+ $X2=34.695 $Y2=2.225
r160 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=38.37 $Y=1.665
+ $X2=38.37 $Y2=2.225
r161 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=38.37 $Y=1.665
+ $X2=38.37 $Y2=1.58
r162 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=37.43 $Y=1.665
+ $X2=37.43 $Y2=2.225
r163 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=37.43 $Y=1.665
+ $X2=37.43 $Y2=1.58
r164 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=36.455 $Y=1.665
+ $X2=36.455 $Y2=1.7
r165 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.595 $Y=1.58
+ $X2=37.43 $Y2=1.58
r166 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=38.205 $Y=1.58
+ $X2=38.37 $Y2=1.58
r167 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=38.205 $Y=1.58
+ $X2=37.595 $Y2=1.58
r168 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=36.605 $Y=1.58
+ $X2=36.455 $Y2=1.665
r169 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.265 $Y=1.58
+ $X2=37.43 $Y2=1.58
r170 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=37.265 $Y=1.58
+ $X2=36.605 $Y2=1.58
r171 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=38.225
+ $Y=1.485 $X2=38.37 $Y2=2.34
r172 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=38.225
+ $Y=1.485 $X2=38.37 $Y2=1.66
r173 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=37.285
+ $Y=1.485 $X2=37.43 $Y2=2.34
r174 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=37.285
+ $Y=1.485 $X2=37.43 $Y2=1.66
r175 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=36.295
+ $Y=1.555 $X2=36.44 $Y2=1.7
r176 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=35.355
+ $Y=1.555 $X2=35.5 $Y2=1.7
r177 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=34.435
+ $Y=1.555 $X2=34.56 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_613# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 49 53 57 61 64 67
c131 57 0 1.3204e-19 $X=35.5 $Y=3.21
c132 49 0 1.97849e-19 $X=38.37 $Y=3.215
c133 34 0 1.97849e-19 $X=37.575 $Y=3.215
c134 33 0 1.91515e-19 $X=38.225 $Y=3.215
c135 32 0 1.97167e-19 $X=36.595 $Y=3.215
c136 31 0 9.57576e-20 $X=37.285 $Y=3.215
c137 29 0 1.87597e-19 $X=36.305 $Y=3.215
c138 28 0 1.97167e-19 $X=34.695 $Y=3.215
c139 27 0 1.87597e-19 $X=35.355 $Y=3.215
r140 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.37 $Y=3.215
+ $X2=38.37 $Y2=3.215
r141 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=37.43 $Y=3.215
+ $X2=37.43 $Y2=3.215
r142 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=36.45 $Y=3.215
+ $X2=36.45 $Y2=3.215
r143 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=35.5 $Y=3.215
+ $X2=35.5 $Y2=3.215
r144 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=34.55 $Y=3.215
+ $X2=34.55 $Y2=3.215
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=37.575 $Y=3.215
+ $X2=37.43 $Y2=3.215
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=38.225 $Y=3.215
+ $X2=38.37 $Y2=3.215
r147 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=38.225 $Y=3.215
+ $X2=37.575 $Y2=3.215
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.595 $Y=3.215
+ $X2=36.45 $Y2=3.215
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=37.285 $Y=3.215
+ $X2=37.43 $Y2=3.215
r150 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=37.285 $Y=3.215
+ $X2=36.595 $Y2=3.215
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.645 $Y=3.215
+ $X2=35.5 $Y2=3.215
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=36.305 $Y=3.215
+ $X2=36.45 $Y2=3.215
r153 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=36.305 $Y=3.215
+ $X2=35.645 $Y2=3.215
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=34.695 $Y=3.215
+ $X2=34.55 $Y2=3.215
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=35.355 $Y=3.215
+ $X2=35.5 $Y2=3.215
r156 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=35.355 $Y=3.215
+ $X2=34.695 $Y2=3.215
r157 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=38.37 $Y=3.775
+ $X2=38.37 $Y2=3.1
r158 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=38.37 $Y=3.775
+ $X2=38.37 $Y2=3.86
r159 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=37.43 $Y=3.775
+ $X2=37.43 $Y2=3.1
r160 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=37.43 $Y=3.775
+ $X2=37.43 $Y2=3.86
r161 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=36.455 $Y=3.775
+ $X2=36.455 $Y2=3.21
r162 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.595 $Y=3.86
+ $X2=37.43 $Y2=3.86
r163 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=38.205 $Y=3.86
+ $X2=38.37 $Y2=3.86
r164 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=38.205 $Y=3.86
+ $X2=37.595 $Y2=3.86
r165 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=36.605 $Y=3.86
+ $X2=36.455 $Y2=3.775
r166 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.265 $Y=3.86
+ $X2=37.43 $Y2=3.86
r167 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=37.265 $Y=3.86
+ $X2=36.605 $Y2=3.86
r168 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=38.225
+ $Y=2.955 $X2=38.37 $Y2=3.1
r169 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=38.225
+ $Y=2.955 $X2=38.37 $Y2=3.78
r170 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=37.285
+ $Y=2.955 $X2=37.43 $Y2=3.1
r171 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=37.285
+ $Y=2.955 $X2=37.43 $Y2=3.78
r172 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=36.295
+ $Y=3.065 $X2=36.44 $Y2=3.21
r173 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=35.355
+ $Y=3.065 $X2=35.5 $Y2=3.21
r174 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=34.435
+ $Y=3.065 $X2=34.56 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_297# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 37 41 49 59 63 68
c128 63 0 1.3204e-19 $X=42.7 $Y=1.7
c129 49 0 1.97167e-19 $X=43.65 $Y=2.225
c130 33 0 1.87597e-19 $X=43.505 $Y=2.225
c131 32 0 1.97167e-19 $X=41.895 $Y=2.225
c132 31 0 1.87597e-19 $X=42.555 $Y=2.225
c133 30 0 1.97849e-19 $X=40.915 $Y=2.225
c134 29 0 9.57576e-20 $X=41.605 $Y=2.225
c135 28 0 1.97849e-19 $X=39.975 $Y=2.225
c136 27 0 1.91515e-19 $X=40.625 $Y=2.225
r137 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=43.655 $Y=2.225
+ $X2=43.655 $Y2=1.73
r138 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=43.65 $Y=2.225
+ $X2=43.65 $Y2=2.225
r139 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=42.7 $Y=2.225
+ $X2=42.7 $Y2=1.7
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=42.7 $Y=2.225
+ $X2=42.7 $Y2=2.225
r141 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=41.745 $Y=2.225
+ $X2=41.745 $Y2=1.7
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=41.75 $Y=2.225
+ $X2=41.75 $Y2=2.225
r143 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=40.77 $Y=2.225
+ $X2=40.77 $Y2=2.225
r144 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.83 $Y=2.225
+ $X2=39.83 $Y2=2.225
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.845 $Y=2.225
+ $X2=42.7 $Y2=2.225
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=43.505 $Y=2.225
+ $X2=43.65 $Y2=2.225
r147 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=43.505 $Y=2.225
+ $X2=42.845 $Y2=2.225
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=41.895 $Y=2.225
+ $X2=41.75 $Y2=2.225
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.555 $Y=2.225
+ $X2=42.7 $Y2=2.225
r150 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=42.555 $Y=2.225
+ $X2=41.895 $Y2=2.225
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=40.915 $Y=2.225
+ $X2=40.77 $Y2=2.225
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=41.605 $Y=2.225
+ $X2=41.75 $Y2=2.225
r153 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=41.605 $Y=2.225
+ $X2=40.915 $Y2=2.225
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=39.975 $Y=2.225
+ $X2=39.83 $Y2=2.225
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=40.625 $Y=2.225
+ $X2=40.77 $Y2=2.225
r156 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=40.625 $Y=2.225
+ $X2=39.975 $Y2=2.225
r157 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=41.745 $Y=1.665
+ $X2=41.745 $Y2=1.7
r158 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=40.77 $Y=1.665
+ $X2=40.77 $Y2=2.225
r159 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=40.77 $Y=1.665
+ $X2=40.77 $Y2=1.58
r160 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=39.83 $Y=1.665
+ $X2=39.83 $Y2=2.225
r161 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=39.83 $Y=1.665
+ $X2=39.83 $Y2=1.58
r162 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.935 $Y=1.58
+ $X2=40.77 $Y2=1.58
r163 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=41.595 $Y=1.58
+ $X2=41.745 $Y2=1.665
r164 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=41.595 $Y=1.58
+ $X2=40.935 $Y2=1.58
r165 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=39.995 $Y=1.58
+ $X2=39.83 $Y2=1.58
r166 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.605 $Y=1.58
+ $X2=40.77 $Y2=1.58
r167 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=40.605 $Y=1.58
+ $X2=39.995 $Y2=1.58
r168 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=43.495
+ $Y=1.555 $X2=43.64 $Y2=1.73
r169 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=42.555
+ $Y=1.555 $X2=42.7 $Y2=1.7
r170 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=41.635
+ $Y=1.555 $X2=41.76 $Y2=1.7
r171 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=40.625
+ $Y=1.485 $X2=40.77 $Y2=2.34
r172 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=40.625
+ $Y=1.485 $X2=40.77 $Y2=1.66
r173 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=39.685
+ $Y=1.485 $X2=39.83 $Y2=2.34
r174 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=39.685
+ $Y=1.485 $X2=39.83 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_591# 1 2 3 4 5 16 18 20 25 27
+ 28 29 30 31 32 33 34 49 53 56 59 62 66
c128 62 0 1.3204e-19 $X=42.7 $Y=3.21
c129 49 0 1.97167e-19 $X=43.65 $Y=3.215
c130 33 0 1.87597e-19 $X=43.505 $Y=3.215
c131 32 0 1.97167e-19 $X=41.895 $Y=3.215
c132 31 0 1.87597e-19 $X=42.555 $Y=3.215
c133 30 0 1.97849e-19 $X=40.915 $Y=3.215
c134 29 0 9.57576e-20 $X=41.605 $Y=3.215
c135 28 0 1.97849e-19 $X=39.975 $Y=3.215
c136 27 0 1.91515e-19 $X=40.625 $Y=3.215
r137 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=43.65 $Y=3.215
+ $X2=43.65 $Y2=3.215
r138 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=42.7 $Y=3.215
+ $X2=42.7 $Y2=3.215
r139 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=41.75 $Y=3.215
+ $X2=41.75 $Y2=3.215
r140 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=40.77 $Y=3.215
+ $X2=40.77 $Y2=3.215
r141 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.83 $Y=3.215
+ $X2=39.83 $Y2=3.215
r142 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.845 $Y=3.215
+ $X2=42.7 $Y2=3.215
r143 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=43.505 $Y=3.215
+ $X2=43.65 $Y2=3.215
r144 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=43.505 $Y=3.215
+ $X2=42.845 $Y2=3.215
r145 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=41.895 $Y=3.215
+ $X2=41.75 $Y2=3.215
r146 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=42.555 $Y=3.215
+ $X2=42.7 $Y2=3.215
r147 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=42.555 $Y=3.215
+ $X2=41.895 $Y2=3.215
r148 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=40.915 $Y=3.215
+ $X2=40.77 $Y2=3.215
r149 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=41.605 $Y=3.215
+ $X2=41.75 $Y2=3.215
r150 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=41.605 $Y=3.215
+ $X2=40.915 $Y2=3.215
r151 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=39.975 $Y=3.215
+ $X2=39.83 $Y2=3.215
r152 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=40.625 $Y=3.215
+ $X2=40.77 $Y2=3.215
r153 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=40.625 $Y=3.215
+ $X2=39.975 $Y2=3.215
r154 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=41.745 $Y=3.775
+ $X2=41.745 $Y2=3.21
r155 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=40.77 $Y=3.775
+ $X2=40.77 $Y2=3.1
r156 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=40.77 $Y=3.775
+ $X2=40.77 $Y2=3.86
r157 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=39.83 $Y=3.775
+ $X2=39.83 $Y2=3.1
r158 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=39.83 $Y=3.775
+ $X2=39.83 $Y2=3.86
r159 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.935 $Y=3.86
+ $X2=40.77 $Y2=3.86
r160 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=41.595 $Y=3.86
+ $X2=41.745 $Y2=3.775
r161 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=41.595 $Y=3.86
+ $X2=40.935 $Y2=3.86
r162 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=39.995 $Y=3.86
+ $X2=39.83 $Y2=3.86
r163 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.605 $Y=3.86
+ $X2=40.77 $Y2=3.86
r164 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=40.605 $Y=3.86
+ $X2=39.995 $Y2=3.86
r165 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=43.495
+ $Y=3.065 $X2=43.64 $Y2=3.21
r166 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=42.555
+ $Y=3.065 $X2=42.7 $Y2=3.21
r167 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=41.635
+ $Y=3.065 $X2=41.76 $Y2=3.21
r168 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=40.625
+ $Y=2.955 $X2=40.77 $Y2=3.1
r169 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=40.625
+ $Y=2.955 $X2=40.77 $Y2=3.78
r170 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=39.685
+ $Y=2.955 $X2=39.83 $Y2=3.1
r171 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=39.685
+ $Y=2.955 $X2=39.83 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_311# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 47 49 50 53 58 63
c119 58 0 1.3204e-19 $X=48.38 $Y=1.7
c120 49 0 1.97849e-19 $X=51.25 $Y=2.225
c121 34 0 1.97849e-19 $X=50.455 $Y=2.225
c122 32 0 1.97167e-19 $X=49.475 $Y=2.225
c123 31 0 1.36925e-19 $X=50.165 $Y=2.225
c124 29 0 1.87597e-19 $X=49.185 $Y=2.225
c125 28 0 1.97167e-19 $X=47.575 $Y=2.225
c126 27 0 1.87597e-19 $X=48.235 $Y=2.225
r127 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.25 $Y=2.225
+ $X2=51.25 $Y2=2.225
r128 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=50.31 $Y=2.225
+ $X2=50.31 $Y2=2.225
r129 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=49.335 $Y=2.225
+ $X2=49.335 $Y2=1.7
r130 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=49.33 $Y=2.225
+ $X2=49.33 $Y2=2.225
r131 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=48.38 $Y=2.225
+ $X2=48.38 $Y2=1.7
r132 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=48.38 $Y=2.225
+ $X2=48.38 $Y2=2.225
r133 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=47.425 $Y=2.225
+ $X2=47.425 $Y2=1.73
r134 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=47.43 $Y=2.225
+ $X2=47.43 $Y2=2.225
r135 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=50.455 $Y=2.225
+ $X2=50.31 $Y2=2.225
r136 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=51.105 $Y=2.225
+ $X2=51.25 $Y2=2.225
r137 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=51.105 $Y=2.225
+ $X2=50.455 $Y2=2.225
r138 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=49.475 $Y=2.225
+ $X2=49.33 $Y2=2.225
r139 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=50.165 $Y=2.225
+ $X2=50.31 $Y2=2.225
r140 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=50.165 $Y=2.225
+ $X2=49.475 $Y2=2.225
r141 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.525 $Y=2.225
+ $X2=48.38 $Y2=2.225
r142 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=49.185 $Y=2.225
+ $X2=49.33 $Y2=2.225
r143 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=49.185 $Y=2.225
+ $X2=48.525 $Y2=2.225
r144 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=47.575 $Y=2.225
+ $X2=47.43 $Y2=2.225
r145 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.235 $Y=2.225
+ $X2=48.38 $Y2=2.225
r146 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=48.235 $Y=2.225
+ $X2=47.575 $Y2=2.225
r147 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=51.25 $Y=1.665
+ $X2=51.25 $Y2=2.225
r148 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=51.25 $Y=1.665
+ $X2=51.25 $Y2=1.58
r149 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=50.31 $Y=1.665
+ $X2=50.31 $Y2=2.225
r150 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=50.31 $Y=1.665
+ $X2=50.31 $Y2=1.58
r151 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=49.335 $Y=1.665
+ $X2=49.335 $Y2=1.7
r152 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.475 $Y=1.58
+ $X2=50.31 $Y2=1.58
r153 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=51.085 $Y=1.58
+ $X2=51.25 $Y2=1.58
r154 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=51.085 $Y=1.58
+ $X2=50.475 $Y2=1.58
r155 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=49.485 $Y=1.58
+ $X2=49.335 $Y2=1.665
r156 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.145 $Y=1.58
+ $X2=50.31 $Y2=1.58
r157 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=50.145 $Y=1.58
+ $X2=49.485 $Y2=1.58
r158 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=51.105
+ $Y=1.485 $X2=51.25 $Y2=2.34
r159 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=51.105
+ $Y=1.485 $X2=51.25 $Y2=1.66
r160 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=50.165
+ $Y=1.485 $X2=50.31 $Y2=2.34
r161 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=50.165
+ $Y=1.485 $X2=50.31 $Y2=1.66
r162 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=49.175
+ $Y=1.555 $X2=49.32 $Y2=1.7
r163 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=48.235
+ $Y=1.555 $X2=48.38 $Y2=1.7
r164 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=47.315
+ $Y=1.555 $X2=47.44 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_613# 1 2 3 4 5 16 17 18 23 24
+ 27 28 29 30 31 32 33 34 49 53 57 61 64 67
c119 57 0 1.3204e-19 $X=48.38 $Y=3.21
c120 49 0 1.97849e-19 $X=51.25 $Y=3.215
c121 34 0 1.97849e-19 $X=50.455 $Y=3.215
c122 32 0 1.97167e-19 $X=49.475 $Y=3.215
c123 31 0 1.36925e-19 $X=50.165 $Y=3.215
c124 29 0 1.87597e-19 $X=49.185 $Y=3.215
c125 28 0 1.97167e-19 $X=47.575 $Y=3.215
c126 27 0 1.87597e-19 $X=48.235 $Y=3.215
r127 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.25 $Y=3.215
+ $X2=51.25 $Y2=3.215
r128 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=50.31 $Y=3.215
+ $X2=50.31 $Y2=3.215
r129 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=49.33 $Y=3.215
+ $X2=49.33 $Y2=3.215
r130 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=48.38 $Y=3.215
+ $X2=48.38 $Y2=3.215
r131 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=47.43 $Y=3.215
+ $X2=47.43 $Y2=3.215
r132 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=50.455 $Y=3.215
+ $X2=50.31 $Y2=3.215
r133 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=51.105 $Y=3.215
+ $X2=51.25 $Y2=3.215
r134 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=51.105 $Y=3.215
+ $X2=50.455 $Y2=3.215
r135 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=49.475 $Y=3.215
+ $X2=49.33 $Y2=3.215
r136 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=50.165 $Y=3.215
+ $X2=50.31 $Y2=3.215
r137 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=50.165 $Y=3.215
+ $X2=49.475 $Y2=3.215
r138 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.525 $Y=3.215
+ $X2=48.38 $Y2=3.215
r139 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=49.185 $Y=3.215
+ $X2=49.33 $Y2=3.215
r140 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=49.185 $Y=3.215
+ $X2=48.525 $Y2=3.215
r141 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=47.575 $Y=3.215
+ $X2=47.43 $Y2=3.215
r142 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=48.235 $Y=3.215
+ $X2=48.38 $Y2=3.215
r143 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=48.235 $Y=3.215
+ $X2=47.575 $Y2=3.215
r144 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=51.25 $Y=3.775
+ $X2=51.25 $Y2=3.1
r145 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=51.25 $Y=3.775
+ $X2=51.25 $Y2=3.86
r146 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=50.31 $Y=3.775
+ $X2=50.31 $Y2=3.1
r147 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=50.31 $Y=3.775
+ $X2=50.31 $Y2=3.86
r148 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=49.335 $Y=3.775
+ $X2=49.335 $Y2=3.21
r149 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.475 $Y=3.86
+ $X2=50.31 $Y2=3.86
r150 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=51.085 $Y=3.86
+ $X2=51.25 $Y2=3.86
r151 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=51.085 $Y=3.86
+ $X2=50.475 $Y2=3.86
r152 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=49.485 $Y=3.86
+ $X2=49.335 $Y2=3.775
r153 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.145 $Y=3.86
+ $X2=50.31 $Y2=3.86
r154 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=50.145 $Y=3.86
+ $X2=49.485 $Y2=3.86
r155 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=51.105
+ $Y=2.955 $X2=51.25 $Y2=3.1
r156 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=51.105
+ $Y=2.955 $X2=51.25 $Y2=3.78
r157 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=50.165
+ $Y=2.955 $X2=50.31 $Y2=3.1
r158 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=50.165
+ $Y=2.955 $X2=50.31 $Y2=3.78
r159 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=49.175
+ $Y=3.065 $X2=49.32 $Y2=3.21
r160 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=48.235
+ $Y=3.065 $X2=48.38 $Y2=3.21
r161 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=47.315
+ $Y=3.065 $X2=47.44 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62 63 64 65 66
+ 67 68 69 70 71 72 73 74 75 76 77 78 79 80 241 243 245 247 251 255 257 259 263
+ 267 271 275 279 283 287 291 295 299 303 307 311 315 319 323 325 327 331 335
+ 339 343 345 347 351 355 359 363 367 371 375 379 383 387 391 395 399 403 407
+ 411 415 419 423 427 429 431 435 439 443 447 451 455 459 463 467 471 475 479
+ 483 487 491 495 497 499 503 507 511 515 517 519 523 527 531 535 539 543 547
+ 551 555 559 563 567 571 575 577 579 581 583 586 587 589 590 592 593 595 596
+ 598 599 601 602 604 605 607 608 610 611 613 614 616 617 619 620 622 623 625
+ 626 628 629 631 632 634 635 637 638 640 641 643 644 646 647 649 650 652 653
+ 655 656 658 659 661 662 664 665 667 668 670 671 673 674 676 677 679 680 682
+ 683 685 686 688 689 691 692 694 695 697 698 700 701 703 704 705 706 707 708
+ 709 710 711 712 713 714 715 716 717 718 719 720 721 722 741 746 795 799 803
+ 808 813 818 867 871 875 880 885 890 895 900 949 953 957 962 967 972 1021 1025
+ 1029 1034 1046 1049 1052 1055 1058 1061 1064 1067 1070 1073 1076 1079 1082
+ 1085 1088 1091 1094 1097 1100 1103 1106 1109 1112 1115 1118 1121 1124 1127
+ 1130 1133 1136 1139 1142 1145 1148 1151
r1360 1151 1152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=50.83 $Y=5.44
+ $X2=50.83 $Y2=5.44
r1361 1148 1149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=50.83 $Y=0
+ $X2=50.83 $Y2=0
r1362 1145 1146 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=41.17 $Y=5.44
+ $X2=41.17 $Y2=5.44
r1363 1142 1143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=41.17 $Y=0
+ $X2=41.17 $Y2=0
r1364 1140 1146 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=40.25 $Y=5.44
+ $X2=41.17 $Y2=5.44
r1365 1139 1140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=40.25 $Y=5.44
+ $X2=40.25 $Y2=5.44
r1366 1137 1143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=40.25 $Y=0
+ $X2=41.17 $Y2=0
r1367 1136 1137 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=40.25 $Y=0
+ $X2=40.25 $Y2=0
r1368 1121 1122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=37.95 $Y=5.44
+ $X2=37.95 $Y2=5.44
r1369 1118 1119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=37.95 $Y=0
+ $X2=37.95 $Y2=0
r1370 1115 1116 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=28.29 $Y=5.44
+ $X2=28.29 $Y2=5.44
r1371 1112 1113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=28.29 $Y=0
+ $X2=28.29 $Y2=0
r1372 1110 1116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=27.37 $Y=5.44
+ $X2=28.29 $Y2=5.44
r1373 1109 1110 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.37 $Y=5.44
+ $X2=27.37 $Y2=5.44
r1374 1107 1113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=27.37 $Y=0
+ $X2=28.29 $Y2=0
r1375 1106 1107 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=27.37 $Y=0
+ $X2=27.37 $Y2=0
r1376 1091 1092 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=5.44
+ $X2=24.61 $Y2=5.44
r1377 1088 1089 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=0
+ $X2=24.61 $Y2=0
r1378 1085 1086 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=5.44
+ $X2=14.95 $Y2=5.44
r1379 1082 1083 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r1380 1080 1086 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=5.44
+ $X2=14.95 $Y2=5.44
r1381 1079 1080 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=5.44
+ $X2=14.03 $Y2=5.44
r1382 1077 1083 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.95 $Y2=0
r1383 1076 1077 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r1384 1061 1062 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=5.44
+ $X2=11.73 $Y2=5.44
r1385 1058 1059 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r1386 1055 1056 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=5.44
+ $X2=2.07 $Y2=5.44
r1387 1052 1053 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r1388 1050 1056 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=5.44
+ $X2=2.07 $Y2=5.44
r1389 1049 1050 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=5.44
+ $X2=1.15 $Y2=5.44
r1390 1047 1053 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r1391 1046 1047 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r1392 1038 1152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.29 $Y=5.44
+ $X2=50.83 $Y2=5.44
r1393 1037 1038 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.29 $Y=5.44
+ $X2=51.29 $Y2=5.44
r1394 1035 1151 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.915 $Y=5.44
+ $X2=50.78 $Y2=5.44
r1395 1035 1037 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=50.915
+ $Y=5.44 $X2=51.29 $Y2=5.44
r1396 1034 1157 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=51.585 $Y=5.44
+ $X2=51.782 $Y2=5.44
r1397 1034 1037 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=51.585 $Y=5.44
+ $X2=51.29 $Y2=5.44
r1398 1033 1149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.29 $Y=0
+ $X2=50.83 $Y2=0
r1399 1032 1033 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.29 $Y=0
+ $X2=51.29 $Y2=0
r1400 1030 1148 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.915 $Y=0
+ $X2=50.78 $Y2=0
r1401 1030 1032 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=50.915 $Y=0
+ $X2=51.29 $Y2=0
r1402 1029 1154 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=51.585 $Y=0
+ $X2=51.782 $Y2=0
r1403 1029 1032 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=51.585 $Y=0
+ $X2=51.29 $Y2=0
r1404 1028 1152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=50.37 $Y=5.44
+ $X2=50.83 $Y2=5.44
r1405 1027 1028 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=50.37 $Y=5.44
+ $X2=50.37 $Y2=5.44
r1406 1025 1151 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.645 $Y=5.44
+ $X2=50.78 $Y2=5.44
r1407 1025 1027 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=50.645
+ $Y=5.44 $X2=50.37 $Y2=5.44
r1408 1024 1149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=50.37 $Y=0
+ $X2=50.83 $Y2=0
r1409 1023 1024 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=50.37 $Y=0
+ $X2=50.37 $Y2=0
r1410 1021 1148 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=50.645 $Y=0
+ $X2=50.78 $Y2=0
r1411 1021 1023 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=50.645 $Y=0
+ $X2=50.37 $Y2=0
r1412 1020 1028 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=49.45 $Y=5.44
+ $X2=50.37 $Y2=5.44
r1413 1019 1020 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=49.45 $Y=5.44
+ $X2=49.45 $Y2=5.44
r1414 1017 1020 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=47.15 $Y=5.44
+ $X2=49.45 $Y2=5.44
r1415 1016 1019 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=47.15 $Y=5.44
+ $X2=49.45 $Y2=5.44
r1416 1016 1017 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=47.15 $Y=5.44
+ $X2=47.15 $Y2=5.44
r1417 1014 1024 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=49.45 $Y=0
+ $X2=50.37 $Y2=0
r1418 1013 1014 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=49.45 $Y=0
+ $X2=49.45 $Y2=0
r1419 1011 1014 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=47.15 $Y=0
+ $X2=49.45 $Y2=0
r1420 1010 1013 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=47.15 $Y=0
+ $X2=49.45 $Y2=0
r1421 1010 1011 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=47.15 $Y=0
+ $X2=47.15 $Y2=0
r1422 1008 1017 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=46.69 $Y=5.44
+ $X2=47.15 $Y2=5.44
r1423 1007 1008 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=46.69 $Y=5.44
+ $X2=46.69 $Y2=5.44
r1424 1005 1011 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=46.69 $Y=0
+ $X2=47.15 $Y2=0
r1425 1004 1005 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=46.69 $Y=0
+ $X2=46.69 $Y2=0
r1426 1002 1008 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=45.77 $Y=5.44
+ $X2=46.69 $Y2=5.44
r1427 1001 1002 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=45.77 $Y=5.44
+ $X2=45.77 $Y2=5.44
r1428 999 1005 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=45.77 $Y=0
+ $X2=46.69 $Y2=0
r1429 998 999 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=45.77 $Y=0
+ $X2=45.77 $Y2=0
r1430 996 1002 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=44.85 $Y=5.44
+ $X2=45.77 $Y2=5.44
r1431 995 996 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=44.85 $Y=5.44
+ $X2=44.85 $Y2=5.44
r1432 993 999 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=44.85 $Y=0
+ $X2=45.77 $Y2=0
r1433 992 993 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=44.85 $Y=0
+ $X2=44.85 $Y2=0
r1434 990 996 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=43.93 $Y=5.44
+ $X2=44.85 $Y2=5.44
r1435 989 990 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=43.93 $Y=5.44
+ $X2=43.93 $Y2=5.44
r1436 987 990 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=41.63 $Y=5.44
+ $X2=43.93 $Y2=5.44
r1437 987 1146 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=41.63 $Y=5.44
+ $X2=41.17 $Y2=5.44
r1438 986 989 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=41.63 $Y=5.44
+ $X2=43.93 $Y2=5.44
r1439 986 987 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=41.63 $Y=5.44
+ $X2=41.63 $Y2=5.44
r1440 984 1145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=41.355 $Y=5.44
+ $X2=41.23 $Y2=5.44
r1441 984 986 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=41.355 $Y=5.44
+ $X2=41.63 $Y2=5.44
r1442 983 993 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=43.93 $Y=0
+ $X2=44.85 $Y2=0
r1443 982 983 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=43.93 $Y=0
+ $X2=43.93 $Y2=0
r1444 980 983 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=41.63 $Y=0
+ $X2=43.93 $Y2=0
r1445 980 1143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=41.63 $Y=0
+ $X2=41.17 $Y2=0
r1446 979 982 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=41.63 $Y=0
+ $X2=43.93 $Y2=0
r1447 979 980 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=41.63 $Y=0
+ $X2=41.63 $Y2=0
r1448 977 1142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=41.355 $Y=0
+ $X2=41.23 $Y2=0
r1449 977 979 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=41.355 $Y=0
+ $X2=41.63 $Y2=0
r1450 976 1140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.79 $Y=5.44
+ $X2=40.25 $Y2=5.44
r1451 975 976 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.79 $Y=5.44
+ $X2=39.79 $Y2=5.44
r1452 973 1133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=39.495 $Y=5.44
+ $X2=39.37 $Y2=5.44
r1453 973 975 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=39.495 $Y=5.44
+ $X2=39.79 $Y2=5.44
r1454 972 1139 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.165 $Y=5.44
+ $X2=40.3 $Y2=5.44
r1455 972 975 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=40.165 $Y=5.44
+ $X2=39.79 $Y2=5.44
r1456 971 1137 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.79 $Y=0
+ $X2=40.25 $Y2=0
r1457 970 971 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.79 $Y=0
+ $X2=39.79 $Y2=0
r1458 968 1130 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=39.495 $Y=0
+ $X2=39.37 $Y2=0
r1459 968 970 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=39.495 $Y=0
+ $X2=39.79 $Y2=0
r1460 967 1136 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.165 $Y=0
+ $X2=40.3 $Y2=0
r1461 967 970 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=40.165 $Y=0
+ $X2=39.79 $Y2=0
r1462 966 1122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.41 $Y=5.44
+ $X2=37.95 $Y2=5.44
r1463 965 966 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.41 $Y=5.44
+ $X2=38.41 $Y2=5.44
r1464 963 1121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=38.035 $Y=5.44
+ $X2=37.9 $Y2=5.44
r1465 963 965 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=38.035 $Y=5.44
+ $X2=38.41 $Y2=5.44
r1466 962 1127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=38.705 $Y=5.44
+ $X2=38.83 $Y2=5.44
r1467 962 965 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=38.705 $Y=5.44
+ $X2=38.41 $Y2=5.44
r1468 961 1119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.41 $Y=0
+ $X2=37.95 $Y2=0
r1469 960 961 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.41 $Y=0
+ $X2=38.41 $Y2=0
r1470 958 1118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=38.035 $Y=0
+ $X2=37.9 $Y2=0
r1471 958 960 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=38.035 $Y=0
+ $X2=38.41 $Y2=0
r1472 957 1124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=38.705 $Y=0
+ $X2=38.83 $Y2=0
r1473 957 960 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=38.705 $Y=0
+ $X2=38.41 $Y2=0
r1474 956 1122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=37.49 $Y=5.44
+ $X2=37.95 $Y2=5.44
r1475 955 956 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=37.49 $Y=5.44
+ $X2=37.49 $Y2=5.44
r1476 953 1121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=37.765 $Y=5.44
+ $X2=37.9 $Y2=5.44
r1477 953 955 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=37.765 $Y=5.44
+ $X2=37.49 $Y2=5.44
r1478 952 1119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=37.49 $Y=0
+ $X2=37.95 $Y2=0
r1479 951 952 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=37.49 $Y=0
+ $X2=37.49 $Y2=0
r1480 949 1118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=37.765 $Y=0
+ $X2=37.9 $Y2=0
r1481 949 951 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=37.765 $Y=0
+ $X2=37.49 $Y2=0
r1482 948 956 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=36.57 $Y=5.44
+ $X2=37.49 $Y2=5.44
r1483 947 948 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=36.57 $Y=5.44
+ $X2=36.57 $Y2=5.44
r1484 945 948 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=34.27 $Y=5.44
+ $X2=36.57 $Y2=5.44
r1485 944 947 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=34.27 $Y=5.44
+ $X2=36.57 $Y2=5.44
r1486 944 945 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=34.27 $Y=5.44
+ $X2=34.27 $Y2=5.44
r1487 942 952 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=36.57 $Y=0
+ $X2=37.49 $Y2=0
r1488 941 942 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=36.57 $Y=0
+ $X2=36.57 $Y2=0
r1489 939 942 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=34.27 $Y=0
+ $X2=36.57 $Y2=0
r1490 938 941 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=34.27 $Y=0
+ $X2=36.57 $Y2=0
r1491 938 939 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=34.27 $Y=0
+ $X2=34.27 $Y2=0
r1492 936 945 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=33.81 $Y=5.44
+ $X2=34.27 $Y2=5.44
r1493 935 936 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=33.81 $Y=5.44
+ $X2=33.81 $Y2=5.44
r1494 933 939 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=33.81 $Y=0
+ $X2=34.27 $Y2=0
r1495 932 933 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=33.81 $Y=0
+ $X2=33.81 $Y2=0
r1496 930 936 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=32.89 $Y=5.44
+ $X2=33.81 $Y2=5.44
r1497 929 930 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=32.89 $Y=5.44
+ $X2=32.89 $Y2=5.44
r1498 927 933 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=32.89 $Y=0
+ $X2=33.81 $Y2=0
r1499 926 927 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=32.89 $Y=0
+ $X2=32.89 $Y2=0
r1500 924 930 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.97 $Y=5.44
+ $X2=32.89 $Y2=5.44
r1501 923 924 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=31.97 $Y=5.44
+ $X2=31.97 $Y2=5.44
r1502 921 927 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.97 $Y=0
+ $X2=32.89 $Y2=0
r1503 920 921 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=31.97 $Y=0
+ $X2=31.97 $Y2=0
r1504 918 924 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.05 $Y=5.44
+ $X2=31.97 $Y2=5.44
r1505 917 918 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=31.05 $Y=5.44
+ $X2=31.05 $Y2=5.44
r1506 915 918 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=28.75 $Y=5.44
+ $X2=31.05 $Y2=5.44
r1507 915 1116 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=28.75 $Y=5.44
+ $X2=28.29 $Y2=5.44
r1508 914 917 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=28.75 $Y=5.44
+ $X2=31.05 $Y2=5.44
r1509 914 915 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=28.75 $Y=5.44
+ $X2=28.75 $Y2=5.44
r1510 912 1115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=28.475 $Y=5.44
+ $X2=28.35 $Y2=5.44
r1511 912 914 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=28.475 $Y=5.44
+ $X2=28.75 $Y2=5.44
r1512 911 921 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=31.05 $Y=0
+ $X2=31.97 $Y2=0
r1513 910 911 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=31.05 $Y=0
+ $X2=31.05 $Y2=0
r1514 908 911 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=28.75 $Y=0
+ $X2=31.05 $Y2=0
r1515 908 1113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=28.75 $Y=0
+ $X2=28.29 $Y2=0
r1516 907 910 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=28.75 $Y=0
+ $X2=31.05 $Y2=0
r1517 907 908 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=28.75 $Y=0
+ $X2=28.75 $Y2=0
r1518 905 1112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=28.475 $Y=0
+ $X2=28.35 $Y2=0
r1519 905 907 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=28.475 $Y=0
+ $X2=28.75 $Y2=0
r1520 904 1110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.91 $Y=5.44
+ $X2=27.37 $Y2=5.44
r1521 903 904 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.91 $Y=5.44
+ $X2=26.91 $Y2=5.44
r1522 901 1103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=26.615 $Y=5.44
+ $X2=26.49 $Y2=5.44
r1523 901 903 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=26.615 $Y=5.44
+ $X2=26.91 $Y2=5.44
r1524 900 1109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.285 $Y=5.44
+ $X2=27.42 $Y2=5.44
r1525 900 903 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=27.285 $Y=5.44
+ $X2=26.91 $Y2=5.44
r1526 899 1107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.91 $Y=0
+ $X2=27.37 $Y2=0
r1527 898 899 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.91 $Y=0
+ $X2=26.91 $Y2=0
r1528 896 1100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=26.615 $Y=0
+ $X2=26.49 $Y2=0
r1529 896 898 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=26.615 $Y=0
+ $X2=26.91 $Y2=0
r1530 895 1106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.285 $Y=0
+ $X2=27.42 $Y2=0
r1531 895 898 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=27.285 $Y=0
+ $X2=26.91 $Y2=0
r1532 891 1097 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=25.615 $Y=5.44
+ $X2=25.49 $Y2=5.44
r1533 891 893 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=25.615 $Y=5.44
+ $X2=25.99 $Y2=5.44
r1534 890 1103 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=26.365 $Y=5.44
+ $X2=26.49 $Y2=5.44
r1535 890 893 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=26.365 $Y=5.44
+ $X2=25.99 $Y2=5.44
r1536 886 1094 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=25.615 $Y=0
+ $X2=25.49 $Y2=0
r1537 886 888 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=25.615 $Y=0
+ $X2=25.99 $Y2=0
r1538 885 1100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=26.365 $Y=0
+ $X2=26.49 $Y2=0
r1539 885 888 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=26.365 $Y=0
+ $X2=25.99 $Y2=0
r1540 884 1092 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.07 $Y=5.44
+ $X2=24.61 $Y2=5.44
r1541 883 884 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=5.44
+ $X2=25.07 $Y2=5.44
r1542 881 1091 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.695 $Y=5.44
+ $X2=24.56 $Y2=5.44
r1543 881 883 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=24.695 $Y=5.44
+ $X2=25.07 $Y2=5.44
r1544 880 1097 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=25.365 $Y=5.44
+ $X2=25.49 $Y2=5.44
r1545 880 883 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.365 $Y=5.44
+ $X2=25.07 $Y2=5.44
r1546 879 1089 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.07 $Y=0
+ $X2=24.61 $Y2=0
r1547 878 879 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=0
+ $X2=25.07 $Y2=0
r1548 876 1088 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.695 $Y=0
+ $X2=24.56 $Y2=0
r1549 876 878 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=24.695 $Y=0
+ $X2=25.07 $Y2=0
r1550 875 1094 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=25.365 $Y=0
+ $X2=25.49 $Y2=0
r1551 875 878 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.365 $Y=0
+ $X2=25.07 $Y2=0
r1552 874 1092 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=5.44
+ $X2=24.61 $Y2=5.44
r1553 873 874 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=5.44
+ $X2=24.15 $Y2=5.44
r1554 871 1091 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.425 $Y=5.44
+ $X2=24.56 $Y2=5.44
r1555 871 873 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=24.425 $Y=5.44
+ $X2=24.15 $Y2=5.44
r1556 870 1089 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=0
+ $X2=24.61 $Y2=0
r1557 869 870 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=0
+ $X2=24.15 $Y2=0
r1558 867 1088 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.425 $Y=0
+ $X2=24.56 $Y2=0
r1559 867 869 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=24.425 $Y=0
+ $X2=24.15 $Y2=0
r1560 866 874 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=5.44
+ $X2=24.15 $Y2=5.44
r1561 865 866 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=5.44
+ $X2=23.23 $Y2=5.44
r1562 863 866 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=5.44
+ $X2=23.23 $Y2=5.44
r1563 862 865 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=5.44
+ $X2=23.23 $Y2=5.44
r1564 862 863 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=5.44
+ $X2=20.93 $Y2=5.44
r1565 860 870 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=0
+ $X2=24.15 $Y2=0
r1566 859 860 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=0
+ $X2=23.23 $Y2=0
r1567 857 860 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r1568 856 859 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r1569 856 857 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=0
+ $X2=20.93 $Y2=0
r1570 854 863 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=5.44
+ $X2=20.93 $Y2=5.44
r1571 853 854 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=5.44
+ $X2=20.47 $Y2=5.44
r1572 851 857 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=20.93 $Y2=0
r1573 850 851 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=0
+ $X2=20.47 $Y2=0
r1574 848 854 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=5.44
+ $X2=20.47 $Y2=5.44
r1575 847 848 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=5.44
+ $X2=19.55 $Y2=5.44
r1576 845 851 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=0
+ $X2=20.47 $Y2=0
r1577 844 845 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=0
+ $X2=19.55 $Y2=0
r1578 842 848 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=18.63 $Y=5.44
+ $X2=19.55 $Y2=5.44
r1579 841 842 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=5.44
+ $X2=18.63 $Y2=5.44
r1580 839 845 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=18.63 $Y=0
+ $X2=19.55 $Y2=0
r1581 838 839 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=0
+ $X2=18.63 $Y2=0
r1582 836 842 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.71 $Y=5.44
+ $X2=18.63 $Y2=5.44
r1583 835 836 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=17.71 $Y=5.44
+ $X2=17.71 $Y2=5.44
r1584 833 836 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=15.41 $Y=5.44
+ $X2=17.71 $Y2=5.44
r1585 833 1086 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=5.44
+ $X2=14.95 $Y2=5.44
r1586 832 835 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=15.41 $Y=5.44
+ $X2=17.71 $Y2=5.44
r1587 832 833 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=15.41 $Y=5.44
+ $X2=15.41 $Y2=5.44
r1588 830 1085 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.135 $Y=5.44
+ $X2=15.01 $Y2=5.44
r1589 830 832 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.135 $Y=5.44
+ $X2=15.41 $Y2=5.44
r1590 829 839 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.71 $Y=0
+ $X2=18.63 $Y2=0
r1591 828 829 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=17.71 $Y=0
+ $X2=17.71 $Y2=0
r1592 826 829 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=17.71 $Y2=0
r1593 826 1083 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=14.95 $Y2=0
r1594 825 828 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=15.41 $Y=0
+ $X2=17.71 $Y2=0
r1595 825 826 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r1596 823 1082 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.135 $Y=0
+ $X2=15.01 $Y2=0
r1597 823 825 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.135 $Y=0
+ $X2=15.41 $Y2=0
r1598 822 1080 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=5.44
+ $X2=14.03 $Y2=5.44
r1599 821 822 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=5.44
+ $X2=13.57 $Y2=5.44
r1600 819 1073 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.275 $Y=5.44
+ $X2=13.15 $Y2=5.44
r1601 819 821 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.275 $Y=5.44
+ $X2=13.57 $Y2=5.44
r1602 818 1079 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.945 $Y=5.44
+ $X2=14.08 $Y2=5.44
r1603 818 821 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.945 $Y=5.44
+ $X2=13.57 $Y2=5.44
r1604 817 1077 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r1605 816 817 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r1606 814 1070 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.275 $Y=0
+ $X2=13.15 $Y2=0
r1607 814 816 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.275 $Y=0
+ $X2=13.57 $Y2=0
r1608 813 1076 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.945 $Y=0
+ $X2=14.08 $Y2=0
r1609 813 816 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.945 $Y=0
+ $X2=13.57 $Y2=0
r1610 812 1062 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=5.44
+ $X2=11.73 $Y2=5.44
r1611 811 812 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=5.44
+ $X2=12.19 $Y2=5.44
r1612 809 1061 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.815 $Y=5.44
+ $X2=11.68 $Y2=5.44
r1613 809 811 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=5.44
+ $X2=12.19 $Y2=5.44
r1614 808 1067 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.485 $Y=5.44
+ $X2=12.61 $Y2=5.44
r1615 808 811 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.485 $Y=5.44
+ $X2=12.19 $Y2=5.44
r1616 807 1059 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r1617 806 807 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r1618 804 1058 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.815 $Y=0
+ $X2=11.68 $Y2=0
r1619 804 806 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=0
+ $X2=12.19 $Y2=0
r1620 803 1064 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.485 $Y=0
+ $X2=12.61 $Y2=0
r1621 803 806 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.485 $Y=0
+ $X2=12.19 $Y2=0
r1622 802 1062 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=5.44
+ $X2=11.73 $Y2=5.44
r1623 801 802 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=5.44
+ $X2=11.27 $Y2=5.44
r1624 799 1061 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.545 $Y=5.44
+ $X2=11.68 $Y2=5.44
r1625 799 801 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.545 $Y=5.44
+ $X2=11.27 $Y2=5.44
r1626 798 1059 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r1627 797 798 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r1628 795 1058 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.68 $Y2=0
r1629 795 797 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.27 $Y2=0
r1630 794 802 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=5.44
+ $X2=11.27 $Y2=5.44
r1631 793 794 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.35 $Y=5.44
+ $X2=10.35 $Y2=5.44
r1632 791 794 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=5.44
+ $X2=10.35 $Y2=5.44
r1633 790 793 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.05 $Y=5.44
+ $X2=10.35 $Y2=5.44
r1634 790 791 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=5.44
+ $X2=8.05 $Y2=5.44
r1635 788 798 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r1636 787 788 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r1637 785 788 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=10.35 $Y2=0
r1638 784 787 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=10.35 $Y2=0
r1639 784 785 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r1640 782 791 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=5.44
+ $X2=8.05 $Y2=5.44
r1641 781 782 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=5.44
+ $X2=7.59 $Y2=5.44
r1642 779 785 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r1643 778 779 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r1644 776 782 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=5.44
+ $X2=7.59 $Y2=5.44
r1645 775 776 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=5.44
+ $X2=6.67 $Y2=5.44
r1646 773 779 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r1647 772 773 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r1648 770 776 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=6.67 $Y2=5.44
r1649 769 770 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=5.44
+ $X2=5.75 $Y2=5.44
r1650 767 773 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r1651 766 767 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r1652 764 770 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=5.44
+ $X2=5.75 $Y2=5.44
r1653 763 764 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r1654 761 764 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=4.83 $Y2=5.44
r1655 761 1056 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=5.44
+ $X2=2.07 $Y2=5.44
r1656 760 763 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=5.44
+ $X2=4.83 $Y2=5.44
r1657 760 761 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=5.44
+ $X2=2.53 $Y2=5.44
r1658 758 1055 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=5.44
+ $X2=2.13 $Y2=5.44
r1659 758 760 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.255 $Y=5.44
+ $X2=2.53 $Y2=5.44
r1660 757 767 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r1661 756 757 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r1662 754 757 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=4.83 $Y2=0
r1663 754 1053 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r1664 753 756 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=4.83 $Y2=0
r1665 753 754 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r1666 751 1052 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.13 $Y2=0
r1667 751 753 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.53 $Y2=0
r1668 750 1050 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=5.44
+ $X2=1.15 $Y2=5.44
r1669 749 750 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=5.44
+ $X2=0.69 $Y2=5.44
r1670 747 1043 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=5.44
+ $X2=0.197 $Y2=5.44
r1671 747 749 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=5.44
+ $X2=0.69 $Y2=5.44
r1672 746 1049 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=5.44
+ $X2=1.2 $Y2=5.44
r1673 746 749 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=5.44
+ $X2=0.69 $Y2=5.44
r1674 745 1047 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r1675 744 745 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r1676 742 1040 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r1677 742 744 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.69 $Y2=0
r1678 741 1046 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=1.2 $Y2=0
r1679 741 744 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=0.69 $Y2=0
r1680 722 1038 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.75 $Y=5.44
+ $X2=51.29 $Y2=5.44
r1681 722 1157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.75 $Y=5.44
+ $X2=51.75 $Y2=5.44
r1682 721 1033 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=51.75 $Y=0
+ $X2=51.29 $Y2=0
r1683 721 1154 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=51.75 $Y=0
+ $X2=51.75 $Y2=0
r1684 720 976 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.33 $Y=5.44
+ $X2=39.79 $Y2=5.44
r1685 720 1133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.33 $Y=5.44
+ $X2=39.33 $Y2=5.44
r1686 719 971 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=39.33 $Y=0
+ $X2=39.79 $Y2=0
r1687 719 1130 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=39.33 $Y=0
+ $X2=39.33 $Y2=0
r1688 718 720 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=5.44
+ $X2=39.33 $Y2=5.44
r1689 718 966 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=5.44
+ $X2=38.41 $Y2=5.44
r1690 718 1127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.87 $Y=5.44
+ $X2=38.87 $Y2=5.44
r1691 717 719 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=0
+ $X2=39.33 $Y2=0
r1692 717 961 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=38.87 $Y=0
+ $X2=38.41 $Y2=0
r1693 717 1124 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=38.87 $Y=0
+ $X2=38.87 $Y2=0
r1694 716 904 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.45 $Y=5.44
+ $X2=26.91 $Y2=5.44
r1695 716 1103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.45 $Y=5.44
+ $X2=26.45 $Y2=5.44
r1696 715 899 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=26.45 $Y=0
+ $X2=26.91 $Y2=0
r1697 715 1100 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=26.45 $Y=0
+ $X2=26.45 $Y2=0
r1698 714 716 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.99 $Y=5.44
+ $X2=26.45 $Y2=5.44
r1699 714 893 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.99 $Y=5.44
+ $X2=25.99 $Y2=5.44
r1700 713 715 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.99 $Y=0
+ $X2=26.45 $Y2=0
r1701 713 888 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.99 $Y=0
+ $X2=25.99 $Y2=0
r1702 712 714 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=5.44
+ $X2=25.99 $Y2=5.44
r1703 712 884 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=5.44
+ $X2=25.07 $Y2=5.44
r1704 712 1097 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=5.44
+ $X2=25.53 $Y2=5.44
r1705 711 713 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=0
+ $X2=25.99 $Y2=0
r1706 711 879 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=0
+ $X2=25.07 $Y2=0
r1707 711 1094 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=0
+ $X2=25.53 $Y2=0
r1708 710 822 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=5.44
+ $X2=13.57 $Y2=5.44
r1709 710 1073 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=5.44
+ $X2=13.11 $Y2=5.44
r1710 709 817 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r1711 709 1070 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r1712 708 710 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=13.11 $Y2=5.44
r1713 708 812 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=12.19 $Y2=5.44
r1714 708 1067 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=5.44
+ $X2=12.65 $Y2=5.44
r1715 707 709 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r1716 707 807 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r1717 707 1064 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r1718 706 750 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=5.44
+ $X2=0.69 $Y2=5.44
r1719 706 1043 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r1720 705 745 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r1721 705 1040 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r1722 703 1019 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=49.725 $Y=5.44
+ $X2=49.45 $Y2=5.44
r1723 703 704 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=49.725 $Y=5.44
+ $X2=49.85 $Y2=5.44
r1724 702 1027 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=49.975 $Y=5.44
+ $X2=50.37 $Y2=5.44
r1725 702 704 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=49.975 $Y=5.44
+ $X2=49.85 $Y2=5.44
r1726 700 1013 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=49.725 $Y=0
+ $X2=49.45 $Y2=0
r1727 700 701 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=49.725 $Y=0
+ $X2=49.85 $Y2=0
r1728 699 1023 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=49.975 $Y=0
+ $X2=50.37 $Y2=0
r1729 699 701 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=49.975 $Y=0
+ $X2=49.85 $Y2=0
r1730 697 1007 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=46.73 $Y=5.44
+ $X2=46.69 $Y2=5.44
r1731 697 698 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=46.73 $Y=5.44
+ $X2=46.875 $Y2=5.44
r1732 696 1016 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=47.02 $Y=5.44
+ $X2=47.15 $Y2=5.44
r1733 696 698 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=47.02 $Y=5.44
+ $X2=46.875 $Y2=5.44
r1734 694 1004 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=46.73 $Y=0
+ $X2=46.69 $Y2=0
r1735 694 695 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=46.73 $Y=0
+ $X2=46.875 $Y2=0
r1736 693 1010 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=47.02 $Y=0
+ $X2=47.15 $Y2=0
r1737 693 695 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=47.02 $Y=0
+ $X2=46.875 $Y2=0
r1738 691 1001 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=45.81 $Y=5.44
+ $X2=45.77 $Y2=5.44
r1739 691 692 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=45.81 $Y=5.44
+ $X2=45.955 $Y2=5.44
r1740 690 1007 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=46.1 $Y=5.44
+ $X2=46.69 $Y2=5.44
r1741 690 692 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=46.1 $Y=5.44
+ $X2=45.955 $Y2=5.44
r1742 688 998 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=45.81 $Y=0
+ $X2=45.77 $Y2=0
r1743 688 689 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=45.81 $Y=0
+ $X2=45.955 $Y2=0
r1744 687 1004 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=46.1 $Y=0
+ $X2=46.69 $Y2=0
r1745 687 689 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=46.1 $Y=0
+ $X2=45.955 $Y2=0
r1746 685 995 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=44.98 $Y=5.44
+ $X2=44.85 $Y2=5.44
r1747 685 686 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.98 $Y=5.44
+ $X2=45.125 $Y2=5.44
r1748 684 1001 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=45.27 $Y=5.44
+ $X2=45.77 $Y2=5.44
r1749 684 686 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=45.27 $Y=5.44
+ $X2=45.125 $Y2=5.44
r1750 682 992 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=44.98 $Y=0
+ $X2=44.85 $Y2=0
r1751 682 683 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.98 $Y=0
+ $X2=45.125 $Y2=0
r1752 681 998 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=45.27 $Y=0
+ $X2=45.77 $Y2=0
r1753 681 683 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=45.27 $Y=0
+ $X2=45.125 $Y2=0
r1754 679 989 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=44.06 $Y=5.44
+ $X2=43.93 $Y2=5.44
r1755 679 680 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.06 $Y=5.44
+ $X2=44.205 $Y2=5.44
r1756 678 995 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=44.35 $Y=5.44
+ $X2=44.85 $Y2=5.44
r1757 678 680 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.35 $Y=5.44
+ $X2=44.205 $Y2=5.44
r1758 676 982 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=44.06 $Y=0
+ $X2=43.93 $Y2=0
r1759 676 677 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.06 $Y=0
+ $X2=44.205 $Y2=0
r1760 675 992 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=44.35 $Y=0
+ $X2=44.85 $Y2=0
r1761 675 677 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=44.35 $Y=0
+ $X2=44.205 $Y2=0
r1762 673 947 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=36.845 $Y=5.44
+ $X2=36.57 $Y2=5.44
r1763 673 674 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=36.845 $Y=5.44
+ $X2=36.97 $Y2=5.44
r1764 672 955 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=37.095 $Y=5.44
+ $X2=37.49 $Y2=5.44
r1765 672 674 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=37.095 $Y=5.44
+ $X2=36.97 $Y2=5.44
r1766 670 941 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=36.845 $Y=0
+ $X2=36.57 $Y2=0
r1767 670 671 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=36.845 $Y=0
+ $X2=36.97 $Y2=0
r1768 669 951 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=37.095 $Y=0
+ $X2=37.49 $Y2=0
r1769 669 671 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=37.095 $Y=0
+ $X2=36.97 $Y2=0
r1770 667 935 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=33.85 $Y=5.44
+ $X2=33.81 $Y2=5.44
r1771 667 668 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=33.85 $Y=5.44
+ $X2=33.995 $Y2=5.44
r1772 666 944 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=34.14 $Y=5.44
+ $X2=34.27 $Y2=5.44
r1773 666 668 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=34.14 $Y=5.44
+ $X2=33.995 $Y2=5.44
r1774 664 932 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=33.85 $Y=0
+ $X2=33.81 $Y2=0
r1775 664 665 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=33.85 $Y=0
+ $X2=33.995 $Y2=0
r1776 663 938 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=34.14 $Y=0
+ $X2=34.27 $Y2=0
r1777 663 665 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=34.14 $Y=0
+ $X2=33.995 $Y2=0
r1778 661 929 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=32.93 $Y=5.44
+ $X2=32.89 $Y2=5.44
r1779 661 662 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.93 $Y=5.44
+ $X2=33.075 $Y2=5.44
r1780 660 935 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=33.22 $Y=5.44
+ $X2=33.81 $Y2=5.44
r1781 660 662 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=33.22 $Y=5.44
+ $X2=33.075 $Y2=5.44
r1782 658 926 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=32.93 $Y=0
+ $X2=32.89 $Y2=0
r1783 658 659 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.93 $Y=0
+ $X2=33.075 $Y2=0
r1784 657 932 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=33.22 $Y=0
+ $X2=33.81 $Y2=0
r1785 657 659 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=33.22 $Y=0
+ $X2=33.075 $Y2=0
r1786 655 923 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=32.1 $Y=5.44
+ $X2=31.97 $Y2=5.44
r1787 655 656 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.1 $Y=5.44
+ $X2=32.245 $Y2=5.44
r1788 654 929 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=32.39 $Y=5.44
+ $X2=32.89 $Y2=5.44
r1789 654 656 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.39 $Y=5.44
+ $X2=32.245 $Y2=5.44
r1790 652 920 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=32.1 $Y=0
+ $X2=31.97 $Y2=0
r1791 652 653 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.1 $Y=0
+ $X2=32.245 $Y2=0
r1792 651 926 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=32.39 $Y=0
+ $X2=32.89 $Y2=0
r1793 651 653 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=32.39 $Y=0
+ $X2=32.245 $Y2=0
r1794 649 917 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=31.18 $Y=5.44
+ $X2=31.05 $Y2=5.44
r1795 649 650 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=31.18 $Y=5.44
+ $X2=31.325 $Y2=5.44
r1796 648 923 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=31.47 $Y=5.44
+ $X2=31.97 $Y2=5.44
r1797 648 650 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=31.47 $Y=5.44
+ $X2=31.325 $Y2=5.44
r1798 646 910 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=31.18 $Y=0
+ $X2=31.05 $Y2=0
r1799 646 647 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=31.18 $Y=0
+ $X2=31.325 $Y2=0
r1800 645 920 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=31.47 $Y=0
+ $X2=31.97 $Y2=0
r1801 645 647 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=31.47 $Y=0
+ $X2=31.325 $Y2=0
r1802 643 865 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=23.505 $Y=5.44
+ $X2=23.23 $Y2=5.44
r1803 643 644 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.505 $Y=5.44
+ $X2=23.63 $Y2=5.44
r1804 642 873 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=23.755 $Y=5.44
+ $X2=24.15 $Y2=5.44
r1805 642 644 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.755 $Y=5.44
+ $X2=23.63 $Y2=5.44
r1806 640 859 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=23.505 $Y=0
+ $X2=23.23 $Y2=0
r1807 640 641 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.505 $Y=0
+ $X2=23.63 $Y2=0
r1808 639 869 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=23.755 $Y=0
+ $X2=24.15 $Y2=0
r1809 639 641 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.755 $Y=0
+ $X2=23.63 $Y2=0
r1810 637 853 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=20.51 $Y=5.44
+ $X2=20.47 $Y2=5.44
r1811 637 638 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.51 $Y=5.44
+ $X2=20.655 $Y2=5.44
r1812 636 862 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=20.8 $Y=5.44
+ $X2=20.93 $Y2=5.44
r1813 636 638 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.8 $Y=5.44
+ $X2=20.655 $Y2=5.44
r1814 634 850 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=20.51 $Y=0
+ $X2=20.47 $Y2=0
r1815 634 635 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.51 $Y=0
+ $X2=20.655 $Y2=0
r1816 633 856 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=20.8 $Y=0
+ $X2=20.93 $Y2=0
r1817 633 635 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.8 $Y=0
+ $X2=20.655 $Y2=0
r1818 631 847 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=19.59 $Y=5.44
+ $X2=19.55 $Y2=5.44
r1819 631 632 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.59 $Y=5.44
+ $X2=19.735 $Y2=5.44
r1820 630 853 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=19.88 $Y=5.44
+ $X2=20.47 $Y2=5.44
r1821 630 632 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.88 $Y=5.44
+ $X2=19.735 $Y2=5.44
r1822 628 844 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=19.59 $Y=0
+ $X2=19.55 $Y2=0
r1823 628 629 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.59 $Y=0
+ $X2=19.735 $Y2=0
r1824 627 850 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=19.88 $Y=0
+ $X2=20.47 $Y2=0
r1825 627 629 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.88 $Y=0
+ $X2=19.735 $Y2=0
r1826 625 841 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=18.76 $Y=5.44
+ $X2=18.63 $Y2=5.44
r1827 625 626 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.76 $Y=5.44
+ $X2=18.905 $Y2=5.44
r1828 624 847 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=19.05 $Y=5.44
+ $X2=19.55 $Y2=5.44
r1829 624 626 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.05 $Y=5.44
+ $X2=18.905 $Y2=5.44
r1830 622 838 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=18.76 $Y=0
+ $X2=18.63 $Y2=0
r1831 622 623 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.76 $Y=0
+ $X2=18.905 $Y2=0
r1832 621 844 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=19.05 $Y=0
+ $X2=19.55 $Y2=0
r1833 621 623 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.05 $Y=0
+ $X2=18.905 $Y2=0
r1834 619 835 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=17.84 $Y=5.44
+ $X2=17.71 $Y2=5.44
r1835 619 620 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=17.84 $Y=5.44
+ $X2=17.985 $Y2=5.44
r1836 618 841 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=18.13 $Y=5.44
+ $X2=18.63 $Y2=5.44
r1837 618 620 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.13 $Y=5.44
+ $X2=17.985 $Y2=5.44
r1838 616 828 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=17.84 $Y=0
+ $X2=17.71 $Y2=0
r1839 616 617 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=17.84 $Y=0
+ $X2=17.985 $Y2=0
r1840 615 838 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=18.13 $Y=0
+ $X2=18.63 $Y2=0
r1841 615 617 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.13 $Y=0
+ $X2=17.985 $Y2=0
r1842 613 793 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.625 $Y=5.44
+ $X2=10.35 $Y2=5.44
r1843 613 614 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.625 $Y=5.44
+ $X2=10.75 $Y2=5.44
r1844 612 801 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.875 $Y=5.44
+ $X2=11.27 $Y2=5.44
r1845 612 614 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.875 $Y=5.44
+ $X2=10.75 $Y2=5.44
r1846 610 787 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.35 $Y2=0
r1847 610 611 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.75 $Y2=0
r1848 609 797 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.875 $Y=0
+ $X2=11.27 $Y2=0
r1849 609 611 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.875 $Y=0
+ $X2=10.75 $Y2=0
r1850 607 781 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=7.63 $Y=5.44
+ $X2=7.59 $Y2=5.44
r1851 607 608 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.63 $Y=5.44
+ $X2=7.775 $Y2=5.44
r1852 606 790 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=5.44
+ $X2=8.05 $Y2=5.44
r1853 606 608 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.92 $Y=5.44
+ $X2=7.775 $Y2=5.44
r1854 604 778 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=7.63 $Y=0 $X2=7.59
+ $Y2=0
r1855 604 605 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.63 $Y=0
+ $X2=7.775 $Y2=0
r1856 603 784 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=8.05 $Y2=0
r1857 603 605 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=7.775 $Y2=0
r1858 601 775 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.71 $Y=5.44
+ $X2=6.67 $Y2=5.44
r1859 601 602 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.71 $Y=5.44
+ $X2=6.855 $Y2=5.44
r1860 600 781 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7 $Y=5.44
+ $X2=7.59 $Y2=5.44
r1861 600 602 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7 $Y=5.44
+ $X2=6.855 $Y2=5.44
r1862 598 772 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.67
+ $Y2=0
r1863 598 599 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.71 $Y=0
+ $X2=6.855 $Y2=0
r1864 597 778 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7 $Y=0 $X2=7.59
+ $Y2=0
r1865 597 599 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.855
+ $Y2=0
r1866 595 769 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=5.44
+ $X2=5.75 $Y2=5.44
r1867 595 596 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.88 $Y=5.44
+ $X2=6.025 $Y2=5.44
r1868 594 775 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.17 $Y=5.44
+ $X2=6.67 $Y2=5.44
r1869 594 596 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.17 $Y=5.44
+ $X2=6.025 $Y2=5.44
r1870 592 766 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=0
+ $X2=5.75 $Y2=0
r1871 592 593 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.88 $Y=0
+ $X2=6.025 $Y2=0
r1872 591 772 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.67
+ $Y2=0
r1873 591 593 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=6.025 $Y2=0
r1874 589 763 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.96 $Y=5.44
+ $X2=4.83 $Y2=5.44
r1875 589 590 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.96 $Y=5.44
+ $X2=5.105 $Y2=5.44
r1876 588 769 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.25 $Y=5.44
+ $X2=5.75 $Y2=5.44
r1877 588 590 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.25 $Y=5.44
+ $X2=5.105 $Y2=5.44
r1878 586 756 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=4.83 $Y2=0
r1879 586 587 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=5.105 $Y2=0
r1880 585 766 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.75
+ $Y2=0
r1881 585 587 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.25 $Y=0
+ $X2=5.105 $Y2=0
r1882 581 1157 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=51.71
+ $Y=5.355 $X2=51.782 $Y2=5.44
r1883 581 583 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=51.71 $Y=5.355
+ $X2=51.71 $Y2=4.72
r1884 577 1154 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=51.71
+ $Y=0.085 $X2=51.782 $Y2=0
r1885 577 579 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=51.71 $Y=0.085
+ $X2=51.71 $Y2=0.38
r1886 573 1151 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=50.78 $Y=5.355
+ $X2=50.78 $Y2=5.44
r1887 573 575 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=50.78 $Y=5.355
+ $X2=50.78 $Y2=5.06
r1888 569 1148 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=50.78 $Y=0.085
+ $X2=50.78 $Y2=0
r1889 569 571 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=50.78 $Y=0.085
+ $X2=50.78 $Y2=0.38
r1890 565 704 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=49.85 $Y=5.355
+ $X2=49.85 $Y2=5.44
r1891 565 567 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=49.85 $Y=5.355
+ $X2=49.85 $Y2=5.06
r1892 561 701 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=49.85 $Y=0.085
+ $X2=49.85 $Y2=0
r1893 561 563 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=49.85 $Y=0.085
+ $X2=49.85 $Y2=0.38
r1894 557 698 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=46.875 $Y=5.355
+ $X2=46.875 $Y2=5.44
r1895 557 559 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=46.875 $Y=5.355
+ $X2=46.875 $Y2=4.995
r1896 553 695 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=46.875 $Y=0.085
+ $X2=46.875 $Y2=0
r1897 553 555 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=46.875 $Y=0.085
+ $X2=46.875 $Y2=0.445
r1898 549 692 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=45.955 $Y=5.355
+ $X2=45.955 $Y2=5.44
r1899 549 551 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=45.955 $Y=5.355
+ $X2=45.955 $Y2=4.995
r1900 545 689 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=45.955 $Y=0.085
+ $X2=45.955 $Y2=0
r1901 545 547 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=45.955 $Y=0.085
+ $X2=45.955 $Y2=0.445
r1902 541 686 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=45.125 $Y=5.355
+ $X2=45.125 $Y2=5.44
r1903 541 543 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=45.125 $Y=5.355
+ $X2=45.125 $Y2=4.995
r1904 537 683 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=45.125 $Y=0.085
+ $X2=45.125 $Y2=0
r1905 537 539 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=45.125 $Y=0.085
+ $X2=45.125 $Y2=0.445
r1906 533 680 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=44.205 $Y=5.355
+ $X2=44.205 $Y2=5.44
r1907 533 535 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=44.205 $Y=5.355
+ $X2=44.205 $Y2=4.995
r1908 529 677 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=44.205 $Y=0.085
+ $X2=44.205 $Y2=0
r1909 529 531 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=44.205 $Y=0.085
+ $X2=44.205 $Y2=0.445
r1910 525 1145 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=41.23
+ $Y=5.355 $X2=41.23 $Y2=5.44
r1911 525 527 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=41.23 $Y=5.355
+ $X2=41.23 $Y2=5.06
r1912 521 1142 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=41.23
+ $Y=0.085 $X2=41.23 $Y2=0
r1913 521 523 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=41.23 $Y=0.085
+ $X2=41.23 $Y2=0.38
r1914 520 1139 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.435 $Y=5.44
+ $X2=40.3 $Y2=5.44
r1915 519 1145 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=41.105 $Y=5.44
+ $X2=41.23 $Y2=5.44
r1916 519 520 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=41.105 $Y=5.44
+ $X2=40.435 $Y2=5.44
r1917 518 1136 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=40.435 $Y=0
+ $X2=40.3 $Y2=0
r1918 517 1142 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=41.105 $Y=0
+ $X2=41.23 $Y2=0
r1919 517 518 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=41.105 $Y=0
+ $X2=40.435 $Y2=0
r1920 513 1139 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=40.3 $Y=5.355
+ $X2=40.3 $Y2=5.44
r1921 513 515 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=40.3 $Y=5.355
+ $X2=40.3 $Y2=5.06
r1922 509 1136 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=40.3 $Y=0.085
+ $X2=40.3 $Y2=0
r1923 509 511 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=40.3 $Y=0.085
+ $X2=40.3 $Y2=0.38
r1924 505 1133 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=39.37
+ $Y=5.355 $X2=39.37 $Y2=5.44
r1925 505 507 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=39.37 $Y=5.355
+ $X2=39.37 $Y2=4.72
r1926 501 1130 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=39.37
+ $Y=0.085 $X2=39.37 $Y2=0
r1927 501 503 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=39.37 $Y=0.085
+ $X2=39.37 $Y2=0.38
r1928 500 1127 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=38.955 $Y=5.44
+ $X2=38.83 $Y2=5.44
r1929 499 1133 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=39.245 $Y=5.44
+ $X2=39.37 $Y2=5.44
r1930 499 500 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=39.245 $Y=5.44
+ $X2=38.955 $Y2=5.44
r1931 498 1124 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=38.955 $Y=0
+ $X2=38.83 $Y2=0
r1932 497 1130 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=39.245 $Y=0
+ $X2=39.37 $Y2=0
r1933 497 498 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=39.245 $Y=0
+ $X2=38.955 $Y2=0
r1934 493 1127 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=38.83
+ $Y=5.355 $X2=38.83 $Y2=5.44
r1935 493 495 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=38.83 $Y=5.355
+ $X2=38.83 $Y2=4.72
r1936 489 1124 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=38.83
+ $Y=0.085 $X2=38.83 $Y2=0
r1937 489 491 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=38.83 $Y=0.085
+ $X2=38.83 $Y2=0.38
r1938 485 1121 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=37.9 $Y=5.355
+ $X2=37.9 $Y2=5.44
r1939 485 487 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=37.9 $Y=5.355
+ $X2=37.9 $Y2=5.06
r1940 481 1118 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=37.9 $Y=0.085
+ $X2=37.9 $Y2=0
r1941 481 483 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=37.9 $Y=0.085
+ $X2=37.9 $Y2=0.38
r1942 477 674 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=36.97 $Y=5.355
+ $X2=36.97 $Y2=5.44
r1943 477 479 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=36.97 $Y=5.355
+ $X2=36.97 $Y2=5.06
r1944 473 671 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=36.97 $Y=0.085
+ $X2=36.97 $Y2=0
r1945 473 475 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=36.97 $Y=0.085
+ $X2=36.97 $Y2=0.38
r1946 469 668 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=33.995 $Y=5.355
+ $X2=33.995 $Y2=5.44
r1947 469 471 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=33.995 $Y=5.355
+ $X2=33.995 $Y2=4.995
r1948 465 665 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=33.995 $Y=0.085
+ $X2=33.995 $Y2=0
r1949 465 467 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=33.995 $Y=0.085
+ $X2=33.995 $Y2=0.445
r1950 461 662 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=33.075 $Y=5.355
+ $X2=33.075 $Y2=5.44
r1951 461 463 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=33.075 $Y=5.355
+ $X2=33.075 $Y2=4.995
r1952 457 659 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=33.075 $Y=0.085
+ $X2=33.075 $Y2=0
r1953 457 459 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=33.075 $Y=0.085
+ $X2=33.075 $Y2=0.445
r1954 453 656 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=32.245 $Y=5.355
+ $X2=32.245 $Y2=5.44
r1955 453 455 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=32.245 $Y=5.355
+ $X2=32.245 $Y2=4.995
r1956 449 653 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=32.245 $Y=0.085
+ $X2=32.245 $Y2=0
r1957 449 451 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=32.245 $Y=0.085
+ $X2=32.245 $Y2=0.445
r1958 445 650 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=31.325 $Y=5.355
+ $X2=31.325 $Y2=5.44
r1959 445 447 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=31.325 $Y=5.355
+ $X2=31.325 $Y2=4.995
r1960 441 647 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=31.325 $Y=0.085
+ $X2=31.325 $Y2=0
r1961 441 443 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=31.325 $Y=0.085
+ $X2=31.325 $Y2=0.445
r1962 437 1115 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=28.35
+ $Y=5.355 $X2=28.35 $Y2=5.44
r1963 437 439 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=28.35 $Y=5.355
+ $X2=28.35 $Y2=5.06
r1964 433 1112 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=28.35
+ $Y=0.085 $X2=28.35 $Y2=0
r1965 433 435 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=28.35 $Y=0.085
+ $X2=28.35 $Y2=0.38
r1966 432 1109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.555 $Y=5.44
+ $X2=27.42 $Y2=5.44
r1967 431 1115 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=28.225 $Y=5.44
+ $X2=28.35 $Y2=5.44
r1968 431 432 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=28.225 $Y=5.44
+ $X2=27.555 $Y2=5.44
r1969 430 1106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=27.555 $Y=0
+ $X2=27.42 $Y2=0
r1970 429 1112 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=28.225 $Y=0
+ $X2=28.35 $Y2=0
r1971 429 430 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=28.225 $Y=0
+ $X2=27.555 $Y2=0
r1972 425 1109 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=27.42 $Y=5.355
+ $X2=27.42 $Y2=5.44
r1973 425 427 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=27.42 $Y=5.355
+ $X2=27.42 $Y2=5.06
r1974 421 1106 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=27.42 $Y=0.085
+ $X2=27.42 $Y2=0
r1975 421 423 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=27.42 $Y=0.085
+ $X2=27.42 $Y2=0.38
r1976 417 1103 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=26.49
+ $Y=5.355 $X2=26.49 $Y2=5.44
r1977 417 419 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=26.49 $Y=5.355
+ $X2=26.49 $Y2=4.72
r1978 413 1100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=26.49
+ $Y=0.085 $X2=26.49 $Y2=0
r1979 413 415 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=26.49 $Y=0.085
+ $X2=26.49 $Y2=0.38
r1980 409 1097 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=25.49
+ $Y=5.355 $X2=25.49 $Y2=5.44
r1981 409 411 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=25.49 $Y=5.355
+ $X2=25.49 $Y2=4.72
r1982 405 1094 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=25.49
+ $Y=0.085 $X2=25.49 $Y2=0
r1983 405 407 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=25.49 $Y=0.085
+ $X2=25.49 $Y2=0.38
r1984 401 1091 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=5.355
+ $X2=24.56 $Y2=5.44
r1985 401 403 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=24.56 $Y=5.355
+ $X2=24.56 $Y2=5.06
r1986 397 1088 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=0.085
+ $X2=24.56 $Y2=0
r1987 397 399 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=24.56 $Y=0.085
+ $X2=24.56 $Y2=0.38
r1988 393 644 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=23.63 $Y=5.355
+ $X2=23.63 $Y2=5.44
r1989 393 395 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=23.63 $Y=5.355
+ $X2=23.63 $Y2=5.06
r1990 389 641 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=23.63 $Y=0.085
+ $X2=23.63 $Y2=0
r1991 389 391 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=23.63 $Y=0.085
+ $X2=23.63 $Y2=0.38
r1992 385 638 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=20.655 $Y=5.355
+ $X2=20.655 $Y2=5.44
r1993 385 387 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=20.655 $Y=5.355
+ $X2=20.655 $Y2=4.995
r1994 381 635 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=20.655 $Y=0.085
+ $X2=20.655 $Y2=0
r1995 381 383 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=20.655 $Y=0.085
+ $X2=20.655 $Y2=0.445
r1996 377 632 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=19.735 $Y=5.355
+ $X2=19.735 $Y2=5.44
r1997 377 379 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=19.735 $Y=5.355
+ $X2=19.735 $Y2=4.995
r1998 373 629 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=19.735 $Y=0.085
+ $X2=19.735 $Y2=0
r1999 373 375 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=19.735 $Y=0.085
+ $X2=19.735 $Y2=0.445
r2000 369 626 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=18.905 $Y=5.355
+ $X2=18.905 $Y2=5.44
r2001 369 371 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=18.905 $Y=5.355
+ $X2=18.905 $Y2=4.995
r2002 365 623 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=18.905 $Y=0.085
+ $X2=18.905 $Y2=0
r2003 365 367 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=18.905 $Y=0.085
+ $X2=18.905 $Y2=0.445
r2004 361 620 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=17.985 $Y=5.355
+ $X2=17.985 $Y2=5.44
r2005 361 363 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=17.985 $Y=5.355
+ $X2=17.985 $Y2=4.995
r2006 357 617 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=17.985 $Y=0.085
+ $X2=17.985 $Y2=0
r2007 357 359 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=17.985 $Y=0.085
+ $X2=17.985 $Y2=0.445
r2008 353 1085 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.01
+ $Y=5.355 $X2=15.01 $Y2=5.44
r2009 353 355 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=15.01 $Y=5.355
+ $X2=15.01 $Y2=5.06
r2010 349 1082 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.01
+ $Y=0.085 $X2=15.01 $Y2=0
r2011 349 351 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=15.01 $Y=0.085
+ $X2=15.01 $Y2=0.38
r2012 348 1079 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.215 $Y=5.44
+ $X2=14.08 $Y2=5.44
r2013 347 1085 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.885 $Y=5.44
+ $X2=15.01 $Y2=5.44
r2014 347 348 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=5.44
+ $X2=14.215 $Y2=5.44
r2015 346 1076 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.215 $Y=0
+ $X2=14.08 $Y2=0
r2016 345 1082 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=15.01 $Y2=0
r2017 345 346 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.215 $Y2=0
r2018 341 1079 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=5.355
+ $X2=14.08 $Y2=5.44
r2019 341 343 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.08 $Y=5.355
+ $X2=14.08 $Y2=5.06
r2020 337 1076 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=0.085
+ $X2=14.08 $Y2=0
r2021 337 339 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.08 $Y=0.085
+ $X2=14.08 $Y2=0.38
r2022 333 1073 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.15
+ $Y=5.355 $X2=13.15 $Y2=5.44
r2023 333 335 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=13.15 $Y=5.355
+ $X2=13.15 $Y2=4.72
r2024 329 1070 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.15
+ $Y=0.085 $X2=13.15 $Y2=0
r2025 329 331 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.15 $Y=0.085
+ $X2=13.15 $Y2=0.38
r2026 328 1067 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.735 $Y=5.44
+ $X2=12.61 $Y2=5.44
r2027 327 1073 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.025 $Y=5.44
+ $X2=13.15 $Y2=5.44
r2028 327 328 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.025 $Y=5.44
+ $X2=12.735 $Y2=5.44
r2029 326 1064 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.735 $Y=0
+ $X2=12.61 $Y2=0
r2030 325 1070 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.025 $Y=0
+ $X2=13.15 $Y2=0
r2031 325 326 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.025 $Y=0
+ $X2=12.735 $Y2=0
r2032 321 1067 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.61
+ $Y=5.355 $X2=12.61 $Y2=5.44
r2033 321 323 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=12.61 $Y=5.355
+ $X2=12.61 $Y2=4.72
r2034 317 1064 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.61
+ $Y=0.085 $X2=12.61 $Y2=0
r2035 317 319 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.61 $Y=0.085
+ $X2=12.61 $Y2=0.38
r2036 313 1061 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=5.355
+ $X2=11.68 $Y2=5.44
r2037 313 315 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.68 $Y=5.355
+ $X2=11.68 $Y2=5.06
r2038 309 1058 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0
r2039 309 311 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0.38
r2040 305 614 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=5.355
+ $X2=10.75 $Y2=5.44
r2041 305 307 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.75 $Y=5.355
+ $X2=10.75 $Y2=5.06
r2042 301 611 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0
r2043 301 303 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0.38
r2044 297 608 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.775 $Y=5.355
+ $X2=7.775 $Y2=5.44
r2045 297 299 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.775 $Y=5.355
+ $X2=7.775 $Y2=4.995
r2046 293 605 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.775 $Y2=0
r2047 293 295 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.775 $Y2=0.445
r2048 289 602 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=5.355
+ $X2=6.855 $Y2=5.44
r2049 289 291 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.855 $Y=5.355
+ $X2=6.855 $Y2=4.995
r2050 285 599 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=0.085
+ $X2=6.855 $Y2=0
r2051 285 287 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.855 $Y=0.085
+ $X2=6.855 $Y2=0.445
r2052 281 596 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=5.355
+ $X2=6.025 $Y2=5.44
r2053 281 283 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.025 $Y=5.355
+ $X2=6.025 $Y2=4.995
r2054 277 593 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=0.085
+ $X2=6.025 $Y2=0
r2055 277 279 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.025 $Y=0.085
+ $X2=6.025 $Y2=0.445
r2056 273 590 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=5.355
+ $X2=5.105 $Y2=5.44
r2057 273 275 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.105 $Y=5.355
+ $X2=5.105 $Y2=4.995
r2058 269 587 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0
r2059 269 271 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0.445
r2060 265 1055 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=5.355
+ $X2=2.13 $Y2=5.44
r2061 265 267 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.13 $Y=5.355
+ $X2=2.13 $Y2=5.06
r2062 261 1052 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0
r2063 261 263 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0.38
r2064 260 1049 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=5.44
+ $X2=1.2 $Y2=5.44
r2065 259 1055 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.005 $Y=5.44
+ $X2=2.13 $Y2=5.44
r2066 259 260 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=5.44
+ $X2=1.335 $Y2=5.44
r2067 258 1046 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0
+ $X2=1.2 $Y2=0
r2068 257 1052 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.13 $Y2=0
r2069 257 258 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.335 $Y2=0
r2070 253 1049 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=5.355
+ $X2=1.2 $Y2=5.44
r2071 253 255 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=5.355
+ $X2=1.2 $Y2=5.06
r2072 249 1046 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r2073 249 251 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.38
r2074 245 1043 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27
+ $Y=5.355 $X2=0.197 $Y2=5.44
r2075 245 247 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.27 $Y=5.355
+ $X2=0.27 $Y2=4.72
r2076 241 1040 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27
+ $Y=0.085 $X2=0.197 $Y2=0
r2077 241 243 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r2078 80 583 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=51.535
+ $Y=4.555 $X2=51.67 $Y2=4.72
r2079 79 579 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=51.535
+ $Y=0.235 $X2=51.67 $Y2=0.38
r2080 78 575 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=50.595 $Y=4.555 $X2=50.78 $Y2=5.06
r2081 77 571 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=50.595 $Y=0.235 $X2=50.78 $Y2=0.38
r2082 76 567 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1
+ $X=49.765 $Y=4.555 $X2=49.89 $Y2=5.06
r2083 75 563 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=49.765 $Y=0.235 $X2=49.89 $Y2=0.38
r2084 74 559 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=46.68
+ $Y=4.785 $X2=46.815 $Y2=4.995
r2085 73 555 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=46.68
+ $Y=0.235 $X2=46.815 $Y2=0.445
r2086 72 551 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=45.85
+ $Y=4.785 $X2=45.975 $Y2=4.995
r2087 71 547 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=45.85
+ $Y=0.235 $X2=45.975 $Y2=0.445
r2088 70 543 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=44.97
+ $Y=4.785 $X2=45.105 $Y2=4.995
r2089 69 539 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=44.97
+ $Y=0.235 $X2=45.105 $Y2=0.445
r2090 68 535 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=44.14
+ $Y=4.785 $X2=44.265 $Y2=4.995
r2091 67 531 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=44.14
+ $Y=0.235 $X2=44.265 $Y2=0.445
r2092 66 527 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1
+ $X=41.055 $Y=4.555 $X2=41.19 $Y2=5.06
r2093 65 523 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1
+ $X=41.055 $Y=0.235 $X2=41.19 $Y2=0.38
r2094 64 515 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=40.115 $Y=4.555 $X2=40.3 $Y2=5.06
r2095 63 511 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=40.115 $Y=0.235 $X2=40.3 $Y2=0.38
r2096 62 507 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=39.235
+ $Y=4.555 $X2=39.41 $Y2=4.72
r2097 61 503 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=39.235
+ $Y=0.235 $X2=39.41 $Y2=0.38
r2098 60 495 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=38.655
+ $Y=4.555 $X2=38.79 $Y2=4.72
r2099 59 491 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=38.655
+ $Y=0.235 $X2=38.79 $Y2=0.38
r2100 58 487 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=37.715 $Y=4.555 $X2=37.9 $Y2=5.06
r2101 57 483 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=37.715 $Y=0.235 $X2=37.9 $Y2=0.38
r2102 56 479 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1
+ $X=36.885 $Y=4.555 $X2=37.01 $Y2=5.06
r2103 55 475 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=36.885 $Y=0.235 $X2=37.01 $Y2=0.38
r2104 54 471 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=33.8
+ $Y=4.785 $X2=33.935 $Y2=4.995
r2105 53 467 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=33.8
+ $Y=0.235 $X2=33.935 $Y2=0.445
r2106 52 463 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=32.97
+ $Y=4.785 $X2=33.095 $Y2=4.995
r2107 51 459 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=32.97
+ $Y=0.235 $X2=33.095 $Y2=0.445
r2108 50 455 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=32.09
+ $Y=4.785 $X2=32.225 $Y2=4.995
r2109 49 451 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=32.09
+ $Y=0.235 $X2=32.225 $Y2=0.445
r2110 48 447 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=31.26
+ $Y=4.785 $X2=31.385 $Y2=4.995
r2111 47 443 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=31.26
+ $Y=0.235 $X2=31.385 $Y2=0.445
r2112 46 439 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1
+ $X=28.175 $Y=4.555 $X2=28.31 $Y2=5.06
r2113 45 435 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1
+ $X=28.175 $Y=0.235 $X2=28.31 $Y2=0.38
r2114 44 427 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=27.235 $Y=4.555 $X2=27.42 $Y2=5.06
r2115 43 423 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=27.235 $Y=0.235 $X2=27.42 $Y2=0.38
r2116 42 419 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=26.355
+ $Y=4.555 $X2=26.53 $Y2=4.72
r2117 41 415 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=26.355
+ $Y=0.235 $X2=26.53 $Y2=0.38
r2118 40 411 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=4.555 $X2=25.45 $Y2=4.72
r2119 39 407 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=0.235 $X2=25.45 $Y2=0.38
r2120 38 403 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=24.375 $Y=4.555 $X2=24.56 $Y2=5.06
r2121 37 399 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=24.375 $Y=0.235 $X2=24.56 $Y2=0.38
r2122 36 395 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1
+ $X=23.545 $Y=4.555 $X2=23.67 $Y2=5.06
r2123 35 391 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=23.545 $Y=0.235 $X2=23.67 $Y2=0.38
r2124 34 387 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.46
+ $Y=4.785 $X2=20.595 $Y2=4.995
r2125 33 383 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.46
+ $Y=0.235 $X2=20.595 $Y2=0.445
r2126 32 379 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=19.63
+ $Y=4.785 $X2=19.755 $Y2=4.995
r2127 31 375 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=19.63
+ $Y=0.235 $X2=19.755 $Y2=0.445
r2128 30 371 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.75
+ $Y=4.785 $X2=18.885 $Y2=4.995
r2129 29 367 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.75
+ $Y=0.235 $X2=18.885 $Y2=0.445
r2130 28 363 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=17.92
+ $Y=4.785 $X2=18.045 $Y2=4.995
r2131 27 359 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=17.92
+ $Y=0.235 $X2=18.045 $Y2=0.445
r2132 26 355 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1
+ $X=14.835 $Y=4.555 $X2=14.97 $Y2=5.06
r2133 25 351 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1
+ $X=14.835 $Y=0.235 $X2=14.97 $Y2=0.38
r2134 24 343 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=13.895 $Y=4.555 $X2=14.08 $Y2=5.06
r2135 23 339 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=13.895 $Y=0.235 $X2=14.08 $Y2=0.38
r2136 22 335 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=4.555 $X2=13.19 $Y2=4.72
r2137 21 331 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=0.235 $X2=13.19 $Y2=0.38
r2138 20 323 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=4.555 $X2=12.57 $Y2=4.72
r2139 19 319 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=0.235 $X2=12.57 $Y2=0.38
r2140 18 315 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1
+ $X=11.495 $Y=4.555 $X2=11.68 $Y2=5.06
r2141 17 311 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1
+ $X=11.495 $Y=0.235 $X2=11.68 $Y2=0.38
r2142 16 307 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1
+ $X=10.665 $Y=4.555 $X2=10.79 $Y2=5.06
r2143 15 303 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=10.665 $Y=0.235 $X2=10.79 $Y2=0.38
r2144 14 299 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.58
+ $Y=4.785 $X2=7.715 $Y2=4.995
r2145 13 295 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.58
+ $Y=0.235 $X2=7.715 $Y2=0.445
r2146 12 291 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=4.785 $X2=6.875 $Y2=4.995
r2147 11 287 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=0.235 $X2=6.875 $Y2=0.445
r2148 10 283 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=4.785 $X2=6.005 $Y2=4.995
r2149 9 279 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.005 $Y2=0.445
r2150 8 275 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=4.785 $X2=5.165 $Y2=4.995
r2151 7 271 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.165 $Y2=0.445
r2152 6 267 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=4.555 $X2=2.09 $Y2=5.06
r2153 5 263 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.09 $Y2=0.38
r2154 4 255 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=4.555 $X2=1.2 $Y2=5.06
r2155 3 251 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r2156 2 247 91 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=4.555 $X2=0.31 $Y2=4.72
r2157 1 243 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=4.29 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0.425
+ $X2=4.33 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=3.45 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.205 $Y=0.34
+ $X2=4.33 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=0.34
+ $X2=3.535 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=3.45 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=2.695 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=0.715
+ $X2=2.56 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.695 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0.8
+ $X2=1.67 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=2.56 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=1.835 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.8
+ $X2=1.67 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=0.8
+ $X2=0.895 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.895 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.73 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.33 $X2=4.29 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.315
+ $Y=0.33 $X2=3.45 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.33 $X2=2.61 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_911# 1 2 3 4 5 18 22 27 28 29 32
+ 34 38 41 43 44
c79 38 0 1.10627e-19 $X=4.29 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=5.015
+ $X2=4.33 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=5.1 $X2=3.45
+ $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.205 $Y=5.1
+ $X2=4.33 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=5.1
+ $X2=3.535 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=5.015
+ $X2=3.45 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=5.015
+ $X2=3.45 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=5.1 $X2=3.45
+ $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=5.1
+ $X2=2.695 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.56 $Y=5.015
+ $X2=2.695 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=5.015
+ $X2=2.56 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=4.725
+ $X2=2.56 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=4.64
+ $X2=1.67 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.425 $Y=4.64
+ $X2=2.56 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.425 $Y=4.64
+ $X2=1.835 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=4.64
+ $X2=0.73 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=4.64
+ $X2=1.67 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=4.64
+ $X2=0.895 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=4.59 $X2=4.29 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.315
+ $Y=4.59 $X2=3.45 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=4.59 $X2=2.61 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=4.555 $X2=1.67 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=4.555 $X2=0.73 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.15 $Y=0.715
+ $X2=12.15 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=0.8
+ $X2=11.21 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.985 $Y=0.8
+ $X2=12.15 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=0.8
+ $X2=11.375 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=0.715
+ $X2=11.21 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.21 $Y=0.715
+ $X2=11.21 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=0.8
+ $X2=11.21 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.045 $Y=0.8
+ $X2=10.455 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.32 $Y=0.715
+ $X2=10.455 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.32 $Y=0.715
+ $X2=10.32 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.32 $Y=0.425
+ $X2=10.32 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=0.34
+ $X2=9.43 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=10.32 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=9.515 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=9.43 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=8.675 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.55 $Y=0.425
+ $X2=8.675 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=0.425
+ $X2=8.55 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.015
+ $Y=0.235 $X2=12.15 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=11.075
+ $Y=0.235 $X2=11.21 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=0.33 $X2=10.27 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.33 $X2=9.43 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.33 $X2=8.59 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_918# 1 2 3 4 5 18 20 21 24 26
+ 31 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=4.64
+ $X2=11.21 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=4.64
+ $X2=12.15 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=4.64
+ $X2=11.375 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=4.64
+ $X2=11.21 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.045 $Y=4.64
+ $X2=10.455 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.32 $Y=5.015
+ $X2=10.32 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.32 $Y=4.725
+ $X2=10.455 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.32 $Y=4.725
+ $X2=10.32 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=5.1 $X2=9.43
+ $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.185 $Y=5.1
+ $X2=10.32 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.185 $Y=5.1
+ $X2=9.515 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=5.015
+ $X2=9.43 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.43 $Y=5.015
+ $X2=9.43 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=5.1 $X2=9.43
+ $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.345 $Y=5.1
+ $X2=8.675 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.55 $Y=5.015
+ $X2=8.675 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=5.015
+ $X2=8.55 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=12.015
+ $Y=4.555 $X2=12.15 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=11.075
+ $Y=4.555 $X2=11.21 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=4.59 $X2=10.27 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=4.59 $X2=9.43 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=4.59 $X2=8.59 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=17.17 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=17.21 $Y=0.425
+ $X2=17.21 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.415 $Y=0.34
+ $X2=16.33 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.085 $Y=0.34
+ $X2=17.21 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.085 $Y=0.34
+ $X2=16.415 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.33 $Y=0.425
+ $X2=16.33 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.33 $Y=0.425
+ $X2=16.33 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.245 $Y=0.34
+ $X2=16.33 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.245 $Y=0.34
+ $X2=15.575 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=15.44 $Y=0.715
+ $X2=15.44 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.44 $Y=0.425
+ $X2=15.575 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.44 $Y=0.425
+ $X2=15.44 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=0.8
+ $X2=14.55 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.305 $Y=0.8
+ $X2=15.44 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.305 $Y=0.8
+ $X2=14.715 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.55 $Y=0.715
+ $X2=14.55 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.55 $Y=0.715
+ $X2=14.55 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=0.8
+ $X2=14.55 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=0.8
+ $X2=13.775 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.61 $Y=0.715
+ $X2=13.775 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.61 $Y=0.715
+ $X2=13.61 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=17.035
+ $Y=0.33 $X2=17.17 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.195
+ $Y=0.33 $X2=16.33 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.365
+ $Y=0.33 $X2=15.49 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=14.415
+ $Y=0.235 $X2=14.55 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=13.475
+ $Y=0.235 $X2=13.61 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_911# 1 2 3 4 5 18 22 27 28 29
+ 32 34 38 41 43 44
c79 38 0 1.10627e-19 $X=17.17 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=17.21 $Y=5.015
+ $X2=17.21 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.415 $Y=5.1
+ $X2=16.33 $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.085 $Y=5.1
+ $X2=17.21 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.085 $Y=5.1
+ $X2=16.415 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.33 $Y=5.015
+ $X2=16.33 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.33 $Y=5.015
+ $X2=16.33 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.245 $Y=5.1
+ $X2=16.33 $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.245 $Y=5.1
+ $X2=15.575 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.44 $Y=5.015
+ $X2=15.575 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.44 $Y=5.015
+ $X2=15.44 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=15.44 $Y=4.725
+ $X2=15.44 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=4.64
+ $X2=14.55 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.305 $Y=4.64
+ $X2=15.44 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.305 $Y=4.64
+ $X2=14.715 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.775 $Y=4.64
+ $X2=13.61 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=4.64
+ $X2=14.55 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=4.64
+ $X2=13.775 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=17.035
+ $Y=4.59 $X2=17.17 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.195
+ $Y=4.59 $X2=16.33 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.365
+ $Y=4.59 $X2=15.49 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=14.415
+ $Y=4.555 $X2=14.55 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=13.475
+ $Y=4.555 $X2=13.61 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=25.03 $Y=0.715
+ $X2=25.03 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=0.8
+ $X2=24.09 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=24.865 $Y=0.8
+ $X2=25.03 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=0.8
+ $X2=24.255 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=24.09 $Y=0.715
+ $X2=24.09 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=24.09 $Y=0.715
+ $X2=24.09 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=0.8
+ $X2=24.09 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=23.925 $Y=0.8
+ $X2=23.335 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.2 $Y=0.715
+ $X2=23.335 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=23.2 $Y=0.715
+ $X2=23.2 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=23.2 $Y=0.425
+ $X2=23.2 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.395 $Y=0.34
+ $X2=22.31 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.065 $Y=0.34
+ $X2=23.2 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=23.065 $Y=0.34
+ $X2=22.395 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.31 $Y=0.425
+ $X2=22.31 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=22.31 $Y=0.425
+ $X2=22.31 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.225 $Y=0.34
+ $X2=22.31 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.225 $Y=0.34
+ $X2=21.555 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=21.43 $Y=0.425
+ $X2=21.555 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=21.43 $Y=0.425
+ $X2=21.43 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=24.895
+ $Y=0.235 $X2=25.03 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=23.955
+ $Y=0.235 $X2=24.09 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=23.015
+ $Y=0.33 $X2=23.15 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.175
+ $Y=0.33 $X2=22.31 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.345
+ $Y=0.33 $X2=21.47 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_918# 1 2 3 4 5 18 20 21 24 26
+ 31 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=4.64
+ $X2=24.09 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.865 $Y=4.64
+ $X2=25.03 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=4.64
+ $X2=24.255 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=4.64
+ $X2=24.09 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=23.925 $Y=4.64
+ $X2=23.335 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=23.2 $Y=5.015
+ $X2=23.2 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.2 $Y=4.725
+ $X2=23.335 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=23.2 $Y=4.725
+ $X2=23.2 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.395 $Y=5.1
+ $X2=22.31 $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.065 $Y=5.1
+ $X2=23.2 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=23.065 $Y=5.1
+ $X2=22.395 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.31 $Y=5.015
+ $X2=22.31 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=22.31 $Y=5.015
+ $X2=22.31 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.225 $Y=5.1
+ $X2=22.31 $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.225 $Y=5.1
+ $X2=21.555 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=21.43 $Y=5.015
+ $X2=21.555 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=21.43 $Y=5.015
+ $X2=21.43 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=24.895
+ $Y=4.555 $X2=25.03 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=23.955
+ $Y=4.555 $X2=24.09 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=23.015
+ $Y=4.59 $X2=23.15 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.175
+ $Y=4.59 $X2=22.31 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.345
+ $Y=4.59 $X2=21.47 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=30.51 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=30.55 $Y=0.425
+ $X2=30.55 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.755 $Y=0.34
+ $X2=29.67 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=30.425 $Y=0.34
+ $X2=30.55 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=30.425 $Y=0.34
+ $X2=29.755 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.67 $Y=0.425
+ $X2=29.67 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=29.67 $Y=0.425
+ $X2=29.67 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.585 $Y=0.34
+ $X2=29.67 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=29.585 $Y=0.34
+ $X2=28.915 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=28.78 $Y=0.715
+ $X2=28.78 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=28.78 $Y=0.425
+ $X2=28.915 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=28.78 $Y=0.425
+ $X2=28.78 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=28.055 $Y=0.8
+ $X2=27.89 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=28.645 $Y=0.8
+ $X2=28.78 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=28.645 $Y=0.8
+ $X2=28.055 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=27.89 $Y=0.715
+ $X2=27.89 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=27.89 $Y=0.715
+ $X2=27.89 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.725 $Y=0.8
+ $X2=27.89 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=27.725 $Y=0.8
+ $X2=27.115 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=26.95 $Y=0.715
+ $X2=27.115 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=26.95 $Y=0.715
+ $X2=26.95 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=30.375
+ $Y=0.33 $X2=30.51 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=29.535
+ $Y=0.33 $X2=29.67 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=28.705
+ $Y=0.33 $X2=28.83 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=27.755
+ $Y=0.235 $X2=27.89 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=26.815
+ $Y=0.235 $X2=26.95 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_911# 1 2 3 4 5 18 22 27 28 29
+ 32 34 38 41 43 44
c79 38 0 1.10627e-19 $X=30.51 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=30.55 $Y=5.015
+ $X2=30.55 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.755 $Y=5.1
+ $X2=29.67 $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=30.425 $Y=5.1
+ $X2=30.55 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=30.425 $Y=5.1
+ $X2=29.755 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.67 $Y=5.015
+ $X2=29.67 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=29.67 $Y=5.015
+ $X2=29.67 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=29.585 $Y=5.1
+ $X2=29.67 $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=29.585 $Y=5.1
+ $X2=28.915 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=28.78 $Y=5.015
+ $X2=28.915 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=28.78 $Y=5.015
+ $X2=28.78 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=28.78 $Y=4.725
+ $X2=28.78 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=28.055 $Y=4.64
+ $X2=27.89 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=28.645 $Y=4.64
+ $X2=28.78 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=28.645 $Y=4.64
+ $X2=28.055 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.115 $Y=4.64
+ $X2=26.95 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=27.725 $Y=4.64
+ $X2=27.89 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=27.725 $Y=4.64
+ $X2=27.115 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=30.375
+ $Y=4.59 $X2=30.51 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=29.535
+ $Y=4.59 $X2=29.67 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=28.705
+ $Y=4.59 $X2=28.83 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=27.755
+ $Y=4.555 $X2=27.89 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=26.815
+ $Y=4.555 $X2=26.95 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=38.37 $Y=0.715
+ $X2=38.37 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.595 $Y=0.8
+ $X2=37.43 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=38.205 $Y=0.8
+ $X2=38.37 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=38.205 $Y=0.8
+ $X2=37.595 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=37.43 $Y=0.715
+ $X2=37.43 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=37.43 $Y=0.715
+ $X2=37.43 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.265 $Y=0.8
+ $X2=37.43 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=37.265 $Y=0.8
+ $X2=36.675 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=36.54 $Y=0.715
+ $X2=36.675 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=36.54 $Y=0.715
+ $X2=36.54 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=36.54 $Y=0.425
+ $X2=36.54 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.735 $Y=0.34
+ $X2=35.65 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=36.405 $Y=0.34
+ $X2=36.54 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=36.405 $Y=0.34
+ $X2=35.735 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.65 $Y=0.425
+ $X2=35.65 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=35.65 $Y=0.425
+ $X2=35.65 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.565 $Y=0.34
+ $X2=35.65 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=35.565 $Y=0.34
+ $X2=34.895 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=34.77 $Y=0.425
+ $X2=34.895 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=34.77 $Y=0.425
+ $X2=34.77 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=38.235
+ $Y=0.235 $X2=38.37 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=37.295
+ $Y=0.235 $X2=37.43 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=36.355
+ $Y=0.33 $X2=36.49 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=35.515
+ $Y=0.33 $X2=35.65 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=34.685
+ $Y=0.33 $X2=34.81 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_918# 1 2 3 4 5 18 20 21 24 26
+ 31 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.595 $Y=4.64
+ $X2=37.43 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=38.205 $Y=4.64
+ $X2=38.37 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=38.205 $Y=4.64
+ $X2=37.595 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=37.265 $Y=4.64
+ $X2=37.43 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=37.265 $Y=4.64
+ $X2=36.675 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=36.54 $Y=5.015
+ $X2=36.54 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=36.54 $Y=4.725
+ $X2=36.675 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=36.54 $Y=4.725
+ $X2=36.54 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.735 $Y=5.1
+ $X2=35.65 $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=36.405 $Y=5.1
+ $X2=36.54 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=36.405 $Y=5.1
+ $X2=35.735 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.65 $Y=5.015
+ $X2=35.65 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=35.65 $Y=5.015
+ $X2=35.65 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=35.565 $Y=5.1
+ $X2=35.65 $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=35.565 $Y=5.1
+ $X2=34.895 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=34.77 $Y=5.015
+ $X2=34.895 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=34.77 $Y=5.015
+ $X2=34.77 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=38.235
+ $Y=4.555 $X2=38.37 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=37.295
+ $Y=4.555 $X2=37.43 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=36.355
+ $Y=4.59 $X2=36.49 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=35.515
+ $Y=4.59 $X2=35.65 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=34.685
+ $Y=4.59 $X2=34.81 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=43.39 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=43.43 $Y=0.425
+ $X2=43.43 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.635 $Y=0.34
+ $X2=42.55 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=43.305 $Y=0.34
+ $X2=43.43 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=43.305 $Y=0.34
+ $X2=42.635 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.55 $Y=0.425
+ $X2=42.55 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=42.55 $Y=0.425
+ $X2=42.55 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.465 $Y=0.34
+ $X2=42.55 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=42.465 $Y=0.34
+ $X2=41.795 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=41.66 $Y=0.715
+ $X2=41.66 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=41.66 $Y=0.425
+ $X2=41.795 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=41.66 $Y=0.425
+ $X2=41.66 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.935 $Y=0.8
+ $X2=40.77 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=41.525 $Y=0.8
+ $X2=41.66 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=41.525 $Y=0.8
+ $X2=40.935 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=40.77 $Y=0.715
+ $X2=40.77 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=40.77 $Y=0.715
+ $X2=40.77 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.605 $Y=0.8
+ $X2=40.77 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=40.605 $Y=0.8
+ $X2=39.995 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=39.83 $Y=0.715
+ $X2=39.995 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=39.83 $Y=0.715
+ $X2=39.83 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=43.255
+ $Y=0.33 $X2=43.39 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=42.415
+ $Y=0.33 $X2=42.55 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=41.585
+ $Y=0.33 $X2=41.71 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=40.635
+ $Y=0.235 $X2=40.77 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=39.695
+ $Y=0.235 $X2=39.83 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_911# 1 2 3 4 5 18 22 27 28 29
+ 32 34 38 41 43 44
c79 38 0 1.10627e-19 $X=43.39 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=43.43 $Y=5.015
+ $X2=43.43 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.635 $Y=5.1
+ $X2=42.55 $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=43.305 $Y=5.1
+ $X2=43.43 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=43.305 $Y=5.1
+ $X2=42.635 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.55 $Y=5.015
+ $X2=42.55 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=42.55 $Y=5.015
+ $X2=42.55 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=42.465 $Y=5.1
+ $X2=42.55 $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=42.465 $Y=5.1
+ $X2=41.795 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=41.66 $Y=5.015
+ $X2=41.795 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=41.66 $Y=5.015
+ $X2=41.66 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=41.66 $Y=4.725
+ $X2=41.66 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.935 $Y=4.64
+ $X2=40.77 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=41.525 $Y=4.64
+ $X2=41.66 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=41.525 $Y=4.64
+ $X2=40.935 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=39.995 $Y=4.64
+ $X2=39.83 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=40.605 $Y=4.64
+ $X2=40.77 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=40.605 $Y=4.64
+ $X2=39.995 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=43.255
+ $Y=4.59 $X2=43.39 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=42.415
+ $Y=4.59 $X2=42.55 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=41.585
+ $Y=4.59 $X2=41.71 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=40.635
+ $Y=4.555 $X2=40.77 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=39.695
+ $Y=4.555 $X2=39.83 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=51.25 $Y=0.715
+ $X2=51.25 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.475 $Y=0.8
+ $X2=50.31 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=51.085 $Y=0.8
+ $X2=51.25 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=51.085 $Y=0.8
+ $X2=50.475 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=50.31 $Y=0.715
+ $X2=50.31 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=50.31 $Y=0.715
+ $X2=50.31 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.145 $Y=0.8
+ $X2=50.31 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=50.145 $Y=0.8
+ $X2=49.555 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=49.42 $Y=0.715
+ $X2=49.555 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=49.42 $Y=0.715
+ $X2=49.42 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=49.42 $Y=0.425
+ $X2=49.42 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.615 $Y=0.34
+ $X2=48.53 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=49.285 $Y=0.34
+ $X2=49.42 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=49.285 $Y=0.34
+ $X2=48.615 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.53 $Y=0.425
+ $X2=48.53 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=48.53 $Y=0.425
+ $X2=48.53 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.445 $Y=0.34
+ $X2=48.53 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=48.445 $Y=0.34
+ $X2=47.775 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=47.65 $Y=0.425
+ $X2=47.775 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=47.65 $Y=0.425
+ $X2=47.65 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=51.115
+ $Y=0.235 $X2=51.25 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=50.175
+ $Y=0.235 $X2=50.31 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=49.235
+ $Y=0.33 $X2=49.37 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=48.395
+ $Y=0.33 $X2=48.53 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=47.565
+ $Y=0.33 $X2=47.69 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_918# 1 2 3 4 5 18 20 21 24 26
+ 31 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.475 $Y=4.64
+ $X2=50.31 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=51.085 $Y=4.64
+ $X2=51.25 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=51.085 $Y=4.64
+ $X2=50.475 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=50.145 $Y=4.64
+ $X2=50.31 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=50.145 $Y=4.64
+ $X2=49.555 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=49.42 $Y=5.015
+ $X2=49.42 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=49.42 $Y=4.725
+ $X2=49.555 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=49.42 $Y=4.725
+ $X2=49.42 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.615 $Y=5.1
+ $X2=48.53 $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=49.285 $Y=5.1
+ $X2=49.42 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=49.285 $Y=5.1
+ $X2=48.615 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.53 $Y=5.015
+ $X2=48.53 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=48.53 $Y=5.015
+ $X2=48.53 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=48.445 $Y=5.1
+ $X2=48.53 $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=48.445 $Y=5.1
+ $X2=47.775 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=47.65 $Y=5.015
+ $X2=47.775 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=47.65 $Y=5.015
+ $X2=47.65 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=51.115
+ $Y=4.555 $X2=51.25 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=50.175
+ $Y=4.555 $X2=50.31 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=49.235
+ $Y=4.59 $X2=49.37 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=48.395
+ $Y=4.59 $X2=48.53 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=47.565
+ $Y=4.59 $X2=47.69 $Y2=4.85
.ends

