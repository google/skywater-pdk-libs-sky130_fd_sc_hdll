* File: sky130_fd_sc_hdll__a32oi_1.spice
* Created: Wed Sep  2 08:20:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a32oi_1  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1005 A_119_47# N_B2_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=5.532 M=1 R=4.33333 SA=75000.2
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.17225
+ AS=0.08775 PD=1.18 PS=0.92 NRD=4.608 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1009 A_339_47# N_A1_M1009_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.17225 PD=0.92 PS=1.18 NRD=14.76 NRS=41.532 M=1 R=4.33333 SA=75001.3
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 A_423_47# N_A2_M1004_g A_339_47# VNB NSHORT L=0.15 W=0.65 AD=0.10725
+ AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=14.76 M=1 R=4.33333 SA=75001.8
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g A_423_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.10725 PD=1.92 PS=0.98 NRD=8.304 NRS=20.304 M=1 R=4.33333 SA=75002.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_B2_M1002_g N_A_27_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1000 N_A_27_297#_M1000_d N_B1_M1000_g N_Y_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.225 AS=0.145 PD=1.45 PS=1.29 NRD=32.4853 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_27_297#_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.225 PD=1.29 PS=1.45 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.3 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1003_d N_A2_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.145 PD=1.3 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A3_M1008_g N_A_27_297#_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.15 PD=2.54 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90002.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hdll__a32oi_1.pxi.spice"
*
.ends
*
*
