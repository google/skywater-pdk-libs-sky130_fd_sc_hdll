* File: sky130_fd_sc_hdll__and2_1.spice
* Created: Wed Sep  2 08:21:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2_1.pex.spice"
.subckt sky130_fd_sc_hdll__and2_1  VNB VPB A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 A_123_75# N_A_M1005_g N_A_27_75#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1386 PD=0.69 PS=1.5 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75000.3
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g A_123_75# VNB NSHORT L=0.15 W=0.42
+ AD=0.0944411 AS=0.0567 PD=0.828224 PS=0.69 NRD=28.56 NRS=22.848 M=1 R=2.8
+ SA=75000.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_75#_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.23725 AS=0.146159 PD=2.03 PS=1.28178 NRD=14.76 NRS=5.532 M=1 R=4.33333
+ SA=75000.9 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1000 N_A_27_75#_M1000_d N_A_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1218 PD=0.71 PS=1.42 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_B_M1004_g N_A_27_75#_M1000_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0957866 AS=0.0609 PD=0.81338 PS=0.71 NRD=31.6579 NRS=2.3443 M=1 R=2.33333
+ SA=90000.7 SB=90001 A=0.0756 P=1.2 MULT=1
MM1002 N_X_M1002_d N_A_27_75#_M1002_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.52 AS=0.228063 PD=3.04 PS=1.93662 NRD=27.5603 NRS=5.8903 M=1 R=5.55556
+ SA=90000.6 SB=90000.4 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_10 A A PROBETYPE=1
pX8_noxref noxref_11 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and2_1.pxi.spice"
*
.ends
*
*
