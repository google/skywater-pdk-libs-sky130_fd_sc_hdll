* File: sky130_fd_sc_hdll__o31ai_1.pxi.spice
* Created: Thu Aug 27 19:22:25 2020
* 
x_PM_SKY130_FD_SC_HDLL__O31AI_1%A1 N_A1_c_45_n N_A1_M1000_g N_A1_c_42_n
+ N_A1_M1005_g A1 N_A1_c_44_n PM_SKY130_FD_SC_HDLL__O31AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O31AI_1%A2 N_A2_c_66_n N_A2_M1006_g N_A2_c_67_n
+ N_A2_M1001_g A2 A2 A2 A2 N_A2_c_68_n PM_SKY130_FD_SC_HDLL__O31AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O31AI_1%A3 N_A3_c_99_n N_A3_M1004_g N_A3_c_100_n
+ N_A3_M1003_g A3 A3 N_A3_c_104_n PM_SKY130_FD_SC_HDLL__O31AI_1%A3
x_PM_SKY130_FD_SC_HDLL__O31AI_1%B1 N_B1_c_135_n N_B1_M1002_g N_B1_c_138_n
+ N_B1_M1007_g B1 N_B1_c_137_n B1 PM_SKY130_FD_SC_HDLL__O31AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O31AI_1%VPWR N_VPWR_M1000_s N_VPWR_M1007_d
+ N_VPWR_c_164_n N_VPWR_c_165_n N_VPWR_c_166_n N_VPWR_c_167_n VPWR
+ N_VPWR_c_168_n N_VPWR_c_163_n PM_SKY130_FD_SC_HDLL__O31AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O31AI_1%Y N_Y_M1002_d N_Y_M1003_d Y Y Y Y Y Y Y
+ N_Y_c_205_n PM_SKY130_FD_SC_HDLL__O31AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O31AI_1%VGND N_VGND_M1005_s N_VGND_M1001_d
+ N_VGND_c_224_n N_VGND_c_225_n N_VGND_c_226_n N_VGND_c_227_n VGND
+ N_VGND_c_228_n N_VGND_c_229_n N_VGND_c_230_n
+ PM_SKY130_FD_SC_HDLL__O31AI_1%VGND
x_PM_SKY130_FD_SC_HDLL__O31AI_1%A_119_47# N_A_119_47#_M1005_d
+ N_A_119_47#_M1004_d N_A_119_47#_c_262_n N_A_119_47#_c_260_n
+ N_A_119_47#_c_261_n N_A_119_47#_c_269_n
+ PM_SKY130_FD_SC_HDLL__O31AI_1%A_119_47#
cc_1 VNB N_A1_c_42_n 0.0221197f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB A1 0.00930364f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A1_c_44_n 0.0445819f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A2_c_66_n 0.0199196f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_A2_c_67_n 0.0167728f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_A2_c_68_n 0.00512542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A3_c_99_n 0.0179319f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A3_c_100_n 0.0218949f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB A3 0.00408954f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_10 VNB N_B1_c_135_n 0.0212279f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB B1 0.0154163f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_B1_c_137_n 0.0440124f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_13 VNB N_VPWR_c_163_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB Y 0.00760184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_224_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_VGND_c_225_n 0.00655427f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_17 VNB N_VGND_c_226_n 0.0202127f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_18 VNB N_VGND_c_227_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_228_n 0.0408342f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_229_n 0.168894f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_230_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_119_47#_c_260_n 0.0102862f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_23 VNB N_A_119_47#_c_261_n 0.00283849f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_24 VPB N_A1_c_45_n 0.0205019f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_25 VPB A1 0.0035502f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_26 VPB N_A1_c_44_n 0.0184112f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_27 VPB N_A2_c_66_n 0.0234198f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_28 VPB N_A2_c_68_n 0.00325558f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A3_c_100_n 0.0270709f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_30 VPB A3 0.00156123f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_31 VPB N_A3_c_104_n 0.00136794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_B1_c_138_n 0.0225344f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_33 VPB B1 0.00462051f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_34 VPB N_B1_c_137_n 0.0217639f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_35 VPB N_VPWR_c_164_n 0.0160252f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_36 VPB N_VPWR_c_165_n 0.0420814f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_37 VPB N_VPWR_c_166_n 0.0129411f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_38 VPB N_VPWR_c_167_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_168_n 0.0509427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_163_n 0.040104f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB Y 0.00122593f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 N_A1_c_45_n N_A2_c_66_n 0.0458229f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_43 N_A1_c_44_n N_A2_c_66_n 0.0253274f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_44 N_A1_c_42_n N_A2_c_67_n 0.0100769f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_45 N_A1_c_45_n N_A2_c_68_n 0.00722107f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_46 A1 N_A2_c_68_n 0.0205196f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A1_c_44_n N_A2_c_68_n 0.00481954f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_48 N_A1_c_45_n N_VPWR_c_165_n 0.0164394f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_49 A1 N_VPWR_c_165_n 0.02421f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A1_c_44_n N_VPWR_c_165_n 0.00211327f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_51 N_A1_c_45_n N_VPWR_c_168_n 0.00642146f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A1_c_45_n N_VPWR_c_163_n 0.0108369f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A1_c_42_n N_VGND_c_225_n 0.00634941f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 A1 N_VGND_c_225_n 0.0139721f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A1_c_44_n N_VGND_c_225_n 0.00431028f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_56 N_A1_c_42_n N_VGND_c_226_n 0.00465454f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A1_c_42_n N_VGND_c_229_n 0.00894173f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 N_A1_c_42_n N_A_119_47#_c_262_n 0.00753207f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A1_c_42_n N_A_119_47#_c_261_n 0.00674737f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A2_c_67_n N_A3_c_99_n 0.0228372f $X=1 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_61 N_A2_c_66_n N_A3_c_100_n 0.0722321f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A2_c_68_n N_A3_c_100_n 0.00518269f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A2_c_66_n A3 8.70257e-19 $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A2_c_68_n A3 0.0186386f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A2_c_66_n N_A3_c_104_n 0.00114408f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A2_c_68_n N_A3_c_104_n 0.0258749f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A2_c_66_n N_VPWR_c_165_n 0.00166661f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A2_c_66_n N_VPWR_c_168_n 0.00429201f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A2_c_68_n N_VPWR_c_168_n 0.0300356f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_70 N_A2_c_66_n N_VPWR_c_163_n 0.00618266f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A2_c_68_n N_VPWR_c_163_n 0.0183557f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A2_c_68_n A_117_297# 0.00511952f $X=0.94 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_73 N_A2_c_67_n N_VGND_c_226_n 0.00439206f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A2_c_67_n N_VGND_c_227_n 0.00268723f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A2_c_67_n N_VGND_c_229_n 0.0061063f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A2_c_66_n N_A_119_47#_c_260_n 8.65373e-19 $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A2_c_67_n N_A_119_47#_c_260_n 0.01036f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A2_c_68_n N_A_119_47#_c_260_n 0.0162351f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A2_c_66_n N_A_119_47#_c_261_n 0.00235664f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A2_c_68_n N_A_119_47#_c_261_n 0.0265777f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A2_c_67_n N_A_119_47#_c_269_n 4.78929e-19 $X=1 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A3_c_99_n N_B1_c_135_n 0.014496f $X=1.42 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_83 N_A3_c_100_n N_B1_c_138_n 0.0130857f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A3_c_104_n N_B1_c_138_n 0.00192598f $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_85 N_A3_c_100_n N_B1_c_137_n 0.0115296f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_86 A3 N_B1_c_137_n 7.69841e-19 $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A3_c_104_n N_B1_c_137_n 2.1198e-19 $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_88 N_A3_c_100_n N_VPWR_c_168_n 0.00588982f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A3_c_104_n N_VPWR_c_168_n 0.010519f $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_90 N_A3_c_100_n N_VPWR_c_163_n 0.0104679f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A3_c_104_n N_VPWR_c_163_n 0.00851311f $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_92 N_A3_c_104_n N_Y_M1003_d 0.010084f $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_93 N_A3_c_99_n Y 0.00169875f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A3_c_100_n Y 0.00687413f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_95 A3 Y 0.0190908f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_96 N_A3_c_104_n Y 0.0772104f $X=1.575 $Y=1.2 $X2=0 $Y2=0
cc_97 N_A3_c_99_n N_Y_c_205_n 0.00269062f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A3_c_99_n N_VGND_c_227_n 0.00268723f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A3_c_99_n N_VGND_c_228_n 0.00431995f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A3_c_99_n N_VGND_c_229_n 0.00633994f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A3_c_99_n N_A_119_47#_c_260_n 0.0104435f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A3_c_100_n N_A_119_47#_c_260_n 0.00322034f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_103 A3 N_A_119_47#_c_260_n 0.0292401f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A3_c_99_n N_A_119_47#_c_269_n 0.00467733f $X=1.42 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_c_138_n N_VPWR_c_167_n 0.00779274f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_106 B1 N_VPWR_c_167_n 0.0138735f $X=2.475 $Y=1.105 $X2=0 $Y2=0
cc_107 N_B1_c_137_n N_VPWR_c_167_n 0.00391367f $X=2.205 $Y=1.202 $X2=0 $Y2=0
cc_108 N_B1_c_138_n N_VPWR_c_168_n 0.00643255f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B1_c_138_n N_VPWR_c_163_n 0.0126309f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B1_c_135_n Y 0.00559581f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B1_c_138_n Y 0.0218758f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_112 B1 Y 0.0243399f $X=2.475 $Y=1.105 $X2=0 $Y2=0
cc_113 N_B1_c_137_n Y 0.0212137f $X=2.205 $Y=1.202 $X2=0 $Y2=0
cc_114 N_B1_c_135_n N_Y_c_205_n 0.0149275f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_115 B1 N_Y_c_205_n 0.0137505f $X=2.475 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B1_c_137_n N_Y_c_205_n 0.0109591f $X=2.205 $Y=1.202 $X2=0 $Y2=0
cc_117 N_B1_c_135_n N_VGND_c_228_n 0.00358715f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_135_n N_VGND_c_229_n 0.00683346f $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B1_c_135_n N_A_119_47#_c_260_n 6.17616e-19 $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B1_c_135_n N_A_119_47#_c_269_n 8.43697e-19 $X=2.06 $Y=0.995 $X2=0 $Y2=0
cc_121 N_VPWR_c_163_n A_117_297# 0.003138f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_122 N_VPWR_c_163_n A_213_297# 0.0110423f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_123 N_VPWR_c_163_n N_Y_M1003_d 0.0113781f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_124 N_VPWR_c_167_n Y 0.0622152f $X=2.44 $Y=1.66 $X2=0 $Y2=0
cc_125 N_VPWR_c_168_n Y 0.0167439f $X=2.355 $Y=2.72 $X2=0 $Y2=0
cc_126 N_VPWR_c_163_n Y 0.0100703f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_127 N_Y_c_205_n N_VGND_c_228_n 0.0369619f $X=2.33 $Y=0.4 $X2=0 $Y2=0
cc_128 N_Y_M1002_d N_VGND_c_229_n 0.00423707f $X=2.135 $Y=0.235 $X2=0 $Y2=0
cc_129 N_Y_c_205_n N_VGND_c_229_n 0.022536f $X=2.33 $Y=0.4 $X2=0 $Y2=0
cc_130 Y N_A_119_47#_M1004_d 5.44209e-19 $X=2.045 $Y=0.85 $X2=0 $Y2=0
cc_131 N_Y_c_205_n N_A_119_47#_M1004_d 0.00713875f $X=2.33 $Y=0.4 $X2=0 $Y2=0
cc_132 N_Y_c_205_n N_A_119_47#_c_260_n 0.0147555f $X=2.33 $Y=0.4 $X2=0 $Y2=0
cc_133 N_Y_c_205_n N_A_119_47#_c_269_n 0.0226284f $X=2.33 $Y=0.4 $X2=0 $Y2=0
cc_134 N_VGND_c_229_n N_A_119_47#_M1005_d 0.00277427f $X=2.53 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_135 N_VGND_c_229_n N_A_119_47#_M1004_d 0.0102227f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_136 N_VGND_c_225_n N_A_119_47#_c_262_n 0.0357963f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_137 N_VGND_c_226_n N_A_119_47#_c_262_n 0.0234201f $X=1.125 $Y=0 $X2=0 $Y2=0
cc_138 N_VGND_c_229_n N_A_119_47#_c_262_n 0.0141066f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_139 N_VGND_M1001_d N_A_119_47#_c_260_n 0.00162006f $X=1.075 $Y=0.235 $X2=0
+ $Y2=0
cc_140 N_VGND_c_226_n N_A_119_47#_c_260_n 0.00255762f $X=1.125 $Y=0 $X2=0 $Y2=0
cc_141 N_VGND_c_227_n N_A_119_47#_c_260_n 0.0122414f $X=1.21 $Y=0.4 $X2=0 $Y2=0
cc_142 N_VGND_c_228_n N_A_119_47#_c_260_n 0.00193763f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_143 N_VGND_c_229_n N_A_119_47#_c_260_n 0.00963293f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_144 N_VGND_c_225_n N_A_119_47#_c_261_n 0.0133879f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_145 N_VGND_c_228_n N_A_119_47#_c_269_n 0.00639221f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_146 N_VGND_c_229_n N_A_119_47#_c_269_n 0.00815833f $X=2.53 $Y=0 $X2=0 $Y2=0
