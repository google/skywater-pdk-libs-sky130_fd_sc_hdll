* File: sky130_fd_sc_hdll__and4_1.pxi.spice
* Created: Wed Sep  2 08:22:53 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4_1%A N_A_c_65_n N_A_c_66_n N_A_M1001_g N_A_M1007_g A
+ N_A_c_64_n PM_SKY130_FD_SC_HDLL__AND4_1%A
x_PM_SKY130_FD_SC_HDLL__AND4_1%B N_B_M1002_g N_B_c_99_n N_B_c_100_n N_B_M1008_g
+ B B N_B_c_98_n PM_SKY130_FD_SC_HDLL__AND4_1%B
x_PM_SKY130_FD_SC_HDLL__AND4_1%C N_C_M1006_g N_C_c_137_n N_C_c_138_n N_C_M1004_g
+ C C C N_C_c_136_n PM_SKY130_FD_SC_HDLL__AND4_1%C
x_PM_SKY130_FD_SC_HDLL__AND4_1%D N_D_M1000_g N_D_c_176_n N_D_c_177_n N_D_M1009_g
+ D N_D_c_175_n D PM_SKY130_FD_SC_HDLL__AND4_1%D
x_PM_SKY130_FD_SC_HDLL__AND4_1%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1001_d
+ N_A_27_47#_M1004_d N_A_27_47#_c_216_n N_A_27_47#_M1003_g N_A_27_47#_c_217_n
+ N_A_27_47#_M1005_g N_A_27_47#_c_218_n N_A_27_47#_c_222_n N_A_27_47#_c_223_n
+ N_A_27_47#_c_224_n N_A_27_47#_c_225_n N_A_27_47#_c_219_n N_A_27_47#_c_236_n
+ N_A_27_47#_c_227_n N_A_27_47#_c_228_n PM_SKY130_FD_SC_HDLL__AND4_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4_1%VPWR N_VPWR_M1001_s N_VPWR_M1008_d N_VPWR_M1009_d
+ N_VPWR_c_301_n N_VPWR_c_302_n N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_305_n
+ VPWR N_VPWR_c_306_n N_VPWR_c_307_n N_VPWR_c_300_n N_VPWR_c_309_n
+ N_VPWR_c_310_n PM_SKY130_FD_SC_HDLL__AND4_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4_1%X N_X_M1005_d N_X_M1003_d X X X X X X X
+ N_X_c_350_n X PM_SKY130_FD_SC_HDLL__AND4_1%X
x_PM_SKY130_FD_SC_HDLL__AND4_1%VGND N_VGND_M1000_d N_VGND_c_375_n VGND
+ N_VGND_c_376_n N_VGND_c_377_n N_VGND_c_378_n N_VGND_c_379_n
+ PM_SKY130_FD_SC_HDLL__AND4_1%VGND
cc_1 VNB N_A_M1007_g 0.0332287f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.0241287f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_c_64_n 0.038823f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_B_M1002_g 0.0258854f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_5 VNB B 0.00818964f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_6 VNB N_B_c_98_n 0.019473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_C_M1006_g 0.0289615f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_8 VNB C 0.00436785f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_9 VNB N_C_c_136_n 0.021187f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_10 VNB N_D_M1000_g 0.0311155f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_11 VNB D 0.00411023f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_12 VNB N_D_c_175_n 0.0205719f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_13 VNB N_A_27_47#_c_216_n 0.0250521f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_14 VNB N_A_27_47#_c_217_n 0.0210597f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_15 VNB N_A_27_47#_c_218_n 0.00393054f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_16 VNB N_A_27_47#_c_219_n 0.00402475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_300_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 0.0258943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_X_c_350_n 0.0207068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_375_n 0.00530675f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_21 VNB N_VGND_c_376_n 0.0570647f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_22 VNB N_VGND_c_377_n 0.0269301f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_23 VNB N_VGND_c_378_n 0.183059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_379_n 0.00516539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A_c_65_n 0.0328685f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_26 VPB N_A_c_66_n 0.0252865f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_27 VPB A 0.0376224f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_28 VPB N_A_c_64_n 0.0117539f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_29 VPB N_B_c_99_n 0.0312978f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_30 VPB N_B_c_100_n 0.0221274f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_31 VPB B 0.0019121f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_B_c_98_n 0.00303637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_C_c_137_n 0.0317669f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_34 VPB N_C_c_138_n 0.0224081f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_35 VPB C 0.00151418f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_36 VPB N_C_c_136_n 0.00340421f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_37 VPB N_D_c_176_n 0.0330594f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_38 VPB N_D_c_177_n 0.0230033f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_39 VPB D 6.7738e-19 $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_40 VPB N_D_c_175_n 0.00278754f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_41 VPB N_A_27_47#_c_216_n 0.028895f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_42 VPB N_A_27_47#_c_218_n 0.00177669f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_43 VPB N_A_27_47#_c_222_n 0.00797266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_223_n 0.00905617f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_224_n 0.00826901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_225_n 0.0028031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_219_n 0.00174064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_47#_c_227_n 0.00733094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_47#_c_228_n 0.00576943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_301_n 0.0101963f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_51 VPB N_VPWR_c_302_n 0.0120831f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_52 VPB N_VPWR_c_303_n 0.00322578f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_53 VPB N_VPWR_c_304_n 0.0158757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_305_n 0.00357129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_306_n 0.0148955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_307_n 0.0253827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_300_n 0.0452452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_309_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_310_n 0.0059074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB X 0.0371346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.010718f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 N_A_M1007_g N_B_M1002_g 0.0214332f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_63 N_A_c_65_n N_B_c_99_n 0.0214332f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_64 N_A_c_66_n N_B_c_100_n 0.0316411f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_65 N_A_M1007_g B 0.00197508f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_c_64_n N_B_c_98_n 0.0214332f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_c_65_n N_A_27_47#_c_218_n 0.00381342f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_68 N_A_M1007_g N_A_27_47#_c_218_n 0.0149243f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_218_n 0.0527162f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_64_n N_A_27_47#_c_218_n 0.00944629f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_c_65_n N_A_27_47#_c_222_n 0.00324092f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_72 N_A_c_66_n N_A_27_47#_c_222_n 9.33038e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_73 A N_A_27_47#_c_222_n 0.0226704f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_M1007_g N_A_27_47#_c_236_n 0.0104144f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_75 A N_A_27_47#_c_236_n 0.0123303f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_64_n N_A_27_47#_c_236_n 0.00373141f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_65_n N_A_27_47#_c_227_n 0.0099466f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_227_n 0.0139295f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_79 A N_VPWR_M1001_s 0.00226849f $X=0.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_80 N_A_c_66_n N_VPWR_c_302_n 0.00839181f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_81 A N_VPWR_c_302_n 0.0188536f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_66_n N_VPWR_c_303_n 5.61609e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_83 N_A_c_66_n N_VPWR_c_306_n 0.00643335f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_84 N_A_c_66_n N_VPWR_c_300_n 0.0106848f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_85 A N_VPWR_c_300_n 0.00141964f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_M1007_g N_VGND_c_376_n 0.00357877f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_M1007_g N_VGND_c_378_n 0.00625228f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_88 A N_VGND_c_378_n 0.0038518f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_89 N_B_M1002_g N_C_M1006_g 0.0308651f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_90 B N_C_M1006_g 0.00673563f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_91 N_B_c_99_n N_C_c_137_n 0.0152209f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_92 N_B_c_100_n N_C_c_138_n 0.0269479f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_93 N_B_M1002_g C 5.62228e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_94 B C 0.0760247f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_95 N_B_c_98_n C 3.08958e-19 $X=1 $Y=1.16 $X2=0 $Y2=0
cc_96 N_B_c_98_n N_C_c_136_n 0.0202062f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_M1002_g N_A_27_47#_c_218_n 0.00230131f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_98 N_B_c_99_n N_A_27_47#_c_218_n 0.00354637f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_99 B N_A_27_47#_c_218_n 0.0566787f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_100 N_B_c_99_n N_A_27_47#_c_222_n 0.00743591f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_101 N_B_c_100_n N_A_27_47#_c_222_n 8.10032e-19 $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_102 N_B_c_99_n N_A_27_47#_c_223_n 0.0177813f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_103 B N_A_27_47#_c_223_n 0.0299509f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_104 N_B_c_98_n N_A_27_47#_c_223_n 4.93463e-19 $X=1 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B_M1002_g N_A_27_47#_c_236_n 0.00346086f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_106 N_B_c_100_n N_VPWR_c_302_n 4.91947e-19 $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_107 N_B_c_100_n N_VPWR_c_303_n 0.0137616f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_108 N_B_c_100_n N_VPWR_c_306_n 0.00643335f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_109 N_B_c_100_n N_VPWR_c_300_n 0.0106848f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_110 B A_203_47# 0.00495335f $X=0.98 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_111 N_B_M1002_g N_VGND_c_376_n 0.0037867f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_112 B N_VGND_c_376_n 0.014225f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_113 N_B_M1002_g N_VGND_c_378_n 0.00553827f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_114 B N_VGND_c_378_n 0.0130234f $X=0.98 $Y=0.425 $X2=0 $Y2=0
cc_115 N_C_M1006_g N_D_M1000_g 0.0296336f $X=1.42 $Y=0.445 $X2=0 $Y2=0
cc_116 C N_D_M1000_g 0.00995552f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_117 N_C_c_137_n N_D_c_176_n 0.0136234f $X=1.445 $Y=1.89 $X2=0 $Y2=0
cc_118 N_C_c_138_n N_D_c_177_n 0.0230234f $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_119 N_C_M1006_g D 2.48137e-19 $X=1.42 $Y=0.445 $X2=0 $Y2=0
cc_120 C D 0.0434507f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_121 N_C_c_136_n D 3.3448e-19 $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_122 N_C_c_136_n N_D_c_175_n 0.0202302f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_123 N_C_c_137_n N_A_27_47#_c_223_n 0.0200404f $X=1.445 $Y=1.89 $X2=0 $Y2=0
cc_124 C N_A_27_47#_c_223_n 0.0117493f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_125 N_C_c_137_n N_A_27_47#_c_224_n 0.00750433f $X=1.445 $Y=1.89 $X2=0 $Y2=0
cc_126 N_C_c_138_n N_A_27_47#_c_224_n 8.5324e-19 $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_127 C N_A_27_47#_c_228_n 0.0122602f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_128 N_C_c_136_n N_A_27_47#_c_228_n 5.14458e-19 $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_129 N_C_c_138_n N_VPWR_c_303_n 0.0131783f $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_130 N_C_c_138_n N_VPWR_c_304_n 0.00682361f $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_131 N_C_c_138_n N_VPWR_c_305_n 5.66644e-19 $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_132 N_C_c_138_n N_VPWR_c_300_n 0.011346f $X=1.445 $Y=1.99 $X2=0 $Y2=0
cc_133 C A_299_47# 0.00556334f $X=1.505 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_134 C N_VGND_c_375_n 0.00838236f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_135 N_C_M1006_g N_VGND_c_376_n 0.00462167f $X=1.42 $Y=0.445 $X2=0 $Y2=0
cc_136 C N_VGND_c_376_n 0.0109654f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_137 N_C_M1006_g N_VGND_c_378_n 0.00793053f $X=1.42 $Y=0.445 $X2=0 $Y2=0
cc_138 C N_VGND_c_378_n 0.0100776f $X=1.505 $Y=0.425 $X2=0 $Y2=0
cc_139 N_D_c_176_n N_A_27_47#_c_216_n 0.019082f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_140 N_D_c_177_n N_A_27_47#_c_216_n 0.0120955f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_141 D N_A_27_47#_c_216_n 0.00185033f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_142 N_D_c_175_n N_A_27_47#_c_216_n 0.0202587f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_143 N_D_M1000_g N_A_27_47#_c_217_n 0.017432f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_144 D N_A_27_47#_c_217_n 0.00346115f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_145 N_D_c_176_n N_A_27_47#_c_224_n 0.00591977f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_146 N_D_c_177_n N_A_27_47#_c_224_n 8.35495e-19 $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_147 N_D_c_176_n N_A_27_47#_c_225_n 0.0197748f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_148 D N_A_27_47#_c_225_n 0.0217124f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_149 N_D_c_175_n N_A_27_47#_c_225_n 0.00156944f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_150 N_D_c_176_n N_A_27_47#_c_219_n 0.00323014f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_151 D N_A_27_47#_c_219_n 0.0249117f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_152 N_D_c_175_n N_A_27_47#_c_219_n 3.54436e-19 $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_153 N_D_c_177_n N_VPWR_c_303_n 5.5092e-19 $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_154 N_D_c_177_n N_VPWR_c_304_n 0.00643335f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_155 N_D_c_176_n N_VPWR_c_305_n 0.00177603f $X=1.935 $Y=1.89 $X2=0 $Y2=0
cc_156 N_D_c_177_n N_VPWR_c_305_n 0.0189027f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_157 N_D_c_177_n N_VPWR_c_300_n 0.0107317f $X=1.935 $Y=1.99 $X2=0 $Y2=0
cc_158 D X 0.00425138f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_159 D N_X_c_350_n 0.00306477f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_160 D N_VGND_M1000_d 0.00357417f $X=1.98 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_161 N_D_M1000_g N_VGND_c_375_n 0.00650113f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_162 D N_VGND_c_375_n 0.00843009f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_163 N_D_M1000_g N_VGND_c_376_n 0.00486119f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_164 D N_VGND_c_376_n 0.00285157f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_165 N_D_M1000_g N_VGND_c_378_n 0.00816509f $X=1.91 $Y=0.445 $X2=0 $Y2=0
cc_166 D N_VGND_c_378_n 0.00499623f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_225_n N_VPWR_M1009_d 0.00891095f $X=2.335 $Y=1.58 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_222_n N_VPWR_c_303_n 0.0253855f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_223_n N_VPWR_c_303_n 0.0207344f $X=1.56 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_224_n N_VPWR_c_303_n 0.0238526f $X=1.685 $Y=2.3 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_224_n N_VPWR_c_304_n 0.0156279f $X=1.685 $Y=2.3 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_216_n N_VPWR_c_305_n 0.00330487f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_224_n N_VPWR_c_305_n 0.0297788f $X=1.685 $Y=2.3 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_225_n N_VPWR_c_305_n 0.0268128f $X=2.335 $Y=1.58 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_222_n N_VPWR_c_306_n 0.0149311f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_216_n N_VPWR_c_307_n 0.00702461f $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_M1001_d N_VPWR_c_300_n 0.00328334f $X=0.585 $Y=2.065 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_M1004_d N_VPWR_c_300_n 0.00413826f $X=1.535 $Y=2.065 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_216_n N_VPWR_c_300_n 0.013802f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_222_n N_VPWR_c_300_n 0.00955092f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_224_n N_VPWR_c_300_n 0.00955092f $X=1.685 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_216_n X 0.0174445f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_217_n X 0.0118959f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_225_n X 0.0091161f $X=2.335 $Y=1.58 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_219_n X 0.0251221f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_217_n N_X_c_350_n 0.015204f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_216_n X 0.0061818f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_218_n A_119_47# 6.81697e-19 $X=0.59 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_27_47#_c_236_n A_119_47# 0.00374032f $X=0.59 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_190 N_A_27_47#_c_216_n N_VGND_c_375_n 6.18354e-19 $X=2.485 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_217_n N_VGND_c_375_n 0.00712906f $X=2.51 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_236_n N_VGND_c_376_n 0.0302888f $X=0.59 $Y=0.42 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_217_n N_VGND_c_377_n 0.00585385f $X=2.51 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_M1007_s N_VGND_c_378_n 0.00269774f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_217_n N_VGND_c_378_n 0.0123955f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_236_n N_VGND_c_378_n 0.0187115f $X=0.59 $Y=0.42 $X2=0 $Y2=0
cc_197 N_VPWR_c_300_n N_X_M1003_d 0.00794142f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_307_n X 0.0267545f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_300_n X 0.0148276f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_X_c_350_n N_VGND_c_375_n 0.0115121f $X=2.91 $Y=0.38 $X2=0 $Y2=0
cc_201 N_X_c_350_n N_VGND_c_377_n 0.0216063f $X=2.91 $Y=0.38 $X2=0 $Y2=0
cc_202 N_X_M1005_d N_VGND_c_378_n 0.00754167f $X=2.585 $Y=0.235 $X2=0 $Y2=0
cc_203 N_X_c_350_n N_VGND_c_378_n 0.0146063f $X=2.91 $Y=0.38 $X2=0 $Y2=0
cc_204 A_119_47# N_VGND_c_378_n 0.00810035f $X=0.595 $Y=0.235 $X2=0.73 $Y2=1.665
cc_205 A_203_47# N_VGND_c_378_n 0.00659673f $X=1.015 $Y=0.235 $X2=1 $Y2=1.325
cc_206 A_299_47# N_VGND_c_378_n 0.00770316f $X=1.495 $Y=0.235 $X2=1.49 $Y2=1.16
