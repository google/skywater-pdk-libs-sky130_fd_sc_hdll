* File: sky130_fd_sc_hdll__or2b_2.pxi.spice
* Created: Wed Sep  2 08:48:12 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2B_2%B_N N_B_N_c_66_n N_B_N_M1003_g N_B_N_M1000_g B_N
+ N_B_N_c_65_n B_N PM_SKY130_FD_SC_HDLL__OR2B_2%B_N
x_PM_SKY130_FD_SC_HDLL__OR2B_2%A_27_53# N_A_27_53#_M1000_s N_A_27_53#_M1003_d
+ N_A_27_53#_M1001_g N_A_27_53#_c_90_n N_A_27_53#_M1004_g N_A_27_53#_c_91_n
+ N_A_27_53#_c_92_n N_A_27_53#_c_93_n N_A_27_53#_c_97_n N_A_27_53#_c_94_n
+ PM_SKY130_FD_SC_HDLL__OR2B_2%A_27_53#
x_PM_SKY130_FD_SC_HDLL__OR2B_2%A N_A_c_135_n N_A_M1009_g N_A_c_133_n N_A_c_134_n
+ N_A_c_136_n N_A_M1005_g N_A_c_138_n A N_A_c_140_n A
+ PM_SKY130_FD_SC_HDLL__OR2B_2%A
x_PM_SKY130_FD_SC_HDLL__OR2B_2%A_228_297# N_A_228_297#_M1001_d
+ N_A_228_297#_M1004_s N_A_228_297#_c_188_n N_A_228_297#_M1002_g
+ N_A_228_297#_c_180_n N_A_228_297#_M1006_g N_A_228_297#_c_181_n
+ N_A_228_297#_c_182_n N_A_228_297#_c_191_n N_A_228_297#_M1008_g
+ N_A_228_297#_c_183_n N_A_228_297#_M1007_g N_A_228_297#_c_184_n
+ N_A_228_297#_c_196_n N_A_228_297#_c_243_p N_A_228_297#_c_185_n
+ N_A_228_297#_c_186_n N_A_228_297#_c_187_n N_A_228_297#_c_194_n
+ PM_SKY130_FD_SC_HDLL__OR2B_2%A_228_297#
x_PM_SKY130_FD_SC_HDLL__OR2B_2%VPWR N_VPWR_M1003_s N_VPWR_M1005_d N_VPWR_M1008_d
+ N_VPWR_c_257_n N_VPWR_c_258_n N_VPWR_c_259_n N_VPWR_c_260_n N_VPWR_c_261_n
+ VPWR N_VPWR_c_262_n N_VPWR_c_263_n N_VPWR_c_264_n N_VPWR_c_256_n
+ PM_SKY130_FD_SC_HDLL__OR2B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2B_2%X N_X_M1006_s N_X_M1002_s X N_X_c_297_n
+ PM_SKY130_FD_SC_HDLL__OR2B_2%X
x_PM_SKY130_FD_SC_HDLL__OR2B_2%VGND N_VGND_M1000_d N_VGND_M1009_d N_VGND_M1007_d
+ N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n VGND
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n
+ PM_SKY130_FD_SC_HDLL__OR2B_2%VGND
cc_1 VNB N_B_N_M1000_g 0.0401282f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB B_N 0.00929235f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_B_N_c_65_n 0.0433565f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_27_53#_M1001_g 0.0334724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_53#_c_90_n 0.0381858f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_A_27_53#_c_91_n 0.0206739f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_A_27_53#_c_92_n 0.0164921f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_8 VNB N_A_27_53#_c_93_n 0.00947015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_94_n 0.00459903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_M1009_g 0.0261823f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_11 VNB N_A_c_133_n 0.00697917f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_c_134_n 0.0131969f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB N_A_228_297#_c_180_n 0.0192804f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_14 VNB N_A_228_297#_c_181_n 0.0278921f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_15 VNB N_A_228_297#_c_182_n 0.021025f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_16 VNB N_A_228_297#_c_183_n 0.0223477f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_17 VNB N_A_228_297#_c_184_n 0.0237142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_228_297#_c_185_n 0.00232623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_228_297#_c_186_n 0.00419696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_228_297#_c_187_n 0.00116733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_256_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_297_n 8.88829e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_23 VNB N_VGND_c_317_n 0.0183442f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_24 VNB N_VGND_c_318_n 0.00540513f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_25 VNB N_VGND_c_319_n 0.0118249f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_26 VNB N_VGND_c_320_n 0.0344094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_321_n 0.0268471f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_322_n 0.0188119f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_323_n 0.0227657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_324_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_325_n 0.210932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_B_N_c_66_n 0.0238137f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB B_N 8.86575e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_34 VPB N_B_N_c_65_n 0.0191537f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_35 VPB N_A_27_53#_c_90_n 0.0334732f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_36 VPB N_A_27_53#_c_92_n 0.00329972f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_37 VPB N_A_27_53#_c_97_n 0.00463829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_53#_c_94_n 0.00639431f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_c_135_n 0.0365664f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_40 VPB N_A_c_136_n 0.00637187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_M1005_g 0.011795f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_42 VPB N_A_c_138_n 0.0290475f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_43 VPB A 0.0281685f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_44 VPB N_A_c_140_n 0.0372853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_228_297#_c_188_n 0.0200192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_228_297#_c_181_n 0.0198283f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_47 VPB N_A_228_297#_c_182_n 0.0104802f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_48 VPB N_A_228_297#_c_191_n 0.0213803f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_49 VPB N_A_228_297#_c_184_n 0.00993078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_228_297#_c_187_n 0.00165371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_228_297#_c_194_n 0.00826359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_257_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_53 VPB N_VPWR_c_258_n 0.0557758f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_54 VPB N_VPWR_c_259_n 0.0121493f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_55 VPB N_VPWR_c_260_n 0.0117975f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_56 VPB N_VPWR_c_261_n 0.0464637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_262_n 0.0435097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_263_n 0.0268687f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_264_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_256_n 0.0664461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_X_c_297_n 0.00129626f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_62 N_B_N_c_65_n N_A_27_53#_c_90_n 0.00538165f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_63 N_B_N_M1000_g N_A_27_53#_c_91_n 0.00300496f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_64 N_B_N_M1000_g N_A_27_53#_c_92_n 0.0268605f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_65 B_N N_A_27_53#_c_92_n 0.0162285f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B_N_c_65_n N_A_27_53#_c_92_n 0.00104773f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_67 B_N N_A_27_53#_c_93_n 0.0259349f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_68 N_B_N_c_65_n N_A_27_53#_c_93_n 0.00813455f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_69 N_B_N_c_66_n N_A_27_53#_c_97_n 0.00610416f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B_N_c_65_n N_A_27_53#_c_97_n 0.00648588f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_71 N_B_N_c_66_n A 0.00227571f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_B_N_c_65_n A 2.63734e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_73 N_B_N_c_66_n N_A_228_297#_c_194_n 0.00166429f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B_N_c_66_n N_VPWR_c_258_n 0.00877297f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 B_N N_VPWR_c_258_n 0.0210621f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_B_N_c_65_n N_VPWR_c_258_n 0.00556766f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_77 N_B_N_c_66_n N_VPWR_c_262_n 0.00298464f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B_N_c_66_n N_VPWR_c_256_n 0.0037574f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B_N_M1000_g N_VGND_c_322_n 0.00413798f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_80 N_B_N_M1000_g N_VGND_c_323_n 0.00505351f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_81 N_B_N_M1000_g N_VGND_c_325_n 0.00754515f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_82 N_A_27_53#_c_90_n N_A_c_135_n 0.010421f $X=1.5 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_83 N_A_27_53#_M1001_g N_A_M1009_g 0.0226511f $X=1.465 $Y=0.475 $X2=0 $Y2=0
cc_84 N_A_27_53#_c_90_n N_A_c_133_n 0.0279021f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_27_53#_c_94_n N_A_c_133_n 0.00139464f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_27_53#_c_90_n N_A_M1005_g 0.035907f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_27_53#_c_90_n A 0.00205903f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_27_53#_c_97_n A 0.0124285f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_89 N_A_27_53#_c_90_n N_A_228_297#_c_196_n 0.0126327f $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_90 N_A_27_53#_M1001_g N_A_228_297#_c_186_n 0.00449357f $X=1.465 $Y=0.475
+ $X2=0 $Y2=0
cc_91 N_A_27_53#_c_90_n N_A_228_297#_c_186_n 3.06238e-19 $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_92 N_A_27_53#_c_90_n N_A_228_297#_c_194_n 0.0155597f $X=1.5 $Y=1.41 $X2=0
+ $Y2=0
cc_93 N_A_27_53#_c_97_n N_A_228_297#_c_194_n 0.0257664f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_94 N_A_27_53#_c_94_n N_A_228_297#_c_194_n 0.0267679f $X=1.265 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_27_53#_c_97_n N_VPWR_c_258_n 0.0192564f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_96 N_A_27_53#_M1001_g N_VGND_c_317_n 0.00555245f $X=1.465 $Y=0.475 $X2=0
+ $Y2=0
cc_97 N_A_27_53#_c_91_n N_VGND_c_322_n 0.0196296f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_27_53#_c_92_n N_VGND_c_322_n 0.00299761f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_99 N_A_27_53#_M1001_g N_VGND_c_323_n 0.00367484f $X=1.465 $Y=0.475 $X2=0
+ $Y2=0
cc_100 N_A_27_53#_c_90_n N_VGND_c_323_n 0.004553f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_27_53#_c_92_n N_VGND_c_323_n 0.0210226f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_102 N_A_27_53#_c_94_n N_VGND_c_323_n 0.0194332f $X=1.265 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_27_53#_M1001_g N_VGND_c_325_n 0.0113859f $X=1.465 $Y=0.475 $X2=0
+ $Y2=0
cc_104 N_A_27_53#_c_91_n N_VGND_c_325_n 0.0119774f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_105 N_A_27_53#_c_92_n N_VGND_c_325_n 0.00606676f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_A_228_297#_c_188_n 0.0169236f $X=1.91 $Y=1.695 $X2=0 $Y2=0
cc_107 N_A_M1009_g N_A_228_297#_c_180_n 0.0194393f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_108 N_A_c_133_n N_A_228_297#_c_180_n 9.15481e-19 $X=1.91 $Y=1.06 $X2=0 $Y2=0
cc_109 N_A_c_133_n N_A_228_297#_c_182_n 0.0232287f $X=1.91 $Y=1.06 $X2=0 $Y2=0
cc_110 N_A_c_136_n N_A_228_297#_c_182_n 0.00275812f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_135_n N_A_228_297#_c_196_n 7.85782e-19 $X=1.81 $Y=2.34 $X2=0 $Y2=0
cc_112 N_A_M1005_g N_A_228_297#_c_196_n 0.019663f $X=1.91 $Y=1.695 $X2=0 $Y2=0
cc_113 A N_A_228_297#_c_196_n 0.0127859f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_114 N_A_M1009_g N_A_228_297#_c_185_n 0.0142024f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_115 N_A_c_133_n N_A_228_297#_c_185_n 0.00160903f $X=1.91 $Y=1.06 $X2=0 $Y2=0
cc_116 N_A_M1009_g N_A_228_297#_c_187_n 0.0025127f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_117 N_A_c_133_n N_A_228_297#_c_187_n 0.002704f $X=1.91 $Y=1.06 $X2=0 $Y2=0
cc_118 N_A_c_136_n N_A_228_297#_c_187_n 0.00164174f $X=1.91 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_M1005_g N_A_228_297#_c_187_n 0.00161078f $X=1.91 $Y=1.695 $X2=0 $Y2=0
cc_120 N_A_c_135_n N_A_228_297#_c_194_n 9.83498e-19 $X=1.81 $Y=2.34 $X2=0 $Y2=0
cc_121 N_A_M1005_g N_A_228_297#_c_194_n 0.00115522f $X=1.91 $Y=1.695 $X2=0 $Y2=0
cc_122 A N_A_228_297#_c_194_n 0.0344364f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_123 N_A_c_140_n N_A_228_297#_c_194_n 0.00119166f $X=1.22 $Y=2.28 $X2=0 $Y2=0
cc_124 A N_VPWR_c_258_n 0.0258924f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_125 N_A_c_140_n N_VPWR_c_258_n 9.3247e-19 $X=1.22 $Y=2.28 $X2=0 $Y2=0
cc_126 N_A_M1005_g N_VPWR_c_259_n 0.00443253f $X=1.91 $Y=1.695 $X2=0 $Y2=0
cc_127 N_A_c_138_n N_VPWR_c_259_n 0.00487993f $X=1.91 $Y=2.34 $X2=0 $Y2=0
cc_128 A N_VPWR_c_259_n 0.0216404f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_129 A N_VPWR_c_262_n 0.0634852f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_130 N_A_c_140_n N_VPWR_c_262_n 0.0240252f $X=1.22 $Y=2.28 $X2=0 $Y2=0
cc_131 A N_VPWR_c_256_n 0.0467241f $X=1.115 $Y=2.125 $X2=0 $Y2=0
cc_132 N_A_c_140_n N_VPWR_c_256_n 0.0331114f $X=1.22 $Y=2.28 $X2=0 $Y2=0
cc_133 N_A_M1009_g N_VGND_c_317_n 0.00403348f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_134 N_A_M1009_g N_VGND_c_318_n 0.00431669f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_135 N_A_M1009_g N_VGND_c_325_n 0.00587083f $X=1.885 $Y=0.475 $X2=0 $Y2=0
cc_136 N_A_228_297#_c_196_n N_VPWR_M1005_d 0.00651861f $X=2.27 $Y=1.58 $X2=0
+ $Y2=0
cc_137 N_A_228_297#_c_188_n N_VPWR_c_259_n 0.00482583f $X=2.45 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_228_297#_c_182_n N_VPWR_c_259_n 3.01556e-19 $X=2.55 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_228_297#_c_196_n N_VPWR_c_259_n 0.0198977f $X=2.27 $Y=1.58 $X2=0
+ $Y2=0
cc_140 N_A_228_297#_c_194_n N_VPWR_c_259_n 0.00230358f $X=1.245 $Y=1.58 $X2=0
+ $Y2=0
cc_141 N_A_228_297#_c_191_n N_VPWR_c_261_n 0.00799675f $X=3.11 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_228_297#_c_188_n N_VPWR_c_263_n 0.00702461f $X=2.45 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_228_297#_c_191_n N_VPWR_c_263_n 0.00567349f $X=3.11 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_228_297#_c_188_n N_VPWR_c_256_n 0.0141931f $X=2.45 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_228_297#_c_191_n N_VPWR_c_256_n 0.0107563f $X=3.11 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_228_297#_c_196_n A_318_297# 0.003951f $X=2.27 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_228_297#_c_188_n N_X_c_297_n 0.0124805f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_228_297#_c_180_n N_X_c_297_n 0.00779986f $X=2.475 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_228_297#_c_181_n N_X_c_297_n 0.0231948f $X=3.01 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_228_297#_c_182_n N_X_c_297_n 7.69592e-19 $X=2.55 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_228_297#_c_191_n N_X_c_297_n 0.0234401f $X=3.11 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_228_297#_c_183_n N_X_c_297_n 0.013198f $X=3.135 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_228_297#_c_184_n N_X_c_297_n 0.0220689f $X=3.11 $Y=1.202 $X2=0 $Y2=0
cc_154 N_A_228_297#_c_196_n N_X_c_297_n 0.00800109f $X=2.27 $Y=1.58 $X2=0 $Y2=0
cc_155 N_A_228_297#_c_185_n N_X_c_297_n 0.00800095f $X=2.27 $Y=0.74 $X2=0 $Y2=0
cc_156 N_A_228_297#_c_187_n N_X_c_297_n 0.0279739f $X=2.355 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_228_297#_c_185_n N_VGND_M1009_d 0.00755106f $X=2.27 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_A_228_297#_c_187_n N_VGND_M1009_d 7.65498e-19 $X=2.355 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_228_297#_c_243_p N_VGND_c_317_n 0.00846569f $X=1.675 $Y=0.47 $X2=0
+ $Y2=0
cc_160 N_A_228_297#_c_185_n N_VGND_c_317_n 0.0035399f $X=2.27 $Y=0.74 $X2=0
+ $Y2=0
cc_161 N_A_228_297#_c_180_n N_VGND_c_318_n 0.00510929f $X=2.475 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_228_297#_c_182_n N_VGND_c_318_n 4.00709e-19 $X=2.55 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_228_297#_c_185_n N_VGND_c_318_n 0.0245048f $X=2.27 $Y=0.74 $X2=0
+ $Y2=0
cc_164 N_A_228_297#_c_183_n N_VGND_c_320_n 0.0102136f $X=3.135 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_228_297#_c_180_n N_VGND_c_321_n 0.00543382f $X=2.475 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_228_297#_c_183_n N_VGND_c_321_n 0.00521195f $X=3.135 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_228_297#_c_185_n N_VGND_c_321_n 0.00104987f $X=2.27 $Y=0.74 $X2=0
+ $Y2=0
cc_168 N_A_228_297#_c_180_n N_VGND_c_325_n 0.0105119f $X=2.475 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_228_297#_c_183_n N_VGND_c_325_n 0.0104625f $X=3.135 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_228_297#_c_243_p N_VGND_c_325_n 0.00625722f $X=1.675 $Y=0.47 $X2=0
+ $Y2=0
cc_171 N_A_228_297#_c_185_n N_VGND_c_325_n 0.0104309f $X=2.27 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_256_n N_X_M1002_s 0.0125882f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_261_n N_X_c_297_n 0.0741971f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_174 N_VPWR_c_263_n N_X_c_297_n 0.0201856f $X=3.285 $Y=2.72 $X2=0 $Y2=0
cc_175 N_VPWR_c_256_n N_X_c_297_n 0.0118397f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_176 N_VPWR_c_261_n N_VGND_c_320_n 0.00980968f $X=3.37 $Y=1.65 $X2=0 $Y2=0
cc_177 N_X_c_297_n N_VGND_c_320_n 0.0376908f $X=2.875 $Y=0.59 $X2=0 $Y2=0
cc_178 N_X_c_297_n N_VGND_c_321_n 0.00990218f $X=2.875 $Y=0.59 $X2=0 $Y2=0
cc_179 N_X_M1006_s N_VGND_c_325_n 0.012724f $X=2.55 $Y=0.235 $X2=0 $Y2=0
cc_180 N_X_c_297_n N_VGND_c_325_n 0.0109165f $X=2.875 $Y=0.59 $X2=0 $Y2=0
