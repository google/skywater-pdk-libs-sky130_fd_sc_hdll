* NGSPICE file created from sky130_fd_sc_hdll__nand2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nand2_1 A B VGND VNB VPB VPWR Y
M1000 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=5.4e+11p ps=5.08e+06u
M1001 Y A a_123_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.755e+11p ps=1.84e+06u
M1002 a_123_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1003 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

