* File: sky130_fd_sc_hdll__nand3_1.pxi.spice
* Created: Wed Sep  2 08:37:33 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3_1%C N_C_c_37_n N_C_M1003_g N_C_c_34_n N_C_M1005_g
+ C C N_C_c_36_n PM_SKY130_FD_SC_HDLL__NAND3_1%C
x_PM_SKY130_FD_SC_HDLL__NAND3_1%B N_B_c_63_n N_B_M1001_g N_B_c_64_n N_B_M1000_g
+ B B PM_SKY130_FD_SC_HDLL__NAND3_1%B
x_PM_SKY130_FD_SC_HDLL__NAND3_1%A N_A_c_96_n N_A_M1002_g N_A_c_97_n N_A_M1004_g
+ A A PM_SKY130_FD_SC_HDLL__NAND3_1%A
x_PM_SKY130_FD_SC_HDLL__NAND3_1%VPWR N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_c_123_n N_VPWR_c_124_n N_VPWR_c_125_n N_VPWR_c_126_n VPWR
+ N_VPWR_c_127_n N_VPWR_c_122_n N_VPWR_c_129_n
+ PM_SKY130_FD_SC_HDLL__NAND3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3_1%Y N_Y_M1002_d N_Y_M1003_d N_Y_M1004_d
+ N_Y_c_158_n N_Y_c_166_n N_Y_c_155_n N_Y_c_156_n N_Y_c_153_n N_Y_c_163_n
+ N_Y_c_154_n N_Y_c_175_n Y PM_SKY130_FD_SC_HDLL__NAND3_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND3_1%VGND N_VGND_M1005_s N_VGND_c_213_n
+ N_VGND_c_214_n VGND N_VGND_c_215_n N_VGND_c_216_n
+ PM_SKY130_FD_SC_HDLL__NAND3_1%VGND
cc_1 VNB N_C_c_34_n 0.0187992f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB C 0.00980239f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_C_c_36_n 0.0484134f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_c_63_n 0.0167612f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_c_64_n 0.0243902f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B 0.00302998f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_7 VNB N_A_c_96_n 0.0231188f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A_c_97_n 0.0358518f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB A 0.0128127f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_10 VNB N_VPWR_c_122_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_153_n 0.00248617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_154_n 0.0230706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_213_n 0.00994635f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB N_VGND_c_214_n 0.0188667f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_VGND_c_215_n 0.0509608f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_16 VNB N_VGND_c_216_n 0.155149f $X=-0.19 $Y=-0.24 $X2=0.22 $Y2=0.85
cc_17 VPB N_C_c_37_n 0.020812f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_18 VPB C 0.00203753f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_19 VPB N_C_c_36_n 0.0193798f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_20 VPB N_B_c_64_n 0.0274153f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_21 VPB B 0.00216641f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_22 VPB N_A_c_97_n 0.0376718f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_23 VPB A 0.00161459f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_24 VPB N_VPWR_c_123_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_25 VPB N_VPWR_c_124_n 0.0433665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_VPWR_c_125_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_27 VPB N_VPWR_c_126_n 0.00503731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_VPWR_c_127_n 0.0288381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_122_n 0.0561169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_129_n 0.00439477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_Y_c_155_n 0.00752809f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=0.85
cc_32 VPB N_Y_c_156_n 0.0317329f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_33 VPB N_Y_c_153_n 0.00166906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 N_C_c_34_n N_B_c_63_n 0.029569f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_35 N_C_c_37_n N_B_c_64_n 0.00921322f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_36 N_C_c_36_n N_B_c_64_n 0.029569f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_37 N_C_c_34_n B 5.08222e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_38 N_C_c_37_n N_VPWR_c_124_n 0.00777002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_39 C N_VPWR_c_124_n 0.0188755f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_40 N_C_c_36_n N_VPWR_c_124_n 0.00239203f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_41 N_C_c_37_n N_VPWR_c_125_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_42 N_C_c_37_n N_VPWR_c_122_n 0.0109312f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_43 N_C_c_37_n N_Y_c_158_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_C_c_37_n N_Y_c_153_n 0.00437338f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_45 N_C_c_34_n N_Y_c_153_n 0.0134206f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_46 C N_Y_c_153_n 0.0391002f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_47 N_C_c_36_n N_Y_c_153_n 0.0144417f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_48 N_C_c_37_n N_Y_c_163_n 0.0024721f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_49 N_C_c_34_n Y 0.0101899f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_50 C N_VGND_M1005_s 0.00404081f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_51 N_C_c_34_n N_VGND_c_214_n 0.00536202f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_52 C N_VGND_c_214_n 0.0188142f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_53 N_C_c_36_n N_VGND_c_214_n 0.00148721f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_54 N_C_c_34_n N_VGND_c_215_n 0.00463936f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_55 N_C_c_34_n N_VGND_c_216_n 0.00880407f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_56 C N_VGND_c_216_n 8.97811e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B_c_63_n N_A_c_96_n 0.0265056f $X=0.94 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_58 B N_A_c_96_n 0.00746207f $X=1.075 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_59 N_B_c_64_n N_A_c_97_n 0.0520177f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B_c_64_n A 3.0004e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_61 B A 0.0246683f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_62 N_B_c_64_n N_VPWR_c_125_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B_c_64_n N_VPWR_c_126_n 0.00555837f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B_c_64_n N_VPWR_c_122_n 0.0120301f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_65 N_B_c_64_n N_Y_c_158_n 0.0109123f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_66 N_B_c_64_n N_Y_c_166_n 0.0154187f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_67 B N_Y_c_166_n 0.0264942f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_68 N_B_c_64_n N_Y_c_156_n 6.35212e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B_c_63_n N_Y_c_153_n 0.00959072f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B_c_64_n N_Y_c_153_n 0.00191844f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_71 B N_Y_c_153_n 0.04324f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_72 N_B_c_64_n N_Y_c_163_n 0.00129054f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B_c_63_n N_Y_c_154_n 0.00100699f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_74 B N_Y_c_154_n 0.00376447f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_75 N_B_c_63_n N_Y_c_175_n 0.0187176f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_76 N_B_c_64_n N_Y_c_175_n 6.51204e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_77 B N_Y_c_175_n 0.0247727f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_78 N_B_c_63_n N_VGND_c_215_n 0.00357877f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_c_63_n N_VGND_c_216_n 0.00557664f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_80 B A_203_47# 0.00381115f $X=1.075 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_81 N_A_c_97_n N_VPWR_c_126_n 0.00849087f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_97_n N_VPWR_c_127_n 0.00597712f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_97_n N_VPWR_c_122_n 0.0113384f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_97_n N_Y_c_158_n 6.80127e-19 $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_97_n N_Y_c_166_n 0.0125212f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_86 A N_Y_c_166_n 0.00282261f $X=1.54 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A_c_97_n N_Y_c_155_n 0.0076545f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_88 A N_Y_c_155_n 0.0288843f $X=1.54 $Y=1.105 $X2=0 $Y2=0
cc_89 N_A_c_97_n N_Y_c_156_n 0.0133425f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_96_n N_Y_c_154_n 0.00678247f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_97_n N_Y_c_154_n 0.00682953f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_92 A N_Y_c_154_n 0.0284541f $X=1.54 $Y=1.105 $X2=0 $Y2=0
cc_93 N_A_c_96_n N_Y_c_175_n 0.0156479f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_94 A N_Y_c_175_n 0.00150996f $X=1.54 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_c_96_n N_VGND_c_215_n 0.00359354f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_c_96_n N_VGND_c_216_n 0.00682647f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_97 N_VPWR_c_122_n N_Y_M1003_d 0.00231261f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_98 N_VPWR_c_122_n N_Y_M1004_d 0.00217517f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_124_n N_Y_c_158_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_100 N_VPWR_c_125_n N_Y_c_158_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_101 N_VPWR_c_126_n N_Y_c_158_n 0.0394373f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_102 N_VPWR_c_122_n N_Y_c_158_n 0.0140101f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_103 N_VPWR_M1000_d N_Y_c_166_n 0.00652763f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_104 N_VPWR_c_126_n N_Y_c_166_n 0.0185497f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_105 N_VPWR_c_126_n N_Y_c_156_n 0.0480927f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_106 N_VPWR_c_127_n N_Y_c_156_n 0.0244686f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_107 N_VPWR_c_122_n N_Y_c_156_n 0.0141694f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_108 N_VPWR_c_124_n N_Y_c_163_n 0.0137498f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_109 Y N_VGND_c_214_n 0.0258822f $X=0.59 $Y=0.425 $X2=0 $Y2=0
cc_110 N_Y_c_154_n N_VGND_c_215_n 0.0242653f $X=1.73 $Y=0.38 $X2=0 $Y2=0
cc_111 N_Y_c_175_n N_VGND_c_215_n 0.0452714f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_112 Y N_VGND_c_215_n 0.0140166f $X=0.59 $Y=0.425 $X2=0 $Y2=0
cc_113 N_Y_M1002_d N_VGND_c_216_n 0.00250309f $X=1.545 $Y=0.235 $X2=0 $Y2=0
cc_114 N_Y_c_154_n N_VGND_c_216_n 0.0142861f $X=1.73 $Y=0.38 $X2=0 $Y2=0
cc_115 N_Y_c_175_n N_VGND_c_216_n 0.0278897f $X=1.515 $Y=0.425 $X2=0 $Y2=0
cc_116 Y N_VGND_c_216_n 0.00849186f $X=0.59 $Y=0.425 $X2=0 $Y2=0
cc_117 N_Y_c_153_n A_119_47# 0.00297272f $X=0.63 $Y=1.495 $X2=-0.19 $Y2=-0.24
cc_118 N_Y_c_175_n A_119_47# 0.0031671f $X=1.515 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_119 Y A_119_47# 9.09492e-19 $X=0.59 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_120 N_Y_c_175_n A_203_47# 0.00729541f $X=1.515 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_121 N_VGND_c_216_n A_119_47# 0.00216819f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
cc_122 N_VGND_c_216_n A_203_47# 0.00305172f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
