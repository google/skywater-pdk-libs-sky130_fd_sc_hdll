* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
X0 a_1011_47# a_27_47# a_1121_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 a_1568_413# a_1667_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 a_608_369# SCE a_721_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND a_319_47# a_517_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1474_413# a_203_47# a_1568_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 a_1127_47# a_1189_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_1189_183# a_27_47# a_1474_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X8 VPWR a_1667_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_319_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_608_369# a_27_47# a_1011_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X11 a_1189_183# a_203_47# a_1474_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 VGND a_1667_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND a_1667_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_504_369# D a_608_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X15 a_702_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X16 a_517_47# D a_608_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 Q a_1667_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 Q a_1667_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_27_47# a_203_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_721_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1474_413# a_27_47# a_1625_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X22 a_1011_47# a_203_47# a_1127_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 VPWR SCE a_504_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X24 a_1667_315# a_1474_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_1625_47# a_1667_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_1667_315# a_1474_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR a_27_47# a_203_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X28 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 Q a_1667_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 VPWR a_1667_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 Q a_1667_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VPWR a_1011_47# a_1189_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=180000u
X33 a_1121_413# a_1189_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X34 VGND a_1011_47# a_1189_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X35 a_319_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X36 a_608_369# a_319_47# a_702_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X37 a_608_369# a_203_47# a_1011_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
