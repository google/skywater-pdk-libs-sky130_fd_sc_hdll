# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a32o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.680000 1.075000 5.575000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.635000 1.075000 4.430000 1.325000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.410000 1.075000 3.405000 1.295000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.120000 1.075000 7.140000 1.625000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.440000 1.075000 8.170000 1.295000 ;
        RECT 7.440000 1.295000 7.635000 1.635000 ;
    END
  END B2
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.635000 1.755000 0.805000 ;
        RECT 0.120000 0.805000 0.340000 1.495000 ;
        RECT 0.120000 1.495000 1.755000 1.665000 ;
        RECT 0.645000 0.255000 0.815000 0.635000 ;
        RECT 0.645000 1.665000 0.815000 2.465000 ;
        RECT 1.585000 0.255000 1.755000 0.635000 ;
        RECT 1.585000 1.665000 1.755000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.095000  1.915000 0.425000 2.635000 ;
      RECT 0.620000  0.995000 2.170000 1.325000 ;
      RECT 0.985000  0.085000 1.365000 0.465000 ;
      RECT 0.985000  1.915000 1.365000 2.635000 ;
      RECT 1.925000  0.085000 2.305000 0.465000 ;
      RECT 1.925000  1.915000 2.305000 2.635000 ;
      RECT 1.950000  1.325000 2.170000 1.495000 ;
      RECT 1.950000  1.495000 5.950000 1.665000 ;
      RECT 2.525000  0.255000 2.695000 0.655000 ;
      RECT 2.525000  0.655000 4.235000 0.825000 ;
      RECT 2.525000  1.915000 5.565000 2.085000 ;
      RECT 2.525000  2.085000 2.695000 2.465000 ;
      RECT 2.865000  0.085000 3.245000 0.465000 ;
      RECT 2.865000  2.255000 3.245000 2.635000 ;
      RECT 3.435000  0.295000 5.645000 0.465000 ;
      RECT 3.515000  2.085000 3.685000 2.465000 ;
      RECT 3.855000  2.255000 4.235000 2.635000 ;
      RECT 4.455000  2.085000 4.625000 2.465000 ;
      RECT 4.795000  0.635000 6.735000 0.805000 ;
      RECT 4.795000  2.255000 5.175000 2.635000 ;
      RECT 5.395000  2.085000 5.565000 2.255000 ;
      RECT 5.395000  2.255000 8.185000 2.425000 ;
      RECT 5.780000  0.805000 5.950000 1.495000 ;
      RECT 5.780000  1.665000 5.950000 1.905000 ;
      RECT 5.780000  1.905000 6.510000 1.915000 ;
      RECT 5.780000  1.915000 7.715000 2.075000 ;
      RECT 5.930000  0.295000 7.165000 0.465000 ;
      RECT 6.445000  2.075000 7.715000 2.085000 ;
      RECT 6.995000  0.255000 7.165000 0.295000 ;
      RECT 6.995000  0.465000 7.165000 0.645000 ;
      RECT 6.995000  0.645000 8.105000 0.815000 ;
      RECT 7.335000  0.085000 7.715000 0.465000 ;
      RECT 7.935000  0.255000 8.105000 0.645000 ;
      RECT 7.935000  1.755000 8.185000 2.255000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32o_4
