* File: sky130_fd_sc_hdll__nor2b_2.pxi.spice
* Created: Wed Sep  2 08:39:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%A N_A_c_60_n N_A_M1004_g N_A_c_64_n N_A_M1000_g
+ N_A_c_65_n N_A_M1005_g N_A_c_61_n N_A_M1008_g A N_A_c_63_n A
+ PM_SKY130_FD_SC_HDLL__NOR2B_2%A
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%A_271_21# N_A_271_21#_M1009_s
+ N_A_271_21#_M1002_s N_A_271_21#_c_97_n N_A_271_21#_M1006_g N_A_271_21#_c_105_n
+ N_A_271_21#_M1001_g N_A_271_21#_c_98_n N_A_271_21#_M1007_g N_A_271_21#_c_106_n
+ N_A_271_21#_M1003_g N_A_271_21#_c_99_n N_A_271_21#_c_100_n N_A_271_21#_c_101_n
+ N_A_271_21#_c_102_n N_A_271_21#_c_103_n N_A_271_21#_c_104_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_2%A_271_21#
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%B_N N_B_N_M1009_g N_B_N_c_167_n N_B_N_c_168_n
+ N_B_N_M1002_g N_B_N_c_162_n N_B_N_c_163_n B_N B_N B_N N_B_N_c_166_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_2%B_N
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1005_s N_A_27_297#_M1003_d N_A_27_297#_c_194_n
+ N_A_27_297#_c_195_n N_A_27_297#_c_196_n N_A_27_297#_c_197_n
+ N_A_27_297#_c_216_p N_A_27_297#_c_206_n N_A_27_297#_c_198_n
+ N_A_27_297#_c_199_n PM_SKY130_FD_SC_HDLL__NOR2B_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%VPWR N_VPWR_M1000_d N_VPWR_M1002_d
+ N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n VPWR N_VPWR_c_237_n
+ N_VPWR_c_238_n N_VPWR_c_233_n VPWR PM_SKY130_FD_SC_HDLL__NOR2B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%Y N_Y_M1004_d N_Y_M1006_s N_Y_M1001_s
+ N_Y_c_278_n N_Y_c_273_n N_Y_c_274_n N_Y_c_275_n N_Y_c_276_n Y N_Y_c_286_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR2B_2%VGND N_VGND_M1004_s N_VGND_M1008_s
+ N_VGND_M1007_d N_VGND_M1009_d N_VGND_c_318_n N_VGND_c_319_n N_VGND_c_320_n
+ N_VGND_c_321_n N_VGND_c_322_n N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n
+ N_VGND_c_326_n VGND N_VGND_c_327_n N_VGND_c_328_n N_VGND_c_329_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_2%VGND
cc_1 VNB N_A_c_60_n 0.0225874f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_61_n 0.0169958f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB A 0.00473824f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_A_c_63_n 0.0481664f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_A_271_21#_c_97_n 0.0165539f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_6 VNB N_A_271_21#_c_98_n 0.0204716f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_7 VNB N_A_271_21#_c_99_n 0.0348031f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_8 VNB N_A_271_21#_c_100_n 0.0130416f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_9 VNB N_A_271_21#_c_101_n 0.0348055f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_271_21#_c_102_n 0.00748545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_271_21#_c_103_n 0.00139127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_271_21#_c_104_n 0.00216451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B_N_c_162_n 0.00266859f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_14 VNB N_B_N_c_163_n 0.0350842f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.56
cc_15 VNB B_N 0.0138864f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB B_N 0.00109931f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_17 VNB N_B_N_c_166_n 0.0442166f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.17
cc_18 VNB N_VPWR_c_233_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_273_n 0.0032419f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_274_n 0.00281417f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_21 VNB N_Y_c_275_n 0.00188026f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_22 VNB N_Y_c_276_n 0.00282996f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_23 VNB N_VGND_c_318_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_24 VNB N_VGND_c_319_n 0.0350705f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_25 VNB N_VGND_c_320_n 0.0198175f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.202
cc_26 VNB N_VGND_c_321_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_27 VNB N_VGND_c_322_n 0.00601139f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.17
cc_28 VNB N_VGND_c_323_n 0.0147615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_324_n 0.0315251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_325_n 0.0200006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_326_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_327_n 0.02876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_328_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_329_n 0.229865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_c_64_n 0.0201091f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_36 VPB N_A_c_65_n 0.016004f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_37 VPB N_A_c_63_n 0.0226591f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_38 VPB N_A_271_21#_c_105_n 0.0164039f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_39 VPB N_A_271_21#_c_106_n 0.0194069f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_40 VPB N_A_271_21#_c_99_n 0.0229536f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_41 VPB N_A_271_21#_c_101_n 0.0128045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_271_21#_c_103_n 0.0189329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_N_c_167_n 0.0376757f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_44 VPB N_B_N_c_168_n 0.0321748f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_45 VPB N_B_N_c_163_n 0.007858f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_46 VPB B_N 0.0372721f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_47 VPB N_A_27_297#_c_194_n 0.0151236f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_48 VPB N_A_27_297#_c_195_n 0.0318598f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_49 VPB N_A_27_297#_c_196_n 0.00226265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_297#_c_197_n 0.00325848f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_51 VPB N_A_27_297#_c_198_n 0.00215223f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_52 VPB N_A_27_297#_c_199_n 0.0115428f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.17
cc_53 VPB N_VPWR_c_234_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_54 VPB N_VPWR_c_235_n 0.0144505f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_55 VPB N_VPWR_c_236_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_56 VPB N_VPWR_c_237_n 0.060023f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_57 VPB N_VPWR_c_238_n 0.0238232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_233_n 0.0570632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_Y_c_275_n 0.0027542f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_60 N_A_c_61_n N_A_271_21#_c_97_n 0.0235436f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A_c_65_n N_A_271_21#_c_105_n 0.00943295f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_62 A N_A_271_21#_c_99_n 0.00236897f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_c_63_n N_A_271_21#_c_99_n 0.0235436f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_64 N_A_c_64_n N_A_27_297#_c_196_n 0.0191894f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_65_n N_A_27_297#_c_196_n 0.0170544f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_66 A N_A_27_297#_c_196_n 0.0442545f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_c_63_n N_A_27_297#_c_196_n 0.00820898f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_68 A N_A_27_297#_c_197_n 0.0141395f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A_c_64_n N_VPWR_c_234_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_65_n N_VPWR_c_234_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_c_65_n N_VPWR_c_237_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_64_n N_VPWR_c_238_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_c_64_n N_VPWR_c_233_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_65_n N_VPWR_c_233_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_60_n N_Y_c_278_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_76 N_A_c_61_n N_Y_c_273_n 0.0100733f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_77 A N_Y_c_273_n 0.0236938f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A_c_60_n N_Y_c_274_n 0.00243049f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_79 A N_Y_c_274_n 0.0324228f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_c_63_n N_Y_c_274_n 0.00480108f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_81 A N_Y_c_275_n 0.011141f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_63_n N_Y_c_275_n 7.60995e-19 $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_83 N_A_c_61_n N_Y_c_286_n 5.27946e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_c_60_n N_VGND_c_319_n 0.0047492f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_c_60_n N_VGND_c_320_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_c_61_n N_VGND_c_320_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_c_61_n N_VGND_c_321_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_c_60_n N_VGND_c_329_n 0.0107167f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_c_61_n N_VGND_c_329_n 0.00615622f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_90 N_A_271_21#_c_103_n N_B_N_c_168_n 0.0117794f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_91 N_A_271_21#_c_101_n N_B_N_c_162_n 4.42171e-19 $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_271_21#_c_102_n N_B_N_c_162_n 6.45958e-19 $X=2.68 $Y=0.68 $X2=0 $Y2=0
cc_93 N_A_271_21#_c_103_n N_B_N_c_162_n 0.00215764f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_94 N_A_271_21#_c_104_n N_B_N_c_162_n 0.0142805f $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_271_21#_c_101_n N_B_N_c_163_n 0.00497665f $X=2.24 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_271_21#_c_103_n N_B_N_c_163_n 0.0159974f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_97 N_A_271_21#_c_104_n N_B_N_c_163_n 7.92131e-19 $X=2.68 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_271_21#_c_103_n B_N 0.0248956f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_99 N_A_271_21#_c_102_n N_B_N_c_166_n 0.014856f $X=2.68 $Y=0.68 $X2=0 $Y2=0
cc_100 N_A_271_21#_c_105_n N_A_27_297#_c_197_n 4.00176e-19 $X=1.455 $Y=1.41
+ $X2=0 $Y2=0
cc_101 N_A_271_21#_c_105_n N_A_27_297#_c_206_n 0.0143578f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_102 N_A_271_21#_c_106_n N_A_27_297#_c_206_n 0.0143578f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_271_21#_c_103_n N_A_27_297#_c_198_n 0.00984622f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_104 N_A_271_21#_c_106_n N_A_27_297#_c_199_n 9.96901e-19 $X=1.925 $Y=1.41
+ $X2=0 $Y2=0
cc_105 N_A_271_21#_c_100_n N_A_27_297#_c_199_n 0.0177877f $X=2.595 $Y=1.16 $X2=0
+ $Y2=0
cc_106 N_A_271_21#_c_101_n N_A_27_297#_c_199_n 0.00812764f $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_271_21#_c_103_n N_A_27_297#_c_199_n 0.0479968f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_108 N_A_271_21#_c_105_n N_VPWR_c_237_n 0.00429453f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_109 N_A_271_21#_c_106_n N_VPWR_c_237_n 0.00429453f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_110 N_A_271_21#_c_103_n N_VPWR_c_237_n 0.0114468f $X=2.68 $Y=2.28 $X2=0 $Y2=0
cc_111 N_A_271_21#_M1002_s N_VPWR_c_233_n 0.0123591f $X=2.555 $Y=2.065 $X2=0
+ $Y2=0
cc_112 N_A_271_21#_c_105_n N_VPWR_c_233_n 0.00609021f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_113 N_A_271_21#_c_106_n N_VPWR_c_233_n 0.00734734f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_114 N_A_271_21#_c_103_n N_VPWR_c_233_n 0.00645481f $X=2.68 $Y=2.28 $X2=0
+ $Y2=0
cc_115 N_A_271_21#_c_97_n N_Y_c_273_n 0.0120386f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_271_21#_c_97_n N_Y_c_275_n 0.00257856f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_271_21#_c_105_n N_Y_c_275_n 0.00130217f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_271_21#_c_98_n N_Y_c_275_n 0.00274923f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_271_21#_c_106_n N_Y_c_275_n 0.00130282f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_271_21#_c_99_n N_Y_c_275_n 0.036848f $X=2.025 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_271_21#_c_100_n N_Y_c_275_n 0.00935835f $X=2.595 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_271_21#_c_97_n N_Y_c_276_n 0.00208031f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_271_21#_c_98_n N_Y_c_276_n 0.00368409f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_271_21#_c_97_n N_Y_c_286_n 0.00639345f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_271_21#_c_98_n N_Y_c_286_n 0.00600712f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_271_21#_c_97_n N_VGND_c_321_n 0.00268723f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_127 N_A_271_21#_c_98_n N_VGND_c_322_n 0.00656994f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_271_21#_c_100_n N_VGND_c_322_n 0.0129839f $X=2.595 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_271_21#_c_101_n N_VGND_c_322_n 0.00429275f $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_271_21#_c_102_n N_VGND_c_322_n 0.0192831f $X=2.68 $Y=0.68 $X2=0 $Y2=0
cc_131 N_A_271_21#_c_102_n N_VGND_c_324_n 0.0154184f $X=2.68 $Y=0.68 $X2=0 $Y2=0
cc_132 N_A_271_21#_c_97_n N_VGND_c_325_n 0.00423334f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_133 N_A_271_21#_c_98_n N_VGND_c_325_n 0.00541359f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_271_21#_c_102_n N_VGND_c_327_n 0.00542302f $X=2.68 $Y=0.68 $X2=0
+ $Y2=0
cc_135 N_A_271_21#_c_97_n N_VGND_c_329_n 0.00587047f $X=1.43 $Y=0.995 $X2=0
+ $Y2=0
cc_136 N_A_271_21#_c_98_n N_VGND_c_329_n 0.0110773f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_271_21#_c_102_n N_VGND_c_329_n 0.00578545f $X=2.68 $Y=0.68 $X2=0
+ $Y2=0
cc_138 N_B_N_c_168_n N_A_27_297#_c_198_n 4.49502e-19 $X=3.075 $Y=1.99 $X2=0
+ $Y2=0
cc_139 B_N N_VPWR_c_235_n 0.00159942f $X=3.32 $Y=1.445 $X2=0 $Y2=0
cc_140 N_B_N_c_168_n N_VPWR_c_236_n 0.00479105f $X=3.075 $Y=1.99 $X2=0 $Y2=0
cc_141 B_N N_VPWR_c_236_n 0.0137828f $X=3.32 $Y=1.445 $X2=0 $Y2=0
cc_142 N_B_N_c_168_n N_VPWR_c_237_n 0.00743866f $X=3.075 $Y=1.99 $X2=0 $Y2=0
cc_143 N_B_N_c_168_n N_VPWR_c_233_n 0.015347f $X=3.075 $Y=1.99 $X2=0 $Y2=0
cc_144 B_N N_VPWR_c_233_n 0.00343698f $X=3.32 $Y=1.445 $X2=0 $Y2=0
cc_145 N_B_N_c_162_n N_VGND_c_324_n 0.00548538f $X=3.27 $Y=1.17 $X2=0 $Y2=0
cc_146 N_B_N_c_163_n N_VGND_c_324_n 0.00306356f $X=3.125 $Y=1.16 $X2=0 $Y2=0
cc_147 B_N N_VGND_c_324_n 0.0127012f $X=3.32 $Y=1.105 $X2=0 $Y2=0
cc_148 N_B_N_c_166_n N_VGND_c_324_n 0.0162897f $X=3.142 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B_N_c_166_n N_VGND_c_327_n 0.00585385f $X=3.142 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B_N_c_166_n N_VGND_c_329_n 0.0132084f $X=3.142 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_27_297#_c_196_n N_VPWR_M1000_d 0.00188315f $X=1.095 $Y=1.55 $X2=-0.19
+ $Y2=1.305
cc_152 N_A_27_297#_c_196_n N_VPWR_c_234_n 0.0145257f $X=1.095 $Y=1.55 $X2=0
+ $Y2=0
cc_153 N_A_27_297#_c_216_p N_VPWR_c_237_n 0.015002f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_154 N_A_27_297#_c_206_n N_VPWR_c_237_n 0.0386815f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_155 N_A_27_297#_c_198_n N_VPWR_c_237_n 0.0191589f $X=2.18 $Y=2.295 $X2=0
+ $Y2=0
cc_156 N_A_27_297#_c_195_n N_VPWR_c_238_n 0.0211751f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_157 N_A_27_297#_M1000_s N_VPWR_c_233_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_158 N_A_27_297#_M1005_s N_VPWR_c_233_n 0.00297222f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_159 N_A_27_297#_M1003_d N_VPWR_c_233_n 0.00217519f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_160 N_A_27_297#_c_195_n N_VPWR_c_233_n 0.0122467f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_161 N_A_27_297#_c_216_p N_VPWR_c_233_n 0.00962794f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_162 N_A_27_297#_c_206_n N_VPWR_c_233_n 0.0239144f $X=2.035 $Y=2.38 $X2=0
+ $Y2=0
cc_163 N_A_27_297#_c_198_n N_VPWR_c_233_n 0.0111632f $X=2.18 $Y=2.295 $X2=0
+ $Y2=0
cc_164 N_A_27_297#_c_206_n N_Y_M1001_s 0.00352392f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_165 N_A_27_297#_c_197_n N_Y_c_273_n 0.00317178f $X=1.22 $Y=1.655 $X2=0 $Y2=0
cc_166 N_A_27_297#_c_197_n N_Y_c_275_n 0.00281802f $X=1.22 $Y=1.655 $X2=0 $Y2=0
cc_167 N_A_27_297#_c_206_n N_Y_c_275_n 0.0134104f $X=2.035 $Y=2.38 $X2=0 $Y2=0
cc_168 N_A_27_297#_c_199_n N_Y_c_275_n 0.00262601f $X=2.16 $Y=1.63 $X2=0 $Y2=0
cc_169 N_A_27_297#_c_194_n N_VGND_c_319_n 0.0114749f $X=0.245 $Y=1.655 $X2=0
+ $Y2=0
cc_170 N_VPWR_c_233_n N_Y_M1001_s 0.00232895f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_171 N_Y_c_273_n N_VGND_M1008_s 0.00161804f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_172 N_Y_c_274_n N_VGND_c_319_n 0.00752789f $X=0.935 $Y=0.81 $X2=0 $Y2=0
cc_173 N_Y_c_278_n N_VGND_c_320_n 0.0238677f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_174 N_Y_c_273_n N_VGND_c_320_n 0.00238269f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_175 N_Y_c_273_n N_VGND_c_321_n 0.0122105f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_176 N_Y_c_276_n N_VGND_c_322_n 0.0109535f $X=1.665 $Y=0.81 $X2=0 $Y2=0
cc_177 N_Y_c_286_n N_VGND_c_322_n 0.0287371f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_178 N_Y_c_273_n N_VGND_c_325_n 0.00198102f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_179 N_Y_c_286_n N_VGND_c_325_n 0.0224022f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_180 N_Y_M1004_d N_VGND_c_329_n 0.002955f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_181 N_Y_M1006_s N_VGND_c_329_n 0.0025535f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_182 N_Y_c_278_n N_VGND_c_329_n 0.0150984f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_183 N_Y_c_273_n N_VGND_c_329_n 0.00896169f $X=1.475 $Y=0.81 $X2=0 $Y2=0
cc_184 N_Y_c_286_n N_VGND_c_329_n 0.0141397f $X=1.69 $Y=0.39 $X2=0 $Y2=0
