* File: sky130_fd_sc_hdll__sdfxtp_1.pex.spice
* Created: Thu Aug 27 19:27:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%CLK 1 2 3 5 6 8 13
c38 1 0 2.71124e-20 $X=0.31 $Y=1.325
r39 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r40 6 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.5 $Y=1.665 $X2=0.31
+ $Y2=1.665
r41 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=1.74 $X2=0.5
+ $Y2=2.135
r42 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r43 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r44 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r45 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r46 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_27_47# 1 2 9 12 13 15 18 20 21 23 24 26
+ 28 29 31 32 36 40 44 45 46 49 51 54 63 66 67 68 70 72 77 82 86
c231 82 0 1.69827e-19 $X=7.315 $Y=1.32
c232 66 0 1.55016e-19 $X=5.75 $Y=1.825
c233 46 0 1.76957e-19 $X=0.665 $Y=1.88
r234 85 87 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.315 $Y=1.41
+ $X2=7.315 $Y2=1.575
r235 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.315
+ $Y=1.41 $X2=7.315 $Y2=1.41
r236 82 85 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.315 $Y=1.32
+ $X2=7.315 $Y2=1.41
r237 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.74 $X2=5.55 $Y2=1.74
r238 76 77 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=0.94 $Y=1.235
+ $X2=0.97 $Y2=1.235
r239 71 86 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=7.35 $Y=1.825
+ $X2=7.35 $Y2=1.41
r240 70 72 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.325 $Y=1.825
+ $X2=7.13 $Y2=1.825
r241 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.325 $Y=1.825
+ $X2=7.325 $Y2=1.825
r242 68 72 1.52846 $w=1.4e-07 $l=1.235e-06 $layer=MET1_cond $X=5.895 $Y=1.87
+ $X2=7.13 $Y2=1.87
r243 66 81 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=5.75 $Y=1.832
+ $X2=5.55 $Y2=1.832
r244 65 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.895 $Y2=1.825
r245 65 67 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.555 $Y2=1.825
r246 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.825
+ $X2=5.75 $Y2=1.825
r247 63 67 5.76732 $w=1.4e-07 $l=4.66e-06 $layer=MET1_cond $X=0.895 $Y=1.87
+ $X2=5.555 $Y2=1.87
r248 60 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.75 $Y=1.825
+ $X2=0.895 $Y2=1.825
r249 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.75 $Y=1.825
+ $X2=0.75 $Y2=1.825
r250 52 76 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r251 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r252 49 61 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.88
r253 49 51 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.235
r254 48 51 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.805
+ $X2=0.78 $Y2=1.235
r255 47 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r256 46 61 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.78 $Y2=1.88
r257 46 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.35 $Y2=1.88
r258 44 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.78 $Y2=0.805
r259 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.345 $Y2=0.72
r260 38 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r261 38 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r262 34 36 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=7.83 $Y=1.245
+ $X2=7.83 $Y2=0.415
r263 33 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.45 $Y=1.32
+ $X2=7.315 $Y2=1.32
r264 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.755 $Y=1.32
+ $X2=7.83 $Y2=1.245
r265 32 33 156.394 $w=1.5e-07 $l=3.05e-07 $layer=POLY_cond $X=7.755 $Y=1.32
+ $X2=7.45 $Y2=1.32
r266 29 31 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.28 $Y=1.99
+ $X2=7.28 $Y2=2.275
r267 28 29 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.28 $Y=1.89 $X2=7.28
+ $Y2=1.99
r268 28 87 104.447 $w=2e-07 $l=3.15e-07 $layer=POLY_cond $X=7.28 $Y=1.89
+ $X2=7.28 $Y2=1.575
r269 24 80 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.575 $Y2=1.74
r270 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.515 $Y2=2.275
r271 23 80 31.9848 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.515 $Y=1.575
+ $X2=5.575 $Y2=1.74
r272 22 23 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=5.515 $Y=1.395
+ $X2=5.515 $Y2=1.575
r273 20 22 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.515 $Y2=1.395
r274 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.055 $Y2=1.32
r275 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=5.055 $Y2=1.32
r276 16 18 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=4.98 $Y2=0.415
r277 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.97 $Y=1.74
+ $X2=0.97 $Y2=2.135
r278 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.97 $Y=1.64 $X2=0.97
+ $Y2=1.74
r279 11 77 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.37
+ $X2=0.97 $Y2=1.235
r280 11 12 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.97 $Y=1.37 $X2=0.97
+ $Y2=1.64
r281 7 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r282 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r283 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r284 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCE 1 3 6 8 10 13 15 19 22 28 33 35 37
c96 28 0 7.84804e-20 $X=2.025 $Y=1.52
c97 15 0 1.59107e-19 $X=3.335 $Y=0.7
c98 6 0 1.74476e-19 $X=2.01 $Y=0.445
r99 35 37 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.047 $Y=0.785
+ $X2=2.047 $Y2=0.84
r100 28 30 70.4729 $w=2.77e-07 $l=4.05e-07 $layer=POLY_cond $X=2.025 $Y=1.577
+ $X2=2.43 $Y2=1.577
r101 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.025
+ $Y=1.52 $X2=2.025 $Y2=1.52
r102 26 28 2.61011 $w=2.77e-07 $l=1.5e-08 $layer=POLY_cond $X=2.01 $Y=1.577
+ $X2=2.025 $Y2=1.577
r103 25 26 8.70036 $w=2.77e-07 $l=5e-08 $layer=POLY_cond $X=1.96 $Y=1.577
+ $X2=2.01 $Y2=1.577
r104 22 35 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=0.7
+ $X2=2.047 $Y2=0.785
r105 22 29 22.8081 $w=3.33e-07 $l=6.63e-07 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=1.52
r106 22 37 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=0.84
r107 20 33 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.42 $Y=0.95
+ $X2=3.53 $Y2=0.95
r108 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=0.95 $X2=3.42 $Y2=0.95
r109 17 19 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0.785
+ $X2=3.42 $Y2=0.95
r110 16 22 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.215 $Y=0.7
+ $X2=2.047 $Y2=0.7
r111 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=3.42 $Y2=0.785
r112 15 16 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=2.215 $Y2=0.7
r113 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.95
r114 11 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.445
r115 8 30 12.8788 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=1.577
r116 8 10 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=2.165
r117 4 26 17.1008 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.01 $Y=1.385
+ $X2=2.01 $Y2=1.577
r118 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=2.01 $Y=1.385 $X2=2.01
+ $Y2=0.445
r119 1 25 12.8788 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=1.577
r120 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_319_47# 1 2 9 11 13 15 18 20 23 24 28
+ 34 36 39 40 42
c115 39 0 2.52956e-19 $X=2.55 $Y=1.04
c116 28 0 1.76415e-19 $X=3.455 $Y=1.52
r117 40 44 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.55 $Y=1.04
+ $X2=2.55 $Y2=0.875
r118 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.04 $X2=2.55 $Y2=1.04
r119 31 34 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.62 $Y=0.36
+ $X2=1.74 $Y2=0.36
r120 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.455
+ $Y=1.52 $X2=3.455 $Y2=1.52
r121 26 28 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=3.435 $Y=1.86
+ $X2=3.435 $Y2=1.52
r122 25 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=1.967
+ $X2=2.47 $Y2=1.967
r123 24 26 6.81772 $w=2.15e-07 $l=1.50612e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=3.435 $Y2=1.86
r124 24 25 41.5415 $w=2.13e-07 $l=7.75e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=2.555 $Y2=1.967
r125 23 42 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.47 $Y=1.86
+ $X2=2.47 $Y2=1.967
r126 22 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.04
r127 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.86
r128 21 36 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.81 $Y=1.967
+ $X2=1.672 $Y2=1.967
r129 20 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=2.47 $Y2=1.967
r130 20 21 30.8211 $w=2.13e-07 $l=5.75e-07 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=1.81 $Y2=1.967
r131 16 36 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=1.967
r132 16 18 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=2.175
r133 15 36 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.62 $Y=1.86
+ $X2=1.672 $Y2=1.967
r134 14 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=0.36
r135 14 15 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=1.86
r136 11 29 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.455 $Y2=1.52
r137 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.42 $Y2=2.165
r138 9 44 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.46 $Y=0.445
+ $X2=2.46 $Y2=0.875
r139 2 18 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.845 $X2=1.725 $Y2=2.175
r140 1 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.74 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%D 1 3 6 8 15
r40 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.52 $X2=2.91 $Y2=1.52
r41 8 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.99 $Y=1.52 $X2=2.91
+ $Y2=1.52
r42 4 11 33.7441 $w=3.01e-07 $l=1.74284e-07 $layer=POLY_cond $X=3 $Y=1.385
+ $X2=2.91 $Y2=1.52
r43 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=3 $Y=1.385 $X2=3 $Y2=0.445
r44 1 11 47.761 $w=3.01e-07 $l=2.69258e-07 $layer=POLY_cond $X=2.95 $Y=1.77
+ $X2=2.91 $Y2=1.52
r45 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.95 $Y=1.77 $X2=2.95
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%SCD 3 6 7 9 10 13
c53 6 0 1.76415e-19 $X=3.935 $Y=1.67
c54 3 0 1.59107e-19 $X=3.91 $Y=0.445
r55 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.52
r56 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.19
r57 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.97
+ $Y=1.355 $X2=3.97 $Y2=1.355
r58 10 14 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=1.19
+ $X2=3.91 $Y2=1.355
r59 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.935 $Y=1.77
+ $X2=3.935 $Y2=2.165
r60 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.77
r61 6 16 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.52
r62 3 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.91 $Y=0.445
+ $X2=3.91 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_203_47# 1 2 7 9 12 15 16 18 21 26 29 38
+ 42 43 45 47 51 52 53 56 58 62
c201 45 0 5.35254e-21 $X=7.395 $Y=0.805
c202 43 0 1.7664e-19 $X=5.385 $Y=0.805
r203 56 58 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=7.365 $Y=0.87
+ $X2=7.365 $Y2=0.705
r204 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.365
+ $Y=0.87 $X2=7.365 $Y2=0.87
r205 51 53 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.45 $Y=0.87
+ $X2=5.45 $Y2=0.705
r206 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=0.87 $X2=5.45 $Y2=0.87
r207 45 47 0.128299 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=7.395 $Y=0.805
+ $X2=7.23 $Y2=0.805
r208 45 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.395 $Y=0.805
+ $X2=7.395 $Y2=0.805
r209 43 47 2.28341 $w=1.4e-07 $l=1.845e-06 $layer=MET1_cond $X=5.385 $Y=0.85
+ $X2=7.23 $Y2=0.85
r210 41 52 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.45 $Y2=0.87
r211 41 70 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.05 $Y2=0.87
r212 40 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.385 $Y2=0.805
r213 40 42 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.045 $Y2=0.805
r214 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=0.805
+ $X2=5.24 $Y2=0.805
r215 38 42 4.52969 $w=1.4e-07 $l=3.66e-06 $layer=MET1_cond $X=1.385 $Y=0.85
+ $X2=5.045 $Y2=0.85
r216 36 66 57.8727 $w=2.28e-07 $l=1.155e-06 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=1.96
r217 36 62 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=0.51
r218 35 38 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.24 $Y=0.805
+ $X2=1.385 $Y2=0.805
r219 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.24 $Y=0.805
+ $X2=1.24 $Y2=0.805
r220 29 57 12.9213 $w=3.28e-07 $l=3.7e-07 $layer=LI1_cond $X=7.735 $Y=0.87
+ $X2=7.365 $Y2=0.87
r221 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.825
+ $Y=1.74 $X2=7.825 $Y2=1.74
r222 24 29 7.26367 $w=3.3e-07 $l=2.11069e-07 $layer=LI1_cond $X=7.84 $Y=1.035
+ $X2=7.735 $Y2=0.87
r223 24 26 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=7.84 $Y=1.035
+ $X2=7.84 $Y2=1.74
r224 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.74 $X2=4.99 $Y2=1.74
r225 19 70 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=0.87
r226 19 21 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=1.74
r227 16 27 48.3784 $w=2.91e-07 $l=2.80624e-07 $layer=POLY_cond $X=7.76 $Y=1.99
+ $X2=7.825 $Y2=1.74
r228 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.76 $Y=1.99
+ $X2=7.76 $Y2=2.275
r229 15 58 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.305 $Y=0.415
+ $X2=7.305 $Y2=0.705
r230 12 53 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.51 $Y=0.415
+ $X2=5.51 $Y2=0.705
r231 7 22 46.5577 $w=3.26e-07 $l=2.57391e-07 $layer=POLY_cond $X=5 $Y=1.99
+ $X2=5.015 $Y2=1.74
r232 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5 $Y=1.99 $X2=5
+ $Y2=2.275
r233 2 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.815 $X2=1.205 $Y2=1.96
r234 1 62 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1189_21# 1 2 9 12 13 15 16 19 22 25 30
+ 32
c92 13 0 1.55016e-19 $X=6.045 $Y=1.99
r93 23 32 6.56857 $w=2.45e-07 $l=1.83916e-07 $layer=LI1_cond $X=6.957 $Y=1.095
+ $X2=6.917 $Y2=0.93
r94 23 25 65.1929 $w=2.03e-07 $l=1.205e-06 $layer=LI1_cond $X=6.957 $Y=1.095
+ $X2=6.957 $Y2=2.3
r95 22 32 6.56857 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=6.917 $Y=0.765
+ $X2=6.917 $Y2=0.93
r96 21 30 11.6128 $w=1.68e-07 $l=1.78e-07 $layer=LI1_cond $X=6.917 $Y=0.45
+ $X2=7.095 $Y2=0.45
r97 21 22 9.30042 $w=2.83e-07 $l=2.3e-07 $layer=LI1_cond $X=6.917 $Y=0.535
+ $X2=6.917 $Y2=0.765
r98 19 35 32.7676 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.12 $Y=0.93
+ $X2=6.12 $Y2=1.065
r99 19 34 41.4854 $w=3.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.12 $Y=0.93
+ $X2=6.12 $Y2=0.795
r100 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.13
+ $Y=0.93 $X2=6.13 $Y2=0.93
r101 16 32 0.295496 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=6.775 $Y=0.93
+ $X2=6.917 $Y2=0.93
r102 16 18 22.525 $w=3.28e-07 $l=6.45e-07 $layer=LI1_cond $X=6.775 $Y=0.93
+ $X2=6.13 $Y2=0.93
r103 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.045 $Y=1.99
+ $X2=6.045 $Y2=2.275
r104 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.045 $Y=1.89 $X2=6.045
+ $Y2=1.99
r105 12 35 273.551 $w=2e-07 $l=8.25e-07 $layer=POLY_cond $X=6.045 $Y=1.89
+ $X2=6.045 $Y2=1.065
r106 9 34 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.02 $Y=0.445
+ $X2=6.02 $Y2=0.795
r107 2 25 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=6.83
+ $Y=1.735 $X2=6.975 $Y2=2.3
r108 1 30 182 $w=1.7e-07 $l=3.46194e-07 $layer=licon1_NDIFF $count=1 $X=6.84
+ $Y=0.235 $X2=7.095 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1011_47# 1 2 7 9 12 14 15 16 20 25 27
+ 28 30
c103 25 0 1.79445e-19 $X=5.79 $Y=1.315
r104 33 34 21.0617 $w=2.01e-07 $l=3.47e-07 $layer=LI1_cond $X=5.79 $Y=1.445
+ $X2=6.137 $Y2=1.445
r105 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.52
+ $Y=1.41 $X2=6.52 $Y2=1.41
r106 28 34 5.0239 $w=2.6e-07 $l=9.3e-08 $layer=LI1_cond $X=6.23 $Y=1.445
+ $X2=6.137 $Y2=1.445
r107 28 30 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=6.23 $Y=1.445
+ $X2=6.52 $Y2=1.445
r108 26 34 1.24766 $w=1.85e-07 $l=1.3e-07 $layer=LI1_cond $X=6.137 $Y=1.575
+ $X2=6.137 $Y2=1.445
r109 26 27 36.8698 $w=1.83e-07 $l=6.15e-07 $layer=LI1_cond $X=6.137 $Y=1.575
+ $X2=6.137 $Y2=2.19
r110 25 33 1.71937 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=5.79 $Y=1.315
+ $X2=5.79 $Y2=1.445
r111 24 25 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.79 $Y=0.535
+ $X2=5.79 $Y2=1.315
r112 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.705 $Y=0.45
+ $X2=5.79 $Y2=0.535
r113 20 22 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=5.705 $Y=0.45
+ $X2=5.3 $Y2=0.45
r114 16 27 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=6.137 $Y2=2.19
r115 16 18 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=5.26 $Y2=2.275
r116 14 31 26.6608 $w=2.7e-07 $l=1.2e-07 $layer=POLY_cond $X=6.64 $Y=1.41
+ $X2=6.52 $Y2=1.41
r117 14 15 1.40033 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=6.64 $Y=1.41
+ $X2=6.74 $Y2=1.467
r118 10 15 30.0832 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=6.765 $Y=1.275
+ $X2=6.74 $Y2=1.467
r119 10 12 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=6.765 $Y=1.275
+ $X2=6.765 $Y2=0.555
r120 7 15 30.0832 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=6.74 $Y=1.66
+ $X2=6.74 $Y2=1.467
r121 7 9 120.5 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.74 $Y=1.66 $X2=6.74
+ $Y2=2.11
r122 2 18 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=2.065 $X2=5.26 $Y2=2.275
r123 1 22 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.3 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1647_21# 1 2 9 11 13 14 16 17 19 20 27
+ 30 32 35 39 42 43
r84 39 41 16.9646 $w=3.58e-07 $l=4.4e-07 $layer=LI1_cond $X=9.22 $Y=0.385
+ $X2=9.22 $Y2=0.825
r85 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.945
+ $Y=1.16 $X2=9.945 $Y2=1.16
r86 33 43 0.674692 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=9.405 $Y=1.16
+ $X2=9.312 $Y2=1.16
r87 33 35 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.405 $Y=1.16
+ $X2=9.945 $Y2=1.16
r88 32 42 6.7841 $w=2.35e-07 $l=1.88348e-07 $layer=LI1_cond $X=9.312 $Y=1.575
+ $X2=9.262 $Y2=1.74
r89 31 43 8.18839 $w=1.82e-07 $l=1.65e-07 $layer=LI1_cond $X=9.312 $Y=1.325
+ $X2=9.312 $Y2=1.16
r90 31 32 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=9.312 $Y=1.325
+ $X2=9.312 $Y2=1.575
r91 30 43 8.18839 $w=1.82e-07 $l=1.65997e-07 $layer=LI1_cond $X=9.31 $Y=0.995
+ $X2=9.312 $Y2=1.16
r92 30 41 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=9.31 $Y=0.995
+ $X2=9.31 $Y2=0.825
r93 25 42 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=9.262 $Y=1.905
+ $X2=9.262 $Y2=1.74
r94 25 27 1.81965 $w=2.83e-07 $l=4.5e-08 $layer=LI1_cond $X=9.262 $Y=1.905
+ $X2=9.262 $Y2=1.95
r95 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.54
+ $Y=1.74 $X2=8.54 $Y2=1.74
r96 20 42 0.153733 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=9.12 $Y=1.74
+ $X2=9.262 $Y2=1.74
r97 20 22 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=9.12 $Y=1.74
+ $X2=8.54 $Y2=1.74
r98 17 36 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=9.91 $Y=1.41
+ $X2=9.945 $Y2=1.16
r99 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.91 $Y=1.41
+ $X2=9.91 $Y2=1.985
r100 14 36 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=9.885 $Y=0.995
+ $X2=9.945 $Y2=1.16
r101 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.885 $Y=0.995
+ $X2=9.885 $Y2=0.56
r102 11 23 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=8.335 $Y=1.99
+ $X2=8.455 $Y2=1.74
r103 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.335 $Y=1.99
+ $X2=8.335 $Y2=2.275
r104 7 23 39.3952 $w=3.9e-07 $l=2.26164e-07 $layer=POLY_cond $X=8.31 $Y=1.575
+ $X2=8.455 $Y2=1.74
r105 7 9 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=8.31 $Y=1.575
+ $X2=8.31 $Y2=0.445
r106 2 27 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=9.08
+ $Y=1.485 $X2=9.205 $Y2=1.95
r107 1 39 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=9.08
+ $Y=0.235 $X2=9.205 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_1474_413# 1 2 7 9 10 12 13 14 15 19 24
+ 26 29 32
c85 32 0 1.25162e-19 $X=8.2 $Y=1.16
c86 15 0 1.64475e-19 $X=8.115 $Y=2.25
r87 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.965
+ $Y=1.16 $X2=8.965 $Y2=1.16
r88 27 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.285 $Y=1.16 $X2=8.2
+ $Y2=1.16
r89 27 29 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.285 $Y=1.16
+ $X2=8.965 $Y2=1.16
r90 25 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.2 $Y=1.325 $X2=8.2
+ $Y2=1.16
r91 25 26 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=8.2 $Y=1.325 $X2=8.2
+ $Y2=2.165
r92 24 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.2 $Y=0.995 $X2=8.2
+ $Y2=1.16
r93 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=8.2 $Y=0.535 $X2=8.2
+ $Y2=0.995
r94 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.115 $Y=0.45
+ $X2=8.2 $Y2=0.535
r95 19 21 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.115 $Y=0.45
+ $X2=7.62 $Y2=0.45
r96 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.115 $Y=2.25
+ $X2=8.2 $Y2=2.165
r97 15 17 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=8.115 $Y=2.25
+ $X2=7.515 $Y2=2.25
r98 13 30 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=9.34 $Y=1.16
+ $X2=8.965 $Y2=1.16
r99 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=9.34 $Y=1.16
+ $X2=9.44 $Y2=1.202
r100 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=9.465 $Y=0.995
+ $X2=9.44 $Y2=1.202
r101 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.465 $Y=0.995
+ $X2=9.465 $Y2=0.56
r102 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=9.44 $Y=1.41
+ $X2=9.44 $Y2=1.202
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.44 $Y=1.41
+ $X2=9.44 $Y2=1.985
r104 2 17 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=2.065 $X2=7.515 $Y2=2.25
r105 1 21 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=7.38
+ $Y=0.235 $X2=7.62 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%VPWR 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 52 54 59 77 86 87 90 93 96
c150 1 0 1.76957e-19 $X=0.59 $Y=1.815
r151 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r152 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r153 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r154 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r155 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r156 84 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.51 $Y2=2.72
r157 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r158 81 96 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.77 $Y=2.72
+ $X2=8.617 $Y2=2.72
r159 81 83 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.77 $Y=2.72
+ $X2=9.43 $Y2=2.72
r160 80 97 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r161 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r162 77 96 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.465 $Y=2.72
+ $X2=8.617 $Y2=2.72
r163 77 79 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=8.465 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 76 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r165 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r166 73 76 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r167 72 75 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r168 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r169 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r170 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r171 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r172 67 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r173 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r174 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r175 64 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.17 $Y2=2.72
r176 64 66 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.53 $Y2=2.72
r177 63 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r178 63 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r179 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r180 60 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.9 $Y=2.72 $X2=0.71
+ $Y2=2.72
r181 60 62 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.9 $Y=2.72
+ $X2=1.61 $Y2=2.72
r182 59 93 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.17 $Y2=2.72
r183 59 62 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=1.61 $Y2=2.72
r184 54 90 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.71 $Y2=2.72
r185 54 56 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r186 52 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r187 52 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r188 50 83 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=9.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r189 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.59 $Y=2.72
+ $X2=9.675 $Y2=2.72
r190 49 86 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=10.35 $Y2=2.72
r191 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=2.72
+ $X2=9.675 $Y2=2.72
r192 47 75 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=6.4 $Y=2.72
+ $X2=6.21 $Y2=2.72
r193 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.4 $Y=2.72
+ $X2=6.485 $Y2=2.72
r194 46 79 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=6.57 $Y=2.72 $X2=6.67
+ $Y2=2.72
r195 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=2.72
+ $X2=6.485 $Y2=2.72
r196 44 69 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.11 $Y=2.72 $X2=3.91
+ $Y2=2.72
r197 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=4.195 $Y2=2.72
r198 43 72 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.28 $Y=2.72 $X2=4.37
+ $Y2=2.72
r199 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.72
+ $X2=4.195 $Y2=2.72
r200 39 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.675 $Y=2.635
+ $X2=9.675 $Y2=2.72
r201 39 41 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.675 $Y=2.635
+ $X2=9.675 $Y2=1.79
r202 35 96 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.617 $Y=2.635
+ $X2=8.617 $Y2=2.72
r203 35 37 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.617 $Y=2.635
+ $X2=8.617 $Y2=2.3
r204 31 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=2.635
+ $X2=6.485 $Y2=2.72
r205 31 33 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.485 $Y=2.635
+ $X2=6.485 $Y2=2
r206 27 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.72
r207 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.33
r208 23 93 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.72
r209 23 25 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.33
r210 19 90 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.72
r211 19 21 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.22
r212 6 41 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=9.53
+ $Y=1.485 $X2=9.675 $Y2=1.79
r213 5 37 600 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=2.065 $X2=8.68 $Y2=2.3
r214 4 33 300 $w=1.7e-07 $l=3.81117e-07 $layer=licon1_PDIFF $count=2 $X=6.135
+ $Y=2.065 $X2=6.485 $Y2=2
r215 3 29 600 $w=1.7e-07 $l=5.63627e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.845 $X2=4.195 $Y2=2.33
r216 2 25 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.845 $X2=2.195 $Y2=2.33
r217 1 21 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.815 $X2=0.735 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%A_608_369# 1 2 3 4 13 17 22 24 25 26 27
+ 28 30 32 36 38 39
c113 30 0 1.7664e-19 $X=4.65 $Y=0.695
r114 39 41 21.3062 $w=2.09e-07 $l=3.65e-07 $layer=LI1_cond $X=4.682 $Y=1.91
+ $X2=4.682 $Y2=2.275
r115 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.65 $Y=0.45 $X2=4.75
+ $Y2=0.45
r116 32 39 5.42244 $w=2.09e-07 $l=9.97246e-08 $layer=LI1_cond $X=4.65 $Y=1.825
+ $X2=4.682 $Y2=1.91
r117 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=0.78
r118 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=1.825
r119 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.695
+ $X2=4.65 $Y2=0.78
r120 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.45
r121 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.695
r122 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=4.65 $Y2=0.78
r123 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=3.895 $Y2=0.78
r124 25 39 1.94907 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=4.682 $Y2=1.91
r125 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=3.89 $Y2=1.91
r126 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.695
+ $X2=3.895 $Y2=0.78
r127 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.81 $Y=0.445
+ $X2=3.81 $Y2=0.695
r128 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.89 $Y2=1.91
r129 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.805 $Y2=2.245
r130 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.81 $Y2=0.445
r131 17 19 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.265 $Y2=0.36
r132 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.805 $Y2=2.245
r133 13 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.185 $Y2=2.33
r134 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=2.065 $X2=4.715 $Y2=2.275
r135 3 15 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.845 $X2=3.185 $Y2=2.33
r136 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.75 $Y2=0.45
r137 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.235 $X2=3.265 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%Q 1 2 10 13 18 24 25
r26 24 25 5.62797 $w=5.38e-07 $l=8.5e-08 $layer=LI1_cond $X=10.2 $Y=1.63
+ $X2=10.2 $Y2=1.545
r27 16 18 1.10748 $w=5.38e-07 $l=5e-08 $layer=LI1_cond $X=10.2 $Y=1.815 $X2=10.2
+ $Y2=1.865
r28 13 16 0.55374 $w=5.38e-07 $l=2.5e-08 $layer=LI1_cond $X=10.2 $Y=1.79
+ $X2=10.2 $Y2=1.815
r29 13 24 3.54394 $w=5.38e-07 $l=1.6e-07 $layer=LI1_cond $X=10.2 $Y=1.79
+ $X2=10.2 $Y2=1.63
r30 13 21 9.63508 $w=5.38e-07 $l=4.35e-07 $layer=LI1_cond $X=10.2 $Y=1.875
+ $X2=10.2 $Y2=2.31
r31 13 18 0.221496 $w=5.38e-07 $l=1e-08 $layer=LI1_cond $X=10.2 $Y=1.875
+ $X2=10.2 $Y2=1.865
r32 12 25 34.8134 $w=2.38e-07 $l=7.25e-07 $layer=LI1_cond $X=10.35 $Y=0.82
+ $X2=10.35 $Y2=1.545
r33 10 12 13.1588 $w=5.38e-07 $l=4.25e-07 $layer=LI1_cond $X=10.2 $Y=0.395
+ $X2=10.2 $Y2=0.82
r34 2 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=1.485 $X2=10.145 $Y2=1.63
r35 2 21 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10
+ $Y=1.485 $X2=10.145 $Y2=2.31
r36 1 10 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=9.96
+ $Y=0.235 $X2=10.145 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_1%VGND 1 2 3 4 5 6 21 25 29 33 37 40 41 43
+ 44 46 47 49 50 51 53 77 86 87 91 97
c152 87 0 2.71124e-20 $X=10.35 $Y=0
r153 97 98 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r154 91 94 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r155 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r156 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r157 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r158 84 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.51
+ $Y2=0
r159 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r160 81 97 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=8.77 $Y=0 $X2=8.612
+ $Y2=0
r161 81 83 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.77 $Y=0 $X2=9.43
+ $Y2=0
r162 80 98 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.51 $Y2=0
r163 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r164 77 97 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=8.455 $Y=0
+ $X2=8.612 $Y2=0
r165 77 79 116.455 $w=1.68e-07 $l=1.785e-06 $layer=LI1_cond $X=8.455 $Y=0
+ $X2=6.67 $Y2=0
r166 76 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r167 75 76 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r168 73 76 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.21 $Y2=0
r169 72 75 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=6.21
+ $Y2=0
r170 72 73 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r171 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r172 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r173 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r174 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r175 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r176 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r177 63 64 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r178 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r179 61 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r180 60 63 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r181 60 61 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r182 58 91 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r183 58 60 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r184 53 91 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r185 53 55 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r186 51 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r187 51 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r188 49 83 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=9.59 $Y=0 $X2=9.43
+ $Y2=0
r189 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.59 $Y=0 $X2=9.675
+ $Y2=0
r190 48 86 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=9.76 $Y=0 $X2=10.35
+ $Y2=0
r191 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.76 $Y=0 $X2=9.675
+ $Y2=0
r192 46 75 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.21
+ $Y2=0
r193 46 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.41
+ $Y2=0
r194 45 79 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.67
+ $Y2=0
r195 45 47 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.41
+ $Y2=0
r196 43 69 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=3.91 $Y2=0
r197 43 44 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.215
+ $Y2=0
r198 42 72 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r199 42 44 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.215
+ $Y2=0
r200 40 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r201 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.24
+ $Y2=0
r202 39 66 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.405 $Y=0
+ $X2=2.53 $Y2=0
r203 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=0 $X2=2.24
+ $Y2=0
r204 35 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.675 $Y=0.085
+ $X2=9.675 $Y2=0
r205 35 37 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.675 $Y=0.085
+ $X2=9.675 $Y2=0.53
r206 31 97 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=8.612 $Y=0.085
+ $X2=8.612 $Y2=0
r207 31 33 13.3537 $w=3.13e-07 $l=3.65e-07 $layer=LI1_cond $X=8.612 $Y=0.085
+ $X2=8.612 $Y2=0.45
r208 27 47 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0
r209 27 29 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0.42
r210 23 44 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r211 23 25 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.36
r212 19 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0
r213 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.24 $Y=0.085
+ $X2=2.24 $Y2=0.36
r214 6 37 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=9.54
+ $Y=0.235 $X2=9.675 $Y2=0.53
r215 5 33 182 $w=1.7e-07 $l=3.93065e-07 $layer=licon1_NDIFF $count=1 $X=8.385
+ $Y=0.235 $X2=8.685 $Y2=0.45
r216 4 29 182 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_NDIFF $count=1 $X=6.095
+ $Y=0.235 $X2=6.48 $Y2=0.42
r217 3 25 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.2 $Y2=0.36
r218 2 21 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.24 $Y2=0.36
r219 1 94 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

