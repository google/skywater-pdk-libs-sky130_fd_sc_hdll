* File: sky130_fd_sc_hdll__isobufsrc_1.pxi.spice
* Created: Wed Sep  2 08:33:40 2020
* 
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A N_A_M1004_g N_A_c_44_n N_A_M1005_g
+ N_A_c_41_n N_A_c_42_n A A PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%SLEEP N_SLEEP_c_70_n N_SLEEP_M1002_g
+ N_SLEEP_c_71_n N_SLEEP_M1001_g SLEEP SLEEP
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%SLEEP
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A_74_47# N_A_74_47#_M1004_s
+ N_A_74_47#_M1005_s N_A_74_47#_c_103_n N_A_74_47#_M1000_g N_A_74_47#_c_104_n
+ N_A_74_47#_M1003_g N_A_74_47#_c_112_n N_A_74_47#_c_105_n N_A_74_47#_c_106_n
+ N_A_74_47#_c_110_n N_A_74_47#_c_107_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%A_74_47#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VPWR N_VPWR_M1005_d N_VPWR_c_159_n VPWR
+ N_VPWR_c_160_n N_VPWR_c_161_n N_VPWR_c_158_n N_VPWR_c_163_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VPWR
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%X N_X_M1002_d N_X_M1003_d N_X_c_188_n
+ N_X_c_184_n N_X_c_189_n X N_X_c_186_n N_X_c_185_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%X
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VGND N_VGND_M1004_d N_VGND_M1000_d
+ N_VGND_c_214_n N_VGND_c_215_n N_VGND_c_216_n N_VGND_c_217_n N_VGND_c_218_n
+ VGND N_VGND_c_219_n N_VGND_c_220_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_1%VGND
cc_1 VNB N_A_M1004_g 0.0365595f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.445
cc_2 VNB N_A_c_41_n 0.0413574f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_3 VNB N_A_c_42_n 0.015019f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_4 VNB A 0.0263972f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_5 VNB N_SLEEP_c_70_n 0.0179274f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.995
cc_6 VNB N_SLEEP_c_71_n 0.0268302f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB SLEEP 0.00375062f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.695
cc_8 VNB N_A_74_47#_c_103_n 0.020138f $X=-0.19 $Y=-0.24 $X2=0.735 $Y2=1.695
cc_9 VNB N_A_74_47#_c_104_n 0.0272567f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_A_74_47#_c_105_n 7.40462e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_74_47#_c_106_n 0.00758253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_74_47#_c_107_n 0.00490456f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_158_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_14 VNB N_X_c_184_n 0.00888499f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_15 VNB N_X_c_185_n 0.0227195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_214_n 0.00752718f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.995
cc_17 VNB N_VGND_c_215_n 0.0134731f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_VGND_c_216_n 0.0151623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_217_n 0.0275208f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_20 VNB N_VGND_c_218_n 0.00403597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_219_n 0.017745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_220_n 0.146529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VPB N_A_c_44_n 0.0233261f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.41
cc_24 VPB N_A_c_41_n 0.0183665f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_25 VPB N_A_c_42_n 0.00764078f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=0.995
cc_26 VPB A 0.00949562f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_27 VPB N_SLEEP_c_71_n 0.0294898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB SLEEP 6.05838e-19 $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.695
cc_29 VPB N_A_74_47#_c_104_n 0.0301504f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_30 VPB N_A_74_47#_c_105_n 0.00222785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_74_47#_c_110_n 0.00334815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_74_47#_c_107_n 0.00553539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_159_n 0.0216601f $X=-0.19 $Y=1.305 $X2=0.735 $Y2=1.695
cc_34 VPB N_VPWR_c_160_n 0.0315786f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_35 VPB N_VPWR_c_161_n 0.0299934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_158_n 0.0678959f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_37 VPB N_VPWR_c_163_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_X_c_186_n 0.0270799f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_39 VPB N_X_c_185_n 0.0225034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_A_M1004_g N_SLEEP_c_70_n 0.0152725f $X=0.705 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_41 N_A_c_44_n N_SLEEP_c_71_n 0.0144679f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_42 N_A_c_42_n N_SLEEP_c_71_n 0.0254207f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_43 N_A_c_42_n SLEEP 0.00220881f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_44 N_A_c_44_n N_A_74_47#_c_112_n 0.0181378f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_45 N_A_M1004_g N_A_74_47#_c_106_n 0.0029978f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_46 N_A_c_41_n N_A_74_47#_c_106_n 0.00498936f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_c_44_n N_A_74_47#_c_110_n 0.00641733f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_48 N_A_c_41_n N_A_74_47#_c_110_n 0.00321379f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A_M1004_g N_A_74_47#_c_107_n 0.0127069f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_50 N_A_c_44_n N_A_74_47#_c_107_n 0.00366203f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A_c_41_n N_A_74_47#_c_107_n 0.0146708f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_c_42_n N_A_74_47#_c_107_n 0.00914382f $X=0.63 $Y=0.995 $X2=0 $Y2=0
cc_53 A N_A_74_47#_c_107_n 0.0438196f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_54 N_A_c_44_n N_VPWR_c_159_n 0.00404321f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_c_44_n N_VPWR_c_160_n 0.00393512f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A_c_44_n N_VPWR_c_158_n 0.00500987f $X=0.735 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A_M1004_g N_VGND_c_214_n 0.00999374f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_58 N_A_M1004_g N_VGND_c_217_n 0.00523996f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_59 A N_VGND_c_217_n 0.00375784f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_60 N_A_M1004_g N_VGND_c_220_n 0.0106169f $X=0.705 $Y=0.445 $X2=0 $Y2=0
cc_61 A N_VGND_c_220_n 0.00623997f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 N_SLEEP_c_70_n N_A_74_47#_c_103_n 0.0104455f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_63 N_SLEEP_c_71_n N_A_74_47#_c_104_n 0.0933866f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_64 SLEEP N_A_74_47#_c_104_n 8.93818e-19 $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_65 N_SLEEP_c_71_n N_A_74_47#_c_112_n 0.0211958f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_66 SLEEP N_A_74_47#_c_112_n 0.0256006f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_67 N_SLEEP_c_71_n N_A_74_47#_c_105_n 0.00298692f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_68 SLEEP N_A_74_47#_c_105_n 0.0162172f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_69 N_SLEEP_c_71_n N_A_74_47#_c_110_n 7.45465e-19 $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_70 N_SLEEP_c_70_n N_A_74_47#_c_107_n 5.86455e-19 $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_71 N_SLEEP_c_71_n N_A_74_47#_c_107_n 0.00145125f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_72 SLEEP N_A_74_47#_c_107_n 0.012092f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_73 N_SLEEP_c_71_n N_VPWR_c_159_n 0.0168582f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_74 N_SLEEP_c_71_n N_VPWR_c_161_n 0.00622633f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_75 N_SLEEP_c_71_n N_VPWR_c_158_n 0.0103479f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_76 N_SLEEP_c_70_n N_X_c_188_n 0.00435905f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_77 N_SLEEP_c_70_n N_X_c_189_n 0.00230643f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_78 N_SLEEP_c_71_n N_X_c_189_n 0.00281723f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_79 SLEEP N_X_c_189_n 0.00634126f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_80 N_SLEEP_c_71_n N_X_c_186_n 0.00185364f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_81 N_SLEEP_c_70_n N_VGND_c_214_n 0.00315458f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_82 N_SLEEP_c_71_n N_VGND_c_214_n 0.00174997f $X=1.325 $Y=1.41 $X2=0 $Y2=0
cc_83 SLEEP N_VGND_c_214_n 0.00876939f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_84 N_SLEEP_c_70_n N_VGND_c_219_n 0.00541359f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_85 N_SLEEP_c_70_n N_VGND_c_220_n 0.00993085f $X=1.24 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_74_47#_c_112_n N_VPWR_M1005_d 0.0094087f $X=1.635 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_74_47#_c_104_n N_VPWR_c_159_n 0.00276341f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_74_47#_c_112_n N_VPWR_c_159_n 0.0214349f $X=1.635 $Y=1.595 $X2=0 $Y2=0
cc_89 N_A_74_47#_c_110_n N_VPWR_c_159_n 0.00283786f $X=0.545 $Y=1.595 $X2=0
+ $Y2=0
cc_90 N_A_74_47#_c_104_n N_VPWR_c_161_n 0.00597712f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_74_47#_c_104_n N_VPWR_c_158_n 0.0110093f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_74_47#_c_110_n N_VPWR_c_158_n 0.0100177f $X=0.545 $Y=1.595 $X2=0 $Y2=0
cc_93 N_A_74_47#_c_112_n A_283_297# 0.00885209f $X=1.635 $Y=1.595 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_74_47#_c_103_n N_X_c_184_n 0.0114928f $X=1.71 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_74_47#_c_104_n N_X_c_184_n 0.00409998f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_74_47#_c_105_n N_X_c_184_n 0.0150383f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_74_47#_c_104_n N_X_c_186_n 0.0167848f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_74_47#_c_112_n N_X_c_186_n 0.00576463f $X=1.635 $Y=1.595 $X2=0 $Y2=0
cc_99 N_A_74_47#_c_103_n N_X_c_185_n 0.00547424f $X=1.71 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_74_47#_c_104_n N_X_c_185_n 0.0156545f $X=1.735 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_74_47#_c_105_n N_X_c_185_n 0.0381477f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_74_47#_c_112_n N_VGND_c_214_n 0.00342128f $X=1.635 $Y=1.595 $X2=0
+ $Y2=0
cc_103 N_A_74_47#_c_106_n N_VGND_c_214_n 0.0103589f $X=0.585 $Y=0.457 $X2=0
+ $Y2=0
cc_104 N_A_74_47#_c_107_n N_VGND_c_214_n 0.0199064f $X=0.545 $Y=1.51 $X2=0 $Y2=0
cc_105 N_A_74_47#_c_103_n N_VGND_c_216_n 0.00482545f $X=1.71 $Y=0.995 $X2=0
+ $Y2=0
cc_106 N_A_74_47#_c_106_n N_VGND_c_217_n 0.011702f $X=0.585 $Y=0.457 $X2=0 $Y2=0
cc_107 N_A_74_47#_c_103_n N_VGND_c_219_n 0.00426565f $X=1.71 $Y=0.995 $X2=0
+ $Y2=0
cc_108 N_A_74_47#_M1004_s N_VGND_c_220_n 0.00223287f $X=0.37 $Y=0.235 $X2=0
+ $Y2=0
cc_109 N_A_74_47#_c_103_n N_VGND_c_220_n 0.00681333f $X=1.71 $Y=0.995 $X2=0
+ $Y2=0
cc_110 N_A_74_47#_c_106_n N_VGND_c_220_n 0.0117059f $X=0.585 $Y=0.457 $X2=0
+ $Y2=0
cc_111 N_VPWR_c_158_n A_283_297# 0.00983149f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_112 N_VPWR_c_158_n N_X_M1003_d 0.00217517f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_113 N_VPWR_c_159_n N_X_c_186_n 0.019448f $X=1.09 $Y=2 $X2=0 $Y2=0
cc_114 N_VPWR_c_161_n N_X_c_186_n 0.0293798f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_c_158_n N_X_c_186_n 0.0168383f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_116 N_X_c_184_n N_VGND_M1000_d 0.00773123f $X=2.025 $Y=0.73 $X2=0 $Y2=0
cc_117 N_X_c_185_n N_VGND_M1000_d 0.00108192f $X=1.98 $Y=1.85 $X2=0 $Y2=0
cc_118 N_X_c_184_n N_VGND_c_215_n 0.00139619f $X=2.025 $Y=0.73 $X2=0 $Y2=0
cc_119 N_X_c_184_n N_VGND_c_216_n 0.0233163f $X=2.025 $Y=0.73 $X2=0 $Y2=0
cc_120 N_X_c_188_n N_VGND_c_219_n 0.0202096f $X=1.47 $Y=0.39 $X2=0 $Y2=0
cc_121 N_X_c_184_n N_VGND_c_219_n 0.00257305f $X=2.025 $Y=0.73 $X2=0 $Y2=0
cc_122 N_X_M1002_d N_VGND_c_220_n 0.0025535f $X=1.315 $Y=0.235 $X2=0 $Y2=0
cc_123 N_X_c_188_n N_VGND_c_220_n 0.0131301f $X=1.47 $Y=0.39 $X2=0 $Y2=0
cc_124 N_X_c_184_n N_VGND_c_220_n 0.00759144f $X=2.025 $Y=0.73 $X2=0 $Y2=0
