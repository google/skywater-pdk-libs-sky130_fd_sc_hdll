* File: sky130_fd_sc_hdll__inputiso1p_1.spice
* Created: Wed Sep  2 08:32:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__inputiso1p_1.pex.spice"
.subckt sky130_fd_sc_hdll__inputiso1p_1  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_A_44_297#_M1000_d N_A_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_SLEEP_M1003_g N_A_44_297#_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0869439 AS=0.0567 PD=0.812523 PS=0.69 NRD=30 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_44_297#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2405 AS=0.134556 PD=2.04 PS=1.25748 NRD=19.38 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1004 A_134_297# N_A_M1004_g N_A_44_297#_M1004_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=42.1974 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1001_d N_SLEEP_M1001_g A_134_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.0609 PD=0.801549 PS=0.71 NRD=35.1645 NRS=42.1974 M=1
+ R=2.33333 SA=90000.6 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1005 N_X_M1005_d N_A_44_297#_M1005_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.41 AS=0.215282 PD=2.82 PS=1.90845 NRD=28.565 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.3 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
c_136 A_134_297# 0 1.05122e-19 $X=0.67 $Y=1.485
*
.include "sky130_fd_sc_hdll__inputiso1p_1.pxi.spice"
*
.ends
*
*
