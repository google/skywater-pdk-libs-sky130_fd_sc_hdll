* File: sky130_fd_sc_hdll__a2bb2oi_4.pex.spice
* Created: Wed Sep  2 08:19:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 26 27 28 29 31 36 48 52
c127 48 0 1.66018e-19 $X=1.435 $Y=1.202
c128 31 0 1.41039e-20 $X=3.76 $Y=1.16
c129 19 0 1.43816e-19 $X=3.785 $Y=1.41
c130 16 0 8.27827e-20 $X=1.46 $Y=0.995
r131 48 49 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r132 46 48 12.8877 $w=3.74e-07 $l=1e-07 $layer=POLY_cond $X=1.335 $Y=1.202
+ $X2=1.435 $Y2=1.202
r133 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.335
+ $Y=1.16 $X2=1.335 $Y2=1.16
r134 44 46 47.6845 $w=3.74e-07 $l=3.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.335 $Y2=1.202
r135 43 44 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r136 42 47 41.1948 $w=2.08e-07 $l=7.8e-07 $layer=LI1_cond $X=0.555 $Y=1.18
+ $X2=1.335 $Y2=1.18
r137 41 43 49.6176 $w=3.74e-07 $l=3.85e-07 $layer=POLY_cond $X=0.555 $Y=1.202
+ $X2=0.94 $Y2=1.202
r138 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.555
+ $Y=1.16 $X2=0.555 $Y2=1.16
r139 39 41 7.73262 $w=3.74e-07 $l=6e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.555 $Y2=1.202
r140 38 39 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r141 36 42 16.9004 $w=2.08e-07 $l=3.2e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.555 $Y2=1.18
r142 36 52 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.23 $Y2=1.18
r143 31 34 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.785 $Y=1.16
+ $X2=3.785 $Y2=1.53
r144 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.76
+ $Y=1.16 $X2=3.76 $Y2=1.16
r145 29 47 10.5628 $w=2.08e-07 $l=2e-07 $layer=LI1_cond $X=1.535 $Y=1.18
+ $X2=1.335 $Y2=1.18
r146 27 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.595 $Y=1.53
+ $X2=3.785 $Y2=1.53
r147 27 28 123.305 $w=1.68e-07 $l=1.89e-06 $layer=LI1_cond $X=3.595 $Y=1.53
+ $X2=1.705 $Y2=1.53
r148 26 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.62 $Y=1.445
+ $X2=1.705 $Y2=1.53
r149 25 29 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.62 $Y=1.285
+ $X2=1.535 $Y2=1.18
r150 25 26 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.62 $Y=1.285
+ $X2=1.62 $Y2=1.445
r151 22 32 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.785 $Y2=1.16
r152 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r153 19 32 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.16
r154 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r155 16 49 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r156 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r157 13 48 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r158 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r159 10 44 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r160 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r161 7 43 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r162 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r163 4 39 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r164 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r165 1 38 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r166 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 42
c67 38 0 1.66018e-19 $X=3.21 $Y=1.16
c68 1 0 1.79953e-19 $X=1.88 $Y=0.995
r69 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.34 $Y2=1.202
r70 37 39 13.6048 $w=3.72e-07 $l=1.05e-07 $layer=POLY_cond $X=3.21 $Y=1.202
+ $X2=3.315 $Y2=1.202
r71 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.21
+ $Y=1.16 $X2=3.21 $Y2=1.16
r72 35 37 47.293 $w=3.72e-07 $l=3.65e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.21 $Y2=1.202
r73 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r74 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r75 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r76 30 32 33.6882 $w=3.72e-07 $l=2.6e-07 $layer=POLY_cond $X=2.09 $Y=1.202
+ $X2=2.35 $Y2=1.202
r77 30 42 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.09
+ $Y=1.16 $X2=2.09 $Y2=1.16
r78 28 30 23.9704 $w=3.72e-07 $l=1.85e-07 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=2.09 $Y2=1.202
r79 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r80 25 38 37.4318 $w=1.98e-07 $l=6.75e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=3.21 $Y2=1.175
r81 25 42 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.075 $Y2=1.175
r82 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r83 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r84 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r85 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r86 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r87 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r88 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r89 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r90 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r91 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r92 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r93 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995 $X2=2.35
+ $Y2=0.56
r94 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r95 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r96 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r97 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995 $X2=1.88
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_831_21# 1 2 3 4 5 6 19 21 22 24 25 27
+ 28 30 31 33 34 36 37 39 40 42 43 52 53 54 57 59 63 65 69 73 75 79 83 85 88 89
+ 90 91 93 94 96 105
c214 28 0 1.0864e-19 $X=4.725 $Y=1.41
r215 105 106 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.69 $Y2=1.202
r216 102 103 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.202
+ $X2=5.195 $Y2=1.202
r217 101 102 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=5.17 $Y2=1.202
r218 98 99 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.7 $Y2=1.202
r219 97 98 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r220 87 88 19.5029 $w=3.23e-07 $l=5.5e-07 $layer=LI1_cond $X=10.297 $Y=0.905
+ $X2=10.297 $Y2=1.455
r221 86 94 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=9.875 $Y=0.82
+ $X2=9.685 $Y2=0.815
r222 85 87 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=10.135 $Y=0.82
+ $X2=10.297 $Y2=0.905
r223 85 86 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=10.135 $Y=0.82
+ $X2=9.875 $Y2=0.82
r224 84 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.835 $Y=1.54
+ $X2=9.71 $Y2=1.54
r225 83 88 7.72402 $w=1.7e-07 $l=2.00035e-07 $layer=LI1_cond $X=10.135 $Y=1.54
+ $X2=10.297 $Y2=1.455
r226 83 84 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=10.135 $Y=1.54
+ $X2=9.835 $Y2=1.54
r227 77 94 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=9.685 $Y=0.725
+ $X2=9.685 $Y2=0.815
r228 77 79 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.685 $Y=0.725
+ $X2=9.685 $Y2=0.39
r229 76 91 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.935 $Y=0.815
+ $X2=8.745 $Y2=0.815
r230 75 94 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=9.495 $Y=0.815
+ $X2=9.685 $Y2=0.815
r231 75 76 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=9.495 $Y=0.815
+ $X2=8.935 $Y2=0.815
r232 74 93 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.895 $Y=1.54
+ $X2=8.77 $Y2=1.54
r233 73 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.585 $Y=1.54
+ $X2=9.71 $Y2=1.54
r234 73 74 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.585 $Y=1.54
+ $X2=8.895 $Y2=1.54
r235 67 91 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=8.745 $Y=0.725
+ $X2=8.745 $Y2=0.815
r236 67 69 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.745 $Y=0.725
+ $X2=8.745 $Y2=0.39
r237 66 90 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.995 $Y=0.815
+ $X2=7.805 $Y2=0.815
r238 65 91 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.555 $Y=0.815
+ $X2=8.745 $Y2=0.815
r239 65 66 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.555 $Y=0.815
+ $X2=7.995 $Y2=0.815
r240 61 90 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.805 $Y=0.725
+ $X2=7.805 $Y2=0.815
r241 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.805 $Y=0.725
+ $X2=7.805 $Y2=0.39
r242 60 89 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=6.865 $Y2=0.815
r243 59 90 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.615 $Y=0.815
+ $X2=7.805 $Y2=0.815
r244 59 60 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.615 $Y=0.815
+ $X2=7.055 $Y2=0.815
r245 55 89 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.815
r246 55 57 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.39
r247 53 89 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=6.675 $Y=0.82
+ $X2=6.865 $Y2=0.815
r248 53 54 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=6.675 $Y=0.82
+ $X2=6.325 $Y2=0.82
r249 51 54 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.24 $Y=0.905
+ $X2=6.325 $Y2=0.82
r250 51 52 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.24 $Y=0.905
+ $X2=6.24 $Y2=1.075
r251 50 105 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=5.495 $Y=1.202
+ $X2=5.665 $Y2=1.202
r252 50 103 38.871 $w=3.72e-07 $l=3e-07 $layer=POLY_cond $X=5.495 $Y=1.202
+ $X2=5.195 $Y2=1.202
r253 49 50 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.16 $X2=5.495 $Y2=1.16
r254 46 101 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=4.715 $Y=1.202
+ $X2=4.725 $Y2=1.202
r255 46 99 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=4.715 $Y=1.202
+ $X2=4.7 $Y2=1.202
r256 45 49 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.715 $Y=1.16
+ $X2=5.495 $Y2=1.16
r257 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.715
+ $Y=1.16 $X2=4.715 $Y2=1.16
r258 43 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.155 $Y=1.16
+ $X2=6.24 $Y2=1.075
r259 43 49 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=6.155 $Y=1.16
+ $X2=5.495 $Y2=1.16
r260 40 106 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r261 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r262 37 105 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r263 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r264 34 103 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r265 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r266 31 102 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.202
r267 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.56
r268 28 101 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r269 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r270 25 99 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=1.202
r271 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=0.56
r272 22 98 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r273 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r274 19 97 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r275 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.56
r276 6 96 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.565
+ $Y=1.485 $X2=9.71 $Y2=1.62
r277 5 93 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.625
+ $Y=1.485 $X2=8.77 $Y2=1.62
r278 4 79 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.525
+ $Y=0.235 $X2=9.71 $Y2=0.39
r279 3 69 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.585
+ $Y=0.235 $X2=8.77 $Y2=0.39
r280 2 63 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.645
+ $Y=0.235 $X2=7.83 $Y2=0.39
r281 1 57 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A1_N 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 36 39 42
r81 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.065 $Y=1.202
+ $X2=8.09 $Y2=1.202
r82 38 39 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=7.595 $Y=1.202
+ $X2=8.065 $Y2=1.202
r83 37 38 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.57 $Y=1.202
+ $X2=7.595 $Y2=1.202
r84 35 37 7.12634 $w=3.72e-07 $l=5.5e-08 $layer=POLY_cond $X=7.515 $Y=1.202
+ $X2=7.57 $Y2=1.202
r85 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.515
+ $Y=1.16 $X2=7.515 $Y2=1.16
r86 33 35 50.5323 $w=3.72e-07 $l=3.9e-07 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.515 $Y2=1.202
r87 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r88 30 32 47.293 $w=3.72e-07 $l=3.65e-07 $layer=POLY_cond $X=6.735 $Y=1.202
+ $X2=7.1 $Y2=1.202
r89 30 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.735
+ $Y=1.16 $X2=6.735 $Y2=1.16
r90 28 30 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.735 $Y2=1.202
r91 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r92 25 36 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=7.13 $Y=1.175
+ $X2=7.515 $Y2=1.175
r93 25 42 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=7.13 $Y=1.175
+ $X2=6.695 $Y2=1.175
r94 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.09 $Y=0.995
+ $X2=8.09 $Y2=1.202
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.09 $Y=0.995
+ $X2=8.09 $Y2=0.56
r96 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.202
r97 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.065 $Y=1.41
+ $X2=8.065 $Y2=1.985
r98 16 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.202
r99 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.595 $Y=1.41
+ $X2=7.595 $Y2=1.985
r100 13 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r101 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r102 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r103 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r104 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r105 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995 $X2=7.1
+ $Y2=0.56
r106 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r107 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r108 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r109 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A2_N 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 44
r76 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.945 $Y=1.202
+ $X2=9.97 $Y2=1.202
r77 37 39 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=9.775 $Y=1.202
+ $X2=9.945 $Y2=1.202
r78 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.775
+ $Y=1.16 $X2=9.775 $Y2=1.16
r79 35 37 38.871 $w=3.72e-07 $l=3e-07 $layer=POLY_cond $X=9.475 $Y=1.202
+ $X2=9.775 $Y2=1.202
r80 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.45 $Y=1.202
+ $X2=9.475 $Y2=1.202
r81 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=9.005 $Y=1.202
+ $X2=9.45 $Y2=1.202
r82 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.98 $Y=1.202
+ $X2=9.005 $Y2=1.202
r83 31 44 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=8.605 $Y=1.175
+ $X2=8.725 $Y2=1.175
r84 30 32 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=8.605 $Y=1.202
+ $X2=8.98 $Y2=1.202
r85 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.605
+ $Y=1.16 $X2=8.605 $Y2=1.16
r86 28 30 9.06989 $w=3.72e-07 $l=7e-08 $layer=POLY_cond $X=8.535 $Y=1.202
+ $X2=8.605 $Y2=1.202
r87 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.51 $Y=1.202
+ $X2=8.535 $Y2=1.202
r88 25 38 43.2545 $w=1.98e-07 $l=7.8e-07 $layer=LI1_cond $X=8.995 $Y=1.175
+ $X2=9.775 $Y2=1.175
r89 25 44 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=8.995 $Y=1.175
+ $X2=8.725 $Y2=1.175
r90 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.97 $Y=0.995
+ $X2=9.97 $Y2=1.202
r91 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.97 $Y=0.995
+ $X2=9.97 $Y2=0.56
r92 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.202
r93 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.985
r94 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.202
r95 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.985
r96 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.45 $Y=0.995
+ $X2=9.45 $Y2=1.202
r97 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.45 $Y=0.995
+ $X2=9.45 $Y2=0.56
r98 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.202
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.985
r100 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.98 $Y=0.995
+ $X2=8.98 $Y2=1.202
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.98 $Y=0.995
+ $X2=8.98 $Y2=0.56
r102 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.202
r103 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.985
r104 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.51 $Y=0.995
+ $X2=8.51 $Y2=1.202
r105 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.51 $Y=0.995
+ $X2=8.51 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_27_297# 1 2 3 4 5 6 7 24 28 29 30 34
+ 38 42 44 46 47 50 52 54 56 61 63 65 68
c101 44 0 1.43816e-19 $X=4.02 $Y=1.965
r102 54 70 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.875 $Y=2.295
+ $X2=5.875 $Y2=2.38
r103 54 56 19.5612 $w=3.78e-07 $l=6.45e-07 $layer=LI1_cond $X=5.875 $Y=2.295
+ $X2=5.875 $Y2=1.65
r104 53 68 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.075 $Y=2.38
+ $X2=4.955 $Y2=2.38
r105 52 70 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.685 $Y=2.38
+ $X2=5.875 $Y2=2.38
r106 52 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.685 $Y=2.38
+ $X2=5.075 $Y2=2.38
r107 48 68 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.955 $Y=2.295
+ $X2=4.955 $Y2=2.38
r108 48 50 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=4.955 $Y=2.295
+ $X2=4.955 $Y2=1.96
r109 46 68 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=4.835 $Y=2.38
+ $X2=4.955 $Y2=2.38
r110 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.835 $Y=2.38
+ $X2=4.145 $Y2=2.38
r111 45 47 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.02 $Y=2.295
+ $X2=4.145 $Y2=2.38
r112 44 67 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=1.965
+ $X2=4.02 $Y2=1.88
r113 44 45 15.2122 $w=2.48e-07 $l=3.3e-07 $layer=LI1_cond $X=4.02 $Y=1.965
+ $X2=4.02 $Y2=2.295
r114 43 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=1.88
+ $X2=3.08 $Y2=1.88
r115 42 67 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=1.88
+ $X2=4.02 $Y2=1.88
r116 42 43 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=1.88
+ $X2=3.205 $Y2=1.88
r117 39 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=1.88
+ $X2=2.14 $Y2=1.88
r118 38 65 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=1.88
+ $X2=3.08 $Y2=1.88
r119 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=1.88
+ $X2=2.265 $Y2=1.88
r120 35 61 2.60907 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.315 $Y=1.88
+ $X2=1.195 $Y2=1.88
r121 34 63 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=1.88
+ $X2=2.14 $Y2=1.88
r122 34 35 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.015 $Y=1.88
+ $X2=1.315 $Y2=1.88
r123 31 61 3.84343 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=1.795
+ $X2=1.195 $Y2=1.88
r124 30 59 2.93484 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=1.625
+ $X2=1.195 $Y2=1.54
r125 30 31 8.16314 $w=2.38e-07 $l=1.7e-07 $layer=LI1_cond $X=1.195 $Y=1.625
+ $X2=1.195 $Y2=1.795
r126 28 59 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=1.195 $Y2=1.54
r127 28 29 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=0.425 $Y2=1.54
r128 24 26 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.65
+ $X2=0.255 $Y2=2.33
r129 22 29 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.425 $Y2=1.54
r130 22 24 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=0.255 $Y=1.625
+ $X2=0.255 $Y2=1.65
r131 7 70 400 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2.33
r132 7 56 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.65
r133 6 50 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.96
r134 5 67 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.96
r135 4 65 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.96
r136 3 63 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r137 2 61 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r138 2 59 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.62
r139 1 26 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.33
r140 1 24 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VPWR 1 2 3 4 5 6 23 25 29 31 35 37 41 45
+ 49 52 53 55 56 57 73 74 77 80 83 86 89
r146 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r147 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r148 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r149 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r150 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r151 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r152 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r153 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r154 71 74 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r155 70 73 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r156 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r157 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r158 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r159 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r160 64 65 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r161 62 65 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=6.67 $Y2=2.72
r162 62 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r163 61 64 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=6.67 $Y2=2.72
r164 61 62 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r165 59 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.55 $Y2=2.72
r166 59 61 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.91 $Y2=2.72
r167 57 78 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r168 57 89 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r169 55 67 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.59 $Y2=2.72
r170 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.705 $Y=2.72
+ $X2=7.83 $Y2=2.72
r171 54 70 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.955 $Y=2.72
+ $X2=8.05 $Y2=2.72
r172 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.955 $Y=2.72
+ $X2=7.83 $Y2=2.72
r173 52 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.67 $Y2=2.72
r174 52 53 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.805 $Y=2.72
+ $X2=6.91 $Y2=2.72
r175 51 67 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=7.59 $Y2=2.72
r176 51 53 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.015 $Y=2.72
+ $X2=6.91 $Y2=2.72
r177 47 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.83 $Y=2.635
+ $X2=7.83 $Y2=2.72
r178 47 49 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=7.83 $Y=2.635
+ $X2=7.83 $Y2=1.96
r179 43 53 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=2.635
+ $X2=6.91 $Y2=2.72
r180 43 45 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=6.91 $Y=2.635
+ $X2=6.91 $Y2=1.96
r181 39 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r182 39 41 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.3
r183 38 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=2.61 $Y2=2.72
r184 37 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.55 $Y2=2.72
r185 37 38 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=2.735 $Y2=2.72
r186 33 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.72
r187 33 35 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.3
r188 32 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.67 $Y2=2.72
r189 31 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.61 $Y2=2.72
r190 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=1.795 $Y2=2.72
r191 27 80 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r192 27 29 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.3
r193 26 77 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.75 $Y2=2.72
r194 25 80 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=1.67 $Y2=2.72
r195 25 26 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=0.855 $Y2=2.72
r196 21 77 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r197 21 23 35.6493 $w=2.08e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r198 6 49 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.685
+ $Y=1.485 $X2=7.83 $Y2=1.96
r199 5 45 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.96
r200 4 41 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.3
r201 3 35 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r202 2 29 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r203 1 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%Y 1 2 3 4 5 6 19 25 28 31 35 37 38 40 42
+ 46 48 49 53 54 60
c97 28 0 9.45358e-20 $X=4.255 $Y=1.415
c98 19 0 8.27827e-20 $X=3.165 $Y=0.775
r99 54 60 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=5.38 $Y=1.87
+ $X2=5.38 $Y2=1.62
r100 53 60 1.83974 $w=4.38e-07 $l=5e-09 $layer=LI1_cond $X=5.38 $Y=1.615
+ $X2=5.38 $Y2=1.62
r101 44 46 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.405 $Y=0.725
+ $X2=5.405 $Y2=0.39
r102 43 49 4.73265 $w=1.8e-07 $l=2.55e-07 $layer=LI1_cond $X=4.655 $Y=0.815
+ $X2=4.4 $Y2=0.815
r103 42 44 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.215 $Y=0.815
+ $X2=5.405 $Y2=0.725
r104 42 43 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=0.815
+ $X2=4.655 $Y2=0.815
r105 38 40 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=4.615 $Y=1.515
+ $X2=4.835 $Y2=1.515
r106 37 53 4.0299 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=5.245 $Y=1.515
+ $X2=5.38 $Y2=1.515
r107 37 40 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=5.245 $Y=1.515
+ $X2=4.835 $Y2=1.515
r108 33 38 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=4.49 $Y=1.515
+ $X2=4.615 $Y2=1.515
r109 33 50 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=4.49 $Y=1.515
+ $X2=4.255 $Y2=1.515
r110 33 35 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.62
r111 29 49 1.65197 $w=3.8e-07 $l=1.1811e-07 $layer=LI1_cond $X=4.465 $Y=0.725
+ $X2=4.4 $Y2=0.815
r112 29 31 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.465 $Y=0.725
+ $X2=4.465 $Y2=0.39
r113 28 50 0.126616 $w=2.2e-07 $l=1e-07 $layer=LI1_cond $X=4.255 $Y=1.415
+ $X2=4.255 $Y2=1.515
r114 27 49 1.65197 $w=2.2e-07 $l=1.84594e-07 $layer=LI1_cond $X=4.255 $Y=0.905
+ $X2=4.4 $Y2=0.815
r115 27 28 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=4.255 $Y=0.905
+ $X2=4.255 $Y2=1.415
r116 25 49 4.73265 $w=1.8e-07 $l=2.55e-07 $layer=LI1_cond $X=4.145 $Y=0.815
+ $X2=4.4 $Y2=0.815
r117 25 48 52.3737 $w=1.78e-07 $l=8.5e-07 $layer=LI1_cond $X=4.145 $Y=0.815
+ $X2=3.295 $Y2=0.815
r118 21 24 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=0.775
+ $X2=3.08 $Y2=0.775
r119 19 48 6.86404 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=3.165 $Y=0.775
+ $X2=3.295 $Y2=0.775
r120 19 24 3.7676 $w=2.58e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0.775
+ $X2=3.08 $Y2=0.775
r121 6 60 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.62
r122 5 35 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
r123 4 46 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.39
r124 3 31 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.39
r125 2 24 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.73
r126 1 21 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_1259_297# 1 2 3 4 5 18 22 23 26 28 30
+ 31 32 36 40 43 49
r68 38 40 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.185 $Y=2.295
+ $X2=10.185 $Y2=1.96
r69 37 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.365 $Y=2.38
+ $X2=9.24 $Y2=2.38
r70 36 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.06 $Y=2.38
+ $X2=10.185 $Y2=2.295
r71 36 37 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=10.06 $Y=2.38
+ $X2=9.365 $Y2=2.38
r72 33 47 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.425 $Y=2.38
+ $X2=8.3 $Y2=2.38
r73 32 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.115 $Y=2.38
+ $X2=9.24 $Y2=2.38
r74 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.115 $Y=2.38
+ $X2=8.425 $Y2=2.38
r75 31 47 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=2.295 $X2=8.3
+ $Y2=2.38
r76 30 45 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=1.625 $X2=8.3
+ $Y2=1.54
r77 30 31 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.3 $Y=1.625 $X2=8.3
+ $Y2=2.295
r78 29 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.48 $Y=1.54 $X2=7.36
+ $Y2=1.54
r79 28 45 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.175 $Y=1.54
+ $X2=8.3 $Y2=1.54
r80 28 29 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.175 $Y=1.54
+ $X2=7.48 $Y2=1.54
r81 24 43 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=1.625
+ $X2=7.36 $Y2=1.54
r82 24 26 32.4125 $w=2.38e-07 $l=6.75e-07 $layer=LI1_cond $X=7.36 $Y=1.625
+ $X2=7.36 $Y2=2.3
r83 22 43 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=7.24 $Y=1.54 $X2=7.36
+ $Y2=1.54
r84 22 23 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=7.24 $Y=1.54
+ $X2=6.585 $Y2=1.54
r85 18 20 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.42 $Y=1.65
+ $X2=6.42 $Y2=2.33
r86 16 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.42 $Y=1.625
+ $X2=6.585 $Y2=1.54
r87 16 18 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=6.42 $Y=1.625
+ $X2=6.42 $Y2=1.65
r88 5 40 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.035
+ $Y=1.485 $X2=10.18 $Y2=1.96
r89 4 49 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.095
+ $Y=1.485 $X2=9.24 $Y2=2.3
r90 3 47 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=2.3
r91 3 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.155
+ $Y=1.485 $X2=8.3 $Y2=1.62
r92 2 43 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.62
r93 2 26 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.3
r94 1 20 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.485 $X2=6.42 $Y2=2.33
r95 1 18 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.485 $X2=6.42 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VGND 1 2 3 4 5 6 7 8 9 28 30 32 36 40 44
+ 48 52 56 60 63 64 66 67 69 70 72 73 75 76 78 79 80 110 111 117 122 125
r165 124 125 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.235
+ $X2=6.505 $Y2=0.235
r166 120 124 3.92463 $w=6.38e-07 $l=2.1e-07 $layer=LI1_cond $X=6.21 $Y=0.235
+ $X2=6.42 $Y2=0.235
r167 120 122 14.7153 $w=6.38e-07 $l=3.95e-07 $layer=LI1_cond $X=6.21 $Y=0.235
+ $X2=5.815 $Y2=0.235
r168 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r169 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r170 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r171 108 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r172 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r173 105 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r174 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r175 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r176 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r177 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r178 99 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r179 98 125 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=7.13 $Y=0
+ $X2=6.505 $Y2=0
r180 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r181 95 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r182 94 122 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=5.815 $Y2=0
r183 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r184 91 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r185 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r186 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r187 87 88 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r188 85 88 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r189 85 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=1.15 $Y2=0
r190 84 87 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=3.91
+ $Y2=0
r191 84 85 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r192 82 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r193 82 84 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.285 $Y=0
+ $X2=1.61 $Y2=0
r194 80 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r195 80 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r196 78 107 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=9.89 $Y2=0
r197 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.095 $Y=0
+ $X2=10.18 $Y2=0
r198 77 110 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=0
+ $X2=10.35 $Y2=0
r199 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=0
+ $X2=10.18 $Y2=0
r200 75 104 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.155 $Y=0
+ $X2=8.97 $Y2=0
r201 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.155 $Y=0 $X2=9.24
+ $Y2=0
r202 74 107 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=9.325 $Y=0
+ $X2=9.89 $Y2=0
r203 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.325 $Y=0 $X2=9.24
+ $Y2=0
r204 72 101 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.215 $Y=0
+ $X2=8.05 $Y2=0
r205 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.215 $Y=0 $X2=8.3
+ $Y2=0
r206 71 104 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=8.385 $Y=0
+ $X2=8.97 $Y2=0
r207 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.385 $Y=0 $X2=8.3
+ $Y2=0
r208 69 98 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r209 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.36
+ $Y2=0
r210 68 101 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=8.05 $Y2=0
r211 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.36
+ $Y2=0
r212 66 90 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=0 $X2=4.83
+ $Y2=0
r213 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0 $X2=4.96
+ $Y2=0
r214 65 94 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.75 $Y2=0
r215 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0 $X2=4.96
+ $Y2=0
r216 63 87 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=3.91
+ $Y2=0
r217 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=4.02
+ $Y2=0
r218 62 90 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.105 $Y=0
+ $X2=4.83 $Y2=0
r219 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.02
+ $Y2=0
r220 58 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0
r221 58 60 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0.39
r222 54 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0
r223 54 56 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0.39
r224 50 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.3 $Y=0.085 $X2=8.3
+ $Y2=0
r225 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.3 $Y=0.085
+ $X2=8.3 $Y2=0.39
r226 46 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r227 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.39
r228 42 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r229 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.39
r230 38 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r231 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.39
r232 34 117 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r233 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r234 33 114 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r235 32 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r236 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.345 $Y2=0
r237 28 114 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r238 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.39
r239 9 60 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=10.045
+ $Y=0.235 $X2=10.18 $Y2=0.39
r240 8 56 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.235 $X2=9.24 $Y2=0.39
r241 7 52 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.165
+ $Y=0.235 $X2=8.3 $Y2=0.39
r242 6 48 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.39
r243 5 124 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=6.42 $Y2=0.39
r244 4 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.39
r245 3 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.39
r246 2 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.39
r247 1 30 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_109_47# 1 2 3 4 15 17 18 19 20 25
c50 20 0 1.79953e-19 $X=1.605 $Y=0.725
r51 23 25 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=2.61 $Y=0.365
+ $X2=3.55 $Y2=0.365
r52 21 28 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=1.755 $Y=0.365
+ $X2=1.605 $Y2=0.365
r53 21 23 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=1.755 $Y=0.365
+ $X2=2.61 $Y2=0.365
r54 20 30 2.76965 $w=3e-07 $l=9e-08 $layer=LI1_cond $X=1.605 $Y=0.725 $X2=1.605
+ $Y2=0.815
r55 19 28 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=1.605 $Y=0.475
+ $X2=1.605 $Y2=0.365
r56 19 20 9.60369 $w=2.98e-07 $l=2.5e-07 $layer=LI1_cond $X=1.605 $Y=0.475
+ $X2=1.605 $Y2=0.725
r57 17 30 4.61608 $w=1.8e-07 $l=1.5e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=1.605 $Y2=0.815
r58 17 18 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=0.815
+ $X2=0.895 $Y2=0.815
r59 13 18 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.895 $Y2=0.815
r60 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.705 $Y=0.725
+ $X2=0.705 $Y2=0.39
r61 4 25 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.39
r62 3 23 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.39
r63 2 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.73
r64 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.39
r65 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

