* File: sky130_fd_sc_hdll__mux2_12.pxi.spice
* Created: Wed Sep  2 08:34:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A1 N_A1_c_209_n N_A1_M1002_g N_A1_c_204_n
+ N_A1_M1016_g N_A1_c_205_n N_A1_M1040_g N_A1_c_210_n N_A1_M1026_g N_A1_c_211_n
+ N_A1_M1035_g N_A1_c_206_n N_A1_M1051_g N_A1_c_207_n N_A1_M1058_g N_A1_c_212_n
+ N_A1_M1048_g A1 N_A1_c_227_p N_A1_c_208_n PM_SKY130_FD_SC_HDLL__MUX2_12%A1
x_PM_SKY130_FD_SC_HDLL__MUX2_12%S N_S_c_299_n N_S_M1006_g N_S_c_292_n
+ N_S_M1000_g N_S_c_293_n N_S_M1020_g N_S_c_300_n N_S_M1015_g N_S_c_301_n
+ N_S_M1042_g N_S_c_294_n N_S_M1023_g N_S_c_295_n N_S_M1054_g N_S_c_302_n
+ N_S_M1056_g N_S_c_303_n N_S_M1012_g N_S_c_296_n N_S_M1038_g N_S_c_297_n
+ N_S_M1039_g N_S_c_304_n N_S_M1032_g S N_S_c_305_n N_S_c_298_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%S
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_973_297# N_A_973_297#_M1038_d
+ N_A_973_297#_M1012_s N_A_973_297#_c_422_n N_A_973_297#_M1005_g
+ N_A_973_297#_c_416_n N_A_973_297#_M1001_g N_A_973_297#_c_417_n
+ N_A_973_297#_M1009_g N_A_973_297#_c_423_n N_A_973_297#_M1029_g
+ N_A_973_297#_c_424_n N_A_973_297#_M1036_g N_A_973_297#_c_418_n
+ N_A_973_297#_M1024_g N_A_973_297#_c_419_n N_A_973_297#_M1044_g
+ N_A_973_297#_c_425_n N_A_973_297#_M1049_g N_A_973_297#_c_430_n
+ N_A_973_297#_c_434_n N_A_973_297#_c_420_n N_A_973_297#_c_439_n
+ N_A_973_297#_c_421_n PM_SKY130_FD_SC_HDLL__MUX2_12%A_973_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A0 N_A0_c_543_n N_A0_M1008_g N_A0_c_538_n
+ N_A0_M1004_g N_A0_c_539_n N_A0_M1011_g N_A0_c_544_n N_A0_M1010_g N_A0_c_545_n
+ N_A0_M1018_g N_A0_c_540_n N_A0_M1041_g N_A0_c_541_n N_A0_M1046_g N_A0_c_546_n
+ N_A0_M1030_g A0 N_A0_c_559_p N_A0_c_542_n PM_SKY130_FD_SC_HDLL__MUX2_12%A0
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_27_47# N_A_27_47#_M1016_d N_A_27_47#_M1040_d
+ N_A_27_47#_M1058_d N_A_27_47#_M1004_d N_A_27_47#_M1011_d N_A_27_47#_M1046_d
+ N_A_27_47#_M1002_d N_A_27_47#_M1026_d N_A_27_47#_M1048_d N_A_27_47#_M1008_s
+ N_A_27_47#_M1010_s N_A_27_47#_M1030_s N_A_27_47#_c_652_n N_A_27_47#_M1003_g
+ N_A_27_47#_c_630_n N_A_27_47#_M1014_g N_A_27_47#_c_631_n N_A_27_47#_M1017_g
+ N_A_27_47#_c_653_n N_A_27_47#_M1007_g N_A_27_47#_c_654_n N_A_27_47#_M1013_g
+ N_A_27_47#_c_632_n N_A_27_47#_M1021_g N_A_27_47#_c_633_n N_A_27_47#_M1025_g
+ N_A_27_47#_c_655_n N_A_27_47#_M1019_g N_A_27_47#_c_656_n N_A_27_47#_M1022_g
+ N_A_27_47#_c_634_n N_A_27_47#_M1027_g N_A_27_47#_c_635_n N_A_27_47#_M1033_g
+ N_A_27_47#_c_657_n N_A_27_47#_M1028_g N_A_27_47#_c_658_n N_A_27_47#_M1031_g
+ N_A_27_47#_c_636_n N_A_27_47#_M1034_g N_A_27_47#_c_637_n N_A_27_47#_M1043_g
+ N_A_27_47#_c_659_n N_A_27_47#_M1037_g N_A_27_47#_c_660_n N_A_27_47#_M1045_g
+ N_A_27_47#_c_638_n N_A_27_47#_M1047_g N_A_27_47#_c_639_n N_A_27_47#_M1052_g
+ N_A_27_47#_c_661_n N_A_27_47#_M1050_g N_A_27_47#_c_662_n N_A_27_47#_M1053_g
+ N_A_27_47#_c_640_n N_A_27_47#_M1055_g N_A_27_47#_c_641_n N_A_27_47#_M1059_g
+ N_A_27_47#_c_663_n N_A_27_47#_M1057_g N_A_27_47#_c_675_n N_A_27_47#_c_736_p
+ N_A_27_47#_c_677_n N_A_27_47#_c_664_n N_A_27_47#_c_665_n N_A_27_47#_c_666_n
+ N_A_27_47#_c_667_n N_A_27_47#_c_710_n N_A_27_47#_c_829_p N_A_27_47#_c_712_n
+ N_A_27_47#_c_715_n N_A_27_47#_c_668_n N_A_27_47#_c_669_n N_A_27_47#_c_642_n
+ N_A_27_47#_c_643_n N_A_27_47#_c_671_n N_A_27_47#_c_679_n N_A_27_47#_c_1004_p
+ N_A_27_47#_c_784_p N_A_27_47#_c_644_n N_A_27_47#_c_682_n N_A_27_47#_c_645_n
+ N_A_27_47#_c_719_n N_A_27_47#_c_1108_p N_A_27_47#_c_779_p N_A_27_47#_c_646_n
+ N_A_27_47#_c_647_n N_A_27_47#_c_648_n N_A_27_47#_c_690_n N_A_27_47#_c_649_n
+ N_A_27_47#_c_729_n N_A_27_47#_c_650_n N_A_27_47#_c_651_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_117_297# N_A_117_297#_M1002_s
+ N_A_117_297#_M1035_s N_A_117_297#_M1005_d N_A_117_297#_M1036_d
+ N_A_117_297#_c_1111_n N_A_117_297#_c_1145_n N_A_117_297#_c_1115_n
+ N_A_117_297#_c_1119_n N_A_117_297#_c_1149_n N_A_117_297#_c_1153_n
+ N_A_117_297#_c_1123_n N_A_117_297#_c_1126_n N_A_117_297#_c_1110_n
+ N_A_117_297#_c_1130_n N_A_117_297#_c_1161_n N_A_117_297#_c_1164_n
+ N_A_117_297#_c_1131_n N_A_117_297#_c_1134_n N_A_117_297#_c_1165_n
+ N_A_117_297#_c_1168_n N_A_117_297#_c_1169_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%A_117_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_12%VPWR N_VPWR_M1006_d N_VPWR_M1015_d
+ N_VPWR_M1056_d N_VPWR_M1032_d N_VPWR_M1029_s N_VPWR_M1049_s N_VPWR_M1003_d
+ N_VPWR_M1007_d N_VPWR_M1019_d N_VPWR_M1028_d N_VPWR_M1037_d N_VPWR_M1050_d
+ N_VPWR_M1057_d N_VPWR_c_1242_n N_VPWR_c_1243_n N_VPWR_c_1244_n N_VPWR_c_1245_n
+ N_VPWR_c_1246_n N_VPWR_c_1247_n N_VPWR_c_1248_n N_VPWR_c_1249_n
+ N_VPWR_c_1250_n N_VPWR_c_1251_n N_VPWR_c_1252_n N_VPWR_c_1253_n
+ N_VPWR_c_1254_n N_VPWR_c_1255_n N_VPWR_c_1256_n N_VPWR_c_1257_n
+ N_VPWR_c_1258_n N_VPWR_c_1259_n N_VPWR_c_1260_n N_VPWR_c_1261_n
+ N_VPWR_c_1262_n N_VPWR_c_1263_n N_VPWR_c_1264_n N_VPWR_c_1265_n
+ N_VPWR_c_1266_n VPWR N_VPWR_c_1267_n N_VPWR_c_1268_n N_VPWR_c_1269_n
+ N_VPWR_c_1270_n N_VPWR_c_1271_n N_VPWR_c_1272_n N_VPWR_c_1273_n
+ N_VPWR_c_1274_n N_VPWR_c_1241_n N_VPWR_c_1276_n N_VPWR_c_1277_n
+ N_VPWR_c_1278_n N_VPWR_c_1279_n N_VPWR_c_1280_n N_VPWR_c_1281_n
+ N_VPWR_c_1282_n VPWR PM_SKY130_FD_SC_HDLL__MUX2_12%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_597_297# N_A_597_297#_M1006_s
+ N_A_597_297#_M1042_s N_A_597_297#_M1008_d N_A_597_297#_M1018_d
+ N_A_597_297#_c_1518_n N_A_597_297#_c_1546_n N_A_597_297#_c_1522_n
+ N_A_597_297#_c_1526_n N_A_597_297#_c_1550_n N_A_597_297#_c_1554_n
+ N_A_597_297#_c_1530_n N_A_597_297#_c_1599_n N_A_597_297#_c_1514_n
+ N_A_597_297#_c_1606_n N_A_597_297#_c_1515_n N_A_597_297#_c_1516_n
+ N_A_597_297#_c_1517_n N_A_597_297#_c_1561_n N_A_597_297#_c_1564_n
+ N_A_597_297#_c_1535_n N_A_597_297#_c_1538_n N_A_597_297#_c_1565_n
+ N_A_597_297#_c_1568_n N_A_597_297#_c_1569_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%A_597_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_12%X N_X_M1014_d N_X_M1021_d N_X_M1027_d
+ N_X_M1034_d N_X_M1047_d N_X_M1055_d N_X_M1003_s N_X_M1013_s N_X_M1022_s
+ N_X_M1031_s N_X_M1045_s N_X_M1053_s N_X_c_1662_n N_X_c_1665_n N_X_c_1669_n
+ N_X_c_1652_n N_X_c_1653_n N_X_c_1680_n N_X_c_1684_n N_X_c_1688_n N_X_c_1654_n
+ N_X_c_1696_n N_X_c_1700_n N_X_c_1704_n N_X_c_1655_n N_X_c_1712_n N_X_c_1716_n
+ N_X_c_1720_n N_X_c_1656_n N_X_c_1728_n N_X_c_1732_n N_X_c_1736_n N_X_c_1657_n
+ N_X_c_1744_n N_X_c_1748_n N_X_c_1751_n N_X_c_1658_n N_X_c_1758_n N_X_c_1659_n
+ N_X_c_1766_n N_X_c_1660_n N_X_c_1774_n N_X_c_1661_n N_X_c_1782_n N_X_c_1786_n
+ N_X_c_1788_n X PM_SKY130_FD_SC_HDLL__MUX2_12%X
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_119_47# N_A_119_47#_M1016_s
+ N_A_119_47#_M1051_s N_A_119_47#_M1000_d N_A_119_47#_M1023_d
+ N_A_119_47#_c_1871_n N_A_119_47#_c_1894_n N_A_119_47#_c_1872_n
+ N_A_119_47#_c_1902_n N_A_119_47#_c_1873_n N_A_119_47#_c_1874_n
+ N_A_119_47#_c_1875_n N_A_119_47#_c_1876_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%A_119_47#
x_PM_SKY130_FD_SC_HDLL__MUX2_12%VGND N_VGND_M1000_s N_VGND_M1020_s
+ N_VGND_M1054_s N_VGND_M1039_s N_VGND_M1009_d N_VGND_M1044_d N_VGND_M1014_s
+ N_VGND_M1017_s N_VGND_M1025_s N_VGND_M1033_s N_VGND_M1043_s N_VGND_M1052_s
+ N_VGND_M1059_s N_VGND_c_1954_n N_VGND_c_1955_n N_VGND_c_1956_n N_VGND_c_1957_n
+ N_VGND_c_1958_n N_VGND_c_1959_n N_VGND_c_1960_n N_VGND_c_1961_n
+ N_VGND_c_1962_n N_VGND_c_1963_n N_VGND_c_1964_n N_VGND_c_1965_n
+ N_VGND_c_1966_n N_VGND_c_1967_n N_VGND_c_1968_n N_VGND_c_1969_n
+ N_VGND_c_1970_n N_VGND_c_1971_n N_VGND_c_1972_n N_VGND_c_1973_n
+ N_VGND_c_1974_n N_VGND_c_1975_n N_VGND_c_1976_n N_VGND_c_1977_n
+ N_VGND_c_1978_n VGND N_VGND_c_1979_n N_VGND_c_1980_n N_VGND_c_1981_n
+ N_VGND_c_1982_n N_VGND_c_1983_n N_VGND_c_1984_n N_VGND_c_1985_n
+ N_VGND_c_1986_n N_VGND_c_1987_n N_VGND_c_1988_n N_VGND_c_1989_n
+ N_VGND_c_1990_n N_VGND_c_1991_n N_VGND_c_1992_n N_VGND_c_1993_n
+ N_VGND_c_1994_n VGND PM_SKY130_FD_SC_HDLL__MUX2_12%VGND
x_PM_SKY130_FD_SC_HDLL__MUX2_12%A_1163_47# N_A_1163_47#_M1001_s
+ N_A_1163_47#_M1024_s N_A_1163_47#_M1004_s N_A_1163_47#_M1041_s
+ N_A_1163_47#_c_2225_n N_A_1163_47#_c_2218_n N_A_1163_47#_c_2219_n
+ N_A_1163_47#_c_2236_n N_A_1163_47#_c_2220_n N_A_1163_47#_c_2221_n
+ N_A_1163_47#_c_2222_n N_A_1163_47#_c_2223_n N_A_1163_47#_c_2224_n
+ PM_SKY130_FD_SC_HDLL__MUX2_12%A_1163_47#
cc_1 VNB N_A1_c_204_n 0.0190697f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A1_c_205_n 0.0167216f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A1_c_206_n 0.0167255f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_A1_c_207_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_5 VNB N_A1_c_208_n 0.0893795f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.202
cc_6 VNB N_S_c_292_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_7 VNB N_S_c_293_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_8 VNB N_S_c_294_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_9 VNB N_S_c_295_n 0.0168138f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_10 VNB N_S_c_296_n 0.0164489f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_11 VNB N_S_c_297_n 0.0166412f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_12 VNB N_S_c_298_n 0.124445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_973_297#_c_416_n 0.0170055f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_14 VNB N_A_973_297#_c_417_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_15 VNB N_A_973_297#_c_418_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_16 VNB N_A_973_297#_c_419_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_17 VNB N_A_973_297#_c_420_n 0.00229688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_973_297#_c_421_n 0.086498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A0_c_538_n 0.0214938f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_20 VNB N_A0_c_539_n 0.0167255f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_21 VNB N_A0_c_540_n 0.0167216f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_22 VNB N_A0_c_541_n 0.0190697f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_23 VNB N_A0_c_542_n 0.0902349f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.202
cc_24 VNB N_A_27_47#_c_630_n 0.0197572f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_25 VNB N_A_27_47#_c_631_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.2
cc_26 VNB N_A_27_47#_c_632_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_633_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_634_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_635_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_636_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_637_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_638_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_27_47#_c_639_n 0.0166924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_27_47#_c_640_n 0.0163356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_27_47#_c_641_n 0.020979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_642_n 0.0130155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_27_47#_c_643_n 0.00746643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_644_n 0.00282197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_645_n 0.00282197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_27_47#_c_646_n 0.00192418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_27_47#_c_647_n 0.00246701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_27_47#_c_648_n 0.00575554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_27_47#_c_649_n 0.0406332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_27_47#_c_650_n 0.0106396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_27_47#_c_651_n 0.243613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VPWR_c_1241_n 0.687231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_1652_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.2
cc_48 VNB N_X_c_1653_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_1654_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_1655_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_X_c_1656_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_X_c_1657_n 0.00392349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_1658_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_X_c_1659_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_X_c_1660_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_X_c_1661_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_119_47#_c_1871_n 0.0224565f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_58 VNB N_A_119_47#_c_1872_n 0.00498055f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_59 VNB N_A_119_47#_c_1873_n 0.00220135f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_60 VNB N_A_119_47#_c_1874_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_61 VNB N_A_119_47#_c_1875_n 0.00220135f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_62 VNB N_A_119_47#_c_1876_n 0.00222096f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.202
cc_63 VNB N_VGND_c_1954_n 0.00711369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1955_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1956_n 0.00758642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1957_n 0.00698018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1958_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1959_n 0.00711369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1960_n 0.0129285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1961_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1962_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1963_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1964_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1965_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1966_n 0.0338358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1967_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1968_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1969_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1970_n 0.00518673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1971_n 0.017949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1972_n 0.00518673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1973_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1974_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1975_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1976_n 0.00516228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1977_n 0.0621464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1978_n 0.00519006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1979_n 0.0603756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1980_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1981_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1982_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1983_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1984_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1985_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1986_n 0.0182134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1987_n 0.762505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1988_n 0.00516228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1989_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1990_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1991_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1992_n 0.00515895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1993_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1994_n 0.00519006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_1163_47#_c_2218_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_105 VNB N_A_1163_47#_c_2219_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_106 VNB N_A_1163_47#_c_2220_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=1.202
cc_107 VNB N_A_1163_47#_c_2221_n 0.0224565f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_108 VNB N_A_1163_47#_c_2222_n 0.00220135f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_109 VNB N_A_1163_47#_c_2223_n 0.00220135f $X=-0.19 $Y=-0.24 $X2=0.965
+ $Y2=1.202
cc_110 VNB N_A_1163_47#_c_2224_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=1.435
+ $Y2=1.202
cc_111 VPB N_A1_c_209_n 0.0191324f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_112 VPB N_A1_c_210_n 0.0162599f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_113 VPB N_A1_c_211_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_114 VPB N_A1_c_212_n 0.0210879f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_115 VPB N_A1_c_208_n 0.0497146f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.202
cc_116 VPB N_S_c_299_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_117 VPB N_S_c_300_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_118 VPB N_S_c_301_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_119 VPB N_S_c_302_n 0.0162591f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_120 VPB N_S_c_303_n 0.0159384f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_121 VPB N_S_c_304_n 0.0161199f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_122 VPB N_S_c_305_n 0.00687561f $X=-0.19 $Y=1.305 $X2=1.15 $Y2=1.2
cc_123 VPB N_S_c_298_n 0.0781467f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_973_297#_c_422_n 0.0164402f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.995
cc_125 VPB N_A_973_297#_c_423_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_126 VPB N_A_973_297#_c_424_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.995
cc_127 VPB N_A_973_297#_c_425_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_128 VPB N_A_973_297#_c_420_n 0.0022837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_973_297#_c_421_n 0.0492207f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A0_c_543_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_131 VPB N_A0_c_544_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_132 VPB N_A0_c_545_n 0.0162599f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_133 VPB N_A0_c_546_n 0.0191324f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_134 VPB N_A0_c_542_n 0.049789f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.202
cc_135 VPB N_A_27_47#_c_652_n 0.0196666f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_136 VPB N_A_27_47#_c_653_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_27_47#_c_654_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_27_47#_c_655_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_27_47#_c_656_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_27_47#_c_657_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_27_47#_c_658_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_27_47#_c_659_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_27_47#_c_660_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_27_47#_c_661_n 0.0162591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_27_47#_c_662_n 0.0159384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_27_47#_c_663_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_27_47#_c_664_n 0.00189756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_27_47#_c_665_n 0.007574f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_27_47#_c_666_n 0.00189756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_27_47#_c_667_n 0.00695839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_27_47#_c_668_n 0.00189756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_27_47#_c_669_n 0.0129953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_27_47#_c_642_n 0.0106155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_27_47#_c_671_n 0.00745915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_27_47#_c_647_n 2.14522e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_27_47#_c_649_n 0.0411682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_27_47#_c_651_n 0.154379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_117_297#_c_1110_n 0.0107269f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_159 VPB N_VPWR_c_1242_n 0.0126709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_1243_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_1244_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1245_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1246_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1247_n 0.0120377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1248_n 0.0131235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1249_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1250_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1251_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1252_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1253_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1254_n 0.0410796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1255_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1256_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1257_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1258_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1259_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1260_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1261_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1262_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1263_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1264_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1265_n 0.0629219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1266_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1267_n 0.0611443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1268_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1269_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1270_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1271_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1272_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1273_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1274_n 0.0182134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1241_n 0.0779009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1276_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1277_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1278_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1279_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1280_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1281_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1282_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_597_297#_c_1514_n 0.00287217f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_201 VPB N_A_597_297#_c_1515_n 0.00271682f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.202
cc_202 VPB N_A_597_297#_c_1516_n 0.00263789f $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=1.202
cc_203 VPB N_A_597_297#_c_1517_n 0.00660038f $X=-0.19 $Y=1.305 $X2=1.75
+ $Y2=1.202
cc_204 N_A1_c_209_n N_A_27_47#_c_675_n 0.0137768f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_210_n N_A_27_47#_c_675_n 0.0108728f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A1_c_211_n N_A_27_47#_c_677_n 0.0108728f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A1_c_212_n N_A_27_47#_c_677_n 0.00974411f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A1_c_204_n N_A_27_47#_c_679_n 0.00767088f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A1_c_205_n N_A_27_47#_c_679_n 0.00836606f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A1_c_208_n N_A_27_47#_c_679_n 8.08246e-19 $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_211 N_A1_c_206_n N_A_27_47#_c_682_n 0.00836606f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A1_c_207_n N_A_27_47#_c_682_n 0.00801464f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A1_c_204_n N_A_27_47#_c_648_n 0.00729564f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A1_c_205_n N_A_27_47#_c_648_n 0.00375115f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A1_c_206_n N_A_27_47#_c_648_n 0.00375115f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A1_c_207_n N_A_27_47#_c_648_n 0.00347927f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A1_c_227_p N_A_27_47#_c_648_n 0.00322221f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A1_c_208_n N_A_27_47#_c_648_n 9.46745e-19 $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A1_c_208_n N_A_27_47#_c_690_n 2.2806e-19 $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_220 N_A1_c_209_n N_A_27_47#_c_649_n 0.00329518f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A1_c_204_n N_A_27_47#_c_649_n 0.00519414f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A1_c_227_p N_A_27_47#_c_649_n 0.0206594f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_223 N_A1_c_208_n N_A_27_47#_c_649_n 0.0163098f $X=1.88 $Y=1.202 $X2=0 $Y2=0
cc_224 N_A1_c_210_n N_A_117_297#_c_1111_n 0.0106503f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A1_c_211_n N_A_117_297#_c_1111_n 0.0106503f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A1_c_227_p N_A_117_297#_c_1111_n 0.0374055f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A1_c_208_n N_A_117_297#_c_1111_n 0.00616252f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_228 N_A1_c_209_n N_A_117_297#_c_1115_n 0.00214429f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A1_c_210_n N_A_117_297#_c_1115_n 5.6422e-19 $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A1_c_227_p N_A_117_297#_c_1115_n 0.0203246f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A1_c_208_n N_A_117_297#_c_1115_n 0.00669726f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_232 N_A1_c_211_n N_A_117_297#_c_1119_n 5.6422e-19 $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A1_c_212_n N_A_117_297#_c_1119_n 0.00214429f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A1_c_227_p N_A_117_297#_c_1119_n 0.0202695f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A1_c_208_n N_A_117_297#_c_1119_n 0.00669726f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_236 N_A1_c_210_n N_A_117_297#_c_1123_n 0.00313189f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_237 N_A1_c_211_n N_A_117_297#_c_1123_n 0.00313189f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A1_c_227_p N_A_117_297#_c_1123_n 0.00107383f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_239 N_A1_c_227_p N_A_117_297#_c_1126_n 0.00117983f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_240 N_A1_c_212_n N_A_117_297#_c_1110_n 0.00600932f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A1_c_227_p N_A_117_297#_c_1110_n 0.00233931f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A1_c_208_n N_A_117_297#_c_1110_n 2.02467e-19 $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_243 N_A1_c_227_p N_A_117_297#_c_1130_n 0.00117983f $X=1.75 $Y=1.16 $X2=0
+ $Y2=0
cc_244 N_A1_c_209_n N_A_117_297#_c_1131_n 0.00532302f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A1_c_210_n N_A_117_297#_c_1131_n 0.00606957f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A1_c_211_n N_A_117_297#_c_1131_n 5.7339e-19 $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A1_c_210_n N_A_117_297#_c_1134_n 5.7339e-19 $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A1_c_211_n N_A_117_297#_c_1134_n 0.00606957f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A1_c_212_n N_A_117_297#_c_1134_n 0.00483111f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A1_c_212_n N_VPWR_c_1242_n 0.0021834f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A1_c_209_n N_VPWR_c_1267_n 0.00429453f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A1_c_210_n N_VPWR_c_1267_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A1_c_211_n N_VPWR_c_1267_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A1_c_212_n N_VPWR_c_1267_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A1_c_209_n N_VPWR_c_1241_n 0.00697643f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A1_c_210_n N_VPWR_c_1241_n 0.00600186f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A1_c_211_n N_VPWR_c_1241_n 0.00600186f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_c_212_n N_VPWR_c_1241_n 0.00728421f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_c_207_n N_A_119_47#_c_1871_n 0.0112292f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A1_c_208_n N_A_119_47#_c_1871_n 0.00224539f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_261 N_A1_c_204_n N_A_119_47#_c_1873_n 0.00440693f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A1_c_205_n N_A_119_47#_c_1873_n 0.00402996f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A1_c_206_n N_A_119_47#_c_1873_n 4.02078e-19 $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A1_c_227_p N_A_119_47#_c_1873_n 0.0974168f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A1_c_208_n N_A_119_47#_c_1873_n 0.00225271f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_266 N_A1_c_205_n N_A_119_47#_c_1874_n 0.00754011f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A1_c_206_n N_A_119_47#_c_1874_n 0.00754011f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A1_c_208_n N_A_119_47#_c_1874_n 0.00468948f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_269 N_A1_c_205_n N_A_119_47#_c_1875_n 4.02078e-19 $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_270 N_A1_c_206_n N_A_119_47#_c_1875_n 0.00402996f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_271 N_A1_c_207_n N_A_119_47#_c_1875_n 0.00716324f $X=1.88 $Y=0.995 $X2=0
+ $Y2=0
cc_272 N_A1_c_208_n N_A_119_47#_c_1875_n 0.00225271f $X=1.88 $Y=1.202 $X2=0
+ $Y2=0
cc_273 N_A1_c_207_n N_VGND_c_1954_n 0.00203215f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A1_c_204_n N_VGND_c_1979_n 0.00357877f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_205_n N_VGND_c_1979_n 0.00357877f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A1_c_206_n N_VGND_c_1979_n 0.00357877f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A1_c_207_n N_VGND_c_1979_n 0.00357877f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A1_c_204_n N_VGND_c_1987_n 0.00572883f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A1_c_205_n N_VGND_c_1987_n 0.00497228f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A1_c_206_n N_VGND_c_1987_n 0.00497228f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A1_c_207_n N_VGND_c_1987_n 0.00605604f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_282 N_S_c_304_n N_A_973_297#_c_422_n 0.00970081f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_283 N_S_c_297_n N_A_973_297#_c_416_n 0.00828698f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_284 N_S_c_295_n N_A_973_297#_c_430_n 6.09671e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_285 N_S_c_296_n N_A_973_297#_c_430_n 0.00968408f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_286 N_S_c_297_n N_A_973_297#_c_430_n 0.00968408f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_287 N_S_c_298_n N_A_973_297#_c_430_n 0.00975822f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_288 N_S_c_302_n N_A_973_297#_c_434_n 7.04702e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_289 N_S_c_303_n N_A_973_297#_c_434_n 0.0119897f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_290 N_S_c_304_n N_A_973_297#_c_434_n 0.0119897f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_291 N_S_c_298_n N_A_973_297#_c_434_n 0.00612724f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_292 N_S_c_298_n N_A_973_297#_c_420_n 0.0143164f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_293 N_S_c_305_n N_A_973_297#_c_439_n 0.00775355f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_294 N_S_c_298_n N_A_973_297#_c_439_n 0.021583f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_295 N_S_c_298_n N_A_973_297#_c_421_n 0.0210988f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_296 N_S_c_292_n N_A_27_47#_c_648_n 0.00187713f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_297 N_S_c_293_n N_A_27_47#_c_648_n 0.00192476f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_298 N_S_c_294_n N_A_27_47#_c_648_n 0.00192476f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_299 N_S_c_295_n N_A_27_47#_c_648_n 0.00465394f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_300 N_S_c_296_n N_A_27_47#_c_648_n 0.00576977f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_301 N_S_c_297_n N_A_27_47#_c_648_n 0.00241086f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_302 N_S_c_305_n N_A_27_47#_c_648_n 0.00449599f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_303 N_S_c_298_n N_A_27_47#_c_648_n 0.00116442f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_304 N_S_c_299_n N_A_117_297#_c_1110_n 0.00808847f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_S_c_300_n N_A_117_297#_c_1110_n 0.00301881f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_S_c_301_n N_A_117_297#_c_1110_n 0.00301881f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_S_c_302_n N_A_117_297#_c_1110_n 0.00705091f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_S_c_303_n N_A_117_297#_c_1110_n 0.00817858f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_309 N_S_c_304_n N_A_117_297#_c_1110_n 0.00365735f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_310 N_S_c_305_n N_A_117_297#_c_1110_n 0.00568194f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_311 N_S_c_298_n N_A_117_297#_c_1110_n 8.5765e-19 $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_312 N_S_c_299_n N_VPWR_c_1242_n 0.00374733f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_313 N_S_c_300_n N_VPWR_c_1243_n 0.00208662f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_314 N_S_c_301_n N_VPWR_c_1243_n 0.00208662f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_315 N_S_c_302_n N_VPWR_c_1244_n 0.00213628f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_316 N_S_c_303_n N_VPWR_c_1244_n 0.00213628f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_317 N_S_c_298_n N_VPWR_c_1244_n 0.00731623f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_318 N_S_c_304_n N_VPWR_c_1245_n 0.00213628f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_319 N_S_c_299_n N_VPWR_c_1255_n 0.00673617f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_320 N_S_c_300_n N_VPWR_c_1255_n 0.00673617f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_321 N_S_c_301_n N_VPWR_c_1257_n 0.00673617f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_322 N_S_c_302_n N_VPWR_c_1257_n 0.00673617f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_323 N_S_c_303_n N_VPWR_c_1259_n 0.00673617f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_324 N_S_c_304_n N_VPWR_c_1259_n 0.00673617f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_325 N_S_c_299_n N_VPWR_c_1241_n 0.00832888f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_326 N_S_c_300_n N_VPWR_c_1241_n 0.0059257f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_327 N_S_c_301_n N_VPWR_c_1241_n 0.0059257f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_328 N_S_c_302_n N_VPWR_c_1241_n 0.0059257f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_329 N_S_c_303_n N_VPWR_c_1241_n 0.0059257f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_330 N_S_c_304_n N_VPWR_c_1241_n 0.00595091f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_331 N_S_c_300_n N_A_597_297#_c_1518_n 0.00916f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_332 N_S_c_301_n N_A_597_297#_c_1518_n 0.00916f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_333 N_S_c_305_n N_A_597_297#_c_1518_n 0.0376251f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_334 N_S_c_298_n N_A_597_297#_c_1518_n 0.00169072f $X=5.22 $Y=1.202 $X2=0
+ $Y2=0
cc_335 N_S_c_299_n N_A_597_297#_c_1522_n 0.00215881f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_336 N_S_c_300_n N_A_597_297#_c_1522_n 5.7874e-19 $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_337 N_S_c_305_n N_A_597_297#_c_1522_n 0.0206325f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_338 N_S_c_298_n N_A_597_297#_c_1522_n 0.00183511f $X=5.22 $Y=1.202 $X2=0
+ $Y2=0
cc_339 N_S_c_301_n N_A_597_297#_c_1526_n 5.7874e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_340 N_S_c_302_n N_A_597_297#_c_1526_n 0.00207067f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_S_c_305_n N_A_597_297#_c_1526_n 0.0206325f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_342 N_S_c_298_n N_A_597_297#_c_1526_n 0.00183511f $X=5.22 $Y=1.202 $X2=0
+ $Y2=0
cc_343 N_S_c_300_n N_A_597_297#_c_1530_n 0.00232817f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_344 N_S_c_301_n N_A_597_297#_c_1530_n 0.00232817f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_345 N_S_c_302_n N_A_597_297#_c_1514_n 0.00272349f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_346 N_S_c_303_n N_A_597_297#_c_1514_n 0.00272349f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_S_c_304_n N_A_597_297#_c_1514_n 0.00272349f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_348 N_S_c_299_n N_A_597_297#_c_1535_n 0.00848227f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_349 N_S_c_300_n N_A_597_297#_c_1535_n 0.00912469f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_350 N_S_c_301_n N_A_597_297#_c_1535_n 7.05028e-19 $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_351 N_S_c_300_n N_A_597_297#_c_1538_n 7.05028e-19 $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_352 N_S_c_301_n N_A_597_297#_c_1538_n 0.00912469f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_353 N_S_c_302_n N_A_597_297#_c_1538_n 0.00772015f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_354 N_S_c_292_n N_A_119_47#_c_1871_n 0.013146f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_355 N_S_c_305_n N_A_119_47#_c_1871_n 0.00261569f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_356 N_S_c_298_n N_A_119_47#_c_1871_n 0.00224539f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_357 N_S_c_292_n N_A_119_47#_c_1894_n 0.0100064f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_358 N_S_c_293_n N_A_119_47#_c_1894_n 0.00627537f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_359 N_S_c_294_n N_A_119_47#_c_1894_n 6.13333e-19 $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_360 N_S_c_293_n N_A_119_47#_c_1872_n 0.00900777f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_361 N_S_c_294_n N_A_119_47#_c_1872_n 0.0101394f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_362 N_S_c_295_n N_A_119_47#_c_1872_n 0.00255406f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_363 N_S_c_305_n N_A_119_47#_c_1872_n 0.0690141f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_364 N_S_c_298_n N_A_119_47#_c_1872_n 0.00698847f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_365 N_S_c_293_n N_A_119_47#_c_1902_n 6.13333e-19 $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_366 N_S_c_294_n N_A_119_47#_c_1902_n 0.00627537f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_367 N_S_c_295_n N_A_119_47#_c_1902_n 0.00473017f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_368 N_S_c_292_n N_A_119_47#_c_1876_n 0.00113159f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_369 N_S_c_293_n N_A_119_47#_c_1876_n 0.00113159f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_370 N_S_c_305_n N_A_119_47#_c_1876_n 0.0262372f $X=3.09 $Y=1.16 $X2=0 $Y2=0
cc_371 N_S_c_298_n N_A_119_47#_c_1876_n 0.00230167f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_372 N_S_c_292_n N_VGND_c_1954_n 0.00336227f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_373 N_S_c_293_n N_VGND_c_1955_n 0.00180171f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_374 N_S_c_294_n N_VGND_c_1955_n 0.00180171f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_375 N_S_c_295_n N_VGND_c_1956_n 0.00201331f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_376 N_S_c_296_n N_VGND_c_1956_n 0.00201363f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_377 N_S_c_298_n N_VGND_c_1956_n 0.00618196f $X=5.22 $Y=1.202 $X2=0 $Y2=0
cc_378 N_S_c_297_n N_VGND_c_1957_n 0.00201363f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_379 N_S_c_292_n N_VGND_c_1967_n 0.00423334f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_380 N_S_c_293_n N_VGND_c_1967_n 0.00423334f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_381 N_S_c_294_n N_VGND_c_1969_n 0.00423334f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_382 N_S_c_295_n N_VGND_c_1969_n 0.00541359f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_383 N_S_c_296_n N_VGND_c_1971_n 0.00541359f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_384 N_S_c_297_n N_VGND_c_1971_n 0.00541359f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_385 N_S_c_292_n N_VGND_c_1987_n 0.00613629f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_386 N_S_c_293_n N_VGND_c_1987_n 0.00505254f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_387 N_S_c_294_n N_VGND_c_1987_n 0.00505254f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_388 N_S_c_295_n N_VGND_c_1987_n 0.00535118f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_389 N_S_c_296_n N_VGND_c_1987_n 0.00535118f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_390 N_S_c_297_n N_VGND_c_1987_n 0.00536223f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A_973_297#_c_416_n N_A_27_47#_c_648_n 0.00242407f $X=5.74 $Y=0.995
+ $X2=0 $Y2=0
cc_392 N_A_973_297#_c_417_n N_A_27_47#_c_648_n 0.00192476f $X=6.16 $Y=0.995
+ $X2=0 $Y2=0
cc_393 N_A_973_297#_c_418_n N_A_27_47#_c_648_n 0.00192476f $X=6.68 $Y=0.995
+ $X2=0 $Y2=0
cc_394 N_A_973_297#_c_419_n N_A_27_47#_c_648_n 0.00187713f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_395 N_A_973_297#_c_430_n N_A_27_47#_c_648_n 0.0267501f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_396 N_A_973_297#_c_420_n N_A_27_47#_c_648_n 0.0141572f $X=6.93 $Y=1.16 $X2=0
+ $Y2=0
cc_397 N_A_973_297#_c_421_n N_A_27_47#_c_648_n 0.00116442f $X=7.1 $Y=1.202 $X2=0
+ $Y2=0
cc_398 N_A_973_297#_c_423_n N_A_117_297#_c_1145_n 0.00916655f $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_399 N_A_973_297#_c_424_n N_A_117_297#_c_1145_n 0.00916655f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_400 N_A_973_297#_c_420_n N_A_117_297#_c_1145_n 0.0374055f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_401 N_A_973_297#_c_421_n N_A_117_297#_c_1145_n 0.00616252f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_402 N_A_973_297#_c_422_n N_A_117_297#_c_1149_n 0.00207151f $X=5.715 $Y=1.41
+ $X2=0 $Y2=0
cc_403 N_A_973_297#_c_423_n N_A_117_297#_c_1149_n 5.79575e-19 $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_404 N_A_973_297#_c_420_n N_A_117_297#_c_1149_n 0.020376f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_405 N_A_973_297#_c_421_n N_A_117_297#_c_1149_n 0.00671335f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_406 N_A_973_297#_c_424_n N_A_117_297#_c_1153_n 5.79575e-19 $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_407 N_A_973_297#_c_425_n N_A_117_297#_c_1153_n 0.00215964f $X=7.125 $Y=1.41
+ $X2=0 $Y2=0
cc_408 N_A_973_297#_c_420_n N_A_117_297#_c_1153_n 0.0204311f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_409 N_A_973_297#_c_421_n N_A_117_297#_c_1153_n 0.00671335f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_410 N_A_973_297#_c_422_n N_A_117_297#_c_1110_n 0.00367026f $X=5.715 $Y=1.41
+ $X2=0 $Y2=0
cc_411 N_A_973_297#_c_434_n N_A_117_297#_c_1110_n 0.0231322f $X=5.01 $Y=1.66
+ $X2=0 $Y2=0
cc_412 N_A_973_297#_c_420_n N_A_117_297#_c_1110_n 0.0107876f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_413 N_A_973_297#_c_421_n N_A_117_297#_c_1110_n 2.02467e-19 $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_414 N_A_973_297#_c_423_n N_A_117_297#_c_1161_n 0.00301881f $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_415 N_A_973_297#_c_424_n N_A_117_297#_c_1161_n 0.00301881f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_416 N_A_973_297#_c_420_n N_A_117_297#_c_1161_n 0.00107383f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_417 N_A_973_297#_c_420_n N_A_117_297#_c_1164_n 0.00117983f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_418 N_A_973_297#_c_422_n N_A_117_297#_c_1165_n 0.00772015f $X=5.715 $Y=1.41
+ $X2=0 $Y2=0
cc_419 N_A_973_297#_c_423_n N_A_117_297#_c_1165_n 0.00912469f $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_420 N_A_973_297#_c_424_n N_A_117_297#_c_1165_n 7.05028e-19 $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_421 N_A_973_297#_c_420_n N_A_117_297#_c_1168_n 0.00117983f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_422 N_A_973_297#_c_423_n N_A_117_297#_c_1169_n 7.05028e-19 $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_423 N_A_973_297#_c_424_n N_A_117_297#_c_1169_n 0.00912469f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_424 N_A_973_297#_c_425_n N_A_117_297#_c_1169_n 0.00845951f $X=7.125 $Y=1.41
+ $X2=0 $Y2=0
cc_425 N_A_973_297#_c_434_n N_VPWR_c_1244_n 0.0400362f $X=5.01 $Y=1.66 $X2=0
+ $Y2=0
cc_426 N_A_973_297#_c_422_n N_VPWR_c_1245_n 0.00213628f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_427 N_A_973_297#_c_434_n N_VPWR_c_1245_n 0.0400362f $X=5.01 $Y=1.66 $X2=0
+ $Y2=0
cc_428 N_A_973_297#_c_420_n N_VPWR_c_1245_n 0.0178233f $X=6.93 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_A_973_297#_c_423_n N_VPWR_c_1246_n 0.00208662f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_430 N_A_973_297#_c_424_n N_VPWR_c_1246_n 0.00208662f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_431 N_A_973_297#_c_425_n N_VPWR_c_1247_n 0.00374733f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_432 N_A_973_297#_c_434_n N_VPWR_c_1259_n 0.0189467f $X=5.01 $Y=1.66 $X2=0
+ $Y2=0
cc_433 N_A_973_297#_c_422_n N_VPWR_c_1261_n 0.00673617f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_434 N_A_973_297#_c_423_n N_VPWR_c_1261_n 0.00673617f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_435 N_A_973_297#_c_424_n N_VPWR_c_1263_n 0.00673617f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_436 N_A_973_297#_c_425_n N_VPWR_c_1263_n 0.00673617f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_437 N_A_973_297#_M1012_s N_VPWR_c_1241_n 0.00130534f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_A_973_297#_c_422_n N_VPWR_c_1241_n 0.00595091f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_439 N_A_973_297#_c_423_n N_VPWR_c_1241_n 0.0059257f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_440 N_A_973_297#_c_424_n N_VPWR_c_1241_n 0.0059257f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_441 N_A_973_297#_c_425_n N_VPWR_c_1241_n 0.00720805f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_442 N_A_973_297#_c_434_n N_VPWR_c_1241_n 0.00347454f $X=5.01 $Y=1.66 $X2=0
+ $Y2=0
cc_443 N_A_973_297#_c_422_n N_A_597_297#_c_1514_n 0.00272349f $X=5.715 $Y=1.41
+ $X2=0 $Y2=0
cc_444 N_A_973_297#_c_423_n N_A_597_297#_c_1514_n 0.00232817f $X=6.185 $Y=1.41
+ $X2=0 $Y2=0
cc_445 N_A_973_297#_c_424_n N_A_597_297#_c_1514_n 0.00232817f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_446 N_A_973_297#_c_425_n N_A_597_297#_c_1514_n 0.00769303f $X=7.125 $Y=1.41
+ $X2=0 $Y2=0
cc_447 N_A_973_297#_c_434_n N_A_597_297#_c_1514_n 0.0166918f $X=5.01 $Y=1.66
+ $X2=0 $Y2=0
cc_448 N_A_973_297#_c_430_n N_VGND_c_1956_n 0.0269761f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_449 N_A_973_297#_c_416_n N_VGND_c_1957_n 0.00201331f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_450 N_A_973_297#_c_430_n N_VGND_c_1957_n 0.0269761f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_451 N_A_973_297#_c_420_n N_VGND_c_1957_n 0.022484f $X=6.93 $Y=1.16 $X2=0
+ $Y2=0
cc_452 N_A_973_297#_c_417_n N_VGND_c_1958_n 0.00180171f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_453 N_A_973_297#_c_418_n N_VGND_c_1958_n 0.00180171f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_454 N_A_973_297#_c_419_n N_VGND_c_1959_n 0.00336227f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_455 N_A_973_297#_c_430_n N_VGND_c_1971_n 0.0189039f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_456 N_A_973_297#_c_416_n N_VGND_c_1973_n 0.00541359f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_457 N_A_973_297#_c_417_n N_VGND_c_1973_n 0.00423334f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A_973_297#_c_418_n N_VGND_c_1975_n 0.00423334f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A_973_297#_c_419_n N_VGND_c_1975_n 0.00423334f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_973_297#_M1038_d N_VGND_c_1987_n 0.00121469f $X=4.875 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_A_973_297#_c_416_n N_VGND_c_1987_n 0.00536223f $X=5.74 $Y=0.995 $X2=0
+ $Y2=0
cc_462 N_A_973_297#_c_417_n N_VGND_c_1987_n 0.00505254f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_463 N_A_973_297#_c_418_n N_VGND_c_1987_n 0.00505254f $X=6.68 $Y=0.995 $X2=0
+ $Y2=0
cc_464 N_A_973_297#_c_419_n N_VGND_c_1987_n 0.00613629f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_465 N_A_973_297#_c_430_n N_VGND_c_1987_n 0.00344927f $X=5.01 $Y=0.42 $X2=0
+ $Y2=0
cc_466 N_A_973_297#_c_416_n N_A_1163_47#_c_2225_n 0.00473017f $X=5.74 $Y=0.995
+ $X2=0 $Y2=0
cc_467 N_A_973_297#_c_417_n N_A_1163_47#_c_2225_n 0.00627537f $X=6.16 $Y=0.995
+ $X2=0 $Y2=0
cc_468 N_A_973_297#_c_418_n N_A_1163_47#_c_2225_n 6.13333e-19 $X=6.68 $Y=0.995
+ $X2=0 $Y2=0
cc_469 N_A_973_297#_c_417_n N_A_1163_47#_c_2218_n 0.00901269f $X=6.16 $Y=0.995
+ $X2=0 $Y2=0
cc_470 N_A_973_297#_c_418_n N_A_1163_47#_c_2218_n 0.00901269f $X=6.68 $Y=0.995
+ $X2=0 $Y2=0
cc_471 N_A_973_297#_c_420_n N_A_1163_47#_c_2218_n 0.0425393f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_472 N_A_973_297#_c_421_n N_A_1163_47#_c_2218_n 0.00468948f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_473 N_A_973_297#_c_416_n N_A_1163_47#_c_2219_n 0.00255533f $X=5.74 $Y=0.995
+ $X2=0 $Y2=0
cc_474 N_A_973_297#_c_417_n N_A_1163_47#_c_2219_n 0.00113286f $X=6.16 $Y=0.995
+ $X2=0 $Y2=0
cc_475 N_A_973_297#_c_420_n N_A_1163_47#_c_2219_n 0.026096f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_476 N_A_973_297#_c_421_n N_A_1163_47#_c_2219_n 0.00230339f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_477 N_A_973_297#_c_417_n N_A_1163_47#_c_2236_n 6.13333e-19 $X=6.16 $Y=0.995
+ $X2=0 $Y2=0
cc_478 N_A_973_297#_c_418_n N_A_1163_47#_c_2236_n 0.00627537f $X=6.68 $Y=0.995
+ $X2=0 $Y2=0
cc_479 N_A_973_297#_c_419_n N_A_1163_47#_c_2236_n 0.0100064f $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_480 N_A_973_297#_c_418_n N_A_1163_47#_c_2220_n 0.00113286f $X=6.68 $Y=0.995
+ $X2=0 $Y2=0
cc_481 N_A_973_297#_c_419_n N_A_1163_47#_c_2220_n 0.00113286f $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_482 N_A_973_297#_c_420_n N_A_1163_47#_c_2220_n 0.026096f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_483 N_A_973_297#_c_421_n N_A_1163_47#_c_2220_n 0.00230339f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_484 N_A_973_297#_c_419_n N_A_1163_47#_c_2221_n 0.0131168f $X=7.1 $Y=0.995
+ $X2=0 $Y2=0
cc_485 N_A_973_297#_c_420_n N_A_1163_47#_c_2221_n 0.00266811f $X=6.93 $Y=1.16
+ $X2=0 $Y2=0
cc_486 N_A_973_297#_c_421_n N_A_1163_47#_c_2221_n 0.00224539f $X=7.1 $Y=1.202
+ $X2=0 $Y2=0
cc_487 N_A0_c_543_n N_A_27_47#_c_710_n 0.00974411f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_488 N_A0_c_544_n N_A_27_47#_c_710_n 0.0108728f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_489 N_A0_c_540_n N_A_27_47#_c_712_n 0.00836606f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_490 N_A0_c_541_n N_A_27_47#_c_712_n 0.00767088f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_491 N_A0_c_542_n N_A_27_47#_c_712_n 8.08246e-19 $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_492 N_A0_c_545_n N_A_27_47#_c_715_n 0.0108728f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A0_c_546_n N_A_27_47#_c_715_n 0.0137768f $X=9.525 $Y=1.41 $X2=0 $Y2=0
cc_494 N_A0_c_546_n N_A_27_47#_c_669_n 0.00329518f $X=9.525 $Y=1.41 $X2=0 $Y2=0
cc_495 N_A0_c_542_n N_A_27_47#_c_669_n 0.00384727f $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_496 N_A0_c_538_n N_A_27_47#_c_719_n 0.00801464f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_497 N_A0_c_539_n N_A_27_47#_c_719_n 0.00836606f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_498 N_A0_c_559_p N_A_27_47#_c_647_n 0.0209934f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_499 N_A0_c_542_n N_A_27_47#_c_647_n 0.00841651f $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_500 N_A0_c_538_n N_A_27_47#_c_648_n 0.00347927f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_501 N_A0_c_539_n N_A_27_47#_c_648_n 0.00375115f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_502 N_A0_c_540_n N_A_27_47#_c_648_n 0.00375115f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_503 N_A0_c_541_n N_A_27_47#_c_648_n 0.00729564f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_504 N_A0_c_559_p N_A_27_47#_c_648_n 0.00322221f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_505 N_A0_c_542_n N_A_27_47#_c_648_n 9.46745e-19 $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_506 N_A0_c_542_n N_A_27_47#_c_729_n 2.2806e-19 $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_507 N_A0_c_541_n N_A_27_47#_c_650_n 0.00519414f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_508 N_A0_c_542_n N_A_27_47#_c_650_n 0.0042097f $X=9.5 $Y=1.202 $X2=0 $Y2=0
cc_509 N_A0_c_543_n N_VPWR_c_1247_n 0.0021834f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_510 N_A0_c_546_n N_VPWR_c_1248_n 0.0021834f $X=9.525 $Y=1.41 $X2=0 $Y2=0
cc_511 N_A0_c_543_n N_VPWR_c_1265_n 0.00429453f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_512 N_A0_c_544_n N_VPWR_c_1265_n 0.00429453f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_513 N_A0_c_545_n N_VPWR_c_1265_n 0.00429453f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_514 N_A0_c_546_n N_VPWR_c_1265_n 0.00429453f $X=9.525 $Y=1.41 $X2=0 $Y2=0
cc_515 N_A0_c_543_n N_VPWR_c_1241_n 0.00728421f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A0_c_544_n N_VPWR_c_1241_n 0.00600186f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A0_c_545_n N_VPWR_c_1241_n 0.00600186f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_518 N_A0_c_546_n N_VPWR_c_1241_n 0.00734734f $X=9.525 $Y=1.41 $X2=0 $Y2=0
cc_519 N_A0_c_544_n N_A_597_297#_c_1546_n 0.0106503f $X=8.585 $Y=1.41 $X2=0
+ $Y2=0
cc_520 N_A0_c_545_n N_A_597_297#_c_1546_n 0.0106503f $X=9.055 $Y=1.41 $X2=0
+ $Y2=0
cc_521 N_A0_c_559_p N_A_597_297#_c_1546_n 0.0374055f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_522 N_A0_c_542_n N_A_597_297#_c_1546_n 0.00616252f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_523 N_A0_c_543_n N_A_597_297#_c_1550_n 0.00214429f $X=8.115 $Y=1.41 $X2=0
+ $Y2=0
cc_524 N_A0_c_544_n N_A_597_297#_c_1550_n 5.6422e-19 $X=8.585 $Y=1.41 $X2=0
+ $Y2=0
cc_525 N_A0_c_559_p N_A_597_297#_c_1550_n 0.0202695f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_526 N_A0_c_542_n N_A_597_297#_c_1550_n 0.00669726f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_527 N_A0_c_545_n N_A_597_297#_c_1554_n 5.6422e-19 $X=9.055 $Y=1.41 $X2=0
+ $Y2=0
cc_528 N_A0_c_546_n N_A_597_297#_c_1554_n 0.00214429f $X=9.525 $Y=1.41 $X2=0
+ $Y2=0
cc_529 N_A0_c_559_p N_A_597_297#_c_1554_n 0.0203246f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_530 N_A0_c_542_n N_A_597_297#_c_1554_n 0.00669726f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_531 N_A0_c_543_n N_A_597_297#_c_1516_n 0.00600932f $X=8.115 $Y=1.41 $X2=0
+ $Y2=0
cc_532 N_A0_c_559_p N_A_597_297#_c_1516_n 0.00233931f $X=9.29 $Y=1.16 $X2=0
+ $Y2=0
cc_533 N_A0_c_542_n N_A_597_297#_c_1516_n 2.02467e-19 $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_534 N_A0_c_544_n N_A_597_297#_c_1561_n 0.00313189f $X=8.585 $Y=1.41 $X2=0
+ $Y2=0
cc_535 N_A0_c_545_n N_A_597_297#_c_1561_n 0.00313189f $X=9.055 $Y=1.41 $X2=0
+ $Y2=0
cc_536 N_A0_c_559_p N_A_597_297#_c_1561_n 0.00107383f $X=9.29 $Y=1.16 $X2=0
+ $Y2=0
cc_537 N_A0_c_559_p N_A_597_297#_c_1564_n 0.00117983f $X=9.29 $Y=1.16 $X2=0
+ $Y2=0
cc_538 N_A0_c_543_n N_A_597_297#_c_1565_n 0.004823f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_539 N_A0_c_544_n N_A_597_297#_c_1565_n 0.00606957f $X=8.585 $Y=1.41 $X2=0
+ $Y2=0
cc_540 N_A0_c_545_n N_A_597_297#_c_1565_n 5.7339e-19 $X=9.055 $Y=1.41 $X2=0
+ $Y2=0
cc_541 N_A0_c_559_p N_A_597_297#_c_1568_n 0.00117983f $X=9.29 $Y=1.16 $X2=0
+ $Y2=0
cc_542 N_A0_c_544_n N_A_597_297#_c_1569_n 5.7339e-19 $X=8.585 $Y=1.41 $X2=0
+ $Y2=0
cc_543 N_A0_c_545_n N_A_597_297#_c_1569_n 0.00606957f $X=9.055 $Y=1.41 $X2=0
+ $Y2=0
cc_544 N_A0_c_546_n N_A_597_297#_c_1569_n 0.00532302f $X=9.525 $Y=1.41 $X2=0
+ $Y2=0
cc_545 N_A0_c_538_n N_VGND_c_1959_n 0.00203215f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A0_c_541_n N_VGND_c_1960_n 0.00202093f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_547 N_A0_c_538_n N_VGND_c_1977_n 0.00357877f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_548 N_A0_c_539_n N_VGND_c_1977_n 0.00357877f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_549 N_A0_c_540_n N_VGND_c_1977_n 0.00357877f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_550 N_A0_c_541_n N_VGND_c_1977_n 0.00357877f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_551 N_A0_c_538_n N_VGND_c_1987_n 0.00605604f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_552 N_A0_c_539_n N_VGND_c_1987_n 0.00497228f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_553 N_A0_c_540_n N_VGND_c_1987_n 0.00497228f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_554 N_A0_c_541_n N_VGND_c_1987_n 0.00605604f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_555 N_A0_c_538_n N_A_1163_47#_c_2221_n 0.0112292f $X=8.14 $Y=0.995 $X2=0
+ $Y2=0
cc_556 N_A0_c_559_p N_A_1163_47#_c_2221_n 0.0974168f $X=9.29 $Y=1.16 $X2=0 $Y2=0
cc_557 N_A0_c_542_n N_A_1163_47#_c_2221_n 0.00224539f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_558 N_A0_c_538_n N_A_1163_47#_c_2222_n 0.00716324f $X=8.14 $Y=0.995 $X2=0
+ $Y2=0
cc_559 N_A0_c_539_n N_A_1163_47#_c_2222_n 0.00402996f $X=8.56 $Y=0.995 $X2=0
+ $Y2=0
cc_560 N_A0_c_540_n N_A_1163_47#_c_2222_n 4.02078e-19 $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_561 N_A0_c_542_n N_A_1163_47#_c_2222_n 0.00225271f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_562 N_A0_c_539_n N_A_1163_47#_c_2223_n 4.02078e-19 $X=8.56 $Y=0.995 $X2=0
+ $Y2=0
cc_563 N_A0_c_540_n N_A_1163_47#_c_2223_n 0.00402996f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_564 N_A0_c_541_n N_A_1163_47#_c_2223_n 0.00440693f $X=9.5 $Y=0.995 $X2=0
+ $Y2=0
cc_565 N_A0_c_542_n N_A_1163_47#_c_2223_n 0.00225271f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_566 N_A0_c_539_n N_A_1163_47#_c_2224_n 0.00754011f $X=8.56 $Y=0.995 $X2=0
+ $Y2=0
cc_567 N_A0_c_540_n N_A_1163_47#_c_2224_n 0.00754011f $X=9.08 $Y=0.995 $X2=0
+ $Y2=0
cc_568 N_A0_c_542_n N_A_1163_47#_c_2224_n 0.00468948f $X=9.5 $Y=1.202 $X2=0
+ $Y2=0
cc_569 N_A_27_47#_c_675_n N_A_117_297#_M1002_s 0.00341977f $X=1.065 $Y=2.38
+ $X2=-0.19 $Y2=-0.24
cc_570 N_A_27_47#_c_677_n N_A_117_297#_M1035_s 0.00341977f $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_571 N_A_27_47#_M1026_d N_A_117_297#_c_1111_n 0.00315544f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_572 N_A_27_47#_c_675_n N_A_117_297#_c_1111_n 0.00144594f $X=1.065 $Y=2.38
+ $X2=0 $Y2=0
cc_573 N_A_27_47#_c_736_p N_A_117_297#_c_1111_n 0.0130853f $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_574 N_A_27_47#_c_677_n N_A_117_297#_c_1111_n 0.00144594f $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_575 N_A_27_47#_M1026_d N_A_117_297#_c_1123_n 0.00234633f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_576 N_A_27_47#_c_675_n N_A_117_297#_c_1123_n 0.00174687f $X=1.065 $Y=2.38
+ $X2=0 $Y2=0
cc_577 N_A_27_47#_c_736_p N_A_117_297#_c_1123_n 0.0135446f $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_c_677_n N_A_117_297#_c_1123_n 0.00174687f $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_579 N_A_27_47#_c_675_n N_A_117_297#_c_1126_n 9.16304e-19 $X=1.065 $Y=2.38
+ $X2=0 $Y2=0
cc_580 N_A_27_47#_c_736_p N_A_117_297#_c_1126_n 3.34135e-19 $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_581 N_A_27_47#_c_649_n N_A_117_297#_c_1126_n 0.00168706f $X=0.26 $Y=0.51
+ $X2=0 $Y2=0
cc_582 N_A_27_47#_M1048_d N_A_117_297#_c_1110_n 2.0128e-19 $X=1.995 $Y=1.485
+ $X2=0 $Y2=0
cc_583 N_A_27_47#_c_677_n N_A_117_297#_c_1110_n 0.00348472f $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_584 N_A_27_47#_c_665_n N_A_117_297#_c_1110_n 0.0302802f $X=2.14 $Y=1.66 $X2=0
+ $Y2=0
cc_585 N_A_27_47#_c_736_p N_A_117_297#_c_1130_n 3.34135e-19 $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_586 N_A_27_47#_c_677_n N_A_117_297#_c_1130_n 9.16304e-19 $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_587 N_A_27_47#_c_665_n N_A_117_297#_c_1130_n 6.74054e-19 $X=2.14 $Y=1.66
+ $X2=0 $Y2=0
cc_588 N_A_27_47#_c_675_n N_A_117_297#_c_1131_n 0.0150323f $X=1.065 $Y=2.38
+ $X2=0 $Y2=0
cc_589 N_A_27_47#_c_736_p N_A_117_297#_c_1131_n 0.0122463f $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_590 N_A_27_47#_c_736_p N_A_117_297#_c_1134_n 0.0122463f $X=1.2 $Y=2 $X2=0
+ $Y2=0
cc_591 N_A_27_47#_c_677_n N_A_117_297#_c_1134_n 0.0149581f $X=2.005 $Y=2.38
+ $X2=0 $Y2=0
cc_592 N_A_27_47#_c_665_n N_A_117_297#_c_1134_n 0.0190508f $X=2.14 $Y=1.66 $X2=0
+ $Y2=0
cc_593 N_A_27_47#_c_664_n N_VPWR_c_1242_n 0.0123662f $X=2.155 $Y=2.295 $X2=0
+ $Y2=0
cc_594 N_A_27_47#_c_665_n N_VPWR_c_1242_n 0.0526296f $X=2.14 $Y=1.66 $X2=0 $Y2=0
cc_595 N_A_27_47#_c_666_n N_VPWR_c_1247_n 0.0123662f $X=7.865 $Y=2.295 $X2=0
+ $Y2=0
cc_596 N_A_27_47#_c_667_n N_VPWR_c_1247_n 0.0453948f $X=7.88 $Y=1.66 $X2=0 $Y2=0
cc_597 N_A_27_47#_c_652_n N_VPWR_c_1248_n 0.00354866f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_598 N_A_27_47#_c_668_n N_VPWR_c_1248_n 0.0123662f $X=9.775 $Y=2.295 $X2=0
+ $Y2=0
cc_599 N_A_27_47#_c_669_n N_VPWR_c_1248_n 0.0543558f $X=9.76 $Y=1.66 $X2=0 $Y2=0
cc_600 N_A_27_47#_c_642_n N_VPWR_c_1248_n 0.0207233f $X=14.66 $Y=1.16 $X2=0
+ $Y2=0
cc_601 N_A_27_47#_c_653_n N_VPWR_c_1249_n 0.00173895f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_602 N_A_27_47#_c_654_n N_VPWR_c_1249_n 0.00173895f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_603 N_A_27_47#_c_655_n N_VPWR_c_1250_n 0.00173895f $X=11.925 $Y=1.41 $X2=0
+ $Y2=0
cc_604 N_A_27_47#_c_656_n N_VPWR_c_1250_n 0.00173895f $X=12.395 $Y=1.41 $X2=0
+ $Y2=0
cc_605 N_A_27_47#_c_657_n N_VPWR_c_1251_n 0.00173895f $X=12.865 $Y=1.41 $X2=0
+ $Y2=0
cc_606 N_A_27_47#_c_658_n N_VPWR_c_1251_n 0.00173895f $X=13.335 $Y=1.41 $X2=0
+ $Y2=0
cc_607 N_A_27_47#_c_659_n N_VPWR_c_1252_n 0.00173895f $X=13.805 $Y=1.41 $X2=0
+ $Y2=0
cc_608 N_A_27_47#_c_660_n N_VPWR_c_1252_n 0.00173895f $X=14.275 $Y=1.41 $X2=0
+ $Y2=0
cc_609 N_A_27_47#_c_661_n N_VPWR_c_1253_n 0.00173895f $X=14.745 $Y=1.41 $X2=0
+ $Y2=0
cc_610 N_A_27_47#_c_662_n N_VPWR_c_1253_n 0.00173895f $X=15.215 $Y=1.41 $X2=0
+ $Y2=0
cc_611 N_A_27_47#_c_663_n N_VPWR_c_1254_n 0.00354866f $X=15.685 $Y=1.41 $X2=0
+ $Y2=0
cc_612 N_A_27_47#_c_666_n N_VPWR_c_1265_n 0.0195137f $X=7.865 $Y=2.295 $X2=0
+ $Y2=0
cc_613 N_A_27_47#_c_710_n N_VPWR_c_1265_n 0.0379761f $X=8.685 $Y=2.38 $X2=0
+ $Y2=0
cc_614 N_A_27_47#_c_715_n N_VPWR_c_1265_n 0.0379761f $X=9.625 $Y=2.38 $X2=0
+ $Y2=0
cc_615 N_A_27_47#_c_668_n N_VPWR_c_1265_n 0.0195137f $X=9.775 $Y=2.295 $X2=0
+ $Y2=0
cc_616 N_A_27_47#_c_779_p N_VPWR_c_1265_n 0.0156426f $X=8.82 $Y=2.38 $X2=0 $Y2=0
cc_617 N_A_27_47#_c_675_n N_VPWR_c_1267_n 0.0379761f $X=1.065 $Y=2.38 $X2=0
+ $Y2=0
cc_618 N_A_27_47#_c_677_n N_VPWR_c_1267_n 0.0379761f $X=2.005 $Y=2.38 $X2=0
+ $Y2=0
cc_619 N_A_27_47#_c_664_n N_VPWR_c_1267_n 0.0195137f $X=2.155 $Y=2.295 $X2=0
+ $Y2=0
cc_620 N_A_27_47#_c_671_n N_VPWR_c_1267_n 0.0194775f $X=0.245 $Y=2.295 $X2=0
+ $Y2=0
cc_621 N_A_27_47#_c_784_p N_VPWR_c_1267_n 0.0156426f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_622 N_A_27_47#_c_652_n N_VPWR_c_1268_n 0.00673617f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_623 N_A_27_47#_c_653_n N_VPWR_c_1268_n 0.00673617f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_624 N_A_27_47#_c_654_n N_VPWR_c_1269_n 0.00673617f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_625 N_A_27_47#_c_655_n N_VPWR_c_1269_n 0.00673617f $X=11.925 $Y=1.41 $X2=0
+ $Y2=0
cc_626 N_A_27_47#_c_656_n N_VPWR_c_1270_n 0.00673617f $X=12.395 $Y=1.41 $X2=0
+ $Y2=0
cc_627 N_A_27_47#_c_657_n N_VPWR_c_1270_n 0.00673617f $X=12.865 $Y=1.41 $X2=0
+ $Y2=0
cc_628 N_A_27_47#_c_658_n N_VPWR_c_1271_n 0.00673617f $X=13.335 $Y=1.41 $X2=0
+ $Y2=0
cc_629 N_A_27_47#_c_659_n N_VPWR_c_1271_n 0.00673617f $X=13.805 $Y=1.41 $X2=0
+ $Y2=0
cc_630 N_A_27_47#_c_660_n N_VPWR_c_1272_n 0.00673617f $X=14.275 $Y=1.41 $X2=0
+ $Y2=0
cc_631 N_A_27_47#_c_661_n N_VPWR_c_1272_n 0.00673617f $X=14.745 $Y=1.41 $X2=0
+ $Y2=0
cc_632 N_A_27_47#_c_662_n N_VPWR_c_1273_n 0.00673617f $X=15.215 $Y=1.41 $X2=0
+ $Y2=0
cc_633 N_A_27_47#_c_663_n N_VPWR_c_1273_n 0.00673617f $X=15.685 $Y=1.41 $X2=0
+ $Y2=0
cc_634 N_A_27_47#_M1002_d N_VPWR_c_1241_n 0.00217518f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_635 N_A_27_47#_M1026_d N_VPWR_c_1241_n 0.00190236f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_636 N_A_27_47#_M1048_d N_VPWR_c_1241_n 0.00179198f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_637 N_A_27_47#_M1008_s N_VPWR_c_1241_n 0.00179198f $X=7.755 $Y=1.485 $X2=0
+ $Y2=0
cc_638 N_A_27_47#_M1010_s N_VPWR_c_1241_n 0.00190236f $X=8.675 $Y=1.485 $X2=0
+ $Y2=0
cc_639 N_A_27_47#_M1030_s N_VPWR_c_1241_n 0.00217518f $X=9.615 $Y=1.485 $X2=0
+ $Y2=0
cc_640 N_A_27_47#_c_652_n N_VPWR_c_1241_n 0.0130007f $X=10.515 $Y=1.41 $X2=0
+ $Y2=0
cc_641 N_A_27_47#_c_653_n N_VPWR_c_1241_n 0.0117184f $X=10.985 $Y=1.41 $X2=0
+ $Y2=0
cc_642 N_A_27_47#_c_654_n N_VPWR_c_1241_n 0.0117184f $X=11.455 $Y=1.41 $X2=0
+ $Y2=0
cc_643 N_A_27_47#_c_655_n N_VPWR_c_1241_n 0.0117184f $X=11.925 $Y=1.41 $X2=0
+ $Y2=0
cc_644 N_A_27_47#_c_656_n N_VPWR_c_1241_n 0.0117184f $X=12.395 $Y=1.41 $X2=0
+ $Y2=0
cc_645 N_A_27_47#_c_657_n N_VPWR_c_1241_n 0.0117184f $X=12.865 $Y=1.41 $X2=0
+ $Y2=0
cc_646 N_A_27_47#_c_658_n N_VPWR_c_1241_n 0.0117184f $X=13.335 $Y=1.41 $X2=0
+ $Y2=0
cc_647 N_A_27_47#_c_659_n N_VPWR_c_1241_n 0.0117184f $X=13.805 $Y=1.41 $X2=0
+ $Y2=0
cc_648 N_A_27_47#_c_660_n N_VPWR_c_1241_n 0.0117184f $X=14.275 $Y=1.41 $X2=0
+ $Y2=0
cc_649 N_A_27_47#_c_661_n N_VPWR_c_1241_n 0.0117184f $X=14.745 $Y=1.41 $X2=0
+ $Y2=0
cc_650 N_A_27_47#_c_662_n N_VPWR_c_1241_n 0.0117184f $X=15.215 $Y=1.41 $X2=0
+ $Y2=0
cc_651 N_A_27_47#_c_663_n N_VPWR_c_1241_n 0.0130007f $X=15.685 $Y=1.41 $X2=0
+ $Y2=0
cc_652 N_A_27_47#_c_675_n N_VPWR_c_1241_n 0.0137178f $X=1.065 $Y=2.38 $X2=0
+ $Y2=0
cc_653 N_A_27_47#_c_677_n N_VPWR_c_1241_n 0.0103607f $X=2.005 $Y=2.38 $X2=0
+ $Y2=0
cc_654 N_A_27_47#_c_664_n N_VPWR_c_1241_n 0.00550351f $X=2.155 $Y=2.295 $X2=0
+ $Y2=0
cc_655 N_A_27_47#_c_666_n N_VPWR_c_1241_n 0.00550351f $X=7.865 $Y=2.295 $X2=0
+ $Y2=0
cc_656 N_A_27_47#_c_710_n N_VPWR_c_1241_n 0.0103607f $X=8.685 $Y=2.38 $X2=0
+ $Y2=0
cc_657 N_A_27_47#_c_715_n N_VPWR_c_1241_n 0.0137178f $X=9.625 $Y=2.38 $X2=0
+ $Y2=0
cc_658 N_A_27_47#_c_668_n N_VPWR_c_1241_n 0.0115483f $X=9.775 $Y=2.295 $X2=0
+ $Y2=0
cc_659 N_A_27_47#_c_671_n N_VPWR_c_1241_n 0.0115431f $X=0.245 $Y=2.295 $X2=0
+ $Y2=0
cc_660 N_A_27_47#_c_784_p N_VPWR_c_1241_n 0.00493251f $X=1.2 $Y=2.38 $X2=0 $Y2=0
cc_661 N_A_27_47#_c_779_p N_VPWR_c_1241_n 0.00493251f $X=8.82 $Y=2.38 $X2=0
+ $Y2=0
cc_662 N_A_27_47#_c_710_n N_A_597_297#_M1008_d 0.00341977f $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_663 N_A_27_47#_c_715_n N_A_597_297#_M1018_d 0.00341977f $X=9.625 $Y=2.38
+ $X2=0 $Y2=0
cc_664 N_A_27_47#_M1010_s N_A_597_297#_c_1546_n 0.00315544f $X=8.675 $Y=1.485
+ $X2=0 $Y2=0
cc_665 N_A_27_47#_c_710_n N_A_597_297#_c_1546_n 0.00144594f $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_666 N_A_27_47#_c_829_p N_A_597_297#_c_1546_n 0.0130853f $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_667 N_A_27_47#_c_715_n N_A_597_297#_c_1546_n 0.00144594f $X=9.625 $Y=2.38
+ $X2=0 $Y2=0
cc_668 N_A_27_47#_c_667_n N_A_597_297#_c_1515_n 0.0108287f $X=7.88 $Y=1.66 $X2=0
+ $Y2=0
cc_669 N_A_27_47#_M1008_s N_A_597_297#_c_1516_n 2.0128e-19 $X=7.755 $Y=1.485
+ $X2=0 $Y2=0
cc_670 N_A_27_47#_c_667_n N_A_597_297#_c_1516_n 0.0299084f $X=7.88 $Y=1.66 $X2=0
+ $Y2=0
cc_671 N_A_27_47#_c_710_n N_A_597_297#_c_1516_n 0.00348472f $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_672 N_A_27_47#_M1010_s N_A_597_297#_c_1561_n 0.00234633f $X=8.675 $Y=1.485
+ $X2=0 $Y2=0
cc_673 N_A_27_47#_c_710_n N_A_597_297#_c_1561_n 0.00174687f $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_674 N_A_27_47#_c_829_p N_A_597_297#_c_1561_n 0.0135446f $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_675 N_A_27_47#_c_715_n N_A_597_297#_c_1561_n 0.00174687f $X=9.625 $Y=2.38
+ $X2=0 $Y2=0
cc_676 N_A_27_47#_c_667_n N_A_597_297#_c_1564_n 5.45688e-19 $X=7.88 $Y=1.66
+ $X2=0 $Y2=0
cc_677 N_A_27_47#_c_710_n N_A_597_297#_c_1564_n 9.16304e-19 $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_678 N_A_27_47#_c_829_p N_A_597_297#_c_1564_n 3.34135e-19 $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_679 N_A_27_47#_c_667_n N_A_597_297#_c_1565_n 0.0186023f $X=7.88 $Y=1.66 $X2=0
+ $Y2=0
cc_680 N_A_27_47#_c_710_n N_A_597_297#_c_1565_n 0.0149581f $X=8.685 $Y=2.38
+ $X2=0 $Y2=0
cc_681 N_A_27_47#_c_829_p N_A_597_297#_c_1565_n 0.0122463f $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_682 N_A_27_47#_c_829_p N_A_597_297#_c_1568_n 3.34135e-19 $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_683 N_A_27_47#_c_715_n N_A_597_297#_c_1568_n 9.16304e-19 $X=9.625 $Y=2.38
+ $X2=0 $Y2=0
cc_684 N_A_27_47#_c_669_n N_A_597_297#_c_1568_n 0.00168706f $X=9.76 $Y=1.66
+ $X2=0 $Y2=0
cc_685 N_A_27_47#_c_829_p N_A_597_297#_c_1569_n 0.0122463f $X=8.82 $Y=2 $X2=0
+ $Y2=0
cc_686 N_A_27_47#_c_715_n N_A_597_297#_c_1569_n 0.0150323f $X=9.625 $Y=2.38
+ $X2=0 $Y2=0
cc_687 N_A_27_47#_c_630_n N_X_c_1662_n 0.00539651f $X=10.54 $Y=0.995 $X2=0 $Y2=0
cc_688 N_A_27_47#_c_631_n N_X_c_1662_n 0.00680665f $X=10.96 $Y=0.995 $X2=0 $Y2=0
cc_689 N_A_27_47#_c_632_n N_X_c_1662_n 5.53497e-19 $X=11.48 $Y=0.995 $X2=0 $Y2=0
cc_690 N_A_27_47#_c_652_n N_X_c_1665_n 0.00215964f $X=10.515 $Y=1.41 $X2=0 $Y2=0
cc_691 N_A_27_47#_c_653_n N_X_c_1665_n 5.79575e-19 $X=10.985 $Y=1.41 $X2=0 $Y2=0
cc_692 N_A_27_47#_c_642_n N_X_c_1665_n 0.0214226f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_693 N_A_27_47#_c_651_n N_X_c_1665_n 0.00671335f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_694 N_A_27_47#_c_652_n N_X_c_1669_n 0.00897418f $X=10.515 $Y=1.41 $X2=0 $Y2=0
cc_695 N_A_27_47#_c_653_n N_X_c_1669_n 0.0100233f $X=10.985 $Y=1.41 $X2=0 $Y2=0
cc_696 N_A_27_47#_c_654_n N_X_c_1669_n 5.91934e-19 $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_697 N_A_27_47#_c_631_n N_X_c_1652_n 0.00929182f $X=10.96 $Y=0.995 $X2=0 $Y2=0
cc_698 N_A_27_47#_c_632_n N_X_c_1652_n 0.00929182f $X=11.48 $Y=0.995 $X2=0 $Y2=0
cc_699 N_A_27_47#_c_642_n N_X_c_1652_n 0.0441201f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_700 N_A_27_47#_c_651_n N_X_c_1652_n 0.00468948f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_701 N_A_27_47#_c_630_n N_X_c_1653_n 0.00262807f $X=10.54 $Y=0.995 $X2=0 $Y2=0
cc_702 N_A_27_47#_c_631_n N_X_c_1653_n 0.00113286f $X=10.96 $Y=0.995 $X2=0 $Y2=0
cc_703 N_A_27_47#_c_642_n N_X_c_1653_n 0.0269421f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_704 N_A_27_47#_c_651_n N_X_c_1653_n 0.00230339f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_705 N_A_27_47#_c_653_n N_X_c_1680_n 0.0137916f $X=10.985 $Y=1.41 $X2=0 $Y2=0
cc_706 N_A_27_47#_c_654_n N_X_c_1680_n 0.0137916f $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_707 N_A_27_47#_c_642_n N_X_c_1680_n 0.0391038f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_708 N_A_27_47#_c_651_n N_X_c_1680_n 0.00616252f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_709 N_A_27_47#_c_631_n N_X_c_1684_n 5.53497e-19 $X=10.96 $Y=0.995 $X2=0 $Y2=0
cc_710 N_A_27_47#_c_632_n N_X_c_1684_n 0.00680665f $X=11.48 $Y=0.995 $X2=0 $Y2=0
cc_711 N_A_27_47#_c_633_n N_X_c_1684_n 0.00680665f $X=11.9 $Y=0.995 $X2=0 $Y2=0
cc_712 N_A_27_47#_c_634_n N_X_c_1684_n 5.53497e-19 $X=12.42 $Y=0.995 $X2=0 $Y2=0
cc_713 N_A_27_47#_c_653_n N_X_c_1688_n 5.91934e-19 $X=10.985 $Y=1.41 $X2=0 $Y2=0
cc_714 N_A_27_47#_c_654_n N_X_c_1688_n 0.0100233f $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_715 N_A_27_47#_c_655_n N_X_c_1688_n 0.0100233f $X=11.925 $Y=1.41 $X2=0 $Y2=0
cc_716 N_A_27_47#_c_656_n N_X_c_1688_n 5.91934e-19 $X=12.395 $Y=1.41 $X2=0 $Y2=0
cc_717 N_A_27_47#_c_633_n N_X_c_1654_n 0.00929182f $X=11.9 $Y=0.995 $X2=0 $Y2=0
cc_718 N_A_27_47#_c_634_n N_X_c_1654_n 0.00929182f $X=12.42 $Y=0.995 $X2=0 $Y2=0
cc_719 N_A_27_47#_c_642_n N_X_c_1654_n 0.0441201f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_720 N_A_27_47#_c_651_n N_X_c_1654_n 0.00468948f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_721 N_A_27_47#_c_655_n N_X_c_1696_n 0.0137916f $X=11.925 $Y=1.41 $X2=0 $Y2=0
cc_722 N_A_27_47#_c_656_n N_X_c_1696_n 0.0137916f $X=12.395 $Y=1.41 $X2=0 $Y2=0
cc_723 N_A_27_47#_c_642_n N_X_c_1696_n 0.0391038f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_724 N_A_27_47#_c_651_n N_X_c_1696_n 0.00616252f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_725 N_A_27_47#_c_633_n N_X_c_1700_n 5.53497e-19 $X=11.9 $Y=0.995 $X2=0 $Y2=0
cc_726 N_A_27_47#_c_634_n N_X_c_1700_n 0.00680665f $X=12.42 $Y=0.995 $X2=0 $Y2=0
cc_727 N_A_27_47#_c_635_n N_X_c_1700_n 0.00680665f $X=12.84 $Y=0.995 $X2=0 $Y2=0
cc_728 N_A_27_47#_c_636_n N_X_c_1700_n 5.53497e-19 $X=13.36 $Y=0.995 $X2=0 $Y2=0
cc_729 N_A_27_47#_c_655_n N_X_c_1704_n 5.91934e-19 $X=11.925 $Y=1.41 $X2=0 $Y2=0
cc_730 N_A_27_47#_c_656_n N_X_c_1704_n 0.0100233f $X=12.395 $Y=1.41 $X2=0 $Y2=0
cc_731 N_A_27_47#_c_657_n N_X_c_1704_n 0.0100233f $X=12.865 $Y=1.41 $X2=0 $Y2=0
cc_732 N_A_27_47#_c_658_n N_X_c_1704_n 5.91934e-19 $X=13.335 $Y=1.41 $X2=0 $Y2=0
cc_733 N_A_27_47#_c_635_n N_X_c_1655_n 0.00929182f $X=12.84 $Y=0.995 $X2=0 $Y2=0
cc_734 N_A_27_47#_c_636_n N_X_c_1655_n 0.00929182f $X=13.36 $Y=0.995 $X2=0 $Y2=0
cc_735 N_A_27_47#_c_642_n N_X_c_1655_n 0.0441201f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_736 N_A_27_47#_c_651_n N_X_c_1655_n 0.00468948f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_737 N_A_27_47#_c_657_n N_X_c_1712_n 0.0137916f $X=12.865 $Y=1.41 $X2=0 $Y2=0
cc_738 N_A_27_47#_c_658_n N_X_c_1712_n 0.0137916f $X=13.335 $Y=1.41 $X2=0 $Y2=0
cc_739 N_A_27_47#_c_642_n N_X_c_1712_n 0.0391038f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_740 N_A_27_47#_c_651_n N_X_c_1712_n 0.00616252f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_741 N_A_27_47#_c_635_n N_X_c_1716_n 5.53497e-19 $X=12.84 $Y=0.995 $X2=0 $Y2=0
cc_742 N_A_27_47#_c_636_n N_X_c_1716_n 0.00680665f $X=13.36 $Y=0.995 $X2=0 $Y2=0
cc_743 N_A_27_47#_c_637_n N_X_c_1716_n 0.00676194f $X=13.78 $Y=0.995 $X2=0 $Y2=0
cc_744 N_A_27_47#_c_638_n N_X_c_1716_n 5.39066e-19 $X=14.3 $Y=0.995 $X2=0 $Y2=0
cc_745 N_A_27_47#_c_657_n N_X_c_1720_n 5.91934e-19 $X=12.865 $Y=1.41 $X2=0 $Y2=0
cc_746 N_A_27_47#_c_658_n N_X_c_1720_n 0.0100233f $X=13.335 $Y=1.41 $X2=0 $Y2=0
cc_747 N_A_27_47#_c_659_n N_X_c_1720_n 0.0100233f $X=13.805 $Y=1.41 $X2=0 $Y2=0
cc_748 N_A_27_47#_c_660_n N_X_c_1720_n 5.91934e-19 $X=14.275 $Y=1.41 $X2=0 $Y2=0
cc_749 N_A_27_47#_c_637_n N_X_c_1656_n 0.00929182f $X=13.78 $Y=0.995 $X2=0 $Y2=0
cc_750 N_A_27_47#_c_638_n N_X_c_1656_n 0.00929182f $X=14.3 $Y=0.995 $X2=0 $Y2=0
cc_751 N_A_27_47#_c_642_n N_X_c_1656_n 0.0441201f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_752 N_A_27_47#_c_651_n N_X_c_1656_n 0.00468948f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_753 N_A_27_47#_c_659_n N_X_c_1728_n 0.0137916f $X=13.805 $Y=1.41 $X2=0 $Y2=0
cc_754 N_A_27_47#_c_660_n N_X_c_1728_n 0.0137916f $X=14.275 $Y=1.41 $X2=0 $Y2=0
cc_755 N_A_27_47#_c_642_n N_X_c_1728_n 0.0391038f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_756 N_A_27_47#_c_651_n N_X_c_1728_n 0.00616252f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_757 N_A_27_47#_c_637_n N_X_c_1732_n 5.39066e-19 $X=13.78 $Y=0.995 $X2=0 $Y2=0
cc_758 N_A_27_47#_c_638_n N_X_c_1732_n 0.00676194f $X=14.3 $Y=0.995 $X2=0 $Y2=0
cc_759 N_A_27_47#_c_639_n N_X_c_1732_n 0.00680665f $X=14.72 $Y=0.995 $X2=0 $Y2=0
cc_760 N_A_27_47#_c_640_n N_X_c_1732_n 5.53497e-19 $X=15.24 $Y=0.995 $X2=0 $Y2=0
cc_761 N_A_27_47#_c_659_n N_X_c_1736_n 5.91934e-19 $X=13.805 $Y=1.41 $X2=0 $Y2=0
cc_762 N_A_27_47#_c_660_n N_X_c_1736_n 0.0100233f $X=14.275 $Y=1.41 $X2=0 $Y2=0
cc_763 N_A_27_47#_c_661_n N_X_c_1736_n 0.0100233f $X=14.745 $Y=1.41 $X2=0 $Y2=0
cc_764 N_A_27_47#_c_662_n N_X_c_1736_n 5.91934e-19 $X=15.215 $Y=1.41 $X2=0 $Y2=0
cc_765 N_A_27_47#_c_639_n N_X_c_1657_n 0.00929182f $X=14.72 $Y=0.995 $X2=0 $Y2=0
cc_766 N_A_27_47#_c_640_n N_X_c_1657_n 0.010806f $X=15.24 $Y=0.995 $X2=0 $Y2=0
cc_767 N_A_27_47#_c_642_n N_X_c_1657_n 0.0106019f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_768 N_A_27_47#_c_651_n N_X_c_1657_n 0.00563654f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_769 N_A_27_47#_c_661_n N_X_c_1744_n 0.0139192f $X=14.745 $Y=1.41 $X2=0 $Y2=0
cc_770 N_A_27_47#_c_662_n N_X_c_1744_n 0.0158202f $X=15.215 $Y=1.41 $X2=0 $Y2=0
cc_771 N_A_27_47#_c_642_n N_X_c_1744_n 0.0104436f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_772 N_A_27_47#_c_651_n N_X_c_1744_n 0.00691238f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_773 N_A_27_47#_c_639_n N_X_c_1748_n 5.53497e-19 $X=14.72 $Y=0.995 $X2=0 $Y2=0
cc_774 N_A_27_47#_c_640_n N_X_c_1748_n 0.00680665f $X=15.24 $Y=0.995 $X2=0 $Y2=0
cc_775 N_A_27_47#_c_641_n N_X_c_1748_n 0.00539651f $X=15.66 $Y=0.995 $X2=0 $Y2=0
cc_776 N_A_27_47#_c_661_n N_X_c_1751_n 5.91934e-19 $X=14.745 $Y=1.41 $X2=0 $Y2=0
cc_777 N_A_27_47#_c_662_n N_X_c_1751_n 0.0100233f $X=15.215 $Y=1.41 $X2=0 $Y2=0
cc_778 N_A_27_47#_c_663_n N_X_c_1751_n 0.00897418f $X=15.685 $Y=1.41 $X2=0 $Y2=0
cc_779 N_A_27_47#_c_632_n N_X_c_1658_n 0.00113286f $X=11.48 $Y=0.995 $X2=0 $Y2=0
cc_780 N_A_27_47#_c_633_n N_X_c_1658_n 0.00113286f $X=11.9 $Y=0.995 $X2=0 $Y2=0
cc_781 N_A_27_47#_c_642_n N_X_c_1658_n 0.0269421f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_782 N_A_27_47#_c_651_n N_X_c_1658_n 0.00230339f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_783 N_A_27_47#_c_654_n N_X_c_1758_n 5.79575e-19 $X=11.455 $Y=1.41 $X2=0 $Y2=0
cc_784 N_A_27_47#_c_655_n N_X_c_1758_n 5.79575e-19 $X=11.925 $Y=1.41 $X2=0 $Y2=0
cc_785 N_A_27_47#_c_642_n N_X_c_1758_n 0.0214226f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_786 N_A_27_47#_c_651_n N_X_c_1758_n 0.00671335f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_787 N_A_27_47#_c_634_n N_X_c_1659_n 0.00113286f $X=12.42 $Y=0.995 $X2=0 $Y2=0
cc_788 N_A_27_47#_c_635_n N_X_c_1659_n 0.00113286f $X=12.84 $Y=0.995 $X2=0 $Y2=0
cc_789 N_A_27_47#_c_642_n N_X_c_1659_n 0.0269421f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_790 N_A_27_47#_c_651_n N_X_c_1659_n 0.00230339f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_791 N_A_27_47#_c_656_n N_X_c_1766_n 5.79575e-19 $X=12.395 $Y=1.41 $X2=0 $Y2=0
cc_792 N_A_27_47#_c_657_n N_X_c_1766_n 5.79575e-19 $X=12.865 $Y=1.41 $X2=0 $Y2=0
cc_793 N_A_27_47#_c_642_n N_X_c_1766_n 0.0214226f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_794 N_A_27_47#_c_651_n N_X_c_1766_n 0.00671335f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_795 N_A_27_47#_c_636_n N_X_c_1660_n 0.00113286f $X=13.36 $Y=0.995 $X2=0 $Y2=0
cc_796 N_A_27_47#_c_637_n N_X_c_1660_n 0.00113286f $X=13.78 $Y=0.995 $X2=0 $Y2=0
cc_797 N_A_27_47#_c_642_n N_X_c_1660_n 0.0269421f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_798 N_A_27_47#_c_651_n N_X_c_1660_n 0.00230339f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_799 N_A_27_47#_c_658_n N_X_c_1774_n 5.79575e-19 $X=13.335 $Y=1.41 $X2=0 $Y2=0
cc_800 N_A_27_47#_c_659_n N_X_c_1774_n 5.79575e-19 $X=13.805 $Y=1.41 $X2=0 $Y2=0
cc_801 N_A_27_47#_c_642_n N_X_c_1774_n 0.0214226f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_802 N_A_27_47#_c_651_n N_X_c_1774_n 0.00671335f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_803 N_A_27_47#_c_638_n N_X_c_1661_n 0.00113286f $X=14.3 $Y=0.995 $X2=0 $Y2=0
cc_804 N_A_27_47#_c_639_n N_X_c_1661_n 0.00113286f $X=14.72 $Y=0.995 $X2=0 $Y2=0
cc_805 N_A_27_47#_c_642_n N_X_c_1661_n 0.0269421f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_806 N_A_27_47#_c_651_n N_X_c_1661_n 0.00230339f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_807 N_A_27_47#_c_660_n N_X_c_1782_n 5.79575e-19 $X=14.275 $Y=1.41 $X2=0 $Y2=0
cc_808 N_A_27_47#_c_661_n N_X_c_1782_n 5.79575e-19 $X=14.745 $Y=1.41 $X2=0 $Y2=0
cc_809 N_A_27_47#_c_642_n N_X_c_1782_n 0.0214226f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_810 N_A_27_47#_c_651_n N_X_c_1782_n 0.00671335f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_811 N_A_27_47#_c_640_n N_X_c_1786_n 7.13294e-19 $X=15.24 $Y=0.995 $X2=0 $Y2=0
cc_812 N_A_27_47#_c_641_n N_X_c_1786_n 0.00220851f $X=15.66 $Y=0.995 $X2=0 $Y2=0
cc_813 N_A_27_47#_c_662_n N_X_c_1788_n 3.04151e-19 $X=15.215 $Y=1.41 $X2=0 $Y2=0
cc_814 N_A_27_47#_c_663_n N_X_c_1788_n 0.00188422f $X=15.685 $Y=1.41 $X2=0 $Y2=0
cc_815 N_A_27_47#_c_639_n X 4.17833e-19 $X=14.72 $Y=0.995 $X2=0 $Y2=0
cc_816 N_A_27_47#_c_661_n X 3.87571e-19 $X=14.745 $Y=1.41 $X2=0 $Y2=0
cc_817 N_A_27_47#_c_662_n X 0.00245231f $X=15.215 $Y=1.41 $X2=0 $Y2=0
cc_818 N_A_27_47#_c_640_n X 0.00278394f $X=15.24 $Y=0.995 $X2=0 $Y2=0
cc_819 N_A_27_47#_c_641_n X 0.00487628f $X=15.66 $Y=0.995 $X2=0 $Y2=0
cc_820 N_A_27_47#_c_663_n X 0.00450039f $X=15.685 $Y=1.41 $X2=0 $Y2=0
cc_821 N_A_27_47#_c_642_n X 0.00880356f $X=14.66 $Y=1.16 $X2=0 $Y2=0
cc_822 N_A_27_47#_c_651_n X 0.0511382f $X=15.66 $Y=1.202 $X2=0 $Y2=0
cc_823 N_A_27_47#_c_679_n N_A_119_47#_M1016_s 0.0028519f $X=1.065 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_824 N_A_27_47#_c_648_n N_A_119_47#_M1016_s 0.00312756f $X=9.615 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_825 N_A_27_47#_c_682_n N_A_119_47#_M1051_s 0.0028519f $X=2.005 $Y=0.402 $X2=0
+ $Y2=0
cc_826 N_A_27_47#_c_648_n N_A_119_47#_M1051_s 0.00312756f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_827 N_A_27_47#_M1058_d N_A_119_47#_c_1871_n 0.00360577f $X=1.955 $Y=0.235
+ $X2=0 $Y2=0
cc_828 N_A_27_47#_c_665_n N_A_119_47#_c_1871_n 0.00930103f $X=2.14 $Y=1.66 $X2=0
+ $Y2=0
cc_829 N_A_27_47#_c_644_n N_A_119_47#_c_1871_n 0.0184232f $X=2.14 $Y=0.385 $X2=0
+ $Y2=0
cc_830 N_A_27_47#_c_682_n N_A_119_47#_c_1871_n 0.0030195f $X=2.005 $Y=0.402
+ $X2=0 $Y2=0
cc_831 N_A_27_47#_c_648_n N_A_119_47#_c_1871_n 0.031319f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_832 N_A_27_47#_c_648_n N_A_119_47#_c_1894_n 0.0181814f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_833 N_A_27_47#_c_648_n N_A_119_47#_c_1872_n 0.0168956f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_834 N_A_27_47#_c_648_n N_A_119_47#_c_1902_n 0.0176612f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_835 N_A_27_47#_c_679_n N_A_119_47#_c_1873_n 0.0124302f $X=1.065 $Y=0.4 $X2=0
+ $Y2=0
cc_836 N_A_27_47#_c_648_n N_A_119_47#_c_1873_n 0.00974243f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_837 N_A_27_47#_c_690_n N_A_119_47#_c_1873_n 8.37317e-19 $X=0.405 $Y=0.51
+ $X2=0 $Y2=0
cc_838 N_A_27_47#_c_649_n N_A_119_47#_c_1873_n 0.0134636f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_839 N_A_27_47#_M1040_d N_A_119_47#_c_1874_n 0.00260599f $X=1.015 $Y=0.235
+ $X2=0 $Y2=0
cc_840 N_A_27_47#_c_679_n N_A_119_47#_c_1874_n 0.00176387f $X=1.065 $Y=0.4 $X2=0
+ $Y2=0
cc_841 N_A_27_47#_c_1004_p N_A_119_47#_c_1874_n 0.0156655f $X=1.335 $Y=0.4 $X2=0
+ $Y2=0
cc_842 N_A_27_47#_c_682_n N_A_119_47#_c_1874_n 0.00176387f $X=2.005 $Y=0.402
+ $X2=0 $Y2=0
cc_843 N_A_27_47#_c_648_n N_A_119_47#_c_1874_n 0.0133851f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_844 N_A_27_47#_c_682_n N_A_119_47#_c_1875_n 0.0124302f $X=2.005 $Y=0.402
+ $X2=0 $Y2=0
cc_845 N_A_27_47#_c_648_n N_A_119_47#_c_1875_n 0.00974243f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_846 N_A_27_47#_c_648_n N_VGND_M1000_s 0.00265275f $X=9.615 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_847 N_A_27_47#_c_648_n N_VGND_M1020_s 0.00339574f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_848 N_A_27_47#_c_648_n N_VGND_M1054_s 0.00419785f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_849 N_A_27_47#_c_648_n N_VGND_M1039_s 0.00166982f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_850 N_A_27_47#_c_648_n N_VGND_M1009_d 0.00339574f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_851 N_A_27_47#_c_648_n N_VGND_M1044_d 0.00265275f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_852 N_A_27_47#_c_644_n N_VGND_c_1954_n 0.0194114f $X=2.14 $Y=0.385 $X2=0
+ $Y2=0
cc_853 N_A_27_47#_c_648_n N_VGND_c_1954_n 0.010655f $X=9.615 $Y=0.51 $X2=0 $Y2=0
cc_854 N_A_27_47#_c_648_n N_VGND_c_1955_n 0.0102455f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_855 N_A_27_47#_c_648_n N_VGND_c_1956_n 0.0195957f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_856 N_A_27_47#_c_648_n N_VGND_c_1957_n 0.0159033f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_857 N_A_27_47#_c_648_n N_VGND_c_1958_n 0.0102455f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_858 N_A_27_47#_c_645_n N_VGND_c_1959_n 0.0194114f $X=8.015 $Y=0.402 $X2=0
+ $Y2=0
cc_859 N_A_27_47#_c_648_n N_VGND_c_1959_n 0.010655f $X=9.615 $Y=0.51 $X2=0 $Y2=0
cc_860 N_A_27_47#_c_630_n N_VGND_c_1960_n 0.00366701f $X=10.54 $Y=0.995 $X2=0
+ $Y2=0
cc_861 N_A_27_47#_c_642_n N_VGND_c_1960_n 0.0232464f $X=14.66 $Y=1.16 $X2=0
+ $Y2=0
cc_862 N_A_27_47#_c_646_n N_VGND_c_1960_n 0.0121207f $X=9.775 $Y=0.425 $X2=0
+ $Y2=0
cc_863 N_A_27_47#_c_729_n N_VGND_c_1960_n 0.00163721f $X=9.76 $Y=0.51 $X2=0
+ $Y2=0
cc_864 N_A_27_47#_c_650_n N_VGND_c_1960_n 0.0309572f $X=9.76 $Y=0.51 $X2=0 $Y2=0
cc_865 N_A_27_47#_c_631_n N_VGND_c_1961_n 0.00166854f $X=10.96 $Y=0.995 $X2=0
+ $Y2=0
cc_866 N_A_27_47#_c_632_n N_VGND_c_1961_n 0.00166854f $X=11.48 $Y=0.995 $X2=0
+ $Y2=0
cc_867 N_A_27_47#_c_633_n N_VGND_c_1962_n 0.00166854f $X=11.9 $Y=0.995 $X2=0
+ $Y2=0
cc_868 N_A_27_47#_c_634_n N_VGND_c_1962_n 0.00166854f $X=12.42 $Y=0.995 $X2=0
+ $Y2=0
cc_869 N_A_27_47#_c_635_n N_VGND_c_1963_n 0.00166854f $X=12.84 $Y=0.995 $X2=0
+ $Y2=0
cc_870 N_A_27_47#_c_636_n N_VGND_c_1963_n 0.00166854f $X=13.36 $Y=0.995 $X2=0
+ $Y2=0
cc_871 N_A_27_47#_c_637_n N_VGND_c_1964_n 0.00166854f $X=13.78 $Y=0.995 $X2=0
+ $Y2=0
cc_872 N_A_27_47#_c_638_n N_VGND_c_1964_n 0.00166854f $X=14.3 $Y=0.995 $X2=0
+ $Y2=0
cc_873 N_A_27_47#_c_639_n N_VGND_c_1965_n 0.00166854f $X=14.72 $Y=0.995 $X2=0
+ $Y2=0
cc_874 N_A_27_47#_c_640_n N_VGND_c_1965_n 0.00166854f $X=15.24 $Y=0.995 $X2=0
+ $Y2=0
cc_875 N_A_27_47#_c_641_n N_VGND_c_1966_n 0.00366701f $X=15.66 $Y=0.995 $X2=0
+ $Y2=0
cc_876 N_A_27_47#_c_648_n N_VGND_c_1967_n 0.00124714f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_877 N_A_27_47#_c_648_n N_VGND_c_1969_n 0.00156886f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_878 N_A_27_47#_c_648_n N_VGND_c_1971_n 0.00189058f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_879 N_A_27_47#_c_648_n N_VGND_c_1973_n 0.00156886f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_880 N_A_27_47#_c_648_n N_VGND_c_1975_n 0.00124714f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_881 N_A_27_47#_c_645_n N_VGND_c_1977_n 0.108576f $X=8.015 $Y=0.402 $X2=0
+ $Y2=0
cc_882 N_A_27_47#_c_646_n N_VGND_c_1977_n 0.0209073f $X=9.775 $Y=0.425 $X2=0
+ $Y2=0
cc_883 N_A_27_47#_c_648_n N_VGND_c_1977_n 0.0015579f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_884 N_A_27_47#_c_643_n N_VGND_c_1979_n 0.0209073f $X=0.245 $Y=0.425 $X2=0
+ $Y2=0
cc_885 N_A_27_47#_c_679_n N_VGND_c_1979_n 0.108576f $X=1.065 $Y=0.4 $X2=0 $Y2=0
cc_886 N_A_27_47#_c_648_n N_VGND_c_1979_n 0.0015579f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_887 N_A_27_47#_c_630_n N_VGND_c_1980_n 0.00541359f $X=10.54 $Y=0.995 $X2=0
+ $Y2=0
cc_888 N_A_27_47#_c_631_n N_VGND_c_1980_n 0.00423334f $X=10.96 $Y=0.995 $X2=0
+ $Y2=0
cc_889 N_A_27_47#_c_632_n N_VGND_c_1981_n 0.00423334f $X=11.48 $Y=0.995 $X2=0
+ $Y2=0
cc_890 N_A_27_47#_c_633_n N_VGND_c_1981_n 0.00423334f $X=11.9 $Y=0.995 $X2=0
+ $Y2=0
cc_891 N_A_27_47#_c_634_n N_VGND_c_1982_n 0.00423334f $X=12.42 $Y=0.995 $X2=0
+ $Y2=0
cc_892 N_A_27_47#_c_635_n N_VGND_c_1982_n 0.00423334f $X=12.84 $Y=0.995 $X2=0
+ $Y2=0
cc_893 N_A_27_47#_c_636_n N_VGND_c_1983_n 0.00423334f $X=13.36 $Y=0.995 $X2=0
+ $Y2=0
cc_894 N_A_27_47#_c_637_n N_VGND_c_1983_n 0.00423334f $X=13.78 $Y=0.995 $X2=0
+ $Y2=0
cc_895 N_A_27_47#_c_638_n N_VGND_c_1984_n 0.00423334f $X=14.3 $Y=0.995 $X2=0
+ $Y2=0
cc_896 N_A_27_47#_c_639_n N_VGND_c_1984_n 0.00423334f $X=14.72 $Y=0.995 $X2=0
+ $Y2=0
cc_897 N_A_27_47#_c_640_n N_VGND_c_1985_n 0.00423334f $X=15.24 $Y=0.995 $X2=0
+ $Y2=0
cc_898 N_A_27_47#_c_641_n N_VGND_c_1985_n 0.00541359f $X=15.66 $Y=0.995 $X2=0
+ $Y2=0
cc_899 N_A_27_47#_M1016_d N_VGND_c_1987_n 0.00133169f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_900 N_A_27_47#_M1040_d N_VGND_c_1987_n 0.00166809f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_901 N_A_27_47#_M1058_d N_VGND_c_1987_n 0.0014225f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_902 N_A_27_47#_M1004_d N_VGND_c_1987_n 0.0014225f $X=7.755 $Y=0.235 $X2=0
+ $Y2=0
cc_903 N_A_27_47#_M1011_d N_VGND_c_1987_n 0.00166809f $X=8.635 $Y=0.235 $X2=0
+ $Y2=0
cc_904 N_A_27_47#_M1046_d N_VGND_c_1987_n 0.00133169f $X=9.575 $Y=0.235 $X2=0
+ $Y2=0
cc_905 N_A_27_47#_c_630_n N_VGND_c_1987_n 0.0108276f $X=10.54 $Y=0.995 $X2=0
+ $Y2=0
cc_906 N_A_27_47#_c_631_n N_VGND_c_1987_n 0.00595861f $X=10.96 $Y=0.995 $X2=0
+ $Y2=0
cc_907 N_A_27_47#_c_632_n N_VGND_c_1987_n 0.00595861f $X=11.48 $Y=0.995 $X2=0
+ $Y2=0
cc_908 N_A_27_47#_c_633_n N_VGND_c_1987_n 0.00595861f $X=11.9 $Y=0.995 $X2=0
+ $Y2=0
cc_909 N_A_27_47#_c_634_n N_VGND_c_1987_n 0.00595861f $X=12.42 $Y=0.995 $X2=0
+ $Y2=0
cc_910 N_A_27_47#_c_635_n N_VGND_c_1987_n 0.00595861f $X=12.84 $Y=0.995 $X2=0
+ $Y2=0
cc_911 N_A_27_47#_c_636_n N_VGND_c_1987_n 0.00595861f $X=13.36 $Y=0.995 $X2=0
+ $Y2=0
cc_912 N_A_27_47#_c_637_n N_VGND_c_1987_n 0.00595861f $X=13.78 $Y=0.995 $X2=0
+ $Y2=0
cc_913 N_A_27_47#_c_638_n N_VGND_c_1987_n 0.00595861f $X=14.3 $Y=0.995 $X2=0
+ $Y2=0
cc_914 N_A_27_47#_c_639_n N_VGND_c_1987_n 0.00595861f $X=14.72 $Y=0.995 $X2=0
+ $Y2=0
cc_915 N_A_27_47#_c_640_n N_VGND_c_1987_n 0.00595861f $X=15.24 $Y=0.995 $X2=0
+ $Y2=0
cc_916 N_A_27_47#_c_641_n N_VGND_c_1987_n 0.0108276f $X=15.66 $Y=0.995 $X2=0
+ $Y2=0
cc_917 N_A_27_47#_c_643_n N_VGND_c_1987_n 0.00348214f $X=0.245 $Y=0.425 $X2=0
+ $Y2=0
cc_918 N_A_27_47#_c_679_n N_VGND_c_1987_n 0.0179106f $X=1.065 $Y=0.4 $X2=0 $Y2=0
cc_919 N_A_27_47#_c_645_n N_VGND_c_1987_n 0.0179106f $X=8.015 $Y=0.402 $X2=0
+ $Y2=0
cc_920 N_A_27_47#_c_646_n N_VGND_c_1987_n 0.00348214f $X=9.775 $Y=0.425 $X2=0
+ $Y2=0
cc_921 N_A_27_47#_c_648_n N_VGND_c_1987_n 0.782671f $X=9.615 $Y=0.51 $X2=0 $Y2=0
cc_922 N_A_27_47#_c_690_n N_VGND_c_1987_n 0.0283252f $X=0.405 $Y=0.51 $X2=0
+ $Y2=0
cc_923 N_A_27_47#_c_729_n N_VGND_c_1987_n 0.0283252f $X=9.76 $Y=0.51 $X2=0 $Y2=0
cc_924 N_A_27_47#_c_719_n N_A_1163_47#_M1004_s 0.0028519f $X=8.685 $Y=0.4 $X2=0
+ $Y2=0
cc_925 N_A_27_47#_c_648_n N_A_1163_47#_M1004_s 0.00312756f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_926 N_A_27_47#_c_712_n N_A_1163_47#_M1041_s 0.0028519f $X=9.625 $Y=0.34 $X2=0
+ $Y2=0
cc_927 N_A_27_47#_c_648_n N_A_1163_47#_M1041_s 0.00312756f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_928 N_A_27_47#_c_648_n N_A_1163_47#_c_2225_n 0.0176673f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_929 N_A_27_47#_c_648_n N_A_1163_47#_c_2218_n 0.0168956f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_930 N_A_27_47#_c_648_n N_A_1163_47#_c_2236_n 0.0181875f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_931 N_A_27_47#_M1004_d N_A_1163_47#_c_2221_n 0.00360577f $X=7.755 $Y=0.235
+ $X2=0 $Y2=0
cc_932 N_A_27_47#_c_667_n N_A_1163_47#_c_2221_n 0.00930103f $X=7.88 $Y=1.66
+ $X2=0 $Y2=0
cc_933 N_A_27_47#_c_645_n N_A_1163_47#_c_2221_n 0.0184232f $X=8.015 $Y=0.402
+ $X2=0 $Y2=0
cc_934 N_A_27_47#_c_719_n N_A_1163_47#_c_2221_n 0.0030195f $X=8.685 $Y=0.4 $X2=0
+ $Y2=0
cc_935 N_A_27_47#_c_648_n N_A_1163_47#_c_2221_n 0.031319f $X=9.615 $Y=0.51 $X2=0
+ $Y2=0
cc_936 N_A_27_47#_c_719_n N_A_1163_47#_c_2222_n 0.0124302f $X=8.685 $Y=0.4 $X2=0
+ $Y2=0
cc_937 N_A_27_47#_c_648_n N_A_1163_47#_c_2222_n 0.00974243f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_938 N_A_27_47#_c_712_n N_A_1163_47#_c_2223_n 0.0124302f $X=9.625 $Y=0.34
+ $X2=0 $Y2=0
cc_939 N_A_27_47#_c_648_n N_A_1163_47#_c_2223_n 0.00974243f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_940 N_A_27_47#_c_729_n N_A_1163_47#_c_2223_n 8.37317e-19 $X=9.76 $Y=0.51
+ $X2=0 $Y2=0
cc_941 N_A_27_47#_c_650_n N_A_1163_47#_c_2223_n 0.0134636f $X=9.76 $Y=0.51 $X2=0
+ $Y2=0
cc_942 N_A_27_47#_M1011_d N_A_1163_47#_c_2224_n 0.00260599f $X=8.635 $Y=0.235
+ $X2=0 $Y2=0
cc_943 N_A_27_47#_c_712_n N_A_1163_47#_c_2224_n 0.00176387f $X=9.625 $Y=0.34
+ $X2=0 $Y2=0
cc_944 N_A_27_47#_c_719_n N_A_1163_47#_c_2224_n 0.00176387f $X=8.685 $Y=0.4
+ $X2=0 $Y2=0
cc_945 N_A_27_47#_c_1108_p N_A_1163_47#_c_2224_n 0.0156655f $X=8.955 $Y=0.4
+ $X2=0 $Y2=0
cc_946 N_A_27_47#_c_648_n N_A_1163_47#_c_2224_n 0.0133851f $X=9.615 $Y=0.51
+ $X2=0 $Y2=0
cc_947 N_A_117_297#_c_1110_n N_VPWR_M1006_d 2.47951e-19 $X=5.805 $Y=1.87
+ $X2=-0.19 $Y2=1.305
cc_948 N_A_117_297#_c_1110_n N_VPWR_M1015_d 0.00235741f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_949 N_A_117_297#_c_1110_n N_VPWR_M1056_d 4.13644e-19 $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_950 N_A_117_297#_c_1110_n N_VPWR_M1032_d 3.27824e-19 $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_951 N_A_117_297#_c_1145_n N_VPWR_M1029_s 0.00315544f $X=6.725 $Y=1.58 $X2=0
+ $Y2=0
cc_952 N_A_117_297#_c_1161_n N_VPWR_M1029_s 0.00235741f $X=6.745 $Y=1.87 $X2=0
+ $Y2=0
cc_953 N_A_117_297#_c_1110_n N_VPWR_c_1242_n 0.0275493f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_954 N_A_117_297#_c_1110_n N_VPWR_c_1243_n 0.0101688f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_955 N_A_117_297#_c_1110_n N_VPWR_c_1244_n 0.0179122f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_956 N_A_117_297#_c_1110_n N_VPWR_c_1245_n 0.0157778f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_957 N_A_117_297#_c_1164_n N_VPWR_c_1245_n 6.68271e-19 $X=6.095 $Y=1.87 $X2=0
+ $Y2=0
cc_958 N_A_117_297#_c_1165_n N_VPWR_c_1245_n 0.0336199f $X=5.95 $Y=1.87 $X2=0
+ $Y2=0
cc_959 N_A_117_297#_c_1145_n N_VPWR_c_1246_n 0.0130979f $X=6.725 $Y=1.58 $X2=0
+ $Y2=0
cc_960 N_A_117_297#_c_1161_n N_VPWR_c_1246_n 0.0101688f $X=6.745 $Y=1.87 $X2=0
+ $Y2=0
cc_961 N_A_117_297#_c_1164_n N_VPWR_c_1246_n 3.34135e-19 $X=6.095 $Y=1.87 $X2=0
+ $Y2=0
cc_962 N_A_117_297#_c_1165_n N_VPWR_c_1246_n 0.0268237f $X=5.95 $Y=1.87 $X2=0
+ $Y2=0
cc_963 N_A_117_297#_c_1168_n N_VPWR_c_1246_n 3.34135e-19 $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_964 N_A_117_297#_c_1169_n N_VPWR_c_1246_n 0.0268237f $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_965 N_A_117_297#_c_1168_n N_VPWR_c_1247_n 0.00114399f $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_966 N_A_117_297#_c_1169_n N_VPWR_c_1247_n 0.0307767f $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_967 N_A_117_297#_c_1165_n N_VPWR_c_1261_n 0.0189467f $X=5.95 $Y=1.87 $X2=0
+ $Y2=0
cc_968 N_A_117_297#_c_1169_n N_VPWR_c_1263_n 0.0189467f $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_969 N_A_117_297#_M1002_s N_VPWR_c_1241_n 0.00184842f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_970 N_A_117_297#_M1035_s N_VPWR_c_1241_n 0.00184842f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_971 N_A_117_297#_M1005_d N_VPWR_c_1241_n 0.00130534f $X=5.805 $Y=1.485 $X2=0
+ $Y2=0
cc_972 N_A_117_297#_M1036_d N_VPWR_c_1241_n 0.00130534f $X=6.745 $Y=1.485 $X2=0
+ $Y2=0
cc_973 N_A_117_297#_c_1123_n N_VPWR_c_1241_n 0.030387f $X=1.525 $Y=1.87 $X2=0
+ $Y2=0
cc_974 N_A_117_297#_c_1126_n N_VPWR_c_1241_n 0.0145656f $X=0.875 $Y=1.87 $X2=0
+ $Y2=0
cc_975 N_A_117_297#_c_1110_n N_VPWR_c_1241_n 0.0547302f $X=5.805 $Y=1.87 $X2=0
+ $Y2=0
cc_976 N_A_117_297#_c_1130_n N_VPWR_c_1241_n 0.0145656f $X=1.815 $Y=1.87 $X2=0
+ $Y2=0
cc_977 N_A_117_297#_c_1165_n N_VPWR_c_1241_n 0.00347454f $X=5.95 $Y=1.87 $X2=0
+ $Y2=0
cc_978 N_A_117_297#_c_1169_n N_VPWR_c_1241_n 0.00347454f $X=6.89 $Y=1.87 $X2=0
+ $Y2=0
cc_979 N_A_117_297#_c_1110_n N_A_597_297#_c_1518_n 0.020688f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_980 N_A_117_297#_c_1110_n N_A_597_297#_c_1530_n 0.0498761f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_981 N_A_117_297#_c_1110_n N_A_597_297#_c_1599_n 0.0249445f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_982 N_A_117_297#_c_1110_n N_A_597_297#_c_1514_n 0.121254f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_983 N_A_117_297#_c_1161_n N_A_597_297#_c_1514_n 0.0498761f $X=6.745 $Y=1.87
+ $X2=0 $Y2=0
cc_984 N_A_117_297#_c_1164_n N_A_597_297#_c_1514_n 0.0249445f $X=6.095 $Y=1.87
+ $X2=0 $Y2=0
cc_985 N_A_117_297#_c_1165_n N_A_597_297#_c_1514_n 0.0160893f $X=5.95 $Y=1.87
+ $X2=0 $Y2=0
cc_986 N_A_117_297#_c_1168_n N_A_597_297#_c_1514_n 0.0249445f $X=6.89 $Y=1.87
+ $X2=0 $Y2=0
cc_987 N_A_117_297#_c_1169_n N_A_597_297#_c_1514_n 0.0168062f $X=6.89 $Y=1.87
+ $X2=0 $Y2=0
cc_988 N_A_117_297#_c_1110_n N_A_597_297#_c_1606_n 0.0249445f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_989 N_A_117_297#_c_1168_n N_A_597_297#_c_1517_n 0.00975633f $X=6.89 $Y=1.87
+ $X2=0 $Y2=0
cc_990 N_A_117_297#_c_1110_n N_A_597_297#_c_1535_n 0.0185376f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_991 N_A_117_297#_c_1110_n N_A_597_297#_c_1538_n 0.0182983f $X=5.805 $Y=1.87
+ $X2=0 $Y2=0
cc_992 N_VPWR_c_1241_n N_A_597_297#_M1006_s 0.00120859f $X=16.33 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_993 N_VPWR_c_1241_n N_A_597_297#_M1042_s 0.00120859f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_994 N_VPWR_c_1241_n N_A_597_297#_M1008_d 0.00184842f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_995 N_VPWR_c_1241_n N_A_597_297#_M1018_d 0.00184842f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_996 N_VPWR_M1015_d N_A_597_297#_c_1518_n 0.0031522f $X=3.455 $Y=1.485 $X2=0
+ $Y2=0
cc_997 N_VPWR_c_1243_n N_A_597_297#_c_1518_n 0.0130979f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_998 N_VPWR_c_1243_n N_A_597_297#_c_1530_n 0.0153241f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_999 N_VPWR_c_1255_n N_A_597_297#_c_1530_n 8.28225e-19 $X=3.465 $Y=2.72 $X2=0
+ $Y2=0
cc_1000 N_VPWR_c_1257_n N_A_597_297#_c_1530_n 8.28225e-19 $X=4.405 $Y=2.72 $X2=0
+ $Y2=0
cc_1001 N_VPWR_c_1241_n N_A_597_297#_c_1530_n 0.0538021f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1002 N_VPWR_c_1242_n N_A_597_297#_c_1599_n 0.00167228f $X=2.66 $Y=1.66 $X2=0
+ $Y2=0
cc_1003 N_VPWR_c_1243_n N_A_597_297#_c_1599_n 6.68271e-19 $X=3.6 $Y=2 $X2=0
+ $Y2=0
cc_1004 N_VPWR_c_1241_n N_A_597_297#_c_1599_n 0.0282533f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1005 N_VPWR_M1056_d N_A_597_297#_c_1514_n 2.3593e-19 $X=4.395 $Y=1.485 $X2=0
+ $Y2=0
cc_1006 N_VPWR_M1032_d N_A_597_297#_c_1514_n 2.3593e-19 $X=5.335 $Y=1.485 $X2=0
+ $Y2=0
cc_1007 N_VPWR_M1049_s N_A_597_297#_c_1514_n 3.49821e-19 $X=7.215 $Y=1.485 $X2=0
+ $Y2=0
cc_1008 N_VPWR_c_1244_n N_A_597_297#_c_1514_n 0.0154913f $X=4.54 $Y=1.66 $X2=0
+ $Y2=0
cc_1009 N_VPWR_c_1245_n N_A_597_297#_c_1514_n 0.0154913f $X=5.48 $Y=1.66 $X2=0
+ $Y2=0
cc_1010 N_VPWR_c_1246_n N_A_597_297#_c_1514_n 0.0153241f $X=6.42 $Y=2 $X2=0
+ $Y2=0
cc_1011 N_VPWR_c_1247_n N_A_597_297#_c_1514_n 0.0254189f $X=7.36 $Y=1.66 $X2=0
+ $Y2=0
cc_1012 N_VPWR_c_1257_n N_A_597_297#_c_1514_n 8.28225e-19 $X=4.405 $Y=2.72 $X2=0
+ $Y2=0
cc_1013 N_VPWR_c_1259_n N_A_597_297#_c_1514_n 0.00185529f $X=5.345 $Y=2.72 $X2=0
+ $Y2=0
cc_1014 N_VPWR_c_1261_n N_A_597_297#_c_1514_n 0.00185529f $X=6.285 $Y=2.72 $X2=0
+ $Y2=0
cc_1015 N_VPWR_c_1263_n N_A_597_297#_c_1514_n 0.00185529f $X=7.225 $Y=2.72 $X2=0
+ $Y2=0
cc_1016 N_VPWR_c_1265_n N_A_597_297#_c_1514_n 9.47375e-19 $X=10.145 $Y=2.72
+ $X2=0 $Y2=0
cc_1017 N_VPWR_c_1241_n N_A_597_297#_c_1514_n 0.288483f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1018 N_VPWR_c_1243_n N_A_597_297#_c_1606_n 6.68271e-19 $X=3.6 $Y=2 $X2=0
+ $Y2=0
cc_1019 N_VPWR_c_1244_n N_A_597_297#_c_1606_n 6.68271e-19 $X=4.54 $Y=1.66 $X2=0
+ $Y2=0
cc_1020 N_VPWR_c_1241_n N_A_597_297#_c_1606_n 0.0282533f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1021 N_VPWR_c_1241_n N_A_597_297#_c_1516_n 0.0256871f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1022 N_VPWR_c_1247_n N_A_597_297#_c_1517_n 0.00800317f $X=7.36 $Y=1.66 $X2=0
+ $Y2=0
cc_1023 N_VPWR_c_1241_n N_A_597_297#_c_1561_n 0.030387f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1024 N_VPWR_c_1241_n N_A_597_297#_c_1564_n 0.0145656f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1025 N_VPWR_c_1242_n N_A_597_297#_c_1535_n 0.0318001f $X=2.66 $Y=1.66 $X2=0
+ $Y2=0
cc_1026 N_VPWR_c_1243_n N_A_597_297#_c_1535_n 0.0268237f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_1027 N_VPWR_c_1255_n N_A_597_297#_c_1535_n 0.0189467f $X=3.465 $Y=2.72 $X2=0
+ $Y2=0
cc_1028 N_VPWR_c_1241_n N_A_597_297#_c_1535_n 0.00325355f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1029 N_VPWR_c_1243_n N_A_597_297#_c_1538_n 0.0268237f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_1030 N_VPWR_c_1244_n N_A_597_297#_c_1538_n 0.0336199f $X=4.54 $Y=1.66 $X2=0
+ $Y2=0
cc_1031 N_VPWR_c_1257_n N_A_597_297#_c_1538_n 0.0189467f $X=4.405 $Y=2.72 $X2=0
+ $Y2=0
cc_1032 N_VPWR_c_1241_n N_A_597_297#_c_1538_n 0.00313501f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1033 N_VPWR_c_1241_n N_A_597_297#_c_1568_n 0.0145656f $X=16.33 $Y=2.72 $X2=0
+ $Y2=0
cc_1034 N_VPWR_c_1241_n N_X_M1003_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1241_n N_X_M1013_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1036 N_VPWR_c_1241_n N_X_M1022_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1241_n N_X_M1031_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1038 N_VPWR_c_1241_n N_X_M1045_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1039 N_VPWR_c_1241_n N_X_M1053_s 0.00231261f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1040 N_VPWR_c_1268_n N_X_c_1669_n 0.0189467f $X=11.085 $Y=2.72 $X2=0 $Y2=0
cc_1041 N_VPWR_c_1241_n N_X_c_1669_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1042 N_VPWR_M1007_d N_X_c_1680_n 0.00334388f $X=11.075 $Y=1.485 $X2=0 $Y2=0
cc_1043 N_VPWR_c_1249_n N_X_c_1680_n 0.0143191f $X=11.22 $Y=2 $X2=0 $Y2=0
cc_1044 N_VPWR_c_1269_n N_X_c_1688_n 0.0189467f $X=12.025 $Y=2.72 $X2=0 $Y2=0
cc_1045 N_VPWR_c_1241_n N_X_c_1688_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1046 N_VPWR_M1019_d N_X_c_1696_n 0.00334388f $X=12.015 $Y=1.485 $X2=0 $Y2=0
cc_1047 N_VPWR_c_1250_n N_X_c_1696_n 0.0143191f $X=12.16 $Y=2 $X2=0 $Y2=0
cc_1048 N_VPWR_c_1270_n N_X_c_1704_n 0.0189467f $X=12.965 $Y=2.72 $X2=0 $Y2=0
cc_1049 N_VPWR_c_1241_n N_X_c_1704_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1050 N_VPWR_M1028_d N_X_c_1712_n 0.00334388f $X=12.955 $Y=1.485 $X2=0 $Y2=0
cc_1051 N_VPWR_c_1251_n N_X_c_1712_n 0.0143191f $X=13.1 $Y=2 $X2=0 $Y2=0
cc_1052 N_VPWR_c_1271_n N_X_c_1720_n 0.0189467f $X=13.905 $Y=2.72 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1241_n N_X_c_1720_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1054 N_VPWR_M1037_d N_X_c_1728_n 0.00334388f $X=13.895 $Y=1.485 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1252_n N_X_c_1728_n 0.0143191f $X=14.04 $Y=2 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1272_n N_X_c_1736_n 0.0189467f $X=14.845 $Y=2.72 $X2=0 $Y2=0
cc_1057 N_VPWR_c_1241_n N_X_c_1736_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1058 N_VPWR_M1050_d N_X_c_1744_n 0.00419277f $X=14.835 $Y=1.485 $X2=0 $Y2=0
cc_1059 N_VPWR_c_1253_n N_X_c_1744_n 0.0143191f $X=14.98 $Y=2 $X2=0 $Y2=0
cc_1060 N_VPWR_c_1273_n N_X_c_1751_n 0.0189467f $X=15.785 $Y=2.72 $X2=0 $Y2=0
cc_1061 N_VPWR_c_1241_n N_X_c_1751_n 0.0123132f $X=16.33 $Y=2.72 $X2=0 $Y2=0
cc_1062 N_VPWR_c_1242_n N_A_119_47#_c_1871_n 0.00823267f $X=2.66 $Y=1.66 $X2=0
+ $Y2=0
cc_1063 N_VPWR_c_1244_n N_VGND_c_1956_n 0.00829786f $X=4.54 $Y=1.66 $X2=0 $Y2=0
cc_1064 N_VPWR_c_1254_n N_VGND_c_1966_n 0.00920291f $X=15.92 $Y=1.66 $X2=0 $Y2=0
cc_1065 N_VPWR_c_1247_n N_A_1163_47#_c_2221_n 0.00823267f $X=7.36 $Y=1.66 $X2=0
+ $Y2=0
cc_1066 N_X_c_1652_n N_VGND_M1017_s 0.00281047f $X=11.525 $Y=0.815 $X2=0 $Y2=0
cc_1067 N_X_c_1654_n N_VGND_M1025_s 0.00281047f $X=12.465 $Y=0.815 $X2=0 $Y2=0
cc_1068 N_X_c_1655_n N_VGND_M1033_s 0.00281047f $X=13.405 $Y=0.815 $X2=0 $Y2=0
cc_1069 N_X_c_1656_n N_VGND_M1043_s 0.00277929f $X=14.345 $Y=0.815 $X2=0 $Y2=0
cc_1070 N_X_c_1657_n N_VGND_M1052_s 0.00281047f $X=15.285 $Y=0.815 $X2=0 $Y2=0
cc_1071 N_X_c_1653_n N_VGND_c_1960_n 0.00835241f $X=10.915 $Y=0.815 $X2=0 $Y2=0
cc_1072 N_X_c_1652_n N_VGND_c_1961_n 0.0191421f $X=11.525 $Y=0.815 $X2=0 $Y2=0
cc_1073 N_X_c_1654_n N_VGND_c_1962_n 0.0191421f $X=12.465 $Y=0.815 $X2=0 $Y2=0
cc_1074 N_X_c_1655_n N_VGND_c_1963_n 0.0191421f $X=13.405 $Y=0.815 $X2=0 $Y2=0
cc_1075 N_X_c_1656_n N_VGND_c_1964_n 0.0196153f $X=14.345 $Y=0.815 $X2=0 $Y2=0
cc_1076 N_X_c_1657_n N_VGND_c_1965_n 0.0191421f $X=15.285 $Y=0.815 $X2=0 $Y2=0
cc_1077 N_X_c_1786_n N_VGND_c_1966_n 0.00835241f $X=15.45 $Y=0.815 $X2=0 $Y2=0
cc_1078 N_X_c_1662_n N_VGND_c_1980_n 0.0188551f $X=10.75 $Y=0.42 $X2=0 $Y2=0
cc_1079 N_X_c_1652_n N_VGND_c_1980_n 0.00198695f $X=11.525 $Y=0.815 $X2=0 $Y2=0
cc_1080 N_X_c_1652_n N_VGND_c_1981_n 0.00198695f $X=11.525 $Y=0.815 $X2=0 $Y2=0
cc_1081 N_X_c_1684_n N_VGND_c_1981_n 0.0188551f $X=11.69 $Y=0.42 $X2=0 $Y2=0
cc_1082 N_X_c_1654_n N_VGND_c_1981_n 0.00198695f $X=12.465 $Y=0.815 $X2=0 $Y2=0
cc_1083 N_X_c_1654_n N_VGND_c_1982_n 0.00198695f $X=12.465 $Y=0.815 $X2=0 $Y2=0
cc_1084 N_X_c_1700_n N_VGND_c_1982_n 0.0188551f $X=12.63 $Y=0.42 $X2=0 $Y2=0
cc_1085 N_X_c_1655_n N_VGND_c_1982_n 0.00198695f $X=13.405 $Y=0.815 $X2=0 $Y2=0
cc_1086 N_X_c_1655_n N_VGND_c_1983_n 0.00198695f $X=13.405 $Y=0.815 $X2=0 $Y2=0
cc_1087 N_X_c_1716_n N_VGND_c_1983_n 0.0188551f $X=13.57 $Y=0.42 $X2=0 $Y2=0
cc_1088 N_X_c_1656_n N_VGND_c_1983_n 0.00198695f $X=14.345 $Y=0.815 $X2=0 $Y2=0
cc_1089 N_X_c_1656_n N_VGND_c_1984_n 0.00198695f $X=14.345 $Y=0.815 $X2=0 $Y2=0
cc_1090 N_X_c_1732_n N_VGND_c_1984_n 0.0188551f $X=14.51 $Y=0.42 $X2=0 $Y2=0
cc_1091 N_X_c_1657_n N_VGND_c_1984_n 0.00198695f $X=15.285 $Y=0.815 $X2=0 $Y2=0
cc_1092 N_X_c_1657_n N_VGND_c_1985_n 0.00198695f $X=15.285 $Y=0.815 $X2=0 $Y2=0
cc_1093 N_X_c_1748_n N_VGND_c_1985_n 0.0189039f $X=15.45 $Y=0.42 $X2=0 $Y2=0
cc_1094 N_X_M1014_d N_VGND_c_1987_n 0.00215201f $X=10.615 $Y=0.235 $X2=0 $Y2=0
cc_1095 N_X_M1021_d N_VGND_c_1987_n 0.00215201f $X=11.555 $Y=0.235 $X2=0 $Y2=0
cc_1096 N_X_M1027_d N_VGND_c_1987_n 0.00215201f $X=12.495 $Y=0.235 $X2=0 $Y2=0
cc_1097 N_X_M1034_d N_VGND_c_1987_n 0.00215201f $X=13.435 $Y=0.235 $X2=0 $Y2=0
cc_1098 N_X_M1047_d N_VGND_c_1987_n 0.00215201f $X=14.375 $Y=0.235 $X2=0 $Y2=0
cc_1099 N_X_M1055_d N_VGND_c_1987_n 0.00215201f $X=15.315 $Y=0.235 $X2=0 $Y2=0
cc_1100 N_X_c_1662_n N_VGND_c_1987_n 0.0122069f $X=10.75 $Y=0.42 $X2=0 $Y2=0
cc_1101 N_X_c_1652_n N_VGND_c_1987_n 0.00876562f $X=11.525 $Y=0.815 $X2=0 $Y2=0
cc_1102 N_X_c_1684_n N_VGND_c_1987_n 0.0122069f $X=11.69 $Y=0.42 $X2=0 $Y2=0
cc_1103 N_X_c_1654_n N_VGND_c_1987_n 0.00876562f $X=12.465 $Y=0.815 $X2=0 $Y2=0
cc_1104 N_X_c_1700_n N_VGND_c_1987_n 0.0122069f $X=12.63 $Y=0.42 $X2=0 $Y2=0
cc_1105 N_X_c_1655_n N_VGND_c_1987_n 0.00876562f $X=13.405 $Y=0.815 $X2=0 $Y2=0
cc_1106 N_X_c_1716_n N_VGND_c_1987_n 0.0122069f $X=13.57 $Y=0.42 $X2=0 $Y2=0
cc_1107 N_X_c_1656_n N_VGND_c_1987_n 0.00875312f $X=14.345 $Y=0.815 $X2=0 $Y2=0
cc_1108 N_X_c_1732_n N_VGND_c_1987_n 0.0122069f $X=14.51 $Y=0.42 $X2=0 $Y2=0
cc_1109 N_X_c_1657_n N_VGND_c_1987_n 0.00876562f $X=15.285 $Y=0.815 $X2=0 $Y2=0
cc_1110 N_X_c_1748_n N_VGND_c_1987_n 0.0122217f $X=15.45 $Y=0.42 $X2=0 $Y2=0
cc_1111 N_A_119_47#_c_1871_n N_VGND_M1000_s 0.00360038f $X=2.965 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_1112 N_A_119_47#_c_1872_n N_VGND_M1020_s 0.00260058f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_1113 N_A_119_47#_c_1871_n N_VGND_c_1954_n 0.0166436f $X=2.965 $Y=0.815 $X2=0
+ $Y2=0
cc_1114 N_A_119_47#_c_1894_n N_VGND_c_1954_n 0.0124989f $X=3.13 $Y=0.42 $X2=0
+ $Y2=0
cc_1115 N_A_119_47#_c_1894_n N_VGND_c_1955_n 0.0122463f $X=3.13 $Y=0.42 $X2=0
+ $Y2=0
cc_1116 N_A_119_47#_c_1872_n N_VGND_c_1955_n 0.015851f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_1117 N_A_119_47#_c_1902_n N_VGND_c_1955_n 0.0122463f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_1118 N_A_119_47#_c_1872_n N_VGND_c_1956_n 0.00835241f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_1119 N_A_119_47#_c_1902_n N_VGND_c_1956_n 0.0194177f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_1120 N_A_119_47#_c_1871_n N_VGND_c_1967_n 0.00178562f $X=2.965 $Y=0.815 $X2=0
+ $Y2=0
cc_1121 N_A_119_47#_c_1894_n N_VGND_c_1967_n 0.0188551f $X=3.13 $Y=0.42 $X2=0
+ $Y2=0
cc_1122 N_A_119_47#_c_1872_n N_VGND_c_1967_n 0.00178562f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_1123 N_A_119_47#_c_1872_n N_VGND_c_1969_n 0.00178562f $X=3.905 $Y=0.815 $X2=0
+ $Y2=0
cc_1124 N_A_119_47#_c_1902_n N_VGND_c_1969_n 0.0188551f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_1125 N_A_119_47#_c_1871_n N_VGND_c_1979_n 0.00286511f $X=2.965 $Y=0.815 $X2=0
+ $Y2=0
cc_1126 N_A_119_47#_M1016_s N_VGND_c_1987_n 0.00122387f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_1127 N_A_119_47#_M1051_s N_VGND_c_1987_n 0.00122387f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_1128 N_A_119_47#_M1000_d N_VGND_c_1987_n 0.00121469f $X=2.995 $Y=0.235 $X2=0
+ $Y2=0
cc_1129 N_A_119_47#_M1023_d N_VGND_c_1987_n 0.00121469f $X=3.935 $Y=0.235 $X2=0
+ $Y2=0
cc_1130 N_A_119_47#_c_1894_n N_VGND_c_1987_n 0.0034345f $X=3.13 $Y=0.42 $X2=0
+ $Y2=0
cc_1131 N_A_119_47#_c_1902_n N_VGND_c_1987_n 0.0034345f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_1132 N_VGND_c_1987_n N_A_1163_47#_M1001_s 0.00121469f $X=16.33 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1133 N_VGND_c_1987_n N_A_1163_47#_M1024_s 0.00121469f $X=16.33 $Y=0 $X2=0
+ $Y2=0
cc_1134 N_VGND_c_1987_n N_A_1163_47#_M1004_s 0.00122387f $X=16.33 $Y=0 $X2=0
+ $Y2=0
cc_1135 N_VGND_c_1987_n N_A_1163_47#_M1041_s 0.00122387f $X=16.33 $Y=0 $X2=0
+ $Y2=0
cc_1136 N_VGND_c_1957_n N_A_1163_47#_c_2225_n 0.0194177f $X=5.48 $Y=0.38 $X2=0
+ $Y2=0
cc_1137 N_VGND_c_1958_n N_A_1163_47#_c_2225_n 0.0122463f $X=6.42 $Y=0.38 $X2=0
+ $Y2=0
cc_1138 N_VGND_c_1973_n N_A_1163_47#_c_2225_n 0.0188551f $X=6.285 $Y=0 $X2=0
+ $Y2=0
cc_1139 N_VGND_c_1987_n N_A_1163_47#_c_2225_n 0.0034345f $X=16.33 $Y=0 $X2=0
+ $Y2=0
cc_1140 N_VGND_M1009_d N_A_1163_47#_c_2218_n 0.00260058f $X=6.235 $Y=0.235 $X2=0
+ $Y2=0
cc_1141 N_VGND_c_1958_n N_A_1163_47#_c_2218_n 0.015851f $X=6.42 $Y=0.38 $X2=0
+ $Y2=0
cc_1142 N_VGND_c_1973_n N_A_1163_47#_c_2218_n 0.00178562f $X=6.285 $Y=0 $X2=0
+ $Y2=0
cc_1143 N_VGND_c_1975_n N_A_1163_47#_c_2218_n 0.00178562f $X=7.225 $Y=0 $X2=0
+ $Y2=0
cc_1144 N_VGND_c_1957_n N_A_1163_47#_c_2219_n 0.00835241f $X=5.48 $Y=0.38 $X2=0
+ $Y2=0
cc_1145 N_VGND_c_1958_n N_A_1163_47#_c_2236_n 0.0122463f $X=6.42 $Y=0.38 $X2=0
+ $Y2=0
cc_1146 N_VGND_c_1959_n N_A_1163_47#_c_2236_n 0.0124989f $X=7.36 $Y=0.385 $X2=0
+ $Y2=0
cc_1147 N_VGND_c_1975_n N_A_1163_47#_c_2236_n 0.0188551f $X=7.225 $Y=0 $X2=0
+ $Y2=0
cc_1148 N_VGND_c_1987_n N_A_1163_47#_c_2236_n 0.0034345f $X=16.33 $Y=0 $X2=0
+ $Y2=0
cc_1149 N_VGND_M1044_d N_A_1163_47#_c_2221_n 0.00360038f $X=7.175 $Y=0.235 $X2=0
+ $Y2=0
cc_1150 N_VGND_c_1959_n N_A_1163_47#_c_2221_n 0.0166436f $X=7.36 $Y=0.385 $X2=0
+ $Y2=0
cc_1151 N_VGND_c_1975_n N_A_1163_47#_c_2221_n 0.00178562f $X=7.225 $Y=0 $X2=0
+ $Y2=0
cc_1152 N_VGND_c_1977_n N_A_1163_47#_c_2221_n 0.00286511f $X=10.145 $Y=0 $X2=0
+ $Y2=0
