* File: sky130_fd_sc_hdll__a21oi_2.spice
* Created: Thu Aug 27 18:53:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21oi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a21oi_2  VNB VPB A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A2_M1003_g A_123_47# VNB NSHORT L=0.15 W=0.65 AD=0.2145
+ AS=0.091 PD=1.96 PS=0.93 NRD=8.304 NRS=15.684 M=1 R=4.33333 SA=75000.3
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1008 A_123_47# N_A1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.091
+ AS=0.1235 PD=0.93 PS=1.03 NRD=15.684 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1005 A_315_47# N_A1_M1005_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.1235 PD=0.86 PS=1.03 NRD=9.228 NRS=9.228 M=1 R=4.33333 SA=75001.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A2_M1007_g A_315_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.06825 PD=1.03 PS=0.86 NRD=9.228 NRS=9.228 M=1 R=4.33333 SA=75001.6
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1007_d N_B1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.104 PD=1.03 PS=0.97 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B1_M1004_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2925 AS=0.104 PD=2.2 PS=0.97 NRD=34.152 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_27_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.29 PD=1.3 PS=2.58 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1000_d N_A1_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A1_M1006_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1006_d N_A2_M1011_g N_A_27_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1011_s N_B1_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_27_297#_M1010_d N_B1_M1010_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.37 AS=0.145 PD=2.74 PS=1.29 NRD=20.685 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX13_noxref noxref_12 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a21oi_2.pxi.spice"
*
.ends
*
*
