* File: sky130_fd_sc_hdll__sedfxbp_1.spice
* Created: Thu Aug 27 19:28:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sedfxbp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sedfxbp_1  VNB VPB CLK D DE SCD SCE VPWR Q_N Q VGND
* 
* VGND	VGND
* Q	Q
* Q_N	Q_N
* VPWR	VPWR
* SCE	SCE
* SCD	SCD
* DE	DE
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1033 N_VGND_M1033_d N_CLK_M1033_g N_A_27_47#_M1033_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_211_363#_M1002_d N_A_27_47#_M1002_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1040 A_413_47# N_D_M1040_g N_A_319_47#_M1040_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1344 PD=0.63 PS=1.48 NRD=14.28 NRS=15.708 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1041 N_VGND_M1041_d N_DE_M1041_g A_413_47# VNB NSHORT L=0.15 W=0.42 AD=0.126
+ AS=0.0441 PD=1.44 PS=0.63 NRD=9.996 NRS=14.28 M=1 R=2.8 SA=75000.6 SB=75000.2
+ A=0.063 P=1.14 MULT=1
MM1030 N_VGND_M1030_d N_DE_M1030_g N_A_455_324#_M1030_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.1302 PD=0.71 PS=1.46 NRD=1.428 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1031 A_779_47# N_A_455_324#_M1031_g N_VGND_M1030_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0966 AS=0.0609 PD=0.88 PS=0.71 NRD=49.992 NRS=1.428 M=1 R=2.8 SA=75000.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1007 N_A_319_47#_M1007_d N_A_851_264#_M1007_g A_779_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.0966 PD=0.69 PS=0.88 NRD=0 NRS=49.992 M=1 R=2.8
+ SA=75001.3 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_A_985_47#_M1015_d N_A_955_21#_M1015_g N_A_319_47#_M1007_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.1302 AS=0.0567 PD=1.46 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75001.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SCE_M1013_g N_A_955_21#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.1092 PD=0.79 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1034 A_1373_119# N_SCD_M1034_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0777 PD=0.63 PS=0.79 NRD=14.28 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1019 N_A_985_47#_M1019_d N_SCE_M1019_g A_1373_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.253777 AS=0.0441 PD=1.67462 PS=0.63 NRD=15.708 NRS=14.28 M=1 R=2.8
+ SA=75001.1 SB=75000.5 A=0.063 P=1.14 MULT=1
MM1011 N_A_1611_413#_M1011_d N_A_27_47#_M1011_g N_A_985_47#_M1019_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0702 AS=0.217523 PD=0.75 PS=1.43538 NRD=14.988 NRS=34.992
+ M=1 R=2.4 SA=75000.6 SB=75001.9 A=0.054 P=1.02 MULT=1
MM1038 A_1738_47# N_A_211_363#_M1038_g N_A_1611_413#_M1011_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0700615 AS=0.0702 PD=0.738462 PS=0.75 NRD=46.536 NRS=21.66 M=1
+ R=2.4 SA=75001.1 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1036 N_VGND_M1036_d N_A_1787_159#_M1036_g A_1738_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.116847 AS=0.0817385 PD=0.939057 PS=0.861538 NRD=14.28 NRS=39.888 M=1
+ R=2.8 SA=75001.4 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1043 N_A_1787_159#_M1043_d N_A_1611_413#_M1043_g N_VGND_M1036_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.178053 PD=1.8 PS=1.43094 NRD=0 NRS=40.308 M=1
+ R=4.26667 SA=75001.5 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1008 A_2181_47# N_A_1787_159#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0730154 AS=0.1302 PD=0.813077 PS=1.46 NRD=33.948 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1010 N_A_2266_413#_M1010_d N_A_211_363#_M1010_g A_2181_47# VNB NSHORT L=0.15
+ W=0.36 AD=0.0747 AS=0.0625846 PD=0.775 PS=0.696923 NRD=19.992 NRS=39.612 M=1
+ R=2.4 SA=75000.7 SB=75001.8 A=0.054 P=1.02 MULT=1
MM1039 A_2391_47# N_A_27_47#_M1039_g N_A_2266_413#_M1010_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0609231 AS=0.0747 PD=0.687692 PS=0.775 NRD=38.076 NRS=24.996 M=1
+ R=2.4 SA=75001.3 SB=75001.2 A=0.054 P=1.02 MULT=1
MM1020 N_VGND_M1020_d N_A_851_264#_M1020_g A_2391_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0910654 AS=0.0710769 PD=0.83215 PS=0.802308 NRD=38.568 NRS=32.628 M=1
+ R=2.8 SA=75001.5 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1027 N_Q_N_M1027_d N_A_851_264#_M1027_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.140935 PD=1.82 PS=1.28785 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_2266_413#_M1014_g N_A_851_264#_M1014_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0997009 AS=0.1092 PD=0.851776 PS=1.36 NRD=31.428 NRS=0 M=1
+ R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1001 N_Q_M1001_d N_A_2266_413#_M1001_g N_VGND_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.154299 PD=1.91 PS=1.31822 NRD=7.38 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1037 N_A_211_363#_M1037_d N_A_27_47#_M1037_g N_VPWR_M1006_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1018 A_409_369# N_D_M1018_g N_A_319_47#_M1018_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.1728 PD=0.87 PS=1.82 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1025 N_VPWR_M1025_d N_A_455_324#_M1025_g A_409_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1728 AS=0.0736 PD=1.82 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1005 N_VPWR_M1005_d N_DE_M1005_g N_A_455_324#_M1005_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0992 AS=0.1728 PD=0.95 PS=1.82 NRD=4.6098 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1021 A_787_369# N_DE_M1021_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1216 AS=0.0992 PD=1.02 PS=0.95 NRD=41.5473 NRS=4.6098 M=1 R=3.55556
+ SA=90000.7 SB=90001.3 A=0.1152 P=1.64 MULT=1
MM1022 N_A_319_47#_M1022_d N_A_851_264#_M1022_g A_787_369# VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1056 AS=0.1216 PD=0.97 PS=1.02 NRD=1.5366 NRS=41.5473 M=1
+ R=3.55556 SA=90001.2 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1026 N_A_985_47#_M1026_d N_SCE_M1026_g N_A_319_47#_M1022_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.2048 AS=0.1056 PD=1.92 PS=0.97 NRD=16.9223 NRS=13.8491 M=1
+ R=3.55556 SA=90001.7 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1017 N_VPWR_M1017_d N_SCE_M1017_g N_A_955_21#_M1017_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1328 AS=0.176 PD=1.055 PS=1.83 NRD=19.9955 NRS=3.0732 M=1
+ R=3.55556 SA=90000.2 SB=90002.9 A=0.1152 P=1.64 MULT=1
MM1032 A_1376_369# N_SCD_M1032_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.112 AS=0.1328 PD=0.99 PS=1.055 NRD=36.9178 NRS=21.5321 M=1 R=3.55556
+ SA=90000.8 SB=90002.3 A=0.1152 P=1.64 MULT=1
MM1012 N_A_985_47#_M1012_d N_A_955_21#_M1012_g A_1376_369# VPB PHIGHVT L=0.18
+ W=0.64 AD=0.168392 AS=0.112 PD=1.33434 PS=0.99 NRD=23.0687 NRS=36.9178 M=1
+ R=3.55556 SA=90001.3 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1023 N_A_1611_413#_M1023_d N_A_211_363#_M1023_g N_A_985_47#_M1012_d VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.06825 AS=0.110508 PD=0.745 PS=0.87566 NRD=9.3772
+ NRS=52.7566 M=1 R=2.33333 SA=90002 SB=90002 A=0.0756 P=1.2 MULT=1
MM1028 A_1712_413# N_A_27_47#_M1028_g N_A_1611_413#_M1023_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.08085 AS=0.06825 PD=0.805 PS=0.745 NRD=64.4781 NRS=11.7215 M=1
+ R=2.33333 SA=90002.5 SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1787_159#_M1024_g A_1712_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.132623 AS=0.08085 PD=0.918974 PS=0.805 NRD=102.007 NRS=64.4781 M=1
+ R=2.33333 SA=90003 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1000 N_A_1787_159#_M1000_d N_A_1611_413#_M1000_g N_VPWR_M1024_d VPB PHIGHVT
+ L=0.18 W=0.75 AD=0.2025 AS=0.236827 PD=2.04 PS=1.64103 NRD=1.3002 NRS=9.1802
+ M=1 R=4.16667 SA=90002.2 SB=90000.2 A=0.135 P=1.86 MULT=1
MM1003 A_2165_413# N_A_1787_159#_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.06825 AS=0.1134 PD=0.745 PS=1.38 NRD=50.4123 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1004 N_A_2266_413#_M1004_d N_A_27_47#_M1004_g A_2165_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.06825 PD=0.71 PS=0.745 NRD=2.3443 NRS=50.4123 M=1
+ R=2.33333 SA=90000.7 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1042 A_2360_413# N_A_211_363#_M1042_g N_A_2266_413#_M1004_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1029 AS=0.0609 PD=0.91 PS=0.71 NRD=89.1031 NRS=2.3443 M=1
+ R=2.33333 SA=90001.2 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1035 N_VPWR_M1035_d N_A_851_264#_M1035_g A_2360_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.1029 PD=0.801549 PS=0.91 NRD=34.0022 NRS=89.1031 M=1
+ R=2.33333 SA=90001.8 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1016 N_Q_N_M1016_d N_A_851_264#_M1016_g N_VPWR_M1035_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.215282 PD=2.54 PS=1.90845 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1029 N_VPWR_M1029_d N_A_2266_413#_M1029_g N_A_851_264#_M1029_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.126595 AS=0.1792 PD=1.05756 PS=1.84 NRD=21.5321 NRS=4.6098
+ M=1 R=3.55556 SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1009 N_Q_M1009_d N_A_2266_413#_M1009_g N_VPWR_M1029_d VPB PHIGHVT L=0.18 W=1
+ AD=0.315 AS=0.197805 PD=2.63 PS=1.65244 NRD=9.8303 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX44_noxref VNB VPB NWDIODE A=24.6228 P=34.59
pX45_noxref noxref_34 DE DE PROBETYPE=1
c_280 VPB 0 1.48265e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sedfxbp_1.pxi.spice"
*
.ends
*
*
