* File: sky130_fd_sc_hdll__nand4_4.spice
* Created: Wed Sep  2 08:38:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4_4.pex.spice"
.subckt sky130_fd_sc_hdll__nand4_4  VNB VPB D C B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1022 N_A_27_47#_M1022_d N_D_M1022_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003 A=0.0975 P=1.6 MULT=1
MM1023 N_A_27_47#_M1022_d N_D_M1023_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1031 N_A_27_47#_M1031_d N_D_M1031_g N_VGND_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1031_d N_C_M1012_g N_A_485_47#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1018 N_A_27_47#_M1018_d N_C_M1018_g N_A_485_47#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1025 N_A_27_47#_M1018_d N_C_M1025_g N_A_485_47#_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1027 N_A_27_47#_M1027_d N_C_M1027_g N_A_485_47#_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_883_47#_M1005_d N_B_M1005_g N_A_485_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1007 N_A_883_47#_M1007_d N_B_M1007_g N_A_485_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1015 N_A_883_47#_M1007_d N_B_M1015_g N_A_485_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1021 N_A_883_47#_M1021_d N_B_M1021_g N_A_485_47#_M1015_s VNB NSHORT L=0.15
+ W=0.65 AD=0.10725 AS=0.104 PD=0.98 PS=0.97 NRD=5.532 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1008 N_A_883_47#_M1021_d N_A_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.104 PD=0.98 PS=0.97 NRD=3.684 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1010 N_A_883_47#_M1010_d N_A_M1010_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1024 N_A_883_47#_M1010_d N_A_M1024_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1026 N_A_883_47#_M1026_d N_A_M1026_g N_Y_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_D_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90007.8 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_D_M1014_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90007.3 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1014_d N_D_M1020_g N_Y_M1020_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90006.9 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_D_M1028_g N_Y_M1020_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90006.4 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1028_d N_C_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90005.9 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90005.5 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1006_d N_C_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003 SB=90005
+ A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1 AD=0.405
+ AS=0.145 PD=1.81 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.405 PD=1.29 PS=1.81 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.5
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1003_d N_B_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.9
+ SB=90003.1 A=0.18 P=2.36 MULT=1
MM1019 N_Y_M1019_d N_B_M1019_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.4
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1029 N_Y_M1019_d N_B_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90005.9
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1004 N_Y_M1004_d N_A_M1004_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.175 PD=1.29 PS=1.35 NRD=0.9653 NRS=5.8903 M=1 R=5.55556 SA=90006.4
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_Y_M1004_d N_A_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.9
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1016 N_Y_M1016_d N_A_M1016_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.3
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1030 N_Y_M1016_d N_A_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=14.6296 P=21.44
pX33_noxref noxref_13 D D PROBETYPE=1
c_49 VNB 0 1.70629e-19 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hdll__nand4_4.pxi.spice"
*
.ends
*
*
