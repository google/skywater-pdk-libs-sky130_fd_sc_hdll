* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o221a_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_117_297# B2 a_305_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR A1 a_785_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_27_47# B1 a_307_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_27_47# B2 a_307_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_307_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR C1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_785_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_305_297# B2 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_117_297# C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_307_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR B1 a_305_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 X a_117_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR a_117_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 X a_117_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_117_297# A2 a_785_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_27_47# C1 a_117_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_307_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_117_297# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND A1 a_307_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_307_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_117_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VGND A2 a_307_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VGND a_117_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_305_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_785_297# A2 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
