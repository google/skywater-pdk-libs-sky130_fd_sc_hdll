* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
X0 a_1126_413# a_27_47# a_1344_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR SET_B a_702_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VPWR a_506_47# a_1044_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X3 a_1244_413# a_1288_261# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X4 Q a_1738_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND SET_B a_866_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_1344_47# a_1288_261# a_1416_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VGND a_1738_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_1126_413# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X9 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 a_636_47# a_702_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VGND a_1738_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VPWR D a_409_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X13 VPWR a_1126_413# a_1288_261# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X14 Q a_1738_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND D a_409_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 a_1738_47# a_1126_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X17 a_506_47# a_211_363# a_636_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X18 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1156_47# a_211_363# a_1126_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VPWR a_1738_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_506_47# a_27_47# a_610_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X22 a_610_413# a_702_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X23 a_1126_413# a_211_363# a_1244_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X24 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X25 VGND a_1738_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_1044_413# a_27_47# a_1126_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X27 a_409_329# a_27_47# a_506_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X28 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X29 a_702_21# a_506_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X30 a_409_329# a_211_363# a_506_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X31 a_866_47# a_506_47# a_702_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1416_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1738_47# a_1126_413# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 VGND a_1126_413# a_1288_261# VNB sky130_fd_pr__nfet_01v8 w=540000u l=150000u
X35 Q a_1738_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VGND a_506_47# a_1156_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 Q a_1738_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VPWR a_1738_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VPWR a_1738_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
