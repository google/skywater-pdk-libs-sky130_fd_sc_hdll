* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0






































































































































































































































































































































.subckt sky130_fd_sc_hdll__tap VGND VPWR
Xsky130_fd_sc_hdll__o22ai_2_0 sky130_fd_sc_hdll__o22ai_2_0/B2 sky130_fd_sc_hdll__o22ai_2_0/B1
+ sky130_fd_sc_hdll__o22ai_2_0/Y sky130_fd_sc_hdll__o22ai_2_0/A1 sky130_fd_sc_hdll__o22ai_2_0/A2
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o22ai_2
Xsky130_fd_sc_hdll__nand2_1_0 sky130_fd_sc_hdll__nand2_1_0/Y sky130_fd_sc_hdll__nand2_1_0/B
+ sky130_fd_sc_hdll__nand2_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_1
Xsky130_fd_sc_hdll__nor3_4_0 sky130_fd_sc_hdll__nor3_4_0/A sky130_fd_sc_hdll__nor3_4_0/C
+ sky130_fd_sc_hdll__nor3_4_0/B sky130_fd_sc_hdll__nor3_4_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_8 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21bo_1_0 sky130_fd_sc_hdll__a21bo_1_0/X sky130_fd_sc_hdll__a21bo_1_0/A1
+ sky130_fd_sc_hdll__a21bo_1_0/B1_N sky130_fd_sc_hdll__a21bo_1_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__a21bo_1
Xsky130_fd_sc_hdll__nand2b_2_0 sky130_fd_sc_hdll__nand2b_2_0/B sky130_fd_sc_hdll__nand2b_2_0/Y
+ sky130_fd_sc_hdll__nand2b_2_0/A_N VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2b_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_305 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_316 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_19 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a31oi_1_0 VGND VPWR sky130_fd_sc_hdll__a31oi_1_0/Y sky130_fd_sc_hdll__a31oi_1_0/B1
+ sky130_fd_sc_hdll__a31oi_1_0/A2 sky130_fd_sc_hdll__a31oi_1_0/A1 sky130_fd_sc_hdll__a31oi_1_0/A3
+ VPWR VGND sky130_fd_sc_hdll__a31oi_1
Xsky130_fd_sc_hdll__mux2i_1_0 sky130_fd_sc_hdll__mux2i_1_0/A1 sky130_fd_sc_hdll__mux2i_1_0/S
+ sky130_fd_sc_hdll__mux2i_1_0/A0 sky130_fd_sc_hdll__mux2i_1_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__mux2i_1
Xsky130_fd_sc_hdll__clkbuf_16_0 sky130_fd_sc_hdll__clkbuf_16_0/X sky130_fd_sc_hdll__clkbuf_16_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkbuf_16
Xsky130_fd_sc_hdll__o211ai_2_0 sky130_fd_sc_hdll__o211ai_2_0/A1 sky130_fd_sc_hdll__o211ai_2_0/A2
+ sky130_fd_sc_hdll__o211ai_2_0/B1 sky130_fd_sc_hdll__o211ai_2_0/Y sky130_fd_sc_hdll__o211ai_2_0/C1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211ai_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_102 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_113 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_124 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_135 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_146 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_157 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_179 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_168 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2b_1_0 sky130_fd_sc_hdll__or2b_1_0/A sky130_fd_sc_hdll__or2b_1_0/B_N
+ sky130_fd_sc_hdll__or2b_1_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2b_1
Xsky130_fd_sc_hdll__dlrtn_1_0 sky130_fd_sc_hdll__dlrtn_1_0/RESET_B sky130_fd_sc_hdll__dlrtn_1_0/D
+ sky130_fd_sc_hdll__dlrtn_1_0/GATE_N sky130_fd_sc_hdll__dlrtn_1_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_1
Xsky130_fd_sc_hdll__clkmux2_2_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_2_0/S sky130_fd_sc_hdll__clkmux2_2_0/A1
+ sky130_fd_sc_hdll__clkmux2_2_0/A0 sky130_fd_sc_hdll__clkmux2_2_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_2
Xsky130_fd_sc_hdll__or2_8_0 sky130_fd_sc_hdll__or2_8_0/X sky130_fd_sc_hdll__or2_8_0/A
+ sky130_fd_sc_hdll__or2_8_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_9 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21ai_2_0 sky130_fd_sc_hdll__o21ai_2_0/B1 sky130_fd_sc_hdll__o21ai_2_0/Y
+ sky130_fd_sc_hdll__o21ai_2_0/A2 sky130_fd_sc_hdll__o21ai_2_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21ai_2
Xsky130_fd_sc_hdll__and3_4_0 sky130_fd_sc_hdll__and3_4_0/A sky130_fd_sc_hdll__and3_4_0/B
+ sky130_fd_sc_hdll__and3_4_0/C sky130_fd_sc_hdll__and3_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__and3_4
Xsky130_fd_sc_hdll__clkbuf_4_0 sky130_fd_sc_hdll__clkbuf_4_0/X sky130_fd_sc_hdll__clkbuf_4_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkbuf_4
Xsky130_fd_sc_hdll__clkinv_4_0 sky130_fd_sc_hdll__clkinv_4_0/A sky130_fd_sc_hdll__clkinv_4_0/Y
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinv_4
Xsky130_fd_sc_hdll__sdfstp_4_0 sky130_fd_sc_hdll__sdfstp_4_0/CLK sky130_fd_sc_hdll__sdfstp_4_0/D
+ sky130_fd_sc_hdll__sdfstp_4_0/SCD sky130_fd_sc_hdll__sdfstp_4_0/Q sky130_fd_sc_hdll__sdfstp_4_0/SCE
+ sky130_fd_sc_hdll__sdfstp_4_0/SET_B VPWR VGND VPWR VGND sky130_fd_sc_hdll__sdfstp_4
Xsky130_fd_sc_hdll__a2bb2oi_1_0 sky130_fd_sc_hdll__a2bb2oi_1_0/A1_N sky130_fd_sc_hdll__a2bb2oi_1_0/Y
+ VGND VPWR sky130_fd_sc_hdll__a2bb2oi_1_0/B2 sky130_fd_sc_hdll__a2bb2oi_1_0/B1 sky130_fd_sc_hdll__a2bb2oi_1_0/A2_N
+ VPWR VGND sky130_fd_sc_hdll__a2bb2oi_1
Xsky130_fd_sc_hdll__nor4bb_2_0 sky130_fd_sc_hdll__nor4bb_2_0/D_N sky130_fd_sc_hdll__nor4bb_2_0/C_N
+ sky130_fd_sc_hdll__nor4bb_2_0/A sky130_fd_sc_hdll__nor4bb_2_0/Y sky130_fd_sc_hdll__nor4bb_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_306 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_317 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_2_0 sky130_fd_sc_hdll__isobufsrc_2_0/A sky130_fd_sc_hdll__isobufsrc_2_0/SLEEP
+ sky130_fd_sc_hdll__isobufsrc_2_0/X VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_2
Xsky130_fd_sc_hdll__sdfxbp_1_0 VGND VPWR sky130_fd_sc_hdll__sdfxbp_1_0/SCD sky130_fd_sc_hdll__sdfxbp_1_0/Q_N
+ sky130_fd_sc_hdll__sdfxbp_1_0/D sky130_fd_sc_hdll__sdfxbp_1_0/SCE sky130_fd_sc_hdll__sdfxbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfxbp_1_0/Q VGND VPWR sky130_fd_sc_hdll__sdfxbp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_103 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_114 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_125 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_136 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_147 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_158 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_169 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2b_1_0 sky130_fd_sc_hdll__nor2b_1_0/B_N sky130_fd_sc_hdll__nor2b_1_0/Y
+ sky130_fd_sc_hdll__nor2b_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2b_1
Xsky130_fd_sc_hdll__a21boi_4_0 sky130_fd_sc_hdll__a21boi_4_0/Y sky130_fd_sc_hdll__a21boi_4_0/A1
+ sky130_fd_sc_hdll__a21boi_4_0/B1_N sky130_fd_sc_hdll__a21boi_4_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__a21boi_4
Xsky130_fd_sc_hdll__nand3_4_0 sky130_fd_sc_hdll__nand3_4_0/Y sky130_fd_sc_hdll__nand3_4_0/A
+ sky130_fd_sc_hdll__nand3_4_0/B sky130_fd_sc_hdll__nand3_4_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3_4
Xsky130_fd_sc_hdll__mux2_4_0 sky130_fd_sc_hdll__mux2_4_0/X sky130_fd_sc_hdll__mux2_4_0/S
+ sky130_fd_sc_hdll__mux2_4_0/A0 sky130_fd_sc_hdll__mux2_4_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__mux2_4
Xsky130_fd_sc_hdll__and2b_4_0 sky130_fd_sc_hdll__and2b_4_0/B sky130_fd_sc_hdll__and2b_4_0/X
+ sky130_fd_sc_hdll__and2b_4_0/A_N VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2b_4
Xsky130_fd_sc_hdll__o22a_2_0 sky130_fd_sc_hdll__o22a_2_0/A2 sky130_fd_sc_hdll__o22a_2_0/X
+ sky130_fd_sc_hdll__o22a_2_0/B1 sky130_fd_sc_hdll__o22a_2_0/A1 sky130_fd_sc_hdll__o22a_2_0/B2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22a_2
Xsky130_fd_sc_hdll__a221oi_2_0 sky130_fd_sc_hdll__a221oi_2_0/B2 sky130_fd_sc_hdll__a221oi_2_0/C1
+ sky130_fd_sc_hdll__a221oi_2_0/A2 sky130_fd_sc_hdll__a221oi_2_0/A1 sky130_fd_sc_hdll__a221oi_2_0/B1
+ sky130_fd_sc_hdll__a221oi_2_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__a221oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_307 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_318 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfrtp_4_0 VPWR VGND sky130_fd_sc_hdll__sdfrtp_4_0/RESET_B VPWR
+ VGND sky130_fd_sc_hdll__sdfrtp_4_0/SCE sky130_fd_sc_hdll__sdfrtp_4_0/SCD sky130_fd_sc_hdll__sdfrtp_4_0/D
+ sky130_fd_sc_hdll__sdfrtp_4_0/CLK sky130_fd_sc_hdll__sdfrtp_4_0/Q sky130_fd_sc_hdll__sdfrtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_104 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_115 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_126 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_137 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_148 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_159 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and4b_1_0 VGND VPWR sky130_fd_sc_hdll__and4b_1_0/C sky130_fd_sc_hdll__and4b_1_0/A_N
+ sky130_fd_sc_hdll__and4b_1_0/X sky130_fd_sc_hdll__and4b_1_0/D sky130_fd_sc_hdll__and4b_1_0/B
+ VPWR VGND sky130_fd_sc_hdll__and4b_1
Xsky130_fd_sc_hdll__probe_p_8_0 sky130_fd_sc_hdll__probe_p_8_0/X sky130_fd_sc_hdll__probe_p_8_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__probe_p_8
Xsky130_fd_sc_hdll__o32ai_4_0 sky130_fd_sc_hdll__o32ai_4_0/A1 sky130_fd_sc_hdll__o32ai_4_0/A2
+ sky130_fd_sc_hdll__o32ai_4_0/A3 sky130_fd_sc_hdll__o32ai_4_0/B1 sky130_fd_sc_hdll__o32ai_4_0/Y
+ sky130_fd_sc_hdll__o32ai_4_0/B2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o32ai_4
Xsky130_fd_sc_hdll__nor3_2_0 sky130_fd_sc_hdll__nor3_2_0/C sky130_fd_sc_hdll__nor3_2_0/Y
+ sky130_fd_sc_hdll__nor3_2_0/A sky130_fd_sc_hdll__nor3_2_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_2
Xsky130_fd_sc_hdll__xor2_4_0 sky130_fd_sc_hdll__xor2_4_0/X sky130_fd_sc_hdll__xor2_4_0/B
+ sky130_fd_sc_hdll__xor2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__xor2_4
Xsky130_fd_sc_hdll__or3b_4_0 sky130_fd_sc_hdll__or3b_4_0/A sky130_fd_sc_hdll__or3b_4_0/B
+ sky130_fd_sc_hdll__or3b_4_0/C_N sky130_fd_sc_hdll__or3b_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__or3b_4
Xsky130_fd_sc_hdll__o21ba_4_0 sky130_fd_sc_hdll__o21ba_4_0/B1_N sky130_fd_sc_hdll__o21ba_4_0/A1
+ sky130_fd_sc_hdll__o21ba_4_0/A2 sky130_fd_sc_hdll__o21ba_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_4
Xsky130_fd_sc_hdll__a31o_1_0 sky130_fd_sc_hdll__a31o_1_0/A2 sky130_fd_sc_hdll__a31o_1_0/B1
+ sky130_fd_sc_hdll__a31o_1_0/A1 sky130_fd_sc_hdll__a31o_1_0/A3 sky130_fd_sc_hdll__a31o_1_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__a31o_1
Xsky130_fd_sc_hdll__xnor3_1_0 sky130_fd_sc_hdll__xnor3_1_0/X sky130_fd_sc_hdll__xnor3_1_0/B
+ sky130_fd_sc_hdll__xnor3_1_0/C sky130_fd_sc_hdll__xnor3_1_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_1
Xsky130_fd_sc_hdll__or4bb_4_0 sky130_fd_sc_hdll__or4bb_4_0/D_N sky130_fd_sc_hdll__or4bb_4_0/B
+ sky130_fd_sc_hdll__or4bb_4_0/A sky130_fd_sc_hdll__or4bb_4_0/C_N sky130_fd_sc_hdll__or4bb_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__or4bb_4
Xsky130_fd_sc_hdll__probec_p_8_0 sky130_fd_sc_hdll__probec_p_8_0/X sky130_fd_sc_hdll__probec_p_8_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__probec_p_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_308 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_319 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_105 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_116 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_127 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_138 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_149 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor3b_4_0 sky130_fd_sc_hdll__nor3b_4_0/A sky130_fd_sc_hdll__nor3b_4_0/C_N
+ sky130_fd_sc_hdll__nor3b_4_0/B sky130_fd_sc_hdll__nor3b_4_0/Y VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_4
Xsky130_fd_sc_hdll__o221ai_4_0 sky130_fd_sc_hdll__o221ai_4_0/B1 sky130_fd_sc_hdll__o221ai_4_0/B2
+ sky130_fd_sc_hdll__o221ai_4_0/A2 sky130_fd_sc_hdll__o221ai_4_0/C1 sky130_fd_sc_hdll__o221ai_4_0/Y
+ sky130_fd_sc_hdll__o221ai_4_0/A1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221ai_4
Xsky130_fd_sc_hdll__or2_6_0 sky130_fd_sc_hdll__or2_6_0/X sky130_fd_sc_hdll__or2_6_0/A
+ sky130_fd_sc_hdll__or2_6_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_6
Xsky130_fd_sc_hdll__o31ai_4_0 sky130_fd_sc_hdll__o31ai_4_0/A3 sky130_fd_sc_hdll__o31ai_4_0/A2
+ sky130_fd_sc_hdll__o31ai_4_0/A1 sky130_fd_sc_hdll__o31ai_4_0/Y sky130_fd_sc_hdll__o31ai_4_0/B1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o31ai_4
Xsky130_fd_sc_hdll__and3_2_0 sky130_fd_sc_hdll__and3_2_0/B sky130_fd_sc_hdll__and3_2_0/X
+ sky130_fd_sc_hdll__and3_2_0/A sky130_fd_sc_hdll__and3_2_0/C VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__and3_2
Xsky130_fd_sc_hdll__clkbuf_2_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__clkbuf_2_0/A
+ sky130_fd_sc_hdll__clkbuf_2_0/X sky130_fd_sc_hdll__clkbuf_2
Xsky130_fd_sc_hdll__clkinv_2_0 sky130_fd_sc_hdll__clkinv_2_0/Y sky130_fd_sc_hdll__clkinv_2_0/A
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinv_2
Xsky130_fd_sc_hdll__sdfstp_2_0 sky130_fd_sc_hdll__sdfstp_2_0/Q sky130_fd_sc_hdll__sdfstp_2_0/SCD
+ sky130_fd_sc_hdll__sdfstp_2_0/D sky130_fd_sc_hdll__sdfstp_2_0/CLK sky130_fd_sc_hdll__sdfstp_2_0/SET_B
+ sky130_fd_sc_hdll__sdfstp_2_0/SCE VGND VPWR VPWR VGND sky130_fd_sc_hdll__sdfstp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_309 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a211o_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_1_0/X sky130_fd_sc_hdll__a211o_1_0/A2
+ sky130_fd_sc_hdll__a211o_1_0/B1 sky130_fd_sc_hdll__a211o_1_0/A1 sky130_fd_sc_hdll__a211o_1_0/C1
+ sky130_fd_sc_hdll__a211o_1
Xsky130_fd_sc_hdll__nor2_8_0 sky130_fd_sc_hdll__nor2_8_0/Y sky130_fd_sc_hdll__nor2_8_0/A
+ sky130_fd_sc_hdll__nor2_8_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_8
Xsky130_fd_sc_hdll__a21o_1_0 sky130_fd_sc_hdll__a21o_1_0/A2 sky130_fd_sc_hdll__a21o_1_0/A1
+ sky130_fd_sc_hdll__a21o_1_0/B1 sky130_fd_sc_hdll__a21o_1_0/X VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__a21o_1
Xsky130_fd_sc_hdll__einvn_4_0 sky130_fd_sc_hdll__einvn_4_0/TE_B sky130_fd_sc_hdll__einvn_4_0/Z
+ sky130_fd_sc_hdll__einvn_4_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_106 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_117 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_128 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_139 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_16_0 sky130_fd_sc_hdll__nand2_16_0/Y sky130_fd_sc_hdll__nand2_16_0/A
+ sky130_fd_sc_hdll__nand2_16_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_16
Xsky130_fd_sc_hdll__buf_16_0 sky130_fd_sc_hdll__buf_16_0/A sky130_fd_sc_hdll__buf_16_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__buf_16
Xsky130_fd_sc_hdll__a21boi_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a21boi_2_0/B1_N
+ sky130_fd_sc_hdll__a21boi_2_0/A2 sky130_fd_sc_hdll__a21boi_2_0/A1 sky130_fd_sc_hdll__a21boi_2_0/Y
+ sky130_fd_sc_hdll__a21boi_2
Xsky130_fd_sc_hdll__nand3_2_0 sky130_fd_sc_hdll__nand3_2_0/A sky130_fd_sc_hdll__nand3_2_0/Y
+ sky130_fd_sc_hdll__nand3_2_0/B sky130_fd_sc_hdll__nand3_2_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3_2
Xsky130_fd_sc_hdll__fill_4_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_4
Xsky130_fd_sc_hdll__einvp_1_0 sky130_fd_sc_hdll__einvp_1_0/TE sky130_fd_sc_hdll__einvp_1_0/A
+ sky130_fd_sc_hdll__einvp_1_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_1
Xsky130_fd_sc_hdll__a32o_4_0 sky130_fd_sc_hdll__a32o_4_0/A3 sky130_fd_sc_hdll__a32o_4_0/X
+ sky130_fd_sc_hdll__a32o_4_0/B1 sky130_fd_sc_hdll__a32o_4_0/B2 sky130_fd_sc_hdll__a32o_4_0/A1
+ sky130_fd_sc_hdll__a32o_4_0/A2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32o_4
Xsky130_fd_sc_hdll__mux2_2_0 VGND VPWR sky130_fd_sc_hdll__mux2_2_0/A1 sky130_fd_sc_hdll__mux2_2_0/A0
+ sky130_fd_sc_hdll__mux2_2_0/S sky130_fd_sc_hdll__mux2_2_0/X VPWR VGND sky130_fd_sc_hdll__mux2_2
Xsky130_fd_sc_hdll__and2b_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__and2b_2_0/X sky130_fd_sc_hdll__and2b_2_0/B
+ sky130_fd_sc_hdll__and2b_2_0/A_N sky130_fd_sc_hdll__and2b_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_107 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_118 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_129 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfrtp_2_0 sky130_fd_sc_hdll__sdfrtp_2_0/RESET_B VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__sdfrtp_2_0/Q sky130_fd_sc_hdll__sdfrtp_2_0/SCE sky130_fd_sc_hdll__sdfrtp_2_0/SCD
+ sky130_fd_sc_hdll__sdfrtp_2_0/D sky130_fd_sc_hdll__sdfrtp_2_0/CLK sky130_fd_sc_hdll__sdfrtp_2
Xsky130_fd_sc_hdll__and2_8_0 sky130_fd_sc_hdll__and2_8_0/X sky130_fd_sc_hdll__and2_8_0/B
+ sky130_fd_sc_hdll__and2_8_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_8
Xsky130_fd_sc_hdll__a22oi_4_0 sky130_fd_sc_hdll__a22oi_4_0/A2 sky130_fd_sc_hdll__a22oi_4_0/B2
+ sky130_fd_sc_hdll__a22oi_4_0/A1 sky130_fd_sc_hdll__a22oi_4_0/B1 sky130_fd_sc_hdll__a22oi_4_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a22oi_4
Xsky130_fd_sc_hdll__muxb4to1_4_0 VPWR VGND VGND VPWR sky130_fd_sc_hdll__muxb4to1_4_0/Z
+ sky130_fd_sc_hdll__muxb4to1_4_0/S[0] sky130_fd_sc_hdll__muxb4to1_4_0/S[1] sky130_fd_sc_hdll__muxb4to1_4_0/D[1]
+ sky130_fd_sc_hdll__muxb4to1_4_0/D[2] sky130_fd_sc_hdll__muxb4to1_4_0/S[2] sky130_fd_sc_hdll__muxb4to1_4_0/S[3]
+ sky130_fd_sc_hdll__muxb4to1_4_0/D[3] sky130_fd_sc_hdll__muxb4to1_4_0/D[0] sky130_fd_sc_hdll__muxb4to1_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_290 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o32ai_2_0 sky130_fd_sc_hdll__o32ai_2_0/A1 sky130_fd_sc_hdll__o32ai_2_0/B1
+ sky130_fd_sc_hdll__o32ai_2_0/A2 sky130_fd_sc_hdll__o32ai_2_0/A3 sky130_fd_sc_hdll__o32ai_2_0/Y
+ sky130_fd_sc_hdll__o32ai_2_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o32ai_2
Xsky130_fd_sc_hdll__o221a_4_0 sky130_fd_sc_hdll__o221a_4_0/C1 sky130_fd_sc_hdll__o221a_4_0/A1
+ sky130_fd_sc_hdll__o221a_4_0/A2 sky130_fd_sc_hdll__o221a_4_0/B1 sky130_fd_sc_hdll__o221a_4_0/B2
+ sky130_fd_sc_hdll__o221a_4_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221a_4
Xsky130_fd_sc_hdll__or3b_2_0 sky130_fd_sc_hdll__or3b_2_0/A sky130_fd_sc_hdll__or3b_2_0/B
+ sky130_fd_sc_hdll__or3b_2_0/C_N sky130_fd_sc_hdll__or3b_2_0/X VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__or3b_2
Xsky130_fd_sc_hdll__xor2_2_0 sky130_fd_sc_hdll__xor2_2_0/B VPWR VGND sky130_fd_sc_hdll__xor2_2_0/X
+ sky130_fd_sc_hdll__xor2_2_0/A VPWR VGND sky130_fd_sc_hdll__xor2_2
Xsky130_fd_sc_hdll__o21ba_2_0 sky130_fd_sc_hdll__o21ba_2_0/B1_N sky130_fd_sc_hdll__o21ba_2_0/A1
+ sky130_fd_sc_hdll__o21ba_2_0/X sky130_fd_sc_hdll__o21ba_2_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_2
Xsky130_fd_sc_hdll__or4bb_2_0 sky130_fd_sc_hdll__or4bb_2_0/A sky130_fd_sc_hdll__or4bb_2_0/X
+ sky130_fd_sc_hdll__or4bb_2_0/B sky130_fd_sc_hdll__or4bb_2_0/D_N sky130_fd_sc_hdll__or4bb_2_0/C_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4bb_2
Xsky130_fd_sc_hdll__dlxtn_4_0 sky130_fd_sc_hdll__dlxtn_4_0/D sky130_fd_sc_hdll__dlxtn_4_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_4_0/Q VGND VPWR VPWR VGND sky130_fd_sc_hdll__dlxtn_4
Xsky130_fd_sc_hdll__nand2_8_0 sky130_fd_sc_hdll__nand2_8_0/A sky130_fd_sc_hdll__nand2_8_0/B
+ sky130_fd_sc_hdll__nand2_8_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_108 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_119 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21bai_4_0 sky130_fd_sc_hdll__o21bai_4_0/Y sky130_fd_sc_hdll__o21bai_4_0/B1_N
+ sky130_fd_sc_hdll__o21bai_4_0/A1 sky130_fd_sc_hdll__o21bai_4_0/A2 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__o21bai_4
Xsky130_fd_sc_hdll__a22o_4_0 sky130_fd_sc_hdll__a22o_4_0/B1 sky130_fd_sc_hdll__a22o_4_0/B2
+ sky130_fd_sc_hdll__a22o_4_0/X sky130_fd_sc_hdll__a22o_4_0/A2 sky130_fd_sc_hdll__a22o_4_0/A1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a22o_4
Xsky130_fd_sc_hdll__dlygate4sd2_1_0 sky130_fd_sc_hdll__dlygate4sd2_1_0/A sky130_fd_sc_hdll__dlygate4sd2_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd2_1
Xsky130_fd_sc_hdll__nand4bb_1_0 sky130_fd_sc_hdll__nand4bb_1_0/C sky130_fd_sc_hdll__nand4bb_1_0/D
+ sky130_fd_sc_hdll__nand4bb_1_0/A_N sky130_fd_sc_hdll__nand4bb_1_0/Y sky130_fd_sc_hdll__nand4bb_1_0/B_N
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__nand4bb_1
Xsky130_fd_sc_hdll__clkbuf_12_0 sky130_fd_sc_hdll__clkbuf_12_0/A sky130_fd_sc_hdll__clkbuf_12_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_12
Xsky130_fd_sc_hdll__nor3b_2_0 sky130_fd_sc_hdll__nor3b_2_0/C_N sky130_fd_sc_hdll__nor3b_2_0/Y
+ sky130_fd_sc_hdll__nor3b_2_0/A sky130_fd_sc_hdll__nor3b_2_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_2
Xsky130_fd_sc_hdll__muxb16to1_1_0 sky130_fd_sc_hdll__muxb16to1_1_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_1_0/D[0] sky130_fd_sc_hdll__muxb16to1_1_0/S[12]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[13] sky130_fd_sc_hdll__muxb16to1_1_0/S[8] sky130_fd_sc_hdll__muxb16to1_1_0/S[9]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[10] sky130_fd_sc_hdll__muxb16to1_1_0/S[11] sky130_fd_sc_hdll__muxb16to1_1_0/S[14]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[12] sky130_fd_sc_hdll__muxb16to1_1_0/D[9]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[10] sky130_fd_sc_hdll__muxb16to1_1_0/D[13] sky130_fd_sc_hdll__muxb16to1_1_0/D[14]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[8] sky130_fd_sc_hdll__muxb16to1_1_0/D[11]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[0] sky130_fd_sc_hdll__muxb16to1_1_0/S[1] sky130_fd_sc_hdll__muxb16to1_1_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[2] sky130_fd_sc_hdll__muxb16to1_1_0/S[2] sky130_fd_sc_hdll__muxb16to1_1_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[4] sky130_fd_sc_hdll__muxb16to1_1_0/S[4] sky130_fd_sc_hdll__muxb16to1_1_0/S[5]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[5] sky130_fd_sc_hdll__muxb16to1_1_0/D[6] sky130_fd_sc_hdll__muxb16to1_1_0/S[6]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[7] sky130_fd_sc_hdll__muxb16to1_1_0/D[7] sky130_fd_sc_hdll__muxb16to1_1_0/D[3]
+ sky130_fd_sc_hdll__muxb16to1_1
Xsky130_fd_sc_hdll__o221ai_2_0 sky130_fd_sc_hdll__o221ai_2_0/B1 sky130_fd_sc_hdll__o221ai_2_0/B2
+ sky130_fd_sc_hdll__o221ai_2_0/Y sky130_fd_sc_hdll__o221ai_2_0/A2 sky130_fd_sc_hdll__o221ai_2_0/A1
+ sky130_fd_sc_hdll__o221ai_2_0/C1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__o221ai_2
Xsky130_fd_sc_hdll__ebufn_1_0 sky130_fd_sc_hdll__ebufn_1_0/Z sky130_fd_sc_hdll__ebufn_1_0/TE_B
+ sky130_fd_sc_hdll__ebufn_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__ebufn_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_291 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_280 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2_4_0 sky130_fd_sc_hdll__or2_4_0/X sky130_fd_sc_hdll__or2_4_0/A
+ sky130_fd_sc_hdll__or2_4_0/B VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2_4
Xsky130_fd_sc_hdll__a21oi_4_0 sky130_fd_sc_hdll__a21oi_4_0/B1 sky130_fd_sc_hdll__a21oi_4_0/A2
+ sky130_fd_sc_hdll__a21oi_4_0/A1 sky130_fd_sc_hdll__a21oi_4_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21oi_4
Xsky130_fd_sc_hdll__o31ai_2_0 sky130_fd_sc_hdll__o31ai_2_0/A1 sky130_fd_sc_hdll__o31ai_2_0/Y
+ sky130_fd_sc_hdll__o31ai_2_0/B1 sky130_fd_sc_hdll__o31ai_2_0/A3 sky130_fd_sc_hdll__o31ai_2_0/A2
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o31ai_2
Xsky130_fd_sc_hdll__o211a_4_0 sky130_fd_sc_hdll__o211a_4_0/A1 sky130_fd_sc_hdll__o211a_4_0/X
+ sky130_fd_sc_hdll__o211a_4_0/C1 sky130_fd_sc_hdll__o211a_4_0/A2 sky130_fd_sc_hdll__o211a_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211a_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_109 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__einvn_2_0 sky130_fd_sc_hdll__einvn_2_0/TE_B sky130_fd_sc_hdll__einvn_2_0/A
+ sky130_fd_sc_hdll__einvn_2_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvn_2
Xsky130_fd_sc_hdll__sdfsbp_1_0 sky130_fd_sc_hdll__sdfsbp_1_0/SCD sky130_fd_sc_hdll__sdfsbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfsbp_1_0/Q_N sky130_fd_sc_hdll__sdfsbp_1_0/D sky130_fd_sc_hdll__sdfsbp_1_0/Q
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_1_0/SET_B sky130_fd_sc_hdll__sdfsbp_1_0/SCE
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_1
Xsky130_fd_sc_hdll__or4_1_0 sky130_fd_sc_hdll__or4_1_0/C sky130_fd_sc_hdll__or4_1_0/A
+ sky130_fd_sc_hdll__or4_1_0/X sky130_fd_sc_hdll__or4_1_0/B sky130_fd_sc_hdll__or4_1_0/D
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_292 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_281 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_270 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inputiso0n_1_0 VPWR VGND sky130_fd_sc_hdll__inputiso0n_1_0/X sky130_fd_sc_hdll__inputiso0n_1_0/SLEEP_B
+ sky130_fd_sc_hdll__inputiso0n_1_0/A VPWR VGND sky130_fd_sc_hdll__inputiso0n_1
Xsky130_fd_sc_hdll__fill_2_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_2
Xsky130_fd_sc_hdll__and4bb_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_1_0/A_N
+ sky130_fd_sc_hdll__and4bb_1_0/D sky130_fd_sc_hdll__and4bb_1_0/X sky130_fd_sc_hdll__and4bb_1_0/C
+ sky130_fd_sc_hdll__and4bb_1_0/B_N sky130_fd_sc_hdll__and4bb_1
Xsky130_fd_sc_hdll__clkinvlp_4_0 sky130_fd_sc_hdll__clkinvlp_4_0/A sky130_fd_sc_hdll__clkinvlp_4_0/Y
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__clkinvlp_4
Xsky130_fd_sc_hdll__a32o_2_0 sky130_fd_sc_hdll__a32o_2_0/B2 sky130_fd_sc_hdll__a32o_2_0/X
+ sky130_fd_sc_hdll__a32o_2_0/A2 sky130_fd_sc_hdll__a32o_2_0/A3 sky130_fd_sc_hdll__a32o_2_0/A1
+ sky130_fd_sc_hdll__a32o_2_0/B1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32o_2
Xsky130_fd_sc_hdll__nand3b_1_0 sky130_fd_sc_hdll__nand3b_1_0/B sky130_fd_sc_hdll__nand3b_1_0/C
+ sky130_fd_sc_hdll__nand3b_1_0/A_N sky130_fd_sc_hdll__nand3b_1_0/Y VPWR VGND VGND
+ VPWR sky130_fd_sc_hdll__nand3b_1
Xsky130_fd_sc_hdll__and2_6_0 sky130_fd_sc_hdll__and2_6_0/X sky130_fd_sc_hdll__and2_6_0/B
+ sky130_fd_sc_hdll__and2_6_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_6
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_293 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_282 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_271 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_260 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a22oi_2_0 sky130_fd_sc_hdll__a22oi_2_0/A1 sky130_fd_sc_hdll__a22oi_2_0/A2
+ sky130_fd_sc_hdll__a22oi_2_0/B1 sky130_fd_sc_hdll__a22oi_2_0/B2 sky130_fd_sc_hdll__a22oi_2_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22oi_2
Xsky130_fd_sc_hdll__muxb4to1_2_0 VGND VPWR sky130_fd_sc_hdll__muxb4to1_2_0/Z VGND
+ VPWR sky130_fd_sc_hdll__muxb4to1_2_0/S[1] sky130_fd_sc_hdll__muxb4to1_2_0/S[2] sky130_fd_sc_hdll__muxb4to1_2_0/S[3]
+ sky130_fd_sc_hdll__muxb4to1_2_0/D[1] sky130_fd_sc_hdll__muxb4to1_2_0/D[0] sky130_fd_sc_hdll__muxb4to1_2_0/D[2]
+ sky130_fd_sc_hdll__muxb4to1_2_0/D[3] sky130_fd_sc_hdll__muxb4to1_2_0/S[0] sky130_fd_sc_hdll__muxb4to1_2
Xsky130_fd_sc_hdll__sdfrbp_1_0 sky130_fd_sc_hdll__sdfrbp_1_0/RESET_B VPWR VGND VGND
+ VPWR sky130_fd_sc_hdll__sdfrbp_1_0/Q_N sky130_fd_sc_hdll__sdfrbp_1_0/D sky130_fd_sc_hdll__sdfrbp_1_0/CLK
+ sky130_fd_sc_hdll__sdfrbp_1_0/Q sky130_fd_sc_hdll__sdfrbp_1_0/SCE sky130_fd_sc_hdll__sdfrbp_1_0/SCD
+ sky130_fd_sc_hdll__sdfrbp_1
Xsky130_fd_sc_hdll__o221a_2_0 sky130_fd_sc_hdll__o221a_2_0/B2 sky130_fd_sc_hdll__o221a_2_0/A2
+ sky130_fd_sc_hdll__o221a_2_0/X sky130_fd_sc_hdll__o221a_2_0/B1 sky130_fd_sc_hdll__o221a_2_0/C1
+ sky130_fd_sc_hdll__o221a_2_0/A1 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221a_2
Xsky130_fd_sc_hdll__dlxtn_2_0 sky130_fd_sc_hdll__dlxtn_2_0/D sky130_fd_sc_hdll__dlxtn_2_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_2_0/Q VGND VPWR VPWR VGND sky130_fd_sc_hdll__dlxtn_2
Xsky130_fd_sc_hdll__a22o_2_0 sky130_fd_sc_hdll__a22o_2_0/A1 sky130_fd_sc_hdll__a22o_2_0/A2
+ sky130_fd_sc_hdll__a22o_2_0/X sky130_fd_sc_hdll__a22o_2_0/B2 sky130_fd_sc_hdll__a22o_2_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22o_2
Xsky130_fd_sc_hdll__nand2_6_0 sky130_fd_sc_hdll__nand2_6_0/Y sky130_fd_sc_hdll__nand2_6_0/A
+ sky130_fd_sc_hdll__nand2_6_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_6
Xsky130_fd_sc_hdll__o21bai_2_0 sky130_fd_sc_hdll__o21bai_2_0/B1_N sky130_fd_sc_hdll__o21bai_2_0/Y
+ sky130_fd_sc_hdll__o21bai_2_0/A2 sky130_fd_sc_hdll__o21bai_2_0/A1 VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__o21bai_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_294 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_283 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_272 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_261 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_250 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21a_4_0 sky130_fd_sc_hdll__o21a_4_0/A1 sky130_fd_sc_hdll__o21a_4_0/A2
+ sky130_fd_sc_hdll__o21a_4_0/B1 sky130_fd_sc_hdll__o21a_4_0/X VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21a_4
Xsky130_fd_sc_hdll__a21oi_2_0 sky130_fd_sc_hdll__a21oi_2_0/B1 sky130_fd_sc_hdll__a21oi_2_0/A2
+ sky130_fd_sc_hdll__a21oi_2_0/A1 sky130_fd_sc_hdll__a21oi_2_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21oi_2
Xsky130_fd_sc_hdll__or2_2_0 sky130_fd_sc_hdll__or2_2_0/B sky130_fd_sc_hdll__or2_2_0/X
+ sky130_fd_sc_hdll__or2_2_0/A VPWR VGND VPWR VGND sky130_fd_sc_hdll__or2_2
Xsky130_fd_sc_hdll__decap_12_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__decap_12
Xsky130_fd_sc_hdll__o211a_2_0 sky130_fd_sc_hdll__o211a_2_0/C1 sky130_fd_sc_hdll__o211a_2_0/B1
+ sky130_fd_sc_hdll__o211a_2_0/A2 sky130_fd_sc_hdll__o211a_2_0/A1 sky130_fd_sc_hdll__o211a_2_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o211a_2
Xsky130_fd_sc_hdll__tapvgnd_1_0 VPWR VGND VPWR sky130_fd_sc_hdll__tapvgnd_1
Xsky130_fd_sc_hdll__nor2_4_0 sky130_fd_sc_hdll__nor2_4_0/Y sky130_fd_sc_hdll__nor2_4_0/A
+ sky130_fd_sc_hdll__nor2_4_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_4
Xsky130_fd_sc_hdll__inputiso1p_1_0 sky130_fd_sc_hdll__inputiso1p_1_0/SLEEP sky130_fd_sc_hdll__inputiso1p_1_0/X
+ sky130_fd_sc_hdll__inputiso1p_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__inputiso1p_1
Xsky130_fd_sc_hdll__dfstp_1_0 sky130_fd_sc_hdll__dfstp_1_0/D VPWR sky130_fd_sc_hdll__dfstp_1_0/CLK
+ VGND sky130_fd_sc_hdll__dfstp_1_0/Q VPWR VGND sky130_fd_sc_hdll__dfstp_1_0/SET_B
+ sky130_fd_sc_hdll__dfstp_1
Xsky130_fd_sc_hdll__nand4b_4_0 sky130_fd_sc_hdll__nand4b_4_0/C sky130_fd_sc_hdll__nand4b_4_0/D
+ sky130_fd_sc_hdll__nand4b_4_0/B sky130_fd_sc_hdll__nand4b_4_0/Y sky130_fd_sc_hdll__nand4b_4_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_295 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_284 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_273 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_262 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_251 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_240 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_12_0 sky130_fd_sc_hdll__nand2_12_0/Y sky130_fd_sc_hdll__nand2_12_0/A
+ sky130_fd_sc_hdll__nand2_12_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_12
Xsky130_fd_sc_hdll__buf_12_0 sky130_fd_sc_hdll__buf_12_0/A sky130_fd_sc_hdll__buf_12_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__buf_12
Xsky130_fd_sc_hdll__a21o_8_0 sky130_fd_sc_hdll__a21o_8_0/A2 sky130_fd_sc_hdll__a21o_8_0/A1
+ sky130_fd_sc_hdll__a21o_8_0/X sky130_fd_sc_hdll__a21o_8_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_8
Xsky130_fd_sc_hdll__sdfrtn_1_0 VPWR VGND sky130_fd_sc_hdll__sdfrtn_1_0/RESET_B VPWR
+ VGND sky130_fd_sc_hdll__sdfrtn_1_0/SCE sky130_fd_sc_hdll__sdfrtn_1_0/SCD sky130_fd_sc_hdll__sdfrtn_1_0/D
+ sky130_fd_sc_hdll__sdfrtn_1_0/CLK_N sky130_fd_sc_hdll__sdfrtn_1_0/Q sky130_fd_sc_hdll__sdfrtn_1
Xsky130_fd_sc_hdll__o2bb2ai_4_0 sky130_fd_sc_hdll__o2bb2ai_4_0/A1_N sky130_fd_sc_hdll__o2bb2ai_4_0/B1
+ sky130_fd_sc_hdll__o2bb2ai_4_0/B2 sky130_fd_sc_hdll__o2bb2ai_4_0/A2_N sky130_fd_sc_hdll__o2bb2ai_4_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o2bb2ai_4
Xsky130_fd_sc_hdll__nor4_1_0 sky130_fd_sc_hdll__nor4_1_0/D sky130_fd_sc_hdll__nor4_1_0/C
+ sky130_fd_sc_hdll__nor4_1_0/Y sky130_fd_sc_hdll__nor4_1_0/A sky130_fd_sc_hdll__nor4_1_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_1
Xsky130_fd_sc_hdll__clkinvlp_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinvlp_2_0/Y
+ sky130_fd_sc_hdll__clkinvlp_2_0/A sky130_fd_sc_hdll__clkinvlp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_263 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_252 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_241 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_230 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__einvp_8_0 sky130_fd_sc_hdll__einvp_8_0/A sky130_fd_sc_hdll__einvp_8_0/Z
+ sky130_fd_sc_hdll__einvp_8_0/TE VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_296 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_285 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and2_4_0 sky130_fd_sc_hdll__and2_4_0/X sky130_fd_sc_hdll__and2_4_0/B
+ sky130_fd_sc_hdll__and2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__and2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_274 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_1_0 sky130_fd_sc_hdll__dfrtp_1_0/RESET_B VGND VPWR sky130_fd_sc_hdll__dfrtp_1_0/Q
+ sky130_fd_sc_hdll__dfrtp_1_0/D sky130_fd_sc_hdll__dfrtp_1_0/CLK VPWR VGND sky130_fd_sc_hdll__dfrtp_1
Xsky130_fd_sc_hdll__sdlclkp_1_0 sky130_fd_sc_hdll__sdlclkp_1_0/CLK VGND VPWR sky130_fd_sc_hdll__sdlclkp_1_0/SCE
+ sky130_fd_sc_hdll__sdlclkp_1_0/GCLK sky130_fd_sc_hdll__sdlclkp_1_0/GATE VPWR VGND
+ sky130_fd_sc_hdll__sdlclkp_1
Xsky130_fd_sc_hdll__a32oi_4_0 sky130_fd_sc_hdll__a32oi_4_0/A3 sky130_fd_sc_hdll__a32oi_4_0/A2
+ sky130_fd_sc_hdll__a32oi_4_0/A1 sky130_fd_sc_hdll__a32oi_4_0/B1 sky130_fd_sc_hdll__a32oi_4_0/Y
+ sky130_fd_sc_hdll__a32oi_4_0/B2 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32oi_4
Xsky130_fd_sc_hdll__and4_1_0 sky130_fd_sc_hdll__and4_1_0/X sky130_fd_sc_hdll__and4_1_0/C
+ sky130_fd_sc_hdll__and4_1_0/A sky130_fd_sc_hdll__and4_1_0/B sky130_fd_sc_hdll__and4_1_0/D
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__and4_1
Xsky130_fd_sc_hdll__nand2_4_0 sky130_fd_sc_hdll__nand2_4_0/Y sky130_fd_sc_hdll__nand2_4_0/A
+ sky130_fd_sc_hdll__nand2_4_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_297 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_286 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_275 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_264 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_253 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_242 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_231 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_220 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21bo_4_0 sky130_fd_sc_hdll__a21bo_4_0/B1_N sky130_fd_sc_hdll__a21bo_4_0/A2
+ sky130_fd_sc_hdll__a21bo_4_0/A1 sky130_fd_sc_hdll__a21bo_4_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21bo_4
Xsky130_fd_sc_hdll__o21a_2_0 sky130_fd_sc_hdll__o21a_2_0/A1 sky130_fd_sc_hdll__o21a_2_0/B1
+ sky130_fd_sc_hdll__o21a_2_0/A2 sky130_fd_sc_hdll__o21a_2_0/X VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21a_2
Xsky130_fd_sc_hdll__a31oi_4_0 sky130_fd_sc_hdll__a31oi_4_0/Y sky130_fd_sc_hdll__a31oi_4_0/B1
+ sky130_fd_sc_hdll__a31oi_4_0/A2 sky130_fd_sc_hdll__a31oi_4_0/A3 sky130_fd_sc_hdll__a31oi_4_0/A1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__a31oi_4
Xsky130_fd_sc_hdll__mux2i_4_0 sky130_fd_sc_hdll__mux2i_4_0/S sky130_fd_sc_hdll__mux2i_4_0/A1
+ sky130_fd_sc_hdll__mux2i_4_0/A0 sky130_fd_sc_hdll__mux2i_4_0/Y VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__mux2i_4
Xsky130_fd_sc_hdll__nand4_1_0 sky130_fd_sc_hdll__nand4_1_0/C sky130_fd_sc_hdll__nand4_1_0/B
+ sky130_fd_sc_hdll__nand4_1_0/Y sky130_fd_sc_hdll__nand4_1_0/D sky130_fd_sc_hdll__nand4_1_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__nand4_1
Xsky130_fd_sc_hdll__and3b_1_0 sky130_fd_sc_hdll__and3b_1_0/A_N sky130_fd_sc_hdll__and3b_1_0/B
+ sky130_fd_sc_hdll__and3b_1_0/X sky130_fd_sc_hdll__and3b_1_0/C VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__and3b_1
Xsky130_fd_sc_hdll__ebufn_8_0 sky130_fd_sc_hdll__ebufn_8_0/A sky130_fd_sc_hdll__ebufn_8_0/Z
+ sky130_fd_sc_hdll__ebufn_8_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_8
Xsky130_fd_sc_hdll__nor2_2_0 sky130_fd_sc_hdll__nor2_2_0/B sky130_fd_sc_hdll__nor2_2_0/Y
+ sky130_fd_sc_hdll__nor2_2_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_298 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlrtn_4_0 sky130_fd_sc_hdll__dlrtn_4_0/RESET_B sky130_fd_sc_hdll__dlrtn_4_0/D
+ sky130_fd_sc_hdll__dlrtn_4_0/GATE_N sky130_fd_sc_hdll__dlrtn_4_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_287 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_276 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_265 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_254 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_243 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_232 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_221 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_210 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4b_2_0 sky130_fd_sc_hdll__nand4b_2_0/D sky130_fd_sc_hdll__nand4b_2_0/C
+ sky130_fd_sc_hdll__nand4b_2_0/B sky130_fd_sc_hdll__nand4b_2_0/Y sky130_fd_sc_hdll__nand4b_2_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4b_2
Xsky130_fd_sc_hdll__or2b_4_0 sky130_fd_sc_hdll__or2b_4_0/A sky130_fd_sc_hdll__or2b_4_0/B_N
+ sky130_fd_sc_hdll__or2b_4_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__or2b_4
Xsky130_fd_sc_hdll__xnor2_1_0 VGND VPWR sky130_fd_sc_hdll__xnor2_1_0/B sky130_fd_sc_hdll__xnor2_1_0/Y
+ sky130_fd_sc_hdll__xnor2_1_0/A VPWR VGND sky130_fd_sc_hdll__xnor2_1
Xsky130_fd_sc_hdll__a21o_6_0 sky130_fd_sc_hdll__a21o_6_0/A2 sky130_fd_sc_hdll__a21o_6_0/A1
+ sky130_fd_sc_hdll__a21o_6_0/X sky130_fd_sc_hdll__a21o_6_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_6
Xsky130_fd_sc_hdll__a2bb2oi_4_0 sky130_fd_sc_hdll__a2bb2oi_4_0/Y sky130_fd_sc_hdll__a2bb2oi_4_0/A2_N
+ sky130_fd_sc_hdll__a2bb2oi_4_0/B2 sky130_fd_sc_hdll__a2bb2oi_4_0/A1_N sky130_fd_sc_hdll__a2bb2oi_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2oi_4
Xsky130_fd_sc_hdll__bufinv_16_0 sky130_fd_sc_hdll__bufinv_16_0/A sky130_fd_sc_hdll__bufinv_16_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufinv_16
Xsky130_fd_sc_hdll__or4b_1_0 sky130_fd_sc_hdll__or4b_1_0/B sky130_fd_sc_hdll__or4b_1_0/D_N
+ sky130_fd_sc_hdll__or4b_1_0/A sky130_fd_sc_hdll__or4b_1_0/X sky130_fd_sc_hdll__or4b_1_0/C
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4b_1
Xsky130_fd_sc_hdll__o2bb2ai_2_0 sky130_fd_sc_hdll__o2bb2ai_2_0/B2 sky130_fd_sc_hdll__o2bb2ai_2_0/Y
+ sky130_fd_sc_hdll__o2bb2ai_2_0/A1_N sky130_fd_sc_hdll__o2bb2ai_2_0/A2_N sky130_fd_sc_hdll__o2bb2ai_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2ai_2
Xsky130_fd_sc_hdll__a2bb2o_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_1_0/B1
+ sky130_fd_sc_hdll__a2bb2o_1_0/A1_N sky130_fd_sc_hdll__a2bb2o_1_0/A2_N sky130_fd_sc_hdll__a2bb2o_1_0/X
+ sky130_fd_sc_hdll__a2bb2o_1_0/B2 sky130_fd_sc_hdll__a2bb2o_1
Xsky130_fd_sc_hdll__xor3_1_0 sky130_fd_sc_hdll__xor3_1_0/X sky130_fd_sc_hdll__xor3_1_0/C
+ sky130_fd_sc_hdll__xor3_1_0/B sky130_fd_sc_hdll__xor3_1_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_1
Xsky130_fd_sc_hdll__dlrtp_1_0 sky130_fd_sc_hdll__dlrtp_1_0/RESET_B sky130_fd_sc_hdll__dlrtp_1_0/D
+ sky130_fd_sc_hdll__dlrtp_1_0/GATE sky130_fd_sc_hdll__dlrtp_1_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_1
Xsky130_fd_sc_hdll__nor2b_4_0 sky130_fd_sc_hdll__nor2b_4_0/B_N sky130_fd_sc_hdll__nor2b_4_0/Y
+ sky130_fd_sc_hdll__nor2b_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor2b_4
Xsky130_fd_sc_hdll__buf_1_0 VGND VPWR sky130_fd_sc_hdll__buf_1_0/X sky130_fd_sc_hdll__buf_1_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_299 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_288 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_277 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_255 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_244 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_233 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_266 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_222 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inv_1_0 sky130_fd_sc_hdll__inv_1_0/Y sky130_fd_sc_hdll__inv_1_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__inv_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_211 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_200 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and2_2_0 VPWR VGND sky130_fd_sc_hdll__and2_2_0/A sky130_fd_sc_hdll__and2_2_0/X
+ sky130_fd_sc_hdll__and2_2_0/B VPWR VGND sky130_fd_sc_hdll__and2_2
Xsky130_fd_sc_hdll__nor4b_1_0 sky130_fd_sc_hdll__nor4b_1_0/C sky130_fd_sc_hdll__nor4b_1_0/B
+ sky130_fd_sc_hdll__nor4b_1_0/A sky130_fd_sc_hdll__nor4b_1_0/D_N sky130_fd_sc_hdll__nor4b_1_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4b_1
Xsky130_fd_sc_hdll__a211oi_1_0 sky130_fd_sc_hdll__a211oi_1_0/A1 sky130_fd_sc_hdll__a211oi_1_0/C1
+ sky130_fd_sc_hdll__a211oi_1_0/B1 sky130_fd_sc_hdll__a211oi_1_0/Y sky130_fd_sc_hdll__a211oi_1_0/A2
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a211oi_1
Xsky130_fd_sc_hdll__sedfxbp_2_0 VPWR VGND sky130_fd_sc_hdll__sedfxbp_2_0/CLK sky130_fd_sc_hdll__sedfxbp_2_0/Q_N
+ sky130_fd_sc_hdll__sedfxbp_2_0/SCD sky130_fd_sc_hdll__sedfxbp_2_0/DE sky130_fd_sc_hdll__sedfxbp_2_0/D
+ sky130_fd_sc_hdll__sedfxbp_2_0/Q sky130_fd_sc_hdll__sedfxbp_2_0/SCE VPWR VGND sky130_fd_sc_hdll__sedfxbp_2
Xsky130_fd_sc_hdll__a32oi_2_0 sky130_fd_sc_hdll__a32oi_2_0/A2 sky130_fd_sc_hdll__a32oi_2_0/B2
+ sky130_fd_sc_hdll__a32oi_2_0/A3 sky130_fd_sc_hdll__a32oi_2_0/A1 sky130_fd_sc_hdll__a32oi_2_0/Y
+ sky130_fd_sc_hdll__a32oi_2_0/B1 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a32oi_2
Xsky130_fd_sc_hdll__and4b_4_0 sky130_fd_sc_hdll__and4b_4_0/X sky130_fd_sc_hdll__and4b_4_0/D
+ sky130_fd_sc_hdll__and4b_4_0/C sky130_fd_sc_hdll__and4b_4_0/B sky130_fd_sc_hdll__and4b_4_0/A_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_289 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_278 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_267 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_256 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_245 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_234 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_223 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_212 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_201 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand2_2_0 sky130_fd_sc_hdll__nand2_2_0/Y sky130_fd_sc_hdll__nand2_2_0/A
+ sky130_fd_sc_hdll__nand2_2_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2_2
Xsky130_fd_sc_hdll__a31o_4_0 sky130_fd_sc_hdll__a31o_4_0/B1 sky130_fd_sc_hdll__a31o_4_0/A2
+ sky130_fd_sc_hdll__a31o_4_0/A3 sky130_fd_sc_hdll__a31o_4_0/A1 sky130_fd_sc_hdll__a31o_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a31o_4
Xsky130_fd_sc_hdll__xnor3_4_0 sky130_fd_sc_hdll__xnor3_4_0/X sky130_fd_sc_hdll__xnor3_4_0/B
+ sky130_fd_sc_hdll__xnor3_4_0/C sky130_fd_sc_hdll__xnor3_4_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_4
Xsky130_fd_sc_hdll__a21bo_2_0 sky130_fd_sc_hdll__a21bo_2_0/B1_N sky130_fd_sc_hdll__a21bo_2_0/A2
+ sky130_fd_sc_hdll__a21bo_2_0/X sky130_fd_sc_hdll__a21bo_2_0/A1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21bo_2
Xsky130_fd_sc_hdll__mux2i_2_0 sky130_fd_sc_hdll__mux2i_2_0/Y sky130_fd_sc_hdll__mux2i_2_0/A1
+ sky130_fd_sc_hdll__mux2i_2_0/A0 sky130_fd_sc_hdll__mux2i_2_0/S VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__mux2i_2
Xsky130_fd_sc_hdll__decap_3_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_3
Xsky130_fd_sc_hdll__a31oi_2_0 sky130_fd_sc_hdll__a31oi_2_0/A3 sky130_fd_sc_hdll__a31oi_2_0/B1
+ sky130_fd_sc_hdll__a31oi_2_0/Y sky130_fd_sc_hdll__a31oi_2_0/A1 sky130_fd_sc_hdll__a31oi_2_0/A2
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__a31oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_279 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_268 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_257 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_246 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_235 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_224 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_213 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_202 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__conb_1_0 sky130_fd_sc_hdll__conb_1_0/LO sky130_fd_sc_hdll__conb_1_0/HI
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__conb_1
Xsky130_fd_sc_hdll__dlrtn_2_0 sky130_fd_sc_hdll__dlrtn_2_0/RESET_B sky130_fd_sc_hdll__dlrtn_2_0/D
+ sky130_fd_sc_hdll__dlrtn_2_0/GATE_N sky130_fd_sc_hdll__dlrtn_2_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtn_2
Xsky130_fd_sc_hdll__or2b_2_0 sky130_fd_sc_hdll__or2b_2_0/A sky130_fd_sc_hdll__or2b_2_0/B_N
+ sky130_fd_sc_hdll__or2b_2_0/X VPWR VGND VGND VPWR sky130_fd_sc_hdll__or2b_2
Xsky130_fd_sc_hdll__diode_8_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__diode_8_0/DIODE
+ sky130_fd_sc_hdll__diode_8
Xsky130_fd_sc_hdll__sdfxtp_1_0 VPWR VGND sky130_fd_sc_hdll__sdfxtp_1_0/CLK sky130_fd_sc_hdll__sdfxtp_1_0/Q
+ sky130_fd_sc_hdll__sdfxtp_1_0/SCD sky130_fd_sc_hdll__sdfxtp_1_0/D sky130_fd_sc_hdll__sdfxtp_1_0/SCE
+ VPWR VGND sky130_fd_sc_hdll__sdfxtp_1
Xsky130_fd_sc_hdll__a211o_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_4_0/C1
+ sky130_fd_sc_hdll__a211o_4_0/B1 sky130_fd_sc_hdll__a211o_4_0/X sky130_fd_sc_hdll__a211o_4_0/A2
+ sky130_fd_sc_hdll__a211o_4_0/A1 sky130_fd_sc_hdll__a211o_4
Xsky130_fd_sc_hdll__a2bb2oi_2_0 sky130_fd_sc_hdll__a2bb2oi_2_0/A2_N sky130_fd_sc_hdll__a2bb2oi_2_0/A1_N
+ sky130_fd_sc_hdll__a2bb2oi_2_0/Y sky130_fd_sc_hdll__a2bb2oi_2_0/B2 sky130_fd_sc_hdll__a2bb2oi_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2oi_2
Xsky130_fd_sc_hdll__a21o_4_0 sky130_fd_sc_hdll__a21o_4_0/A2 sky130_fd_sc_hdll__a21o_4_0/A1
+ sky130_fd_sc_hdll__a21o_4_0/X sky130_fd_sc_hdll__a21o_4_0/B1 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_4
Xsky130_fd_sc_hdll__dlygate4sd1_1_0 sky130_fd_sc_hdll__dlygate4sd1_1_0/A sky130_fd_sc_hdll__dlygate4sd1_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd1_1
Xsky130_fd_sc_hdll__sdfxbp_2_0 VPWR VGND sky130_fd_sc_hdll__sdfxbp_2_0/Q_N sky130_fd_sc_hdll__sdfxbp_2_0/Q
+ sky130_fd_sc_hdll__sdfxbp_2_0/CLK sky130_fd_sc_hdll__sdfxbp_2_0/SCE sky130_fd_sc_hdll__sdfxbp_2_0/D
+ sky130_fd_sc_hdll__sdfxbp_2_0/SCD VGND VPWR sky130_fd_sc_hdll__sdfxbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_269 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_258 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_247 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_236 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_225 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_214 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_203 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2b_2_0 sky130_fd_sc_hdll__nor2b_2_0/B_N sky130_fd_sc_hdll__nor2b_2_0/A
+ sky130_fd_sc_hdll__nor2b_2_0/Y VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2b_2
Xsky130_fd_sc_hdll__nor4_8_0 sky130_fd_sc_hdll__nor4_8_0/A sky130_fd_sc_hdll__nor4_8_0/C
+ sky130_fd_sc_hdll__nor4_8_0/D sky130_fd_sc_hdll__nor4_8_0/B sky130_fd_sc_hdll__nor4_8_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_8
Xsky130_fd_sc_hdll__einvp_4_0 sky130_fd_sc_hdll__einvp_4_0/TE sky130_fd_sc_hdll__einvp_4_0/A
+ sky130_fd_sc_hdll__einvp_4_0/Z VPWR VGND VPWR VGND sky130_fd_sc_hdll__einvp_4
Xsky130_fd_sc_hdll__muxb8to1_1_0 VGND sky130_fd_sc_hdll__muxb8to1_1_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_1_0/D[0] sky130_fd_sc_hdll__muxb8to1_1_0/S[0] sky130_fd_sc_hdll__muxb8to1_1_0/S[1]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[1] sky130_fd_sc_hdll__muxb8to1_1_0/D[2] sky130_fd_sc_hdll__muxb8to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[3] sky130_fd_sc_hdll__muxb8to1_1_0/D[4] sky130_fd_sc_hdll__muxb8to1_1_0/S[4]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[5] sky130_fd_sc_hdll__muxb8to1_1_0/D[5] sky130_fd_sc_hdll__muxb8to1_1_0/D[6]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[6] sky130_fd_sc_hdll__muxb8to1_1_0/S[7] sky130_fd_sc_hdll__muxb8to1_1_0/D[7]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[3] sky130_fd_sc_hdll__muxb8to1_1
Xsky130_fd_sc_hdll__o2bb2a_1_0 sky130_fd_sc_hdll__o2bb2a_1_0/A1_N sky130_fd_sc_hdll__o2bb2a_1_0/X
+ sky130_fd_sc_hdll__o2bb2a_1_0/A2_N sky130_fd_sc_hdll__o2bb2a_1_0/B2 sky130_fd_sc_hdll__o2bb2a_1_0/B1
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__o2bb2a_1
Xsky130_fd_sc_hdll__or3_1_0 sky130_fd_sc_hdll__or3_1_0/A sky130_fd_sc_hdll__or3_1_0/X
+ sky130_fd_sc_hdll__or3_1_0/B sky130_fd_sc_hdll__or3_1_0/C VPWR VGND VPWR VGND sky130_fd_sc_hdll__or3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_259 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_248 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_237 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_226 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_215 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_204 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__and4b_2_0 VPWR VGND sky130_fd_sc_hdll__and4b_2_0/X sky130_fd_sc_hdll__and4b_2_0/A_N
+ sky130_fd_sc_hdll__and4b_2_0/D sky130_fd_sc_hdll__and4b_2_0/C sky130_fd_sc_hdll__and4b_2_0/B
+ VGND VPWR sky130_fd_sc_hdll__and4b_2
Xsky130_fd_sc_hdll__o22ai_1_0 sky130_fd_sc_hdll__o22ai_1_0/B2 sky130_fd_sc_hdll__o22ai_1_0/A1
+ sky130_fd_sc_hdll__o22ai_1_0/Y sky130_fd_sc_hdll__o22ai_1_0/B1 sky130_fd_sc_hdll__o22ai_1_0/A2
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__o22ai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_90 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a31o_2_0 sky130_fd_sc_hdll__a31o_2_0/X sky130_fd_sc_hdll__a31o_2_0/B1
+ sky130_fd_sc_hdll__a31o_2_0/A3 sky130_fd_sc_hdll__a31o_2_0/A1 sky130_fd_sc_hdll__a31o_2_0/A2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a31o_2
Xsky130_fd_sc_hdll__xnor3_2_0 sky130_fd_sc_hdll__xnor3_2_0/X sky130_fd_sc_hdll__xnor3_2_0/B
+ sky130_fd_sc_hdll__xnor3_2_0/C sky130_fd_sc_hdll__xnor3_2_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xnor3_2
Xsky130_fd_sc_hdll__nand2b_1_0 sky130_fd_sc_hdll__nand2b_1_0/Y sky130_fd_sc_hdll__nand2b_1_0/A_N
+ sky130_fd_sc_hdll__nand2b_1_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand2b_1
Xsky130_fd_sc_hdll__nand4bb_4_0 sky130_fd_sc_hdll__nand4bb_4_0/B_N sky130_fd_sc_hdll__nand4bb_4_0/A_N
+ sky130_fd_sc_hdll__nand4bb_4_0/C sky130_fd_sc_hdll__nand4bb_4_0/Y sky130_fd_sc_hdll__nand4bb_4_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4bb_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_249 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_238 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_227 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_216 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_205 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o211ai_1_0 sky130_fd_sc_hdll__o211ai_1_0/A1 sky130_fd_sc_hdll__o211ai_1_0/A2
+ sky130_fd_sc_hdll__o211ai_1_0/Y sky130_fd_sc_hdll__o211ai_1_0/C1 sky130_fd_sc_hdll__o211ai_1_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o211ai_1
Xsky130_fd_sc_hdll__muxb16to1_4_0 VGND sky130_fd_sc_hdll__muxb16to1_4_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_4_0/S[6] sky130_fd_sc_hdll__muxb16to1_4_0/S[10]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[12] sky130_fd_sc_hdll__muxb16to1_4_0/D[13] sky130_fd_sc_hdll__muxb16to1_4_0/D[8]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[15] sky130_fd_sc_hdll__muxb16to1_4_0/D[10] sky130_fd_sc_hdll__muxb16to1_4_0/D[9]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[14] sky130_fd_sc_hdll__muxb16to1_4_0/S[14] sky130_fd_sc_hdll__muxb16to1_4_0/D[11]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[11] sky130_fd_sc_hdll__muxb16to1_4_0/S[8] sky130_fd_sc_hdll__muxb16to1_4_0/S[15]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[12] sky130_fd_sc_hdll__muxb16to1_4_0/S[9] sky130_fd_sc_hdll__muxb16to1_4_0/S[13]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[3] sky130_fd_sc_hdll__muxb16to1_4_0/D[0] sky130_fd_sc_hdll__muxb16to1_4_0/D[4]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[5] sky130_fd_sc_hdll__muxb16to1_4_0/D[2] sky130_fd_sc_hdll__muxb16to1_4_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[6] sky130_fd_sc_hdll__muxb16to1_4_0/S[2] sky130_fd_sc_hdll__muxb16to1_4_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[7] sky130_fd_sc_hdll__muxb16to1_4_0/S[0] sky130_fd_sc_hdll__muxb16to1_4_0/S[1]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[4] sky130_fd_sc_hdll__muxb16to1_4_0/S[5] sky130_fd_sc_hdll__muxb16to1_4_0/D[7]
+ sky130_fd_sc_hdll__muxb16to1_4
Xsky130_fd_sc_hdll__ebufn_4_0 sky130_fd_sc_hdll__ebufn_4_0/A sky130_fd_sc_hdll__ebufn_4_0/Z
+ sky130_fd_sc_hdll__ebufn_4_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_4
Xsky130_fd_sc_hdll__clkmux2_1_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_1_0/S sky130_fd_sc_hdll__clkmux2_1_0/A1
+ sky130_fd_sc_hdll__clkmux2_1_0/A0 sky130_fd_sc_hdll__clkmux2_1_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_80 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_91 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o21ai_1_0 VGND VPWR sky130_fd_sc_hdll__o21ai_1_0/A2 sky130_fd_sc_hdll__o21ai_1_0/A1
+ sky130_fd_sc_hdll__o21ai_1_0/B1 sky130_fd_sc_hdll__o21ai_1_0/Y VPWR VGND sky130_fd_sc_hdll__o21ai_1
Xsky130_fd_sc_hdll__a222oi_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a222oi_1_0/C2
+ sky130_fd_sc_hdll__a222oi_1_0/C1 sky130_fd_sc_hdll__a222oi_1_0/B1 sky130_fd_sc_hdll__a222oi_1_0/A2
+ sky130_fd_sc_hdll__a222oi_1_0/A1 sky130_fd_sc_hdll__a222oi_1_0/Y sky130_fd_sc_hdll__a222oi_1_0/B2
+ sky130_fd_sc_hdll__a222oi_1
Xsky130_fd_sc_hdll__diode_6_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__diode_6_0/DIODE
+ sky130_fd_sc_hdll__diode_6
Xsky130_fd_sc_hdll__clkinv_16_0 sky130_fd_sc_hdll__clkinv_16_0/Y sky130_fd_sc_hdll__clkinv_16_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_16
Xsky130_fd_sc_hdll__a21o_2_0 sky130_fd_sc_hdll__a21o_2_0/X sky130_fd_sc_hdll__a21o_2_0/B1
+ sky130_fd_sc_hdll__a21o_2_0/A1 sky130_fd_sc_hdll__a21o_2_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__a21o_2
Xsky130_fd_sc_hdll__a211o_2_0 sky130_fd_sc_hdll__a211o_2_0/X sky130_fd_sc_hdll__a211o_2_0/A2
+ sky130_fd_sc_hdll__a211o_2_0/A1 sky130_fd_sc_hdll__a211o_2_0/B1 sky130_fd_sc_hdll__a211o_2_0/C1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a211o_2
Xsky130_fd_sc_hdll__nor4bb_1_0 sky130_fd_sc_hdll__nor4bb_1_0/A sky130_fd_sc_hdll__nor4bb_1_0/C_N
+ sky130_fd_sc_hdll__nor4bb_1_0/D_N sky130_fd_sc_hdll__nor4bb_1_0/B sky130_fd_sc_hdll__nor4bb_1_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_239 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_228 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_217 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_206 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_1_0 sky130_fd_sc_hdll__isobufsrc_1_0/A sky130_fd_sc_hdll__isobufsrc_1_0/X
+ sky130_fd_sc_hdll__isobufsrc_1_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_1
Xsky130_fd_sc_hdll__or4_4_0 sky130_fd_sc_hdll__or4_4_0/B sky130_fd_sc_hdll__or4_4_0/C
+ sky130_fd_sc_hdll__or4_4_0/A sky130_fd_sc_hdll__or4_4_0/D sky130_fd_sc_hdll__or4_4_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__or4_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_70 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_81 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_92 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor4_6_0 sky130_fd_sc_hdll__nor4_6_0/A sky130_fd_sc_hdll__nor4_6_0/C
+ sky130_fd_sc_hdll__nor4_6_0/D sky130_fd_sc_hdll__nor4_6_0/B sky130_fd_sc_hdll__nor4_6_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_6
Xsky130_fd_sc_hdll__and4bb_4_0 sky130_fd_sc_hdll__and4bb_4_0/C sky130_fd_sc_hdll__and4bb_4_0/A_N
+ sky130_fd_sc_hdll__and4bb_4_0/D sky130_fd_sc_hdll__and4bb_4_0/X sky130_fd_sc_hdll__and4bb_4_0/B_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_4
Xsky130_fd_sc_hdll__einvp_2_0 sky130_fd_sc_hdll__einvp_2_0/A sky130_fd_sc_hdll__einvp_2_0/Z
+ sky130_fd_sc_hdll__einvp_2_0/TE VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvp_2
Xsky130_fd_sc_hdll__a221oi_1_0 sky130_fd_sc_hdll__a221oi_1_0/Y sky130_fd_sc_hdll__a221oi_1_0/C1
+ sky130_fd_sc_hdll__a221oi_1_0/A1 sky130_fd_sc_hdll__a221oi_1_0/A2 sky130_fd_sc_hdll__a221oi_1_0/B2
+ sky130_fd_sc_hdll__a221oi_1_0/B1 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a221oi_1
Xsky130_fd_sc_hdll__buf_8_0 sky130_fd_sc_hdll__buf_8_0/A sky130_fd_sc_hdll__buf_8_0/X
+ VGND VPWR VPWR VGND sky130_fd_sc_hdll__buf_8
Xsky130_fd_sc_hdll__inv_8_0 sky130_fd_sc_hdll__inv_8_0/A sky130_fd_sc_hdll__inv_8_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__inv_8
Xsky130_fd_sc_hdll__o22a_1_0 sky130_fd_sc_hdll__o22a_1_0/A2 sky130_fd_sc_hdll__o22a_1_0/X
+ sky130_fd_sc_hdll__o22a_1_0/B1 sky130_fd_sc_hdll__o22a_1_0/A1 sky130_fd_sc_hdll__o22a_1_0/B2
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o22a_1
Xsky130_fd_sc_hdll__inputiso0p_1_0 sky130_fd_sc_hdll__inputiso0p_1_0/X sky130_fd_sc_hdll__inputiso0p_1_0/SLEEP
+ sky130_fd_sc_hdll__inputiso0p_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__inputiso0p_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_229 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_218 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_207 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand3b_4_0 sky130_fd_sc_hdll__nand3b_4_0/A_N sky130_fd_sc_hdll__nand3b_4_0/Y
+ sky130_fd_sc_hdll__nand3b_4_0/B sky130_fd_sc_hdll__nand3b_4_0/C VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__nand3b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_60 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_71 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_82 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_93 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor3_1_0 sky130_fd_sc_hdll__nor3_1_0/C sky130_fd_sc_hdll__nor3_1_0/Y
+ sky130_fd_sc_hdll__nor3_1_0/A sky130_fd_sc_hdll__nor3_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_219 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_208 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4bb_2_0 sky130_fd_sc_hdll__nand4bb_2_0/D sky130_fd_sc_hdll__nand4bb_2_0/C
+ sky130_fd_sc_hdll__nand4bb_2_0/B_N sky130_fd_sc_hdll__nand4bb_2_0/A_N sky130_fd_sc_hdll__nand4bb_2_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4bb_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_50 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_61 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_72 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_83 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_94 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__muxb16to1_2_0 sky130_fd_sc_hdll__muxb16to1_2_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb16to1_2_0/D[2] sky130_fd_sc_hdll__muxb16to1_2_0/D[1]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[7] sky130_fd_sc_hdll__muxb16to1_2_0/S[6] sky130_fd_sc_hdll__muxb16to1_2_0/S[5]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[9] sky130_fd_sc_hdll__muxb16to1_2_0/D[8] sky130_fd_sc_hdll__muxb16to1_2_0/S[14]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[13] sky130_fd_sc_hdll__muxb16to1_2_0/S[12] sky130_fd_sc_hdll__muxb16to1_2_0/S[11]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[10] sky130_fd_sc_hdll__muxb16to1_2_0/S[9] sky130_fd_sc_hdll__muxb16to1_2_0/S[8]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[15] sky130_fd_sc_hdll__muxb16to1_2_0/D[14] sky130_fd_sc_hdll__muxb16to1_2_0/D[13]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[12] sky130_fd_sc_hdll__muxb16to1_2_0/D[11] sky130_fd_sc_hdll__muxb16to1_2_0/D[10]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[15] sky130_fd_sc_hdll__muxb16to1_2_0/S[4] sky130_fd_sc_hdll__muxb16to1_2_0/S[3]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[2] sky130_fd_sc_hdll__muxb16to1_2_0/S[1] sky130_fd_sc_hdll__muxb16to1_2_0/S[0]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[7] sky130_fd_sc_hdll__muxb16to1_2_0/D[6] sky130_fd_sc_hdll__muxb16to1_2_0/D[5]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[4] sky130_fd_sc_hdll__muxb16to1_2_0/D[3] sky130_fd_sc_hdll__muxb16to1_2_0/D[0]
+ sky130_fd_sc_hdll__muxb16to1_2
Xsky130_fd_sc_hdll__ebufn_2_0 sky130_fd_sc_hdll__ebufn_2_0/Z sky130_fd_sc_hdll__ebufn_2_0/A
+ sky130_fd_sc_hdll__ebufn_2_0/TE_B VGND VPWR VGND VPWR sky130_fd_sc_hdll__ebufn_2
Xsky130_fd_sc_hdll__diode_4_0 sky130_fd_sc_hdll__diode_4_0/DIODE VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__diode_4
Xsky130_fd_sc_hdll__and3_1_0 VGND VPWR sky130_fd_sc_hdll__and3_1_0/X sky130_fd_sc_hdll__and3_1_0/B
+ sky130_fd_sc_hdll__and3_1_0/A sky130_fd_sc_hdll__and3_1_0/C VPWR VGND sky130_fd_sc_hdll__and3_1
Xsky130_fd_sc_hdll__clkbuf_1_0 VGND VPWR sky130_fd_sc_hdll__clkbuf_1_0/X sky130_fd_sc_hdll__clkbuf_1_0/A
+ VPWR sky130_fd_sc_hdll__clkbuf_1_0/VNB VGND sky130_fd_sc_hdll__clkbuf_1
Xsky130_fd_sc_hdll__clkinv_1_0 sky130_fd_sc_hdll__clkinv_1_0/Y sky130_fd_sc_hdll__clkinv_1_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkinv_1
Xsky130_fd_sc_hdll__sdfstp_1_0 sky130_fd_sc_hdll__sdfstp_1_0/SCE sky130_fd_sc_hdll__sdfstp_1_0/SET_B
+ VPWR VGND sky130_fd_sc_hdll__sdfstp_1_0/CLK sky130_fd_sc_hdll__sdfstp_1_0/D sky130_fd_sc_hdll__sdfstp_1_0/SCD
+ sky130_fd_sc_hdll__sdfstp_1_0/Q VPWR VGND sky130_fd_sc_hdll__sdfstp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_209 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfstp_4_0 sky130_fd_sc_hdll__dfstp_4_0/Q sky130_fd_sc_hdll__dfstp_4_0/D
+ VPWR sky130_fd_sc_hdll__dfstp_4_0/CLK VGND VPWR VGND sky130_fd_sc_hdll__dfstp_4_0/SET_B
+ sky130_fd_sc_hdll__dfstp_4
Xsky130_fd_sc_hdll__or4_2_0 sky130_fd_sc_hdll__or4_2_0/B sky130_fd_sc_hdll__or4_2_0/C
+ sky130_fd_sc_hdll__or4_2_0/A sky130_fd_sc_hdll__or4_2_0/X sky130_fd_sc_hdll__or4_2_0/D
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4_2
Xsky130_fd_sc_hdll__sdfsbp_2_0 sky130_fd_sc_hdll__sdfsbp_2_0/Q_N sky130_fd_sc_hdll__sdfsbp_2_0/Q
+ sky130_fd_sc_hdll__sdfsbp_2_0/CLK sky130_fd_sc_hdll__sdfsbp_2_0/D sky130_fd_sc_hdll__sdfsbp_2_0/SCD
+ sky130_fd_sc_hdll__sdfsbp_2_0/SCE sky130_fd_sc_hdll__sdfsbp_2_0/SET_B VGND VPWR
+ VPWR VGND sky130_fd_sc_hdll__sdfsbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_40 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_51 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_62 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_73 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_84 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_95 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a21boi_1_0 sky130_fd_sc_hdll__a21boi_1_0/Y sky130_fd_sc_hdll__a21boi_1_0/A1
+ sky130_fd_sc_hdll__a21boi_1_0/B1_N sky130_fd_sc_hdll__a21boi_1_0/A2 VPWR VGND VPWR
+ VGND sky130_fd_sc_hdll__a21boi_1
Xsky130_fd_sc_hdll__and4bb_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4bb_2_0/A_N
+ sky130_fd_sc_hdll__and4bb_2_0/C sky130_fd_sc_hdll__and4bb_2_0/B_N sky130_fd_sc_hdll__and4bb_2_0/X
+ sky130_fd_sc_hdll__and4bb_2_0/D sky130_fd_sc_hdll__and4bb_2
Xsky130_fd_sc_hdll__nand3_1_0 sky130_fd_sc_hdll__nand3_1_0/Y sky130_fd_sc_hdll__nand3_1_0/A
+ sky130_fd_sc_hdll__nand3_1_0/C sky130_fd_sc_hdll__nand3_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nand3_1
Xsky130_fd_sc_hdll__nor4_4_0 sky130_fd_sc_hdll__nor4_4_0/A sky130_fd_sc_hdll__nor4_4_0/C
+ sky130_fd_sc_hdll__nor4_4_0/Y sky130_fd_sc_hdll__nor4_4_0/D sky130_fd_sc_hdll__nor4_4_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4_4
Xsky130_fd_sc_hdll__mux2_1_0 VGND VPWR sky130_fd_sc_hdll__mux2_1_0/S sky130_fd_sc_hdll__mux2_1_0/A1
+ sky130_fd_sc_hdll__mux2_1_0/A0 sky130_fd_sc_hdll__mux2_1_0/X VPWR VGND sky130_fd_sc_hdll__mux2_1
Xsky130_fd_sc_hdll__and2b_1_0 sky130_fd_sc_hdll__and2b_1_0/X sky130_fd_sc_hdll__and2b_1_0/A_N
+ sky130_fd_sc_hdll__and2b_1_0/B VGND VPWR VPWR VGND sky130_fd_sc_hdll__and2b_1
Xsky130_fd_sc_hdll__buf_6_0 VPWR VGND sky130_fd_sc_hdll__buf_6_0/X sky130_fd_sc_hdll__buf_6_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_6
Xsky130_fd_sc_hdll__inv_16_0 sky130_fd_sc_hdll__inv_16_0/Y sky130_fd_sc_hdll__inv_16_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__inv_16
Xsky130_fd_sc_hdll__inv_6_0 sky130_fd_sc_hdll__inv_6_0/Y sky130_fd_sc_hdll__inv_6_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_6
Xsky130_fd_sc_hdll__tapvgnd2_1_0 VPWR VGND VPWR sky130_fd_sc_hdll__tapvgnd2_1
Xsky130_fd_sc_hdll__nand3b_2_0 sky130_fd_sc_hdll__nand3b_2_0/Y sky130_fd_sc_hdll__nand3b_2_0/C
+ sky130_fd_sc_hdll__nand3b_2_0/A_N sky130_fd_sc_hdll__nand3b_2_0/B VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__nand3b_2
Xsky130_fd_sc_hdll__sdfrtp_1_0 VPWR VGND VGND VPWR sky130_fd_sc_hdll__sdfrtp_1_0/RESET_B
+ sky130_fd_sc_hdll__sdfrtp_1_0/Q sky130_fd_sc_hdll__sdfrtp_1_0/CLK sky130_fd_sc_hdll__sdfrtp_1_0/D
+ sky130_fd_sc_hdll__sdfrtp_1_0/SCD sky130_fd_sc_hdll__sdfrtp_1_0/SCE sky130_fd_sc_hdll__sdfrtp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_30 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_41 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_52 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_63 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_74 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_85 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_96 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_4_0 sky130_fd_sc_hdll__dfrtp_4_0/Q sky130_fd_sc_hdll__dfrtp_4_0/D
+ sky130_fd_sc_hdll__dfrtp_4_0/CLK VGND VPWR sky130_fd_sc_hdll__dfrtp_4_0/RESET_B
+ VPWR VGND sky130_fd_sc_hdll__dfrtp_4
Xsky130_fd_sc_hdll__isobufsrc_16_0 sky130_fd_sc_hdll__isobufsrc_16_0/A sky130_fd_sc_hdll__isobufsrc_16_0/X
+ sky130_fd_sc_hdll__isobufsrc_16_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_16
Xsky130_fd_sc_hdll__sdlclkp_4_0 sky130_fd_sc_hdll__sdlclkp_4_0/SCE sky130_fd_sc_hdll__sdlclkp_4_0/GATE
+ sky130_fd_sc_hdll__sdlclkp_4_0/GCLK VGND VPWR sky130_fd_sc_hdll__sdlclkp_4_0/CLK
+ VPWR VGND sky130_fd_sc_hdll__sdlclkp_4
Xsky130_fd_sc_hdll__sdfrbp_2_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__sdfrbp_2_0/RESET_B
+ sky130_fd_sc_hdll__sdfrbp_2_0/Q_N sky130_fd_sc_hdll__sdfrbp_2_0/Q sky130_fd_sc_hdll__sdfrbp_2_0/SCD
+ sky130_fd_sc_hdll__sdfrbp_2_0/SCE sky130_fd_sc_hdll__sdfrbp_2_0/CLK sky130_fd_sc_hdll__sdfrbp_2_0/D
+ sky130_fd_sc_hdll__sdfrbp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_190 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or3b_1_0 sky130_fd_sc_hdll__or3b_1_0/A sky130_fd_sc_hdll__or3b_1_0/C_N
+ sky130_fd_sc_hdll__or3b_1_0/X sky130_fd_sc_hdll__or3b_1_0/B VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__or3b_1
Xsky130_fd_sc_hdll__o32ai_1_0 sky130_fd_sc_hdll__o32ai_1_0/A2 sky130_fd_sc_hdll__o32ai_1_0/Y
+ sky130_fd_sc_hdll__o32ai_1_0/A1 sky130_fd_sc_hdll__o32ai_1_0/A3 sky130_fd_sc_hdll__o32ai_1_0/B2
+ sky130_fd_sc_hdll__o32ai_1_0/B1 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o32ai_1
Xsky130_fd_sc_hdll__xor2_1_0 sky130_fd_sc_hdll__xor2_1_0/B sky130_fd_sc_hdll__xor2_1_0/X
+ sky130_fd_sc_hdll__xor2_1_0/A VGND VPWR VPWR VGND sky130_fd_sc_hdll__xor2_1
Xsky130_fd_sc_hdll__o21ba_1_0 sky130_fd_sc_hdll__o21ba_1_0/B1_N sky130_fd_sc_hdll__o21ba_1_0/A1
+ sky130_fd_sc_hdll__o21ba_1_0/X sky130_fd_sc_hdll__o21ba_1_0/A2 VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__o21ba_1
Xsky130_fd_sc_hdll__or4bb_1_0 sky130_fd_sc_hdll__or4bb_1_0/A sky130_fd_sc_hdll__or4bb_1_0/X
+ sky130_fd_sc_hdll__or4bb_1_0/B sky130_fd_sc_hdll__or4bb_1_0/D_N sky130_fd_sc_hdll__or4bb_1_0/C_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4bb_1
Xsky130_fd_sc_hdll__and4_4_0 sky130_fd_sc_hdll__and4_4_0/X sky130_fd_sc_hdll__and4_4_0/C
+ sky130_fd_sc_hdll__and4_4_0/A sky130_fd_sc_hdll__and4_4_0/B sky130_fd_sc_hdll__and4_4_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_31 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_42 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_53 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_64 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_75 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_86 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_97 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_20 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o221ai_1_0 sky130_fd_sc_hdll__o221ai_1_0/A2 sky130_fd_sc_hdll__o221ai_1_0/Y
+ sky130_fd_sc_hdll__o221ai_1_0/B1 sky130_fd_sc_hdll__o221ai_1_0/C1 sky130_fd_sc_hdll__o221ai_1_0/A1
+ sky130_fd_sc_hdll__o221ai_1_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221ai_1
Xsky130_fd_sc_hdll__nor3b_1_0 sky130_fd_sc_hdll__nor3b_1_0/C_N sky130_fd_sc_hdll__nor3b_1_0/Y
+ sky130_fd_sc_hdll__nor3b_1_0/A sky130_fd_sc_hdll__nor3b_1_0/B VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__nor3b_1
Xsky130_fd_sc_hdll__mux2_16_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_16_0/X sky130_fd_sc_hdll__mux2_16_0/S
+ sky130_fd_sc_hdll__mux2_16_0/A1 sky130_fd_sc_hdll__mux2_16_0/A0 sky130_fd_sc_hdll__mux2_16
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_191 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_180 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4_4_0 sky130_fd_sc_hdll__nand4_4_0/A sky130_fd_sc_hdll__nand4_4_0/D
+ sky130_fd_sc_hdll__nand4_4_0/C sky130_fd_sc_hdll__nand4_4_0/B sky130_fd_sc_hdll__nand4_4_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__nand4_4
Xsky130_fd_sc_hdll__decap_8_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_8
Xsky130_fd_sc_hdll__diode_2_0 sky130_fd_sc_hdll__diode_2_0/DIODE VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__diode_2
Xsky130_fd_sc_hdll__o31ai_1_0 sky130_fd_sc_hdll__o31ai_1_0/Y sky130_fd_sc_hdll__o31ai_1_0/A2
+ sky130_fd_sc_hdll__o31ai_1_0/A1 sky130_fd_sc_hdll__o31ai_1_0/A3 sky130_fd_sc_hdll__o31ai_1_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__o31ai_1
Xsky130_fd_sc_hdll__clkinv_12_0 sky130_fd_sc_hdll__clkinv_12_0/Y sky130_fd_sc_hdll__clkinv_12_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_12
Xsky130_fd_sc_hdll__and3b_4_0 sky130_fd_sc_hdll__and3b_4_0/A_N sky130_fd_sc_hdll__and3b_4_0/X
+ sky130_fd_sc_hdll__and3b_4_0/C sky130_fd_sc_hdll__and3b_4_0/B VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__and3b_4
Xsky130_fd_sc_hdll__einvn_1_0 sky130_fd_sc_hdll__einvn_1_0/Z sky130_fd_sc_hdll__einvn_1_0/A
+ sky130_fd_sc_hdll__einvn_1_0/TE_B VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_1
Xsky130_fd_sc_hdll__dfstp_2_0 sky130_fd_sc_hdll__dfstp_2_0/Q VGND sky130_fd_sc_hdll__dfstp_2_0/CLK
+ VPWR sky130_fd_sc_hdll__dfstp_2_0/D VPWR VGND sky130_fd_sc_hdll__dfstp_2_0/SET_B
+ sky130_fd_sc_hdll__dfstp_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_32 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_43 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_54 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_65 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_76 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_87 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_98 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_10 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_21 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__xnor2_4_0 sky130_fd_sc_hdll__xnor2_4_0/Y sky130_fd_sc_hdll__xnor2_4_0/B
+ sky130_fd_sc_hdll__xnor2_4_0/A VGND VPWR VGND VPWR sky130_fd_sc_hdll__xnor2_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_192 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_181 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_170 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__fill_1_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__fill_1
Xsky130_fd_sc_hdll__or4b_4_0 sky130_fd_sc_hdll__or4b_4_0/D_N sky130_fd_sc_hdll__or4b_4_0/B
+ sky130_fd_sc_hdll__or4b_4_0/C sky130_fd_sc_hdll__or4b_4_0/A sky130_fd_sc_hdll__or4b_4_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__or4b_4
Xsky130_fd_sc_hdll__a2bb2o_4_0 sky130_fd_sc_hdll__a2bb2o_4_0/X sky130_fd_sc_hdll__a2bb2o_4_0/B1
+ sky130_fd_sc_hdll__a2bb2o_4_0/B2 sky130_fd_sc_hdll__a2bb2o_4_0/A1_N sky130_fd_sc_hdll__a2bb2o_4_0/A2_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_4
Xsky130_fd_sc_hdll__nor4_2_0 sky130_fd_sc_hdll__nor4_2_0/C sky130_fd_sc_hdll__nor4_2_0/D
+ sky130_fd_sc_hdll__nor4_2_0/Y sky130_fd_sc_hdll__nor4_2_0/A sky130_fd_sc_hdll__nor4_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4_2
Xsky130_fd_sc_hdll__xor3_4_0 sky130_fd_sc_hdll__xor3_4_0/X sky130_fd_sc_hdll__xor3_4_0/C
+ sky130_fd_sc_hdll__xor3_4_0/B sky130_fd_sc_hdll__xor3_4_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_4
Xsky130_fd_sc_hdll__dlrtp_4_0 sky130_fd_sc_hdll__dlrtp_4_0/RESET_B sky130_fd_sc_hdll__dlrtp_4_0/D
+ sky130_fd_sc_hdll__dlrtp_4_0/GATE sky130_fd_sc_hdll__dlrtp_4_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_0 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_8_0 sky130_fd_sc_hdll__isobufsrc_8_0/A sky130_fd_sc_hdll__isobufsrc_8_0/X
+ sky130_fd_sc_hdll__isobufsrc_8_0/SLEEP VPWR VGND VGND VPWR sky130_fd_sc_hdll__isobufsrc_8
Xsky130_fd_sc_hdll__a32o_1_0 sky130_fd_sc_hdll__a32o_1_0/X sky130_fd_sc_hdll__a32o_1_0/A3
+ sky130_fd_sc_hdll__a32o_1_0/B2 sky130_fd_sc_hdll__a32o_1_0/B1 sky130_fd_sc_hdll__a32o_1_0/A1
+ sky130_fd_sc_hdll__a32o_1_0/A2 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a32o_1
Xsky130_fd_sc_hdll__buf_4_0 VPWR VGND sky130_fd_sc_hdll__buf_4_0/X sky130_fd_sc_hdll__buf_4_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_4
Xsky130_fd_sc_hdll__inv_4_0 sky130_fd_sc_hdll__inv_4_0/Y sky130_fd_sc_hdll__inv_4_0/A
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_33 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_44 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_55 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_66 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_77 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_88 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_99 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_11 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_22 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dfrtp_2_0 sky130_fd_sc_hdll__dfrtp_2_0/RESET_B VPWR VGND sky130_fd_sc_hdll__dfrtp_2_0/Q
+ sky130_fd_sc_hdll__dfrtp_2_0/CLK sky130_fd_sc_hdll__dfrtp_2_0/D VPWR VGND sky130_fd_sc_hdll__dfrtp_2
Xsky130_fd_sc_hdll__nor4b_4_0 sky130_fd_sc_hdll__nor4b_4_0/B sky130_fd_sc_hdll__nor4b_4_0/A
+ sky130_fd_sc_hdll__nor4b_4_0/D_N sky130_fd_sc_hdll__nor4b_4_0/C sky130_fd_sc_hdll__nor4b_4_0/Y
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor4b_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_160 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a211oi_4_0 sky130_fd_sc_hdll__a211oi_4_0/A2 sky130_fd_sc_hdll__a211oi_4_0/A1
+ sky130_fd_sc_hdll__a211oi_4_0/C1 sky130_fd_sc_hdll__a211oi_4_0/Y sky130_fd_sc_hdll__a211oi_4_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__a211oi_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_193 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_182 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_171 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdlclkp_2_0 sky130_fd_sc_hdll__sdlclkp_2_0/CLK VPWR VGND sky130_fd_sc_hdll__sdlclkp_2_0/GCLK
+ sky130_fd_sc_hdll__sdlclkp_2_0/SCE sky130_fd_sc_hdll__sdlclkp_2_0/GATE VPWR VGND
+ sky130_fd_sc_hdll__sdlclkp_2
Xsky130_fd_sc_hdll__a22oi_1_0 sky130_fd_sc_hdll__a22oi_1_0/B1 sky130_fd_sc_hdll__a22oi_1_0/A1
+ sky130_fd_sc_hdll__a22oi_1_0/B2 sky130_fd_sc_hdll__a22oi_1_0/A2 sky130_fd_sc_hdll__a22oi_1_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22oi_1
Xsky130_fd_sc_hdll__muxb4to1_1_0 sky130_fd_sc_hdll__muxb4to1_1_0/S[0] sky130_fd_sc_hdll__muxb4to1_1_0/D[0]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[2] sky130_fd_sc_hdll__muxb4to1_1_0/D[3] sky130_fd_sc_hdll__muxb4to1_1_0/S[3]
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__muxb4to1_1_0/Z sky130_fd_sc_hdll__muxb4to1_1
Xsky130_fd_sc_hdll__o221a_1_0 sky130_fd_sc_hdll__o221a_1_0/A2 sky130_fd_sc_hdll__o221a_1_0/X
+ sky130_fd_sc_hdll__o221a_1_0/B1 sky130_fd_sc_hdll__o221a_1_0/C1 sky130_fd_sc_hdll__o221a_1_0/A1
+ sky130_fd_sc_hdll__o221a_1_0/B2 VPWR VGND VGND VPWR sky130_fd_sc_hdll__o221a_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_1 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlxtn_1_0 VGND VPWR sky130_fd_sc_hdll__dlxtn_1_0/Q sky130_fd_sc_hdll__dlxtn_1_0/GATE_N
+ sky130_fd_sc_hdll__dlxtn_1_0/D VPWR VGND sky130_fd_sc_hdll__dlxtn_1
Xsky130_fd_sc_hdll__and4_2_0 sky130_fd_sc_hdll__and4_2_0/X sky130_fd_sc_hdll__and4_2_0/C
+ sky130_fd_sc_hdll__and4_2_0/A sky130_fd_sc_hdll__and4_2_0/B sky130_fd_sc_hdll__and4_2_0/D
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__and4_2
Xsky130_fd_sc_hdll__o21bai_1_0 sky130_fd_sc_hdll__o21bai_1_0/A1 sky130_fd_sc_hdll__o21bai_1_0/Y
+ sky130_fd_sc_hdll__o21bai_1_0/B1_N sky130_fd_sc_hdll__o21bai_1_0/A2 VPWR VGND VPWR
+ VGND sky130_fd_sc_hdll__o21bai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_12 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__a22o_1_0 sky130_fd_sc_hdll__a22o_1_0/A1 sky130_fd_sc_hdll__a22o_1_0/A2
+ sky130_fd_sc_hdll__a22o_1_0/X sky130_fd_sc_hdll__a22o_1_0/B2 sky130_fd_sc_hdll__a22o_1_0/B1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a22o_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_23 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_34 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_45 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_56 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_67 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_78 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_89 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_320 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_150 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_161 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_194 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_183 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_172 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfbbp_1_0 sky130_fd_sc_hdll__sdfbbp_1_0/SCD sky130_fd_sc_hdll__sdfbbp_1_0/SCE
+ sky130_fd_sc_hdll__sdfbbp_1_0/RESET_B VGND sky130_fd_sc_hdll__sdfbbp_1_0/CLK sky130_fd_sc_hdll__sdfbbp_1_0/Q
+ VPWR sky130_fd_sc_hdll__sdfbbp_1_0/D sky130_fd_sc_hdll__sdfbbp_1_0/Q_N sky130_fd_sc_hdll__sdfbbp_1_0/SET_B
+ VPWR VGND sky130_fd_sc_hdll__sdfbbp_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_2 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or2_1_0 sky130_fd_sc_hdll__or2_1_0/A sky130_fd_sc_hdll__or2_1_0/X
+ sky130_fd_sc_hdll__or2_1_0/B VPWR VGND VGND VPWR sky130_fd_sc_hdll__or2_1
Xsky130_fd_sc_hdll__a21oi_1_0 sky130_fd_sc_hdll__a21oi_1_0/A1 sky130_fd_sc_hdll__a21oi_1_0/B1
+ sky130_fd_sc_hdll__a21oi_1_0/Y sky130_fd_sc_hdll__a21oi_1_0/A2 VPWR VGND VPWR VGND
+ sky130_fd_sc_hdll__a21oi_1
Xsky130_fd_sc_hdll__nand4_2_0 sky130_fd_sc_hdll__nand4_2_0/B sky130_fd_sc_hdll__nand4_2_0/A
+ sky130_fd_sc_hdll__nand4_2_0/Y sky130_fd_sc_hdll__nand4_2_0/D sky130_fd_sc_hdll__nand4_2_0/C
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand4_2
Xsky130_fd_sc_hdll__decap_6_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__decap_6
Xsky130_fd_sc_hdll__o211a_1_0 sky130_fd_sc_hdll__o211a_1_0/C1 sky130_fd_sc_hdll__o211a_1_0/B1
+ sky130_fd_sc_hdll__o211a_1_0/A2 sky130_fd_sc_hdll__o211a_1_0/A1 sky130_fd_sc_hdll__o211a_1_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211a_1
Xsky130_fd_sc_hdll__and3b_2_0 VGND VPWR sky130_fd_sc_hdll__and3b_2_0/B sky130_fd_sc_hdll__and3b_2_0/X
+ sky130_fd_sc_hdll__and3b_2_0/A_N sky130_fd_sc_hdll__and3b_2_0/C VGND VPWR sky130_fd_sc_hdll__and3b_2
Xsky130_fd_sc_hdll__bufbuf_16_0 sky130_fd_sc_hdll__bufbuf_16_0/A sky130_fd_sc_hdll__bufbuf_16_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufbuf_16
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_35 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_46 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_57 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_68 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_79 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_13 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_310 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_321 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_24 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_140 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_151 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_162 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_195 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_184 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_173 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__xnor2_2_0 VGND VPWR sky130_fd_sc_hdll__xnor2_2_0/Y sky130_fd_sc_hdll__xnor2_2_0/A
+ sky130_fd_sc_hdll__xnor2_2_0/B VPWR VGND sky130_fd_sc_hdll__xnor2_2
Xsky130_fd_sc_hdll__clkbuf_8_0 sky130_fd_sc_hdll__clkbuf_8_0/X sky130_fd_sc_hdll__clkbuf_8_0/A
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_8
Xsky130_fd_sc_hdll__clkinv_8_0 sky130_fd_sc_hdll__clkinv_8_0/Y sky130_fd_sc_hdll__clkinv_8_0/A
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__clkinv_8
Xsky130_fd_sc_hdll__sdfxtp_4_0 VGND VPWR sky130_fd_sc_hdll__sdfxtp_4_0/SCD sky130_fd_sc_hdll__sdfxtp_4_0/D
+ sky130_fd_sc_hdll__sdfxtp_4_0/SCE sky130_fd_sc_hdll__sdfxtp_4_0/CLK sky130_fd_sc_hdll__sdfxtp_4_0/Q
+ VGND VPWR sky130_fd_sc_hdll__sdfxtp_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_3 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or4b_2_0 sky130_fd_sc_hdll__or4b_2_0/C sky130_fd_sc_hdll__or4b_2_0/A
+ sky130_fd_sc_hdll__or4b_2_0/X sky130_fd_sc_hdll__or4b_2_0/B sky130_fd_sc_hdll__or4b_2_0/D_N
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__or4b_2
Xsky130_fd_sc_hdll__a2bb2o_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__a2bb2o_2_0/B1
+ sky130_fd_sc_hdll__a2bb2o_2_0/A1_N sky130_fd_sc_hdll__a2bb2o_2_0/A2_N sky130_fd_sc_hdll__a2bb2o_2_0/X
+ sky130_fd_sc_hdll__a2bb2o_2_0/B2 sky130_fd_sc_hdll__a2bb2o_2
Xsky130_fd_sc_hdll__xor3_2_0 sky130_fd_sc_hdll__xor3_2_0/X sky130_fd_sc_hdll__xor3_2_0/C
+ sky130_fd_sc_hdll__xor3_2_0/B sky130_fd_sc_hdll__xor3_2_0/A VGND VPWR VGND VPWR
+ sky130_fd_sc_hdll__xor3_2
Xsky130_fd_sc_hdll__dlrtp_2_0 sky130_fd_sc_hdll__dlrtp_2_0/RESET_B sky130_fd_sc_hdll__dlrtp_2_0/D
+ sky130_fd_sc_hdll__dlrtp_2_0/GATE sky130_fd_sc_hdll__dlrtp_2_0/Q VGND VPWR VPWR
+ VGND sky130_fd_sc_hdll__dlrtp_2
Xsky130_fd_sc_hdll__buf_2_0 VPWR VGND sky130_fd_sc_hdll__buf_2_0/X sky130_fd_sc_hdll__buf_2_0/A
+ VPWR VGND sky130_fd_sc_hdll__buf_2
Xsky130_fd_sc_hdll__inv_12_0 sky130_fd_sc_hdll__inv_12_0/A sky130_fd_sc_hdll__inv_12_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__inv_12
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_36 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_47 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_58 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_69 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_300 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_14 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_311 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_322 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_25 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inv_2_0 sky130_fd_sc_hdll__inv_2_0/A sky130_fd_sc_hdll__inv_2_0/Y
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__inv_2
Xsky130_fd_sc_hdll__tap_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hdll__tap_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_130 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_141 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_152 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__dlygate4sd3_1_0 sky130_fd_sc_hdll__dlygate4sd3_1_0/A sky130_fd_sc_hdll__dlygate4sd3_1_0/X
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__dlygate4sd3_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_196 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_185 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_174 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_163 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__muxb8to1_4_0 VGND sky130_fd_sc_hdll__muxb8to1_4_0/Z VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_4_0/S[6] sky130_fd_sc_hdll__muxb8to1_4_0/D[3] sky130_fd_sc_hdll__muxb8to1_4_0/D[0]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[4] sky130_fd_sc_hdll__muxb8to1_4_0/D[5] sky130_fd_sc_hdll__muxb8to1_4_0/D[2]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[1] sky130_fd_sc_hdll__muxb8to1_4_0/D[6] sky130_fd_sc_hdll__muxb8to1_4_0/S[2]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[3] sky130_fd_sc_hdll__muxb8to1_4_0/S[7] sky130_fd_sc_hdll__muxb8to1_4_0/S[0]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[1] sky130_fd_sc_hdll__muxb8to1_4_0/S[4] sky130_fd_sc_hdll__muxb8to1_4_0/S[5]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[7] sky130_fd_sc_hdll__muxb8to1_4
Xsky130_fd_sc_hdll__mux2_8_0 sky130_fd_sc_hdll__mux2_8_0/S sky130_fd_sc_hdll__mux2_8_0/A1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_8_0/A0 sky130_fd_sc_hdll__mux2_8_0/X
+ sky130_fd_sc_hdll__mux2_8
Xsky130_fd_sc_hdll__o2bb2a_4_0 sky130_fd_sc_hdll__o2bb2a_4_0/A2_N sky130_fd_sc_hdll__o2bb2a_4_0/A1_N
+ sky130_fd_sc_hdll__o2bb2a_4_0/X sky130_fd_sc_hdll__o2bb2a_4_0/B2 sky130_fd_sc_hdll__o2bb2a_4_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2a_4
Xsky130_fd_sc_hdll__nor4b_2_0 sky130_fd_sc_hdll__nor4b_2_0/D_N sky130_fd_sc_hdll__nor4b_2_0/Y
+ sky130_fd_sc_hdll__nor4b_2_0/C sky130_fd_sc_hdll__nor4b_2_0/A sky130_fd_sc_hdll__nor4b_2_0/B
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4b_2
Xsky130_fd_sc_hdll__a211oi_2_0 sky130_fd_sc_hdll__a211oi_2_0/A2 sky130_fd_sc_hdll__a211oi_2_0/C1
+ sky130_fd_sc_hdll__a211oi_2_0/B1 sky130_fd_sc_hdll__a211oi_2_0/Y sky130_fd_sc_hdll__a211oi_2_0/A1
+ VPWR VGND VPWR VGND sky130_fd_sc_hdll__a211oi_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_4 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__or3_4_0 sky130_fd_sc_hdll__or3_4_0/A sky130_fd_sc_hdll__or3_4_0/X
+ sky130_fd_sc_hdll__or3_4_0/B sky130_fd_sc_hdll__or3_4_0/C VPWR VGND VPWR VGND sky130_fd_sc_hdll__or3_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_26 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_37 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_48 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_59 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_15 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_301 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_312 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_323 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o22ai_4_0 sky130_fd_sc_hdll__o22ai_4_0/A1 sky130_fd_sc_hdll__o22ai_4_0/Y
+ sky130_fd_sc_hdll__o22ai_4_0/A2 sky130_fd_sc_hdll__o22ai_4_0/B1 sky130_fd_sc_hdll__o22ai_4_0/B2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22ai_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_120 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_131 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_142 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_153 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_164 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_197 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_186 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_175 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__mux2_12_0 VPWR VGND VPWR VGND sky130_fd_sc_hdll__mux2_12_0/X sky130_fd_sc_hdll__mux2_12_0/S
+ sky130_fd_sc_hdll__mux2_12_0/A1 sky130_fd_sc_hdll__mux2_12_0/A0 sky130_fd_sc_hdll__mux2_12
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_5 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__inputiso1n_1_0 sky130_fd_sc_hdll__inputiso1n_1_0/A sky130_fd_sc_hdll__inputiso1n_1_0/SLEEP_B
+ sky130_fd_sc_hdll__inputiso1n_1_0/X VGND VPWR VGND VPWR sky130_fd_sc_hdll__inputiso1n_1
Xsky130_fd_sc_hdll__o21a_1_0 sky130_fd_sc_hdll__o21a_1_0/X sky130_fd_sc_hdll__o21a_1_0/A1
+ sky130_fd_sc_hdll__o21a_1_0/B1 sky130_fd_sc_hdll__o21a_1_0/A2 VPWR VGND VGND VPWR
+ sky130_fd_sc_hdll__o21a_1
Xsky130_fd_sc_hdll__nand2b_4_0 sky130_fd_sc_hdll__nand2b_4_0/B sky130_fd_sc_hdll__nand2b_4_0/A_N
+ sky130_fd_sc_hdll__nand2b_4_0/Y VGND VPWR VGND VPWR sky130_fd_sc_hdll__nand2b_4
Xsky130_fd_sc_hdll__decap_4_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__decap_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_27 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_38 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_49 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__o211ai_4_0 sky130_fd_sc_hdll__o211ai_4_0/A1 sky130_fd_sc_hdll__o211ai_4_0/B1
+ sky130_fd_sc_hdll__o211ai_4_0/A2 sky130_fd_sc_hdll__o211ai_4_0/C1 sky130_fd_sc_hdll__o211ai_4_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o211ai_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_16 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_302 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_313 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_324 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_110 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_121 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_132 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_143 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_154 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nor2_1_0 sky130_fd_sc_hdll__nor2_1_0/B sky130_fd_sc_hdll__nor2_1_0/Y
+ sky130_fd_sc_hdll__nor2_1_0/A VPWR VGND VGND VPWR sky130_fd_sc_hdll__nor2_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_198 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_187 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__nand4b_1_0 sky130_fd_sc_hdll__nand4b_1_0/Y sky130_fd_sc_hdll__nand4b_1_0/C
+ sky130_fd_sc_hdll__nand4b_1_0/D sky130_fd_sc_hdll__nand4b_1_0/A_N sky130_fd_sc_hdll__nand4b_1_0/B
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__nand4b_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_176 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_165 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__clkmux2_4_0 VGND VPWR sky130_fd_sc_hdll__clkmux2_4_0/S sky130_fd_sc_hdll__clkmux2_4_0/A1
+ sky130_fd_sc_hdll__clkmux2_4_0/A0 sky130_fd_sc_hdll__clkmux2_4_0/X VPWR VGND sky130_fd_sc_hdll__clkmux2_4
Xsky130_fd_sc_hdll__o21ai_4_0 sky130_fd_sc_hdll__o21ai_4_0/Y sky130_fd_sc_hdll__o21ai_4_0/B1
+ sky130_fd_sc_hdll__o21ai_4_0/A2 sky130_fd_sc_hdll__o21ai_4_0/A1 VGND VPWR VPWR VGND
+ sky130_fd_sc_hdll__o21ai_4
Xsky130_fd_sc_hdll__clkbuf_6_0 sky130_fd_sc_hdll__clkbuf_6_0/A sky130_fd_sc_hdll__clkbuf_6_0/X
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__clkbuf_6
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_6 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sdfxtp_2_0 VPWR VGND sky130_fd_sc_hdll__sdfxtp_2_0/SCE sky130_fd_sc_hdll__sdfxtp_2_0/D
+ sky130_fd_sc_hdll__sdfxtp_2_0/SCD sky130_fd_sc_hdll__sdfxtp_2_0/Q sky130_fd_sc_hdll__sdfxtp_2_0/CLK
+ VGND VPWR sky130_fd_sc_hdll__sdfxtp_2
Xsky130_fd_sc_hdll__einvn_8_0 sky130_fd_sc_hdll__einvn_8_0/A sky130_fd_sc_hdll__einvn_8_0/TE_B
+ sky130_fd_sc_hdll__einvn_8_0/Z VGND VPWR VPWR VGND sky130_fd_sc_hdll__einvn_8
Xsky130_fd_sc_hdll__nor4bb_4_0 sky130_fd_sc_hdll__nor4bb_4_0/D_N sky130_fd_sc_hdll__nor4bb_4_0/Y
+ sky130_fd_sc_hdll__nor4bb_4_0/A sky130_fd_sc_hdll__nor4bb_4_0/B sky130_fd_sc_hdll__nor4bb_4_0/C_N
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__nor4bb_4
Xsky130_fd_sc_hdll__o2bb2ai_1_0 sky130_fd_sc_hdll__o2bb2ai_1_0/Y sky130_fd_sc_hdll__o2bb2ai_1_0/A1_N
+ sky130_fd_sc_hdll__o2bb2ai_1_0/A2_N sky130_fd_sc_hdll__o2bb2ai_1_0/B2 sky130_fd_sc_hdll__o2bb2ai_1_0/B1
+ VPWR VGND VGND VPWR sky130_fd_sc_hdll__o2bb2ai_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_28 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_39 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__isobufsrc_4_0 sky130_fd_sc_hdll__isobufsrc_4_0/A sky130_fd_sc_hdll__isobufsrc_4_0/X
+ sky130_fd_sc_hdll__isobufsrc_4_0/SLEEP VGND VPWR VGND VPWR sky130_fd_sc_hdll__isobufsrc_4
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_17 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_303 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_314 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_325 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__bufbuf_8_0 sky130_fd_sc_hdll__bufbuf_8_0/A sky130_fd_sc_hdll__bufbuf_8_0/X
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufbuf_8
Xsky130_fd_sc_hdll__bufinv_8_0 sky130_fd_sc_hdll__bufinv_8_0/A sky130_fd_sc_hdll__bufinv_8_0/Y
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__bufinv_8
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_100 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_111 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_122 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_133 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_144 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_155 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_199 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_188 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_177 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_166 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__fill_8_0 VGND VPWR VPWR VGND sky130_fd_sc_hdll__fill_8
Xsky130_fd_sc_hdll__muxb8to1_2_0 sky130_fd_sc_hdll__muxb8to1_2_0/Z VGND VPWR VGND
+ VPWR sky130_fd_sc_hdll__muxb8to1_2_0/D[2] sky130_fd_sc_hdll__muxb8to1_2_0/D[1] sky130_fd_sc_hdll__muxb8to1_2_0/S[7]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[6] sky130_fd_sc_hdll__muxb8to1_2_0/S[5] sky130_fd_sc_hdll__muxb8to1_2_0/S[4]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[3] sky130_fd_sc_hdll__muxb8to1_2_0/S[2] sky130_fd_sc_hdll__muxb8to1_2_0/S[1]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[0] sky130_fd_sc_hdll__muxb8to1_2_0/D[7] sky130_fd_sc_hdll__muxb8to1_2_0/D[6]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[5] sky130_fd_sc_hdll__muxb8to1_2_0/D[4] sky130_fd_sc_hdll__muxb8to1_2_0/D[3]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[0] sky130_fd_sc_hdll__muxb8to1_2
Xsky130_fd_sc_hdll__and2_1_0 VPWR VGND sky130_fd_sc_hdll__and2_1_0/X sky130_fd_sc_hdll__and2_1_0/B
+ sky130_fd_sc_hdll__and2_1_0/A VPWR VGND sky130_fd_sc_hdll__and2_1
Xsky130_fd_sc_hdll__o2bb2a_2_0 sky130_fd_sc_hdll__o2bb2a_2_0/A1_N sky130_fd_sc_hdll__o2bb2a_2_0/X
+ sky130_fd_sc_hdll__o2bb2a_2_0/A2_N sky130_fd_sc_hdll__o2bb2a_2_0/B2 sky130_fd_sc_hdll__o2bb2a_2_0/B1
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o2bb2a_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_7 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__sedfxbp_1_0 VGND VPWR sky130_fd_sc_hdll__sedfxbp_1_0/SCE sky130_fd_sc_hdll__sedfxbp_1_0/Q
+ sky130_fd_sc_hdll__sedfxbp_1_0/D sky130_fd_sc_hdll__sedfxbp_1_0/DE sky130_fd_sc_hdll__sedfxbp_1_0/SCD
+ sky130_fd_sc_hdll__sedfxbp_1_0/Q_N sky130_fd_sc_hdll__sedfxbp_1_0/CLK VPWR VGND
+ sky130_fd_sc_hdll__sedfxbp_1
Xsky130_fd_sc_hdll__a221oi_4_0 sky130_fd_sc_hdll__a221oi_4_0/A2 sky130_fd_sc_hdll__a221oi_4_0/Y
+ sky130_fd_sc_hdll__a221oi_4_0/C1 sky130_fd_sc_hdll__a221oi_4_0/A1 sky130_fd_sc_hdll__a221oi_4_0/B2
+ sky130_fd_sc_hdll__a221oi_4_0/B1 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a221oi_4
Xsky130_fd_sc_hdll__o22a_4_0 sky130_fd_sc_hdll__o22a_4_0/B2 sky130_fd_sc_hdll__o22a_4_0/B1
+ sky130_fd_sc_hdll__o22a_4_0/X sky130_fd_sc_hdll__o22a_4_0/A1 sky130_fd_sc_hdll__o22a_4_0/A2
+ VGND VPWR VGND VPWR sky130_fd_sc_hdll__o22a_4
Xsky130_fd_sc_hdll__a32oi_1_0 sky130_fd_sc_hdll__a32oi_1_0/A2 sky130_fd_sc_hdll__a32oi_1_0/Y
+ sky130_fd_sc_hdll__a32oi_1_0/A1 sky130_fd_sc_hdll__a32oi_1_0/B2 sky130_fd_sc_hdll__a32oi_1_0/B1
+ sky130_fd_sc_hdll__a32oi_1_0/A3 VGND VPWR VPWR VGND sky130_fd_sc_hdll__a32oi_1
Xsky130_fd_sc_hdll__or3_2_0 sky130_fd_sc_hdll__or3_2_0/A sky130_fd_sc_hdll__or3_2_0/B
+ sky130_fd_sc_hdll__or3_2_0/X sky130_fd_sc_hdll__or3_2_0/C VGND VPWR VPWR VGND sky130_fd_sc_hdll__or3_2
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_29 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_304 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_315 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_18 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_101 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_112 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_123 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_134 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_145 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_156 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_189 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_178 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
Xsky130_fd_sc_hdll__tapvpwrvgnd_1_167 VPWR VGND sky130_fd_sc_hdll__tapvpwrvgnd_1
.ends
