* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb8to1_2 D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[7]
+ S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
X0 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_2603_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_3891_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X4 VPWR D[5] a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_3891_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X6 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X7 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Z a_4142_265# a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND D[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VGND S[5] a_3277_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 VGND S[7] a_4565_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 a_4688_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND D[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_3421_69# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X27 VPWR D[4] a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_3400_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_3891_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 Z S[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 a_2854_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 a_4142_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X36 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 Z a_4565_47# a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X39 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_2603_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 VPWR S[7] a_4565_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 a_2603_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 Z a_3277_47# a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X51 a_3891_297# a_4142_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X52 Z S[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X53 Z S[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X54 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X55 a_4709_69# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 VPWR S[5] a_3277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_4142_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X59 a_3421_69# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 a_4709_69# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X61 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_2854_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X63 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 VGND D[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X65 Z a_2854_265# a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X66 VPWR D[7] a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X67 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_2603_297# a_2854_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X70 a_4688_333# a_4565_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X71 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 VGND D[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X73 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X74 VPWR D[6] a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 a_3400_333# a_3277_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X77 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 Z S[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X79 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
