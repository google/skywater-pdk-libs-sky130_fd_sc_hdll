* File: sky130_fd_sc_hdll__or4b_1.pxi.spice
* Created: Wed Sep  2 08:49:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4B_1%D_N N_D_N_c_74_n N_D_N_M1004_g N_D_N_M1000_g D_N
+ D_N N_D_N_c_73_n PM_SKY130_FD_SC_HDLL__OR4B_1%D_N
x_PM_SKY130_FD_SC_HDLL__OR4B_1%A_117_297# N_A_117_297#_M1000_d
+ N_A_117_297#_M1004_d N_A_117_297#_c_101_n N_A_117_297#_M1009_g
+ N_A_117_297#_M1001_g N_A_117_297#_c_98_n N_A_117_297#_c_102_n
+ N_A_117_297#_c_99_n N_A_117_297#_c_100_n
+ PM_SKY130_FD_SC_HDLL__OR4B_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__OR4B_1%C N_C_c_138_n N_C_M1010_g N_C_M1008_g C C C C
+ PM_SKY130_FD_SC_HDLL__OR4B_1%C
x_PM_SKY130_FD_SC_HDLL__OR4B_1%B N_B_c_174_n N_B_c_175_n N_B_c_177_n N_B_c_178_n
+ N_B_M1005_g N_B_M1006_g N_B_c_176_n B B B B N_B_c_180_n B B B B
+ PM_SKY130_FD_SC_HDLL__OR4B_1%B
x_PM_SKY130_FD_SC_HDLL__OR4B_1%A N_A_c_216_n N_A_M1007_g N_A_M1003_g A
+ N_A_c_218_n A PM_SKY130_FD_SC_HDLL__OR4B_1%A
x_PM_SKY130_FD_SC_HDLL__OR4B_1%A_225_297# N_A_225_297#_M1001_d
+ N_A_225_297#_M1006_d N_A_225_297#_M1009_s N_A_225_297#_c_254_n
+ N_A_225_297#_M1011_g N_A_225_297#_c_255_n N_A_225_297#_M1002_g
+ N_A_225_297#_c_263_n N_A_225_297#_c_330_p N_A_225_297#_c_256_n
+ N_A_225_297#_c_257_n N_A_225_297#_c_334_p N_A_225_297#_c_258_n
+ N_A_225_297#_c_299_n N_A_225_297#_c_264_n N_A_225_297#_c_265_n
+ N_A_225_297#_c_259_n N_A_225_297#_c_266_n N_A_225_297#_c_260_n
+ N_A_225_297#_c_261_n PM_SKY130_FD_SC_HDLL__OR4B_1%A_225_297#
x_PM_SKY130_FD_SC_HDLL__OR4B_1%VPWR N_VPWR_M1004_s N_VPWR_M1007_d N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n VPWR
+ N_VPWR_c_354_n N_VPWR_c_348_n PM_SKY130_FD_SC_HDLL__OR4B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4B_1%X N_X_M1002_d N_X_M1011_d N_X_c_389_n N_X_c_391_n
+ N_X_c_390_n X PM_SKY130_FD_SC_HDLL__OR4B_1%X
x_PM_SKY130_FD_SC_HDLL__OR4B_1%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1008_d
+ N_VGND_M1003_d N_VGND_c_407_n N_VGND_c_408_n N_VGND_c_409_n N_VGND_c_410_n
+ N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n VGND N_VGND_c_414_n
+ N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n N_VGND_c_418_n
+ PM_SKY130_FD_SC_HDLL__OR4B_1%VGND
cc_1 VNB N_D_N_M1000_g 0.0353378f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB D_N 0.0257888f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_N_c_73_n 0.0432637f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_117_297#_M1001_g 0.0341488f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_5 VNB N_A_117_297#_c_98_n 0.0142777f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_6 VNB N_A_117_297#_c_99_n 0.0127075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_297#_c_100_n 0.0388177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_C_c_138_n 0.0200253f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_C_M1008_g 0.0263738f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_10 VNB C 0.00754447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_174_n 0.00674306f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_B_c_175_n 0.0235704f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_13 VNB N_B_c_176_n 0.0144642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_c_216_n 0.0193174f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_15 VNB N_A_M1003_g 0.0282089f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_16 VNB N_A_c_218_n 0.00548445f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_17 VNB N_A_225_297#_c_254_n 0.0242891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_297#_c_255_n 0.0209439f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_19 VNB N_A_225_297#_c_256_n 0.00554352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_297#_c_257_n 0.00342296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_225_297#_c_258_n 0.00145828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_225_297#_c_259_n 0.00206408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_225_297#_c_260_n 0.00209425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_225_297#_c_261_n 0.00184153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_348_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_389_n 0.0163908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_390_n 0.0276689f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_VGND_c_407_n 0.0114258f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_29 VNB N_VGND_c_408_n 0.0197154f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_30 VNB N_VGND_c_409_n 0.0188657f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=0.85
cc_31 VNB N_VGND_c_410_n 0.00877358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_411_n 0.0158321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_412_n 8.39112e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_413_n 0.0129653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_414_n 0.0236453f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_415_n 0.243934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_416_n 0.00632108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_417_n 0.00544933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_418_n 0.0102719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_D_N_c_74_n 0.0241214f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB D_N 0.00399928f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_42 VPB N_D_N_c_73_n 0.0189781f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_43 VPB N_A_117_297#_c_101_n 0.0197389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_117_297#_c_102_n 0.0121629f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_45 VPB N_A_117_297#_c_99_n 0.00828518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_117_297#_c_100_n 0.0156292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_C_c_138_n 0.0232713f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB C 0.00185559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_B_c_177_n 0.00573755f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_50 VPB N_B_c_178_n 0.0501192f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_51 VPB N_B_M1005_g 0.0107552f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_52 VPB N_B_c_180_n 0.0595604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_c_216_n 0.0270354f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_A_c_218_n 0.00209843f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_55 VPB N_A_225_297#_c_254_n 0.0323205f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_225_297#_c_263_n 0.00630299f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_57 VPB N_A_225_297#_c_264_n 0.00158307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_225_297#_c_265_n 0.00754111f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_225_297#_c_266_n 0.00139551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_349_n 0.0114263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_350_n 0.0551265f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_62 VPB N_VPWR_c_351_n 0.0115426f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_63 VPB N_VPWR_c_352_n 0.0655885f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_64 VPB N_VPWR_c_353_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=0.85
cc_65 VPB N_VPWR_c_354_n 0.0234554f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_348_n 0.0759838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_X_c_391_n 0.00810971f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_68 VPB N_X_c_390_n 0.00992963f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_69 VPB X 0.0349983f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_70 N_D_N_M1000_g N_A_117_297#_c_98_n 0.00836126f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_71 D_N N_A_117_297#_c_98_n 0.0163351f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_72 N_D_N_c_74_n N_A_117_297#_c_102_n 0.00709049f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_D_N_c_73_n N_A_117_297#_c_102_n 0.00356719f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_74 D_N N_A_117_297#_c_99_n 0.0227733f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_75 N_D_N_c_73_n N_A_117_297#_c_99_n 0.00449331f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_76 N_D_N_c_73_n N_A_117_297#_c_100_n 0.00639522f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_77 N_D_N_c_74_n N_A_225_297#_c_265_n 0.00127278f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_78 N_D_N_c_74_n N_VPWR_c_350_n 0.0121354f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_79 D_N N_VPWR_c_350_n 0.0207642f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_80 N_D_N_c_73_n N_VPWR_c_350_n 0.00203685f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_81 N_D_N_c_74_n N_VPWR_c_352_n 0.00349149f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_D_N_c_74_n N_VPWR_c_348_n 0.00448105f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_D_N_M1000_g N_VGND_c_408_n 0.00432572f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_84 D_N N_VGND_c_408_n 0.0280862f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_85 N_D_N_c_73_n N_VGND_c_408_n 0.001395f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_86 N_D_N_M1000_g N_VGND_c_409_n 0.00555245f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_87 N_D_N_M1000_g N_VGND_c_410_n 0.00263598f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_88 N_D_N_M1000_g N_VGND_c_415_n 0.0121732f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_89 D_N N_VGND_c_415_n 0.00136771f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_117_297#_c_101_n N_C_c_138_n 0.0236423f $X=1.485 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_117_297#_c_99_n N_C_c_138_n 2.18501e-19 $X=1.215 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_117_297#_c_100_n N_C_c_138_n 0.0240795f $X=1.485 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_117_297#_M1001_g N_C_M1008_g 0.0166579f $X=1.51 $Y=0.475 $X2=0 $Y2=0
cc_94 N_A_117_297#_c_101_n C 0.00308949f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_117_297#_c_99_n C 0.0181267f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_117_297#_c_100_n C 0.00663347f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_97 N_A_117_297#_c_101_n N_B_c_180_n 0.00528936f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_117_297#_c_102_n N_B_c_180_n 0.0162027f $X=0.73 $Y=1.72 $X2=0 $Y2=0
cc_99 N_A_117_297#_c_101_n N_A_225_297#_c_263_n 0.014523f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_100 N_A_117_297#_M1001_g N_A_225_297#_c_257_n 0.00532403f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_101 N_A_117_297#_c_101_n N_A_225_297#_c_265_n 0.00645992f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_102 N_A_117_297#_c_102_n N_A_225_297#_c_265_n 0.0313055f $X=0.73 $Y=1.72
+ $X2=0 $Y2=0
cc_103 N_A_117_297#_c_99_n N_A_225_297#_c_265_n 0.0176028f $X=1.215 $Y=1.16
+ $X2=0 $Y2=0
cc_104 N_A_117_297#_c_100_n N_A_225_297#_c_265_n 0.00758805f $X=1.485 $Y=1.202
+ $X2=0 $Y2=0
cc_105 N_A_117_297#_c_102_n N_VPWR_c_350_n 0.0224405f $X=0.73 $Y=1.72 $X2=0
+ $Y2=0
cc_106 N_A_117_297#_c_102_n N_VPWR_c_348_n 0.00106784f $X=0.73 $Y=1.72 $X2=0
+ $Y2=0
cc_107 N_A_117_297#_c_98_n N_VGND_c_409_n 0.0128191f $X=0.73 $Y=0.5 $X2=0 $Y2=0
cc_108 N_A_117_297#_M1001_g N_VGND_c_410_n 0.0042334f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_109 N_A_117_297#_c_98_n N_VGND_c_410_n 0.0207056f $X=0.73 $Y=0.5 $X2=0 $Y2=0
cc_110 N_A_117_297#_c_99_n N_VGND_c_410_n 0.00902763f $X=1.215 $Y=1.16 $X2=0
+ $Y2=0
cc_111 N_A_117_297#_c_100_n N_VGND_c_410_n 0.00756977f $X=1.485 $Y=1.202 $X2=0
+ $Y2=0
cc_112 N_A_117_297#_M1001_g N_VGND_c_411_n 0.00555245f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_113 N_A_117_297#_M1001_g N_VGND_c_412_n 5.74535e-19 $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_114 N_A_117_297#_M1001_g N_VGND_c_415_n 0.0115458f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_115 N_A_117_297#_c_98_n N_VGND_c_415_n 0.00912835f $X=0.73 $Y=0.5 $X2=0 $Y2=0
cc_116 N_C_M1008_g N_B_c_174_n 0.0181868f $X=2.015 $Y=0.475 $X2=-0.19 $Y2=-0.24
cc_117 N_C_c_138_n N_B_c_175_n 0.0181868f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_118 C N_B_c_175_n 0.00941954f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_119 C N_B_c_177_n 0.00354894f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_120 N_C_c_138_n N_B_M1005_g 0.0319112f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_121 C N_B_M1005_g 0.00726812f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_122 N_C_M1008_g N_B_c_176_n 0.0125555f $X=2.015 $Y=0.475 $X2=0 $Y2=0
cc_123 N_C_c_138_n N_B_c_180_n 0.00527095f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_124 C N_A_c_216_n 0.00122619f $X=2.135 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_125 C N_A_c_218_n 0.0232376f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_126 N_C_c_138_n N_A_225_297#_c_263_n 0.0109699f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_127 C N_A_225_297#_c_263_n 0.0474955f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_128 N_C_c_138_n N_A_225_297#_c_256_n 0.00252042f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C_M1008_g N_A_225_297#_c_256_n 0.0108447f $X=2.015 $Y=0.475 $X2=0 $Y2=0
cc_130 C N_A_225_297#_c_256_n 0.0455778f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_131 N_C_c_138_n N_A_225_297#_c_257_n 9.23324e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_132 C N_A_225_297#_c_257_n 0.0152593f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_133 N_C_c_138_n N_A_225_297#_c_265_n 9.19411e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_134 C N_A_225_297#_c_266_n 0.00635864f $X=2.135 $Y=1.105 $X2=0 $Y2=0
cc_135 C A_315_297# 0.00278453f $X=2.135 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_136 C A_416_297# 0.00161889f $X=2.135 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_137 N_C_M1008_g N_VGND_c_411_n 0.00187556f $X=2.015 $Y=0.475 $X2=0 $Y2=0
cc_138 N_C_M1008_g N_VGND_c_412_n 0.0100346f $X=2.015 $Y=0.475 $X2=0 $Y2=0
cc_139 N_C_M1008_g N_VGND_c_415_n 0.00267543f $X=2.015 $Y=0.475 $X2=0 $Y2=0
cc_140 N_B_c_175_n N_A_c_216_n 0.0180423f $X=2.43 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_141 N_B_c_177_n N_A_c_216_n 0.00376819f $X=2.43 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_142 N_B_M1005_g N_A_c_216_n 0.0231537f $X=2.43 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_143 N_B_c_180_n N_A_c_216_n 6.03833e-19 $X=2.47 $Y=2.31 $X2=-0.19 $Y2=-0.24
cc_144 N_B_c_176_n N_A_M1003_g 0.0177253f $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_145 N_B_c_175_n N_A_c_218_n 0.00240539f $X=2.43 $Y=1.31 $X2=0 $Y2=0
cc_146 N_B_c_178_n N_A_225_297#_c_263_n 7.51174e-19 $X=2.43 $Y=2.035 $X2=0 $Y2=0
cc_147 N_B_M1005_g N_A_225_297#_c_263_n 0.0144447f $X=2.43 $Y=1.695 $X2=0 $Y2=0
cc_148 N_B_c_180_n N_A_225_297#_c_263_n 0.0953992f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_149 N_B_c_174_n N_A_225_297#_c_256_n 0.0099557f $X=2.43 $Y=0.86 $X2=0 $Y2=0
cc_150 N_B_c_176_n N_A_225_297#_c_256_n 0.00734988f $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_151 N_B_c_180_n N_A_225_297#_c_265_n 0.0261176f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_152 N_B_M1005_g N_A_225_297#_c_266_n 0.00471908f $X=2.43 $Y=1.695 $X2=0 $Y2=0
cc_153 N_B_c_180_n N_A_225_297#_c_266_n 0.0137296f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_154 N_B_c_180_n N_VPWR_c_350_n 0.020342f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_155 N_B_c_178_n N_VPWR_c_351_n 0.00520464f $X=2.43 $Y=2.035 $X2=0 $Y2=0
cc_156 N_B_c_180_n N_VPWR_c_351_n 0.0210034f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_157 N_B_c_178_n N_VPWR_c_352_n 0.00698479f $X=2.43 $Y=2.035 $X2=0 $Y2=0
cc_158 N_B_c_180_n N_VPWR_c_352_n 0.111255f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_159 N_B_c_178_n N_VPWR_c_348_n 0.00955749f $X=2.43 $Y=2.035 $X2=0 $Y2=0
cc_160 N_B_c_180_n N_VPWR_c_348_n 0.0803497f $X=2.47 $Y=2.31 $X2=0 $Y2=0
cc_161 N_B_c_176_n N_VGND_c_412_n 0.00613475f $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_162 N_B_c_176_n N_VGND_c_413_n 0.00375785f $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_163 N_B_c_176_n N_VGND_c_415_n 0.00463104f $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_164 N_B_c_176_n N_VGND_c_418_n 5.6593e-19 $X=2.43 $Y=0.76 $X2=0 $Y2=0
cc_165 N_A_c_216_n N_A_225_297#_c_254_n 0.0349746f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_218_n N_A_225_297#_c_254_n 0.00107624f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_M1003_g N_A_225_297#_c_255_n 0.0175774f $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_168 N_A_c_216_n N_A_225_297#_c_263_n 2.06235e-19 $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_218_n N_A_225_297#_c_263_n 0.00230038f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_216_n N_A_225_297#_c_258_n 0.00240831f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_M1003_g N_A_225_297#_c_258_n 0.0116486f $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_172 N_A_c_218_n N_A_225_297#_c_258_n 0.0217578f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_c_216_n N_A_225_297#_c_299_n 0.0141303f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_218_n N_A_225_297#_c_299_n 0.0136748f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_c_216_n N_A_225_297#_c_264_n 0.00170148f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_216_n N_A_225_297#_c_259_n 5.77159e-19 $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_218_n N_A_225_297#_c_259_n 0.0128912f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_216_n N_A_225_297#_c_266_n 0.0111966f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_218_n N_A_225_297#_c_266_n 0.0112473f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_c_216_n N_A_225_297#_c_260_n 0.00444957f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_218_n N_A_225_297#_c_260_n 0.0275754f $X=2.89 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_M1003_g N_A_225_297#_c_261_n 0.00174468f $X=2.955 $Y=0.475 $X2=0
+ $Y2=0
cc_183 N_A_c_216_n N_VPWR_c_351_n 0.00330158f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_216_n N_VPWR_c_352_n 0.00351268f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_216_n N_VPWR_c_348_n 0.00445321f $X=2.93 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_M1003_g N_VGND_c_412_n 4.90246e-19 $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_187 N_A_M1003_g N_VGND_c_413_n 0.00188229f $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_188 N_A_M1003_g N_VGND_c_415_n 0.00266683f $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_189 N_A_M1003_g N_VGND_c_418_n 0.0100988f $X=2.955 $Y=0.475 $X2=0 $Y2=0
cc_190 N_A_225_297#_c_299_n N_VPWR_M1007_d 0.00593118f $X=3.245 $Y=1.58 $X2=0
+ $Y2=0
cc_191 N_A_225_297#_c_265_n N_VPWR_c_350_n 9.92714e-19 $X=1.25 $Y=1.685 $X2=0
+ $Y2=0
cc_192 N_A_225_297#_c_254_n N_VPWR_c_351_n 0.00505337f $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_225_297#_c_299_n N_VPWR_c_351_n 0.0202939f $X=3.245 $Y=1.58 $X2=0
+ $Y2=0
cc_194 N_A_225_297#_c_266_n N_VPWR_c_351_n 0.00726621f $X=2.775 $Y=1.58 $X2=0
+ $Y2=0
cc_195 N_A_225_297#_c_254_n N_VPWR_c_354_n 0.00702461f $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_225_297#_c_254_n N_VPWR_c_348_n 0.0148476f $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_225_297#_c_263_n A_315_297# 0.00218559f $X=2.69 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_198 N_A_225_297#_c_263_n A_416_297# 0.00155579f $X=2.69 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_199 N_A_225_297#_c_263_n A_504_297# 0.00334472f $X=2.69 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_200 N_A_225_297#_c_266_n A_504_297# 0.00441537f $X=2.775 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_201 N_A_225_297#_c_254_n N_X_c_391_n 0.0124367f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_225_297#_c_299_n N_X_c_391_n 0.0120449f $X=3.245 $Y=1.58 $X2=0 $Y2=0
cc_203 N_A_225_297#_c_254_n N_X_c_390_n 7.5048e-19 $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_225_297#_c_255_n N_X_c_390_n 0.0134968f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A_225_297#_c_264_n N_X_c_390_n 0.00566258f $X=3.33 $Y=1.495 $X2=0 $Y2=0
cc_206 N_A_225_297#_c_260_n N_X_c_390_n 0.0208334f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_225_297#_c_261_n N_X_c_390_n 0.00709789f $X=3.375 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_225_297#_c_256_n N_VGND_M1008_d 0.00180643f $X=2.61 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_225_297#_c_258_n N_VGND_M1003_d 0.00700166f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_210 N_A_225_297#_c_261_n N_VGND_M1003_d 7.06785e-19 $X=3.375 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_225_297#_c_330_p N_VGND_c_411_n 0.00876148f $X=1.75 $Y=0.47 $X2=0
+ $Y2=0
cc_212 N_A_225_297#_c_256_n N_VGND_c_411_n 0.00240437f $X=2.61 $Y=0.74 $X2=0
+ $Y2=0
cc_213 N_A_225_297#_c_330_p N_VGND_c_412_n 0.0131398f $X=1.75 $Y=0.47 $X2=0
+ $Y2=0
cc_214 N_A_225_297#_c_256_n N_VGND_c_412_n 0.0197523f $X=2.61 $Y=0.74 $X2=0
+ $Y2=0
cc_215 N_A_225_297#_c_334_p N_VGND_c_412_n 0.0110176f $X=2.695 $Y=0.47 $X2=0
+ $Y2=0
cc_216 N_A_225_297#_c_256_n N_VGND_c_413_n 0.00307941f $X=2.61 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A_225_297#_c_334_p N_VGND_c_413_n 0.00876148f $X=2.695 $Y=0.47 $X2=0
+ $Y2=0
cc_218 N_A_225_297#_c_258_n N_VGND_c_413_n 0.00232988f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_219 N_A_225_297#_c_255_n N_VGND_c_414_n 0.00585385f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_225_297#_c_255_n N_VGND_c_415_n 0.0123336f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_225_297#_c_330_p N_VGND_c_415_n 0.00625722f $X=1.75 $Y=0.47 $X2=0
+ $Y2=0
cc_222 N_A_225_297#_c_256_n N_VGND_c_415_n 0.0115926f $X=2.61 $Y=0.74 $X2=0
+ $Y2=0
cc_223 N_A_225_297#_c_334_p N_VGND_c_415_n 0.00625722f $X=2.695 $Y=0.47 $X2=0
+ $Y2=0
cc_224 N_A_225_297#_c_258_n N_VGND_c_415_n 0.0073302f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_225 N_A_225_297#_c_254_n N_VGND_c_418_n 3.3049e-19 $X=3.47 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_225_297#_c_255_n N_VGND_c_418_n 0.00498808f $X=3.495 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_225_297#_c_334_p N_VGND_c_418_n 0.0135697f $X=2.695 $Y=0.47 $X2=0
+ $Y2=0
cc_228 N_A_225_297#_c_258_n N_VGND_c_418_n 0.0277382f $X=3.245 $Y=0.74 $X2=0
+ $Y2=0
cc_229 N_VPWR_c_348_n N_X_M1011_d 0.00442383f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_230 N_VPWR_c_354_n X 0.0264344f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_348_n X 0.0143649f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_232 N_X_c_389_n N_VGND_c_414_n 0.0127126f $X=3.705 $Y=0.59 $X2=0 $Y2=0
cc_233 N_X_M1002_d N_VGND_c_415_n 0.00419212f $X=3.57 $Y=0.235 $X2=0 $Y2=0
cc_234 N_X_c_389_n N_VGND_c_415_n 0.0130147f $X=3.705 $Y=0.59 $X2=0 $Y2=0
