* File: sky130_fd_sc_hdll__ebufn_8.pxi.spice
* Created: Wed Sep  2 08:30:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%A N_A_c_137_n N_A_M1005_g N_A_c_133_n
+ N_A_M1013_g N_A_c_138_n N_A_M1033_g N_A_M1026_g A A N_A_c_136_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_8%A
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%TE_B N_TE_B_c_177_n N_TE_B_M1007_g
+ N_TE_B_c_182_n N_TE_B_M1014_g N_TE_B_c_178_n N_TE_B_c_184_n N_TE_B_c_185_n
+ N_TE_B_M1000_g N_TE_B_c_186_n N_TE_B_c_187_n N_TE_B_M1001_g N_TE_B_c_188_n
+ N_TE_B_c_189_n N_TE_B_M1002_g N_TE_B_c_190_n N_TE_B_c_191_n N_TE_B_M1003_g
+ N_TE_B_c_192_n N_TE_B_c_193_n N_TE_B_M1006_g N_TE_B_c_194_n N_TE_B_c_195_n
+ N_TE_B_M1012_g N_TE_B_c_196_n N_TE_B_c_197_n N_TE_B_M1016_g N_TE_B_c_198_n
+ N_TE_B_c_199_n N_TE_B_M1021_g N_TE_B_c_179_n N_TE_B_c_180_n N_TE_B_c_202_n
+ N_TE_B_c_203_n N_TE_B_c_204_n N_TE_B_c_205_n N_TE_B_c_206_n N_TE_B_c_207_n
+ N_TE_B_c_208_n TE_B TE_B PM_SKY130_FD_SC_HDLL__EBUFN_8%TE_B
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%A_321_47# N_A_321_47#_M1007_d
+ N_A_321_47#_M1014_d N_A_321_47#_c_351_n N_A_321_47#_M1009_g
+ N_A_321_47#_c_352_n N_A_321_47#_c_353_n N_A_321_47#_c_354_n
+ N_A_321_47#_M1010_g N_A_321_47#_c_355_n N_A_321_47#_c_356_n
+ N_A_321_47#_M1018_g N_A_321_47#_c_357_n N_A_321_47#_c_358_n
+ N_A_321_47#_M1019_g N_A_321_47#_c_359_n N_A_321_47#_c_360_n
+ N_A_321_47#_M1022_g N_A_321_47#_c_361_n N_A_321_47#_c_362_n
+ N_A_321_47#_M1032_g N_A_321_47#_c_363_n N_A_321_47#_c_364_n
+ N_A_321_47#_M1034_g N_A_321_47#_c_365_n N_A_321_47#_c_366_n
+ N_A_321_47#_M1036_g N_A_321_47#_c_367_n N_A_321_47#_c_368_n
+ N_A_321_47#_c_369_n N_A_321_47#_c_370_n N_A_321_47#_c_371_n
+ N_A_321_47#_c_372_n N_A_321_47#_c_373_n N_A_321_47#_c_378_n
+ N_A_321_47#_c_374_n N_A_321_47#_c_375_n N_A_321_47#_c_376_n
+ N_A_321_47#_c_377_n N_A_321_47#_c_379_n N_A_321_47#_c_380_n
+ N_A_321_47#_c_416_n PM_SKY130_FD_SC_HDLL__EBUFN_8%A_321_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%A_124_297# N_A_124_297#_M1013_d
+ N_A_124_297#_M1005_s N_A_124_297#_M1004_g N_A_124_297#_c_519_n
+ N_A_124_297#_M1008_g N_A_124_297#_M1011_g N_A_124_297#_c_520_n
+ N_A_124_297#_M1015_g N_A_124_297#_M1023_g N_A_124_297#_c_521_n
+ N_A_124_297#_M1017_g N_A_124_297#_M1024_g N_A_124_297#_c_522_n
+ N_A_124_297#_M1020_g N_A_124_297#_M1025_g N_A_124_297#_c_523_n
+ N_A_124_297#_M1028_g N_A_124_297#_M1027_g N_A_124_297#_c_524_n
+ N_A_124_297#_M1030_g N_A_124_297#_M1029_g N_A_124_297#_c_525_n
+ N_A_124_297#_M1031_g N_A_124_297#_c_526_n N_A_124_297#_M1035_g
+ N_A_124_297#_M1037_g N_A_124_297#_c_554_p N_A_124_297#_c_529_n
+ N_A_124_297#_c_591_p N_A_124_297#_c_516_n N_A_124_297#_c_551_n
+ N_A_124_297#_c_517_n N_A_124_297#_c_518_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_8%A_124_297#
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%VPWR N_VPWR_M1005_d N_VPWR_M1033_d
+ N_VPWR_M1000_d N_VPWR_M1002_d N_VPWR_M1006_d N_VPWR_M1016_d N_VPWR_c_647_n
+ N_VPWR_c_648_n N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_651_n N_VPWR_c_652_n
+ VPWR N_VPWR_c_653_n N_VPWR_c_654_n N_VPWR_c_655_n N_VPWR_c_656_n
+ N_VPWR_c_646_n N_VPWR_c_658_n N_VPWR_c_659_n N_VPWR_c_660_n N_VPWR_c_661_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_8%VPWR
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%A_437_309# N_A_437_309#_M1000_s
+ N_A_437_309#_M1001_s N_A_437_309#_M1003_s N_A_437_309#_M1012_s
+ N_A_437_309#_M1021_s N_A_437_309#_M1015_d N_A_437_309#_M1020_d
+ N_A_437_309#_M1030_d N_A_437_309#_M1035_d N_A_437_309#_c_789_n
+ N_A_437_309#_c_793_n N_A_437_309#_c_790_n N_A_437_309#_c_797_n
+ N_A_437_309#_c_799_n N_A_437_309#_c_802_n N_A_437_309#_c_804_n
+ N_A_437_309#_c_807_n N_A_437_309#_c_809_n N_A_437_309#_c_791_n
+ N_A_437_309#_c_810_n N_A_437_309#_c_811_n N_A_437_309#_c_812_n
+ N_A_437_309#_c_813_n PM_SKY130_FD_SC_HDLL__EBUFN_8%A_437_309#
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%Z N_Z_M1004_s N_Z_M1023_s N_Z_M1025_s
+ N_Z_M1029_s N_Z_M1008_s N_Z_M1017_s N_Z_M1028_s N_Z_M1031_s N_Z_c_930_n Z Z Z
+ Z Z Z Z Z Z Z Z Z Z Z Z Z Z N_Z_c_900_n Z Z Z Z Z Z Z Z Z Z Z Z N_Z_c_897_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_8%Z
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%VGND N_VGND_M1013_s N_VGND_M1026_s
+ N_VGND_M1009_s N_VGND_M1018_s N_VGND_M1022_s N_VGND_M1034_s N_VGND_c_1004_n
+ N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n N_VGND_c_1008_n VGND
+ N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n N_VGND_c_1012_n
+ N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n N_VGND_c_1016_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_8%VGND
x_PM_SKY130_FD_SC_HDLL__EBUFN_8%A_485_47# N_A_485_47#_M1009_d
+ N_A_485_47#_M1010_d N_A_485_47#_M1019_d N_A_485_47#_M1032_d
+ N_A_485_47#_M1036_d N_A_485_47#_M1011_d N_A_485_47#_M1024_d
+ N_A_485_47#_M1027_d N_A_485_47#_M1037_d N_A_485_47#_c_1132_n
+ N_A_485_47#_c_1137_n N_A_485_47#_c_1133_n N_A_485_47#_c_1144_n
+ N_A_485_47#_c_1145_n N_A_485_47#_c_1150_n N_A_485_47#_c_1151_n
+ N_A_485_47#_c_1156_n N_A_485_47#_c_1157_n N_A_485_47#_c_1134_n
+ N_A_485_47#_c_1162_n N_A_485_47#_c_1164_n N_A_485_47#_c_1166_n
+ N_A_485_47#_c_1168_n PM_SKY130_FD_SC_HDLL__EBUFN_8%A_485_47#
cc_1 VNB N_A_c_133_n 0.0224185f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_A_M1026_g 0.0175938f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_3 VNB A 0.0148258f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_c_136_n 0.065476f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_5 VNB N_TE_B_c_177_n 0.0201845f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.41
cc_6 VNB N_TE_B_c_178_n 0.0199077f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_7 VNB N_TE_B_c_179_n 0.0249493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_TE_B_c_180_n 0.0203092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB TE_B 0.00267876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_321_47#_c_351_n 0.0184787f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.41
cc_11 VNB N_A_321_47#_c_352_n 0.0137076f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=1.025
cc_12 VNB N_A_321_47#_c_353_n 0.00771506f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_13 VNB N_A_321_47#_c_354_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_14 VNB N_A_321_47#_c_355_n 0.0137061f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_15 VNB N_A_321_47#_c_356_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_321_47#_c_357_n 0.0137076f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_17 VNB N_A_321_47#_c_358_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.202
cc_18 VNB N_A_321_47#_c_359_n 0.0137061f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_19 VNB N_A_321_47#_c_360_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_321_47#_c_361_n 0.0137076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_321_47#_c_362_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_321_47#_c_363_n 0.0137061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_321_47#_c_364_n 0.0155949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_321_47#_c_365_n 0.0153441f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_321_47#_c_366_n 0.0169495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_321_47#_c_367_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_321_47#_c_368_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_321_47#_c_369_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_321_47#_c_370_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_321_47#_c_371_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_321_47#_c_372_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_321_47#_c_373_n 0.0129526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_321_47#_c_374_n 0.0032241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_321_47#_c_375_n 0.0354407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_321_47#_c_376_n 0.0332203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_321_47#_c_377_n 0.0104843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_124_297#_M1004_g 0.0202161f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.985
cc_38 VNB N_A_124_297#_M1011_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_124_297#_M1023_g 0.018595f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_40 VNB N_A_124_297#_M1024_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_124_297#_M1025_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_124_297#_M1027_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_124_297#_M1029_g 0.01909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_124_297#_M1037_g 0.0218603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_124_297#_c_516_n 0.00496447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_124_297#_c_517_n 0.186296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_124_297#_c_518_n 0.00213216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VPWR_c_646_n 0.459507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB Z 0.0226184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Z_c_897_n 0.010637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1004_n 0.0118369f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_52 VNB N_VGND_c_1005_n 0.0287663f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.202
cc_53 VNB N_VGND_c_1006_n 0.013643f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_54 VNB N_VGND_c_1007_n 0.00617769f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.16
cc_55 VNB N_VGND_c_1008_n 0.0135644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1009_n 0.0240083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1010_n 0.0354185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1011_n 0.013643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1012_n 0.106153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1013_n 0.515562f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1014_n 0.006263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1015_n 0.00617769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1016_n 0.006263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_485_47#_c_1132_n 0.00633746f $X=-0.19 $Y=-0.24 $X2=0.257 $Y2=1.53
cc_65 VNB N_A_485_47#_c_1133_n 0.00316415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_485_47#_c_1134_n 0.00882053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VPB N_A_c_137_n 0.018233f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.41
cc_68 VPB N_A_c_138_n 0.0160851f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_69 VPB A 0.0132795f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_70 VPB N_A_c_136_n 0.0219139f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.202
cc_71 VPB N_TE_B_c_182_n 0.01994f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_72 VPB N_TE_B_c_178_n 0.0113386f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_73 VPB N_TE_B_c_184_n 0.0153293f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.985
cc_74 VPB N_TE_B_c_185_n 0.0192205f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_75 VPB N_TE_B_c_186_n 0.0163203f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_76 VPB N_TE_B_c_187_n 0.0162041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_TE_B_c_188_n 0.0155544f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_78 VPB N_TE_B_c_189_n 0.0159249f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_79 VPB N_TE_B_c_190_n 0.0155544f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=1.202
cc_80 VPB N_TE_B_c_191_n 0.0162041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_TE_B_c_192_n 0.0155544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_TE_B_c_193_n 0.0159249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_TE_B_c_194_n 0.0155544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_TE_B_c_195_n 0.0162041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_TE_B_c_196_n 0.0155544f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_TE_B_c_197_n 0.0159249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_TE_B_c_198_n 0.0297161f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_TE_B_c_199_n 0.0194998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_TE_B_c_179_n 0.0143708f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_TE_B_c_180_n 0.0127657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_TE_B_c_202_n 0.00735165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_TE_B_c_203_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_TE_B_c_204_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_TE_B_c_205_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_TE_B_c_206_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_TE_B_c_207_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_TE_B_c_208_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB TE_B 0.00306059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_321_47#_c_378_n 0.00878946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_321_47#_c_379_n 0.00180385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_321_47#_c_380_n 0.002661f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_124_297#_c_519_n 0.0201091f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_103 VPB N_A_124_297#_c_520_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.202
cc_104 VPB N_A_124_297#_c_521_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_105 VPB N_A_124_297#_c_522_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_124_297#_c_523_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_A_124_297#_c_524_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_124_297#_c_525_n 0.0158723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_124_297#_c_526_n 0.0191743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_124_297#_c_517_n 0.0542821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_124_297#_c_518_n 0.00223368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_647_n 0.0107162f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_113 VPB N_VPWR_c_648_n 0.0310119f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_114 VPB N_VPWR_c_649_n 0.00277705f $X=-0.19 $Y=1.305 $X2=0.257 $Y2=1.16
cc_115 VPB N_VPWR_c_650_n 0.0138213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_651_n 0.00614834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_652_n 0.0288739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_653_n 0.0144188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_654_n 0.0138213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_655_n 0.0138213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_VPWR_c_656_n 0.112673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_646_n 0.0540829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_658_n 0.0058967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_VPWR_c_659_n 0.00606303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_660_n 0.00606303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_661_n 0.00614834f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_437_309#_c_789_n 0.00373697f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_437_309#_c_790_n 0.00177027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_437_309#_c_791_n 0.0249987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB Z 0.00715958f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB Z 0.0125444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_Z_c_900_n 0.0215737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 N_A_M1026_g N_TE_B_c_177_n 0.0218642f $X=1.025 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_c_138_n N_TE_B_c_182_n 0.0237928f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_M1026_g N_TE_B_c_178_n 0.0215243f $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_136 N_A_c_136_n N_TE_B_c_178_n 0.00249401f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_c_138_n TE_B 0.00860187f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_M1026_g TE_B 0.0116025f $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_139 N_A_c_136_n TE_B 0.0106198f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A_c_138_n N_A_321_47#_c_378_n 7.25712e-19 $X=1 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_M1026_g N_A_321_47#_c_377_n 7.0951e-19 $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_142 A N_A_124_297#_c_529_n 0.00702447f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_c_136_n N_A_124_297#_c_529_n 0.0144629f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_144 N_A_c_136_n N_A_124_297#_c_516_n 0.0108804f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_145 N_A_c_137_n N_A_124_297#_c_518_n 0.00125661f $X=0.53 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_133_n N_A_124_297#_c_518_n 0.00442767f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_c_138_n N_A_124_297#_c_518_n 0.00884396f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_M1026_g N_A_124_297#_c_518_n 0.00654752f $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_149 A N_A_124_297#_c_518_n 0.0273981f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_c_136_n N_A_124_297#_c_518_n 0.0199975f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_151 A N_VPWR_M1005_d 0.00417858f $X=0.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_152 N_A_c_137_n N_VPWR_c_648_n 0.01278f $X=0.53 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_138_n N_VPWR_c_648_n 6.57033e-19 $X=1 $Y=1.41 $X2=0 $Y2=0
cc_154 A N_VPWR_c_648_n 0.0267675f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A_c_136_n N_VPWR_c_648_n 0.00105323f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_c_137_n N_VPWR_c_649_n 6.97267e-19 $X=0.53 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_138_n N_VPWR_c_649_n 0.0149638f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_137_n N_VPWR_c_653_n 0.00681171f $X=0.53 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_138_n N_VPWR_c_653_n 0.00427505f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_137_n N_VPWR_c_646_n 0.0114004f $X=0.53 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_138_n N_VPWR_c_646_n 0.00740765f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_133_n N_VGND_c_1005_n 0.0147806f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_163 A N_VGND_c_1005_n 0.029924f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A_c_136_n N_VGND_c_1005_n 0.00211088f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_c_133_n N_VGND_c_1009_n 0.00646692f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_M1026_g N_VGND_c_1009_n 0.0124143f $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_167 N_A_c_133_n N_VGND_c_1013_n 0.0118487f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_M1026_g N_VGND_c_1013_n 0.00510095f $X=1.025 $Y=0.56 $X2=0 $Y2=0
cc_169 N_TE_B_c_203_n N_A_321_47#_c_352_n 0.0172028f $X=3.065 $Y=1.395 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_186_n N_A_321_47#_c_353_n 0.0172028f $X=2.975 $Y=1.395 $X2=0
+ $Y2=0
cc_171 N_TE_B_c_180_n N_A_321_47#_c_353_n 0.00251242f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_172 N_TE_B_c_204_n N_A_321_47#_c_355_n 0.0172028f $X=3.585 $Y=1.395 $X2=0
+ $Y2=0
cc_173 N_TE_B_c_205_n N_A_321_47#_c_357_n 0.0172028f $X=4.105 $Y=1.395 $X2=0
+ $Y2=0
cc_174 N_TE_B_c_206_n N_A_321_47#_c_359_n 0.0172028f $X=4.625 $Y=1.395 $X2=0
+ $Y2=0
cc_175 N_TE_B_c_207_n N_A_321_47#_c_361_n 0.0172028f $X=5.145 $Y=1.395 $X2=0
+ $Y2=0
cc_176 N_TE_B_c_208_n N_A_321_47#_c_363_n 0.0172028f $X=5.665 $Y=1.395 $X2=0
+ $Y2=0
cc_177 N_TE_B_c_188_n N_A_321_47#_c_367_n 0.0172028f $X=3.495 $Y=1.395 $X2=0
+ $Y2=0
cc_178 N_TE_B_c_190_n N_A_321_47#_c_368_n 0.0172028f $X=4.015 $Y=1.395 $X2=0
+ $Y2=0
cc_179 N_TE_B_c_192_n N_A_321_47#_c_369_n 0.0172028f $X=4.535 $Y=1.395 $X2=0
+ $Y2=0
cc_180 N_TE_B_c_194_n N_A_321_47#_c_370_n 0.0172028f $X=5.055 $Y=1.395 $X2=0
+ $Y2=0
cc_181 N_TE_B_c_196_n N_A_321_47#_c_371_n 0.0172028f $X=5.575 $Y=1.395 $X2=0
+ $Y2=0
cc_182 N_TE_B_c_198_n N_A_321_47#_c_372_n 0.0172028f $X=6.095 $Y=1.395 $X2=0
+ $Y2=0
cc_183 N_TE_B_c_182_n N_A_321_47#_c_378_n 0.0130979f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_TE_B_c_185_n N_A_321_47#_c_378_n 0.0060647f $X=2.545 $Y=1.47 $X2=0
+ $Y2=0
cc_185 N_TE_B_c_177_n N_A_321_47#_c_374_n 0.00381839f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_TE_B_c_179_n N_A_321_47#_c_374_n 0.00915045f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_187 N_TE_B_c_180_n N_A_321_47#_c_374_n 0.00232001f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_188 TE_B N_A_321_47#_c_374_n 0.00904843f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_189 N_TE_B_c_184_n N_A_321_47#_c_375_n 0.0399692f $X=2.455 $Y=1.395 $X2=0
+ $Y2=0
cc_190 N_TE_B_c_180_n N_A_321_47#_c_375_n 0.0122741f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_191 N_TE_B_c_177_n N_A_321_47#_c_377_n 0.0129331f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_TE_B_c_178_n N_A_321_47#_c_377_n 0.00391179f $X=1.655 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_TE_B_c_182_n N_A_321_47#_c_379_n 0.00445914f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_TE_B_c_179_n N_A_321_47#_c_379_n 0.00237936f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_195 TE_B N_A_321_47#_c_379_n 0.0160149f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_196 N_TE_B_c_182_n N_A_321_47#_c_380_n 0.00103881f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_TE_B_c_178_n N_A_321_47#_c_380_n 9.2802e-19 $X=1.655 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_TE_B_c_185_n N_A_321_47#_c_380_n 9.78685e-19 $X=2.545 $Y=1.47 $X2=0
+ $Y2=0
cc_199 N_TE_B_c_179_n N_A_321_47#_c_380_n 0.00929198f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_200 N_TE_B_c_180_n N_A_321_47#_c_380_n 0.00363129f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_201 TE_B N_A_321_47#_c_380_n 0.0115235f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_202 N_TE_B_c_179_n N_A_321_47#_c_416_n 0.0147346f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_203 N_TE_B_c_180_n N_A_321_47#_c_416_n 0.00445721f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_204 TE_B N_A_321_47#_c_416_n 0.0143613f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_205 TE_B N_A_124_297#_c_529_n 0.00242116f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_206 N_TE_B_c_178_n N_A_124_297#_c_516_n 0.00540404f $X=1.655 $Y=1.16 $X2=0
+ $Y2=0
cc_207 N_TE_B_c_179_n N_A_124_297#_c_516_n 0.00162963f $X=2.07 $Y=1.232 $X2=0
+ $Y2=0
cc_208 TE_B N_A_124_297#_c_516_n 0.0484104f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_209 N_TE_B_c_178_n N_A_124_297#_c_518_n 2.12051e-19 $X=1.655 $Y=1.16 $X2=0
+ $Y2=0
cc_210 TE_B N_A_124_297#_c_518_n 0.0795932f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_211 TE_B N_VPWR_M1033_d 0.00589982f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_212 N_TE_B_c_182_n N_VPWR_c_649_n 0.00889037f $X=1.555 $Y=1.41 $X2=0 $Y2=0
cc_213 N_TE_B_c_178_n N_VPWR_c_649_n 3.44951e-19 $X=1.655 $Y=1.16 $X2=0 $Y2=0
cc_214 TE_B N_VPWR_c_649_n 0.0282994f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_215 N_TE_B_c_195_n N_VPWR_c_650_n 0.00456556f $X=5.145 $Y=1.47 $X2=0 $Y2=0
cc_216 N_TE_B_c_197_n N_VPWR_c_650_n 0.00313882f $X=5.665 $Y=1.47 $X2=0 $Y2=0
cc_217 N_TE_B_c_185_n N_VPWR_c_651_n 0.0115461f $X=2.545 $Y=1.47 $X2=0 $Y2=0
cc_218 N_TE_B_c_187_n N_VPWR_c_651_n 0.0073741f $X=3.065 $Y=1.47 $X2=0 $Y2=0
cc_219 N_TE_B_c_189_n N_VPWR_c_651_n 4.80713e-19 $X=3.585 $Y=1.47 $X2=0 $Y2=0
cc_220 N_TE_B_c_182_n N_VPWR_c_652_n 0.00597712f $X=1.555 $Y=1.41 $X2=0 $Y2=0
cc_221 N_TE_B_c_185_n N_VPWR_c_652_n 0.00313882f $X=2.545 $Y=1.47 $X2=0 $Y2=0
cc_222 N_TE_B_c_187_n N_VPWR_c_654_n 0.00456556f $X=3.065 $Y=1.47 $X2=0 $Y2=0
cc_223 N_TE_B_c_189_n N_VPWR_c_654_n 0.00313882f $X=3.585 $Y=1.47 $X2=0 $Y2=0
cc_224 N_TE_B_c_191_n N_VPWR_c_655_n 0.00456556f $X=4.105 $Y=1.47 $X2=0 $Y2=0
cc_225 N_TE_B_c_193_n N_VPWR_c_655_n 0.00313882f $X=4.625 $Y=1.47 $X2=0 $Y2=0
cc_226 N_TE_B_c_199_n N_VPWR_c_656_n 0.00456556f $X=6.185 $Y=1.47 $X2=0 $Y2=0
cc_227 N_TE_B_c_182_n N_VPWR_c_646_n 0.0115763f $X=1.555 $Y=1.41 $X2=0 $Y2=0
cc_228 N_TE_B_c_185_n N_VPWR_c_646_n 0.00502902f $X=2.545 $Y=1.47 $X2=0 $Y2=0
cc_229 N_TE_B_c_187_n N_VPWR_c_646_n 0.00531152f $X=3.065 $Y=1.47 $X2=0 $Y2=0
cc_230 N_TE_B_c_189_n N_VPWR_c_646_n 0.00386885f $X=3.585 $Y=1.47 $X2=0 $Y2=0
cc_231 N_TE_B_c_191_n N_VPWR_c_646_n 0.00531152f $X=4.105 $Y=1.47 $X2=0 $Y2=0
cc_232 N_TE_B_c_193_n N_VPWR_c_646_n 0.00386885f $X=4.625 $Y=1.47 $X2=0 $Y2=0
cc_233 N_TE_B_c_195_n N_VPWR_c_646_n 0.00531152f $X=5.145 $Y=1.47 $X2=0 $Y2=0
cc_234 N_TE_B_c_197_n N_VPWR_c_646_n 0.00386885f $X=5.665 $Y=1.47 $X2=0 $Y2=0
cc_235 N_TE_B_c_199_n N_VPWR_c_646_n 0.00656631f $X=6.185 $Y=1.47 $X2=0 $Y2=0
cc_236 N_TE_B_c_187_n N_VPWR_c_659_n 5.42676e-19 $X=3.065 $Y=1.47 $X2=0 $Y2=0
cc_237 N_TE_B_c_189_n N_VPWR_c_659_n 0.0103345f $X=3.585 $Y=1.47 $X2=0 $Y2=0
cc_238 N_TE_B_c_191_n N_VPWR_c_659_n 0.0073741f $X=4.105 $Y=1.47 $X2=0 $Y2=0
cc_239 N_TE_B_c_193_n N_VPWR_c_659_n 4.80713e-19 $X=4.625 $Y=1.47 $X2=0 $Y2=0
cc_240 N_TE_B_c_191_n N_VPWR_c_660_n 5.42676e-19 $X=4.105 $Y=1.47 $X2=0 $Y2=0
cc_241 N_TE_B_c_193_n N_VPWR_c_660_n 0.0103345f $X=4.625 $Y=1.47 $X2=0 $Y2=0
cc_242 N_TE_B_c_195_n N_VPWR_c_660_n 0.0073741f $X=5.145 $Y=1.47 $X2=0 $Y2=0
cc_243 N_TE_B_c_197_n N_VPWR_c_660_n 4.80713e-19 $X=5.665 $Y=1.47 $X2=0 $Y2=0
cc_244 N_TE_B_c_195_n N_VPWR_c_661_n 5.42676e-19 $X=5.145 $Y=1.47 $X2=0 $Y2=0
cc_245 N_TE_B_c_197_n N_VPWR_c_661_n 0.0103345f $X=5.665 $Y=1.47 $X2=0 $Y2=0
cc_246 N_TE_B_c_199_n N_VPWR_c_661_n 0.00886456f $X=6.185 $Y=1.47 $X2=0 $Y2=0
cc_247 N_TE_B_c_185_n N_A_437_309#_c_789_n 0.00509617f $X=2.545 $Y=1.47 $X2=0
+ $Y2=0
cc_248 N_TE_B_c_185_n N_A_437_309#_c_793_n 0.0145793f $X=2.545 $Y=1.47 $X2=0
+ $Y2=0
cc_249 N_TE_B_c_186_n N_A_437_309#_c_793_n 6.43855e-19 $X=2.975 $Y=1.395 $X2=0
+ $Y2=0
cc_250 N_TE_B_c_187_n N_A_437_309#_c_793_n 0.0140179f $X=3.065 $Y=1.47 $X2=0
+ $Y2=0
cc_251 N_TE_B_c_180_n N_A_437_309#_c_790_n 0.00110667f $X=2.22 $Y=1.232 $X2=0
+ $Y2=0
cc_252 N_TE_B_c_187_n N_A_437_309#_c_797_n 0.00430831f $X=3.065 $Y=1.47 $X2=0
+ $Y2=0
cc_253 N_TE_B_c_189_n N_A_437_309#_c_797_n 0.00403422f $X=3.585 $Y=1.47 $X2=0
+ $Y2=0
cc_254 N_TE_B_c_189_n N_A_437_309#_c_799_n 0.0135204f $X=3.585 $Y=1.47 $X2=0
+ $Y2=0
cc_255 N_TE_B_c_190_n N_A_437_309#_c_799_n 6.43855e-19 $X=4.015 $Y=1.395 $X2=0
+ $Y2=0
cc_256 N_TE_B_c_191_n N_A_437_309#_c_799_n 0.0140179f $X=4.105 $Y=1.47 $X2=0
+ $Y2=0
cc_257 N_TE_B_c_191_n N_A_437_309#_c_802_n 0.00430831f $X=4.105 $Y=1.47 $X2=0
+ $Y2=0
cc_258 N_TE_B_c_193_n N_A_437_309#_c_802_n 0.00403422f $X=4.625 $Y=1.47 $X2=0
+ $Y2=0
cc_259 N_TE_B_c_193_n N_A_437_309#_c_804_n 0.0135204f $X=4.625 $Y=1.47 $X2=0
+ $Y2=0
cc_260 N_TE_B_c_194_n N_A_437_309#_c_804_n 6.43855e-19 $X=5.055 $Y=1.395 $X2=0
+ $Y2=0
cc_261 N_TE_B_c_195_n N_A_437_309#_c_804_n 0.0140179f $X=5.145 $Y=1.47 $X2=0
+ $Y2=0
cc_262 N_TE_B_c_195_n N_A_437_309#_c_807_n 0.00430831f $X=5.145 $Y=1.47 $X2=0
+ $Y2=0
cc_263 N_TE_B_c_197_n N_A_437_309#_c_807_n 0.00403422f $X=5.665 $Y=1.47 $X2=0
+ $Y2=0
cc_264 N_TE_B_c_199_n N_A_437_309#_c_809_n 0.0136757f $X=6.185 $Y=1.47 $X2=0
+ $Y2=0
cc_265 N_TE_B_c_188_n N_A_437_309#_c_810_n 6.24408e-19 $X=3.495 $Y=1.395 $X2=0
+ $Y2=0
cc_266 N_TE_B_c_192_n N_A_437_309#_c_811_n 6.24408e-19 $X=4.535 $Y=1.395 $X2=0
+ $Y2=0
cc_267 N_TE_B_c_196_n N_A_437_309#_c_812_n 6.24408e-19 $X=5.575 $Y=1.395 $X2=0
+ $Y2=0
cc_268 N_TE_B_c_197_n N_A_437_309#_c_813_n 0.0135204f $X=5.665 $Y=1.47 $X2=0
+ $Y2=0
cc_269 N_TE_B_c_198_n N_A_437_309#_c_813_n 6.43855e-19 $X=6.095 $Y=1.395 $X2=0
+ $Y2=0
cc_270 N_TE_B_c_199_n N_A_437_309#_c_813_n 0.015737f $X=6.185 $Y=1.47 $X2=0
+ $Y2=0
cc_271 N_TE_B_c_184_n N_Z_c_900_n 0.00694639f $X=2.455 $Y=1.395 $X2=0 $Y2=0
cc_272 N_TE_B_c_185_n N_Z_c_900_n 0.0154731f $X=2.545 $Y=1.47 $X2=0 $Y2=0
cc_273 N_TE_B_c_186_n N_Z_c_900_n 0.00647232f $X=2.975 $Y=1.395 $X2=0 $Y2=0
cc_274 N_TE_B_c_187_n N_Z_c_900_n 0.0138785f $X=3.065 $Y=1.47 $X2=0 $Y2=0
cc_275 N_TE_B_c_188_n N_Z_c_900_n 0.00640772f $X=3.495 $Y=1.395 $X2=0 $Y2=0
cc_276 N_TE_B_c_189_n N_Z_c_900_n 0.0138785f $X=3.585 $Y=1.47 $X2=0 $Y2=0
cc_277 N_TE_B_c_190_n N_Z_c_900_n 0.00640772f $X=4.015 $Y=1.395 $X2=0 $Y2=0
cc_278 N_TE_B_c_191_n N_Z_c_900_n 0.0138785f $X=4.105 $Y=1.47 $X2=0 $Y2=0
cc_279 N_TE_B_c_192_n N_Z_c_900_n 0.00640772f $X=4.535 $Y=1.395 $X2=0 $Y2=0
cc_280 N_TE_B_c_193_n N_Z_c_900_n 0.0138785f $X=4.625 $Y=1.47 $X2=0 $Y2=0
cc_281 N_TE_B_c_194_n N_Z_c_900_n 0.00640772f $X=5.055 $Y=1.395 $X2=0 $Y2=0
cc_282 N_TE_B_c_195_n N_Z_c_900_n 0.0138785f $X=5.145 $Y=1.47 $X2=0 $Y2=0
cc_283 N_TE_B_c_196_n N_Z_c_900_n 0.00640772f $X=5.575 $Y=1.395 $X2=0 $Y2=0
cc_284 N_TE_B_c_197_n N_Z_c_900_n 0.0138785f $X=5.665 $Y=1.47 $X2=0 $Y2=0
cc_285 N_TE_B_c_198_n N_Z_c_900_n 0.00906427f $X=6.095 $Y=1.395 $X2=0 $Y2=0
cc_286 N_TE_B_c_199_n N_Z_c_900_n 0.0164674f $X=6.185 $Y=1.47 $X2=0 $Y2=0
cc_287 N_TE_B_c_180_n N_Z_c_900_n 0.0027955f $X=2.22 $Y=1.232 $X2=0 $Y2=0
cc_288 N_TE_B_c_202_n N_Z_c_900_n 0.0018791f $X=2.545 $Y=1.395 $X2=0 $Y2=0
cc_289 N_TE_B_c_203_n N_Z_c_900_n 0.00176164f $X=3.065 $Y=1.395 $X2=0 $Y2=0
cc_290 N_TE_B_c_204_n N_Z_c_900_n 0.00176164f $X=3.585 $Y=1.395 $X2=0 $Y2=0
cc_291 N_TE_B_c_205_n N_Z_c_900_n 0.00176164f $X=4.105 $Y=1.395 $X2=0 $Y2=0
cc_292 N_TE_B_c_206_n N_Z_c_900_n 0.00176164f $X=4.625 $Y=1.395 $X2=0 $Y2=0
cc_293 N_TE_B_c_207_n N_Z_c_900_n 0.00176164f $X=5.145 $Y=1.395 $X2=0 $Y2=0
cc_294 N_TE_B_c_208_n N_Z_c_900_n 0.00176164f $X=5.665 $Y=1.395 $X2=0 $Y2=0
cc_295 TE_B N_VGND_M1026_s 0.00384013f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_296 N_TE_B_c_177_n N_VGND_c_1009_n 0.00414152f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_297 N_TE_B_c_178_n N_VGND_c_1009_n 3.24606e-19 $X=1.655 $Y=1.16 $X2=0 $Y2=0
cc_298 TE_B N_VGND_c_1009_n 0.0256921f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_299 N_TE_B_c_177_n N_VGND_c_1010_n 0.00541359f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_300 N_TE_B_c_177_n N_VGND_c_1013_n 0.0112237f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_301 TE_B N_VGND_c_1013_n 0.00197758f $X=1.165 $Y=1.445 $X2=0 $Y2=0
cc_302 N_TE_B_c_177_n N_A_485_47#_c_1133_n 3.20478e-19 $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_A_321_47#_c_366_n N_A_124_297#_M1004_g 0.0132555f $X=6.45 $Y=0.96 $X2=0
+ $Y2=0
cc_304 N_A_321_47#_c_376_n N_A_124_297#_M1004_g 0.0211819f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_305 N_A_321_47#_c_375_n N_A_124_297#_c_516_n 0.191275f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_306 N_A_321_47#_c_376_n N_A_124_297#_c_516_n 7.54558e-19 $X=6.71 $Y=1.16
+ $X2=0 $Y2=0
cc_307 N_A_321_47#_c_377_n N_A_124_297#_c_516_n 0.00444024f $X=1.79 $Y=0.56
+ $X2=0 $Y2=0
cc_308 N_A_321_47#_c_379_n N_A_124_297#_c_516_n 0.00479555f $X=1.79 $Y=1.63
+ $X2=0 $Y2=0
cc_309 N_A_321_47#_c_416_n N_A_124_297#_c_516_n 0.047079f $X=1.942 $Y=1.15 $X2=0
+ $Y2=0
cc_310 N_A_321_47#_c_375_n N_A_124_297#_c_551_n 0.0127153f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_311 N_A_321_47#_c_376_n N_A_124_297#_c_551_n 4.24061e-19 $X=6.71 $Y=1.16
+ $X2=0 $Y2=0
cc_312 N_A_321_47#_c_375_n N_A_124_297#_c_517_n 0.00100363f $X=6.71 $Y=1.16
+ $X2=0 $Y2=0
cc_313 N_A_321_47#_c_378_n N_VPWR_c_649_n 0.0478069f $X=1.79 $Y=2.31 $X2=0 $Y2=0
cc_314 N_A_321_47#_c_378_n N_VPWR_c_652_n 0.0259025f $X=1.79 $Y=2.31 $X2=0 $Y2=0
cc_315 N_A_321_47#_M1014_d N_VPWR_c_646_n 0.00217517f $X=1.645 $Y=1.485 $X2=0
+ $Y2=0
cc_316 N_A_321_47#_c_378_n N_VPWR_c_646_n 0.0149397f $X=1.79 $Y=2.31 $X2=0 $Y2=0
cc_317 N_A_321_47#_c_378_n N_A_437_309#_c_789_n 0.0330734f $X=1.79 $Y=2.31 $X2=0
+ $Y2=0
cc_318 N_A_321_47#_c_378_n N_A_437_309#_c_790_n 0.0152479f $X=1.79 $Y=2.31 $X2=0
+ $Y2=0
cc_319 N_A_321_47#_c_353_n N_Z_c_900_n 0.00268878f $X=2.885 $Y=1.035 $X2=0 $Y2=0
cc_320 N_A_321_47#_c_365_n N_Z_c_900_n 0.00101952f $X=6.375 $Y=1.035 $X2=0 $Y2=0
cc_321 N_A_321_47#_c_373_n N_Z_c_900_n 0.00895263f $X=6.375 $Y=0.96 $X2=0 $Y2=0
cc_322 N_A_321_47#_c_375_n N_Z_c_900_n 0.32962f $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_321_47#_c_380_n N_Z_c_900_n 0.0245672f $X=1.775 $Y=1.495 $X2=0 $Y2=0
cc_324 N_A_321_47#_c_354_n N_VGND_c_1006_n 0.00342417f $X=3.33 $Y=0.96 $X2=0
+ $Y2=0
cc_325 N_A_321_47#_c_356_n N_VGND_c_1006_n 0.00342417f $X=3.85 $Y=0.96 $X2=0
+ $Y2=0
cc_326 N_A_321_47#_c_358_n N_VGND_c_1007_n 5.32249e-19 $X=4.37 $Y=0.96 $X2=0
+ $Y2=0
cc_327 N_A_321_47#_c_360_n N_VGND_c_1007_n 0.00755398f $X=4.89 $Y=0.96 $X2=0
+ $Y2=0
cc_328 N_A_321_47#_c_362_n N_VGND_c_1007_n 0.00798115f $X=5.41 $Y=0.96 $X2=0
+ $Y2=0
cc_329 N_A_321_47#_c_364_n N_VGND_c_1007_n 6.02788e-19 $X=5.93 $Y=0.96 $X2=0
+ $Y2=0
cc_330 N_A_321_47#_c_358_n N_VGND_c_1008_n 0.00342417f $X=4.37 $Y=0.96 $X2=0
+ $Y2=0
cc_331 N_A_321_47#_c_360_n N_VGND_c_1008_n 0.00342417f $X=4.89 $Y=0.96 $X2=0
+ $Y2=0
cc_332 N_A_321_47#_c_351_n N_VGND_c_1010_n 0.00342417f $X=2.81 $Y=0.96 $X2=0
+ $Y2=0
cc_333 N_A_321_47#_c_377_n N_VGND_c_1010_n 0.0373877f $X=1.79 $Y=0.56 $X2=0
+ $Y2=0
cc_334 N_A_321_47#_c_362_n N_VGND_c_1011_n 0.00342417f $X=5.41 $Y=0.96 $X2=0
+ $Y2=0
cc_335 N_A_321_47#_c_364_n N_VGND_c_1011_n 0.00342417f $X=5.93 $Y=0.96 $X2=0
+ $Y2=0
cc_336 N_A_321_47#_c_366_n N_VGND_c_1012_n 0.00342417f $X=6.45 $Y=0.96 $X2=0
+ $Y2=0
cc_337 N_A_321_47#_M1007_d N_VGND_c_1013_n 0.00251112f $X=1.605 $Y=0.235 $X2=0
+ $Y2=0
cc_338 N_A_321_47#_c_351_n N_VGND_c_1013_n 0.00540331f $X=2.81 $Y=0.96 $X2=0
+ $Y2=0
cc_339 N_A_321_47#_c_354_n N_VGND_c_1013_n 0.00427787f $X=3.33 $Y=0.96 $X2=0
+ $Y2=0
cc_340 N_A_321_47#_c_356_n N_VGND_c_1013_n 0.00427787f $X=3.85 $Y=0.96 $X2=0
+ $Y2=0
cc_341 N_A_321_47#_c_358_n N_VGND_c_1013_n 0.00427787f $X=4.37 $Y=0.96 $X2=0
+ $Y2=0
cc_342 N_A_321_47#_c_360_n N_VGND_c_1013_n 0.00427787f $X=4.89 $Y=0.96 $X2=0
+ $Y2=0
cc_343 N_A_321_47#_c_362_n N_VGND_c_1013_n 0.00427787f $X=5.41 $Y=0.96 $X2=0
+ $Y2=0
cc_344 N_A_321_47#_c_364_n N_VGND_c_1013_n 0.00427787f $X=5.93 $Y=0.96 $X2=0
+ $Y2=0
cc_345 N_A_321_47#_c_366_n N_VGND_c_1013_n 0.00466313f $X=6.45 $Y=0.96 $X2=0
+ $Y2=0
cc_346 N_A_321_47#_c_377_n N_VGND_c_1013_n 0.0213263f $X=1.79 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_A_321_47#_c_351_n N_VGND_c_1014_n 0.00901456f $X=2.81 $Y=0.96 $X2=0
+ $Y2=0
cc_348 N_A_321_47#_c_354_n N_VGND_c_1014_n 0.00798115f $X=3.33 $Y=0.96 $X2=0
+ $Y2=0
cc_349 N_A_321_47#_c_356_n N_VGND_c_1014_n 6.02788e-19 $X=3.85 $Y=0.96 $X2=0
+ $Y2=0
cc_350 N_A_321_47#_c_354_n N_VGND_c_1015_n 5.89906e-19 $X=3.33 $Y=0.96 $X2=0
+ $Y2=0
cc_351 N_A_321_47#_c_356_n N_VGND_c_1015_n 0.00773282f $X=3.85 $Y=0.96 $X2=0
+ $Y2=0
cc_352 N_A_321_47#_c_358_n N_VGND_c_1015_n 0.00782596f $X=4.37 $Y=0.96 $X2=0
+ $Y2=0
cc_353 N_A_321_47#_c_360_n N_VGND_c_1015_n 5.46358e-19 $X=4.89 $Y=0.96 $X2=0
+ $Y2=0
cc_354 N_A_321_47#_c_362_n N_VGND_c_1016_n 5.89906e-19 $X=5.41 $Y=0.96 $X2=0
+ $Y2=0
cc_355 N_A_321_47#_c_364_n N_VGND_c_1016_n 0.00773282f $X=5.93 $Y=0.96 $X2=0
+ $Y2=0
cc_356 N_A_321_47#_c_366_n N_VGND_c_1016_n 0.00930435f $X=6.45 $Y=0.96 $X2=0
+ $Y2=0
cc_357 N_A_321_47#_c_377_n N_A_485_47#_c_1132_n 0.0350095f $X=1.79 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_321_47#_c_351_n N_A_485_47#_c_1137_n 0.0129905f $X=2.81 $Y=0.96 $X2=0
+ $Y2=0
cc_359 N_A_321_47#_c_352_n N_A_485_47#_c_1137_n 0.00393903f $X=3.255 $Y=1.035
+ $X2=0 $Y2=0
cc_360 N_A_321_47#_c_354_n N_A_485_47#_c_1137_n 0.0123018f $X=3.33 $Y=0.96 $X2=0
+ $Y2=0
cc_361 N_A_321_47#_c_355_n N_A_485_47#_c_1137_n 2.04719e-19 $X=3.775 $Y=1.035
+ $X2=0 $Y2=0
cc_362 N_A_321_47#_c_375_n N_A_485_47#_c_1137_n 0.047834f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_363 N_A_321_47#_c_375_n N_A_485_47#_c_1133_n 0.0293764f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_364 N_A_321_47#_c_377_n N_A_485_47#_c_1133_n 0.0182702f $X=1.79 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_321_47#_c_354_n N_A_485_47#_c_1144_n 0.00450849f $X=3.33 $Y=0.96
+ $X2=0 $Y2=0
cc_366 N_A_321_47#_c_356_n N_A_485_47#_c_1145_n 0.0123018f $X=3.85 $Y=0.96 $X2=0
+ $Y2=0
cc_367 N_A_321_47#_c_357_n N_A_485_47#_c_1145_n 0.00393903f $X=4.295 $Y=1.035
+ $X2=0 $Y2=0
cc_368 N_A_321_47#_c_358_n N_A_485_47#_c_1145_n 0.0123018f $X=4.37 $Y=0.96 $X2=0
+ $Y2=0
cc_369 N_A_321_47#_c_359_n N_A_485_47#_c_1145_n 2.04719e-19 $X=4.815 $Y=1.035
+ $X2=0 $Y2=0
cc_370 N_A_321_47#_c_375_n N_A_485_47#_c_1145_n 0.0475999f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_371 N_A_321_47#_c_358_n N_A_485_47#_c_1150_n 0.00467419f $X=4.37 $Y=0.96
+ $X2=0 $Y2=0
cc_372 N_A_321_47#_c_360_n N_A_485_47#_c_1151_n 0.0123018f $X=4.89 $Y=0.96 $X2=0
+ $Y2=0
cc_373 N_A_321_47#_c_361_n N_A_485_47#_c_1151_n 0.00393903f $X=5.335 $Y=1.035
+ $X2=0 $Y2=0
cc_374 N_A_321_47#_c_362_n N_A_485_47#_c_1151_n 0.0123018f $X=5.41 $Y=0.96 $X2=0
+ $Y2=0
cc_375 N_A_321_47#_c_363_n N_A_485_47#_c_1151_n 2.04719e-19 $X=5.855 $Y=1.035
+ $X2=0 $Y2=0
cc_376 N_A_321_47#_c_375_n N_A_485_47#_c_1151_n 0.0475999f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_377 N_A_321_47#_c_362_n N_A_485_47#_c_1156_n 0.00450849f $X=5.41 $Y=0.96
+ $X2=0 $Y2=0
cc_378 N_A_321_47#_c_364_n N_A_485_47#_c_1157_n 0.0122265f $X=5.93 $Y=0.96 $X2=0
+ $Y2=0
cc_379 N_A_321_47#_c_365_n N_A_485_47#_c_1157_n 0.00393903f $X=6.375 $Y=1.035
+ $X2=0 $Y2=0
cc_380 N_A_321_47#_c_366_n N_A_485_47#_c_1157_n 0.0132198f $X=6.45 $Y=0.96 $X2=0
+ $Y2=0
cc_381 N_A_321_47#_c_375_n N_A_485_47#_c_1157_n 0.0476314f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_382 N_A_321_47#_c_376_n N_A_485_47#_c_1157_n 0.00226806f $X=6.71 $Y=1.16
+ $X2=0 $Y2=0
cc_383 N_A_321_47#_c_355_n N_A_485_47#_c_1162_n 0.00386339f $X=3.775 $Y=1.035
+ $X2=0 $Y2=0
cc_384 N_A_321_47#_c_375_n N_A_485_47#_c_1162_n 0.0158845f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_385 N_A_321_47#_c_359_n N_A_485_47#_c_1164_n 0.00386799f $X=4.815 $Y=1.035
+ $X2=0 $Y2=0
cc_386 N_A_321_47#_c_375_n N_A_485_47#_c_1164_n 0.0159243f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_387 N_A_321_47#_c_363_n N_A_485_47#_c_1166_n 0.00386339f $X=5.855 $Y=1.035
+ $X2=0 $Y2=0
cc_388 N_A_321_47#_c_375_n N_A_485_47#_c_1166_n 0.0158845f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_389 N_A_321_47#_c_366_n N_A_485_47#_c_1168_n 0.00821429f $X=6.45 $Y=0.96
+ $X2=0 $Y2=0
cc_390 N_A_321_47#_c_375_n N_A_485_47#_c_1168_n 0.0183192f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_391 N_A_321_47#_c_376_n N_A_485_47#_c_1168_n 0.00625982f $X=6.71 $Y=1.16
+ $X2=0 $Y2=0
cc_392 N_A_124_297#_c_554_p N_VPWR_c_649_n 0.0451172f $X=0.765 $Y=2.22 $X2=0
+ $Y2=0
cc_393 N_A_124_297#_c_516_n N_VPWR_c_649_n 0.00140918f $X=7.52 $Y=1.145 $X2=0
+ $Y2=0
cc_394 N_A_124_297#_c_554_p N_VPWR_c_653_n 0.0124854f $X=0.765 $Y=2.22 $X2=0
+ $Y2=0
cc_395 N_A_124_297#_c_519_n N_VPWR_c_656_n 0.00429453f $X=7.205 $Y=1.41 $X2=0
+ $Y2=0
cc_396 N_A_124_297#_c_520_n N_VPWR_c_656_n 0.00429453f $X=7.675 $Y=1.41 $X2=0
+ $Y2=0
cc_397 N_A_124_297#_c_521_n N_VPWR_c_656_n 0.00429453f $X=8.145 $Y=1.41 $X2=0
+ $Y2=0
cc_398 N_A_124_297#_c_522_n N_VPWR_c_656_n 0.00429453f $X=8.615 $Y=1.41 $X2=0
+ $Y2=0
cc_399 N_A_124_297#_c_523_n N_VPWR_c_656_n 0.00429453f $X=9.085 $Y=1.41 $X2=0
+ $Y2=0
cc_400 N_A_124_297#_c_524_n N_VPWR_c_656_n 0.00429453f $X=9.555 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A_124_297#_c_525_n N_VPWR_c_656_n 0.00429453f $X=10.025 $Y=1.41 $X2=0
+ $Y2=0
cc_402 N_A_124_297#_c_526_n N_VPWR_c_656_n 0.00429453f $X=10.495 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_A_124_297#_M1005_s N_VPWR_c_646_n 0.00604325f $X=0.62 $Y=1.485 $X2=0
+ $Y2=0
cc_404 N_A_124_297#_c_519_n N_VPWR_c_646_n 0.00743756f $X=7.205 $Y=1.41 $X2=0
+ $Y2=0
cc_405 N_A_124_297#_c_520_n N_VPWR_c_646_n 0.00606499f $X=7.675 $Y=1.41 $X2=0
+ $Y2=0
cc_406 N_A_124_297#_c_521_n N_VPWR_c_646_n 0.00606499f $X=8.145 $Y=1.41 $X2=0
+ $Y2=0
cc_407 N_A_124_297#_c_522_n N_VPWR_c_646_n 0.00606499f $X=8.615 $Y=1.41 $X2=0
+ $Y2=0
cc_408 N_A_124_297#_c_523_n N_VPWR_c_646_n 0.00606499f $X=9.085 $Y=1.41 $X2=0
+ $Y2=0
cc_409 N_A_124_297#_c_524_n N_VPWR_c_646_n 0.00606499f $X=9.555 $Y=1.41 $X2=0
+ $Y2=0
cc_410 N_A_124_297#_c_525_n N_VPWR_c_646_n 0.00606499f $X=10.025 $Y=1.41 $X2=0
+ $Y2=0
cc_411 N_A_124_297#_c_526_n N_VPWR_c_646_n 0.00701975f $X=10.495 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_A_124_297#_c_554_p N_VPWR_c_646_n 0.00704765f $X=0.765 $Y=2.22 $X2=0
+ $Y2=0
cc_413 N_A_124_297#_c_519_n N_A_437_309#_c_791_n 0.0345153f $X=7.205 $Y=1.41
+ $X2=0 $Y2=0
cc_414 N_A_124_297#_c_520_n N_A_437_309#_c_791_n 0.0206878f $X=7.675 $Y=1.41
+ $X2=0 $Y2=0
cc_415 N_A_124_297#_c_521_n N_A_437_309#_c_791_n 0.0206878f $X=8.145 $Y=1.41
+ $X2=0 $Y2=0
cc_416 N_A_124_297#_c_522_n N_A_437_309#_c_791_n 0.0206878f $X=8.615 $Y=1.41
+ $X2=0 $Y2=0
cc_417 N_A_124_297#_c_523_n N_A_437_309#_c_791_n 0.0206878f $X=9.085 $Y=1.41
+ $X2=0 $Y2=0
cc_418 N_A_124_297#_c_524_n N_A_437_309#_c_791_n 0.0206878f $X=9.555 $Y=1.41
+ $X2=0 $Y2=0
cc_419 N_A_124_297#_c_525_n N_A_437_309#_c_791_n 0.0206878f $X=10.025 $Y=1.41
+ $X2=0 $Y2=0
cc_420 N_A_124_297#_c_526_n N_A_437_309#_c_791_n 0.0206878f $X=10.495 $Y=1.41
+ $X2=0 $Y2=0
cc_421 N_A_124_297#_M1004_g N_Z_c_930_n 0.00337382f $X=7.18 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A_124_297#_M1011_g N_Z_c_930_n 0.0105488f $X=7.65 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A_124_297#_M1023_g N_Z_c_930_n 0.0106269f $X=8.12 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A_124_297#_M1024_g N_Z_c_930_n 0.0106269f $X=8.59 $Y=0.56 $X2=0 $Y2=0
cc_425 N_A_124_297#_M1025_g N_Z_c_930_n 0.0106269f $X=9.06 $Y=0.56 $X2=0 $Y2=0
cc_426 N_A_124_297#_M1027_g N_Z_c_930_n 0.0106269f $X=9.53 $Y=0.56 $X2=0 $Y2=0
cc_427 N_A_124_297#_M1029_g N_Z_c_930_n 0.0106269f $X=10 $Y=0.56 $X2=0 $Y2=0
cc_428 N_A_124_297#_M1037_g N_Z_c_930_n 0.0140914f $X=10.52 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A_124_297#_c_591_p N_Z_c_930_n 0.00256035f $X=7.715 $Y=1.145 $X2=0
+ $Y2=0
cc_430 N_A_124_297#_c_516_n N_Z_c_930_n 0.00182713f $X=7.52 $Y=1.145 $X2=0 $Y2=0
cc_431 N_A_124_297#_c_551_n N_Z_c_930_n 0.203603f $X=9.99 $Y=1.16 $X2=0 $Y2=0
cc_432 N_A_124_297#_c_517_n N_Z_c_930_n 0.0223478f $X=10.495 $Y=1.217 $X2=0
+ $Y2=0
cc_433 N_A_124_297#_c_526_n Z 0.00135624f $X=10.495 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A_124_297#_M1037_g Z 0.0199297f $X=10.52 $Y=0.56 $X2=0 $Y2=0
cc_435 N_A_124_297#_c_551_n Z 0.0167743f $X=9.99 $Y=1.16 $X2=0 $Y2=0
cc_436 N_A_124_297#_c_519_n N_Z_c_900_n 0.0168513f $X=7.205 $Y=1.41 $X2=0 $Y2=0
cc_437 N_A_124_297#_c_520_n N_Z_c_900_n 0.013509f $X=7.675 $Y=1.41 $X2=0 $Y2=0
cc_438 N_A_124_297#_c_521_n N_Z_c_900_n 0.0136002f $X=8.145 $Y=1.41 $X2=0 $Y2=0
cc_439 N_A_124_297#_c_522_n N_Z_c_900_n 0.0136002f $X=8.615 $Y=1.41 $X2=0 $Y2=0
cc_440 N_A_124_297#_c_523_n N_Z_c_900_n 0.0136002f $X=9.085 $Y=1.41 $X2=0 $Y2=0
cc_441 N_A_124_297#_c_524_n N_Z_c_900_n 0.0136002f $X=9.555 $Y=1.41 $X2=0 $Y2=0
cc_442 N_A_124_297#_c_525_n N_Z_c_900_n 0.0136002f $X=10.025 $Y=1.41 $X2=0 $Y2=0
cc_443 N_A_124_297#_c_526_n N_Z_c_900_n 0.0175577f $X=10.495 $Y=1.41 $X2=0 $Y2=0
cc_444 N_A_124_297#_c_516_n N_Z_c_900_n 0.0491047f $X=7.52 $Y=1.145 $X2=0 $Y2=0
cc_445 N_A_124_297#_c_551_n N_Z_c_900_n 0.244493f $X=9.99 $Y=1.16 $X2=0 $Y2=0
cc_446 N_A_124_297#_c_517_n N_Z_c_900_n 0.0516717f $X=10.495 $Y=1.217 $X2=0
+ $Y2=0
cc_447 N_A_124_297#_c_518_n N_VGND_c_1009_n 0.0234059f $X=0.765 $Y=0.445 $X2=0
+ $Y2=0
cc_448 N_A_124_297#_M1004_g N_VGND_c_1012_n 0.00357877f $X=7.18 $Y=0.56 $X2=0
+ $Y2=0
cc_449 N_A_124_297#_M1011_g N_VGND_c_1012_n 0.00357877f $X=7.65 $Y=0.56 $X2=0
+ $Y2=0
cc_450 N_A_124_297#_M1023_g N_VGND_c_1012_n 0.00357877f $X=8.12 $Y=0.56 $X2=0
+ $Y2=0
cc_451 N_A_124_297#_M1024_g N_VGND_c_1012_n 0.00357877f $X=8.59 $Y=0.56 $X2=0
+ $Y2=0
cc_452 N_A_124_297#_M1025_g N_VGND_c_1012_n 0.00357877f $X=9.06 $Y=0.56 $X2=0
+ $Y2=0
cc_453 N_A_124_297#_M1027_g N_VGND_c_1012_n 0.00357877f $X=9.53 $Y=0.56 $X2=0
+ $Y2=0
cc_454 N_A_124_297#_M1029_g N_VGND_c_1012_n 0.00357877f $X=10 $Y=0.56 $X2=0
+ $Y2=0
cc_455 N_A_124_297#_M1037_g N_VGND_c_1012_n 0.00357877f $X=10.52 $Y=0.56 $X2=0
+ $Y2=0
cc_456 N_A_124_297#_M1013_d N_VGND_c_1013_n 0.006832f $X=0.63 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_124_297#_M1004_g N_VGND_c_1013_n 0.00603279f $X=7.18 $Y=0.56 $X2=0
+ $Y2=0
cc_458 N_A_124_297#_M1011_g N_VGND_c_1013_n 0.00548399f $X=7.65 $Y=0.56 $X2=0
+ $Y2=0
cc_459 N_A_124_297#_M1023_g N_VGND_c_1013_n 0.00548399f $X=8.12 $Y=0.56 $X2=0
+ $Y2=0
cc_460 N_A_124_297#_M1024_g N_VGND_c_1013_n 0.00548399f $X=8.59 $Y=0.56 $X2=0
+ $Y2=0
cc_461 N_A_124_297#_M1025_g N_VGND_c_1013_n 0.00548399f $X=9.06 $Y=0.56 $X2=0
+ $Y2=0
cc_462 N_A_124_297#_M1027_g N_VGND_c_1013_n 0.00548399f $X=9.53 $Y=0.56 $X2=0
+ $Y2=0
cc_463 N_A_124_297#_M1029_g N_VGND_c_1013_n 0.00560377f $X=10 $Y=0.56 $X2=0
+ $Y2=0
cc_464 N_A_124_297#_M1037_g N_VGND_c_1013_n 0.00647566f $X=10.52 $Y=0.56 $X2=0
+ $Y2=0
cc_465 N_A_124_297#_c_518_n N_VGND_c_1013_n 0.00753309f $X=0.765 $Y=0.445 $X2=0
+ $Y2=0
cc_466 N_A_124_297#_c_516_n N_A_485_47#_c_1137_n 0.00492838f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_467 N_A_124_297#_c_516_n N_A_485_47#_c_1133_n 0.00257709f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_468 N_A_124_297#_c_516_n N_A_485_47#_c_1145_n 0.00492838f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_469 N_A_124_297#_c_516_n N_A_485_47#_c_1151_n 0.00492838f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_470 N_A_124_297#_c_516_n N_A_485_47#_c_1157_n 0.0049309f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_471 N_A_124_297#_M1004_g N_A_485_47#_c_1134_n 0.0123142f $X=7.18 $Y=0.56
+ $X2=0 $Y2=0
cc_472 N_A_124_297#_M1011_g N_A_485_47#_c_1134_n 0.00840951f $X=7.65 $Y=0.56
+ $X2=0 $Y2=0
cc_473 N_A_124_297#_M1023_g N_A_485_47#_c_1134_n 0.00847746f $X=8.12 $Y=0.56
+ $X2=0 $Y2=0
cc_474 N_A_124_297#_M1024_g N_A_485_47#_c_1134_n 0.00847746f $X=8.59 $Y=0.56
+ $X2=0 $Y2=0
cc_475 N_A_124_297#_M1025_g N_A_485_47#_c_1134_n 0.00847746f $X=9.06 $Y=0.56
+ $X2=0 $Y2=0
cc_476 N_A_124_297#_M1027_g N_A_485_47#_c_1134_n 0.00847746f $X=9.53 $Y=0.56
+ $X2=0 $Y2=0
cc_477 N_A_124_297#_M1029_g N_A_485_47#_c_1134_n 0.00876725f $X=10 $Y=0.56 $X2=0
+ $Y2=0
cc_478 N_A_124_297#_M1037_g N_A_485_47#_c_1134_n 0.00876725f $X=10.52 $Y=0.56
+ $X2=0 $Y2=0
cc_479 N_A_124_297#_c_551_n N_A_485_47#_c_1134_n 0.0025603f $X=9.99 $Y=1.16
+ $X2=0 $Y2=0
cc_480 N_A_124_297#_c_516_n N_A_485_47#_c_1162_n 0.00148759f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_481 N_A_124_297#_c_516_n N_A_485_47#_c_1164_n 0.00149207f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_482 N_A_124_297#_c_516_n N_A_485_47#_c_1166_n 0.00148759f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_483 N_A_124_297#_c_516_n N_A_485_47#_c_1168_n 0.00699828f $X=7.52 $Y=1.145
+ $X2=0 $Y2=0
cc_484 N_VPWR_c_646_n N_A_437_309#_M1000_s 0.00239949f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_485 N_VPWR_c_646_n N_A_437_309#_M1001_s 0.00335964f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_646_n N_A_437_309#_M1003_s 0.00335964f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_646_n N_A_437_309#_M1012_s 0.00335964f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_646_n N_A_437_309#_M1021_s 0.00706283f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_646_n N_A_437_309#_M1015_d 0.00231289f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_646_n N_A_437_309#_M1020_d 0.00231289f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_646_n N_A_437_309#_M1030_d 0.00231289f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_646_n N_A_437_309#_M1035_d 0.00233941f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_651_n N_A_437_309#_c_789_n 0.0178356f $X=2.78 $Y=2.36 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_652_n N_A_437_309#_c_789_n 0.0172681f $X=2.565 $Y=2.72 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_646_n N_A_437_309#_c_789_n 0.00950719f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_496 N_VPWR_M1000_d N_A_437_309#_c_793_n 0.00450015f $X=2.635 $Y=1.545 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_651_n N_A_437_309#_c_793_n 0.0235907f $X=2.78 $Y=2.36 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_652_n N_A_437_309#_c_793_n 0.00227617f $X=2.565 $Y=2.72 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_654_n N_A_437_309#_c_793_n 0.00305754f $X=3.605 $Y=2.72 $X2=0
+ $Y2=0
cc_500 N_VPWR_c_646_n N_A_437_309#_c_793_n 0.0112842f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_651_n N_A_437_309#_c_797_n 0.0142149f $X=2.78 $Y=2.36 $X2=0
+ $Y2=0
cc_502 N_VPWR_c_654_n N_A_437_309#_c_797_n 0.0116627f $X=3.605 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_646_n N_A_437_309#_c_797_n 0.00644035f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_504 N_VPWR_c_659_n N_A_437_309#_c_797_n 0.0142151f $X=3.82 $Y=2.36 $X2=0
+ $Y2=0
cc_505 N_VPWR_M1002_d N_A_437_309#_c_799_n 0.00450015f $X=3.675 $Y=1.545 $X2=0
+ $Y2=0
cc_506 N_VPWR_c_654_n N_A_437_309#_c_799_n 0.00312887f $X=3.605 $Y=2.72 $X2=0
+ $Y2=0
cc_507 N_VPWR_c_655_n N_A_437_309#_c_799_n 0.00305754f $X=4.645 $Y=2.72 $X2=0
+ $Y2=0
cc_508 N_VPWR_c_646_n N_A_437_309#_c_799_n 0.01269f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_509 N_VPWR_c_659_n N_A_437_309#_c_799_n 0.0235907f $X=3.82 $Y=2.36 $X2=0
+ $Y2=0
cc_510 N_VPWR_c_655_n N_A_437_309#_c_802_n 0.0116627f $X=4.645 $Y=2.72 $X2=0
+ $Y2=0
cc_511 N_VPWR_c_646_n N_A_437_309#_c_802_n 0.00644035f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_512 N_VPWR_c_659_n N_A_437_309#_c_802_n 0.0142149f $X=3.82 $Y=2.36 $X2=0
+ $Y2=0
cc_513 N_VPWR_c_660_n N_A_437_309#_c_802_n 0.0142151f $X=4.86 $Y=2.36 $X2=0
+ $Y2=0
cc_514 N_VPWR_M1006_d N_A_437_309#_c_804_n 0.00450015f $X=4.715 $Y=1.545 $X2=0
+ $Y2=0
cc_515 N_VPWR_c_650_n N_A_437_309#_c_804_n 0.00305754f $X=5.685 $Y=2.72 $X2=0
+ $Y2=0
cc_516 N_VPWR_c_655_n N_A_437_309#_c_804_n 0.00312887f $X=4.645 $Y=2.72 $X2=0
+ $Y2=0
cc_517 N_VPWR_c_646_n N_A_437_309#_c_804_n 0.01269f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_518 N_VPWR_c_660_n N_A_437_309#_c_804_n 0.0235907f $X=4.86 $Y=2.36 $X2=0
+ $Y2=0
cc_519 N_VPWR_c_650_n N_A_437_309#_c_807_n 0.0116627f $X=5.685 $Y=2.72 $X2=0
+ $Y2=0
cc_520 N_VPWR_c_646_n N_A_437_309#_c_807_n 0.00644035f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_521 N_VPWR_c_660_n N_A_437_309#_c_807_n 0.0142149f $X=4.86 $Y=2.36 $X2=0
+ $Y2=0
cc_522 N_VPWR_c_661_n N_A_437_309#_c_807_n 0.0142151f $X=5.9 $Y=2.36 $X2=0 $Y2=0
cc_523 N_VPWR_c_656_n N_A_437_309#_c_809_n 0.282556f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_524 N_VPWR_c_646_n N_A_437_309#_c_809_n 0.168757f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_525 N_VPWR_c_661_n N_A_437_309#_c_809_n 0.0157915f $X=5.9 $Y=2.36 $X2=0 $Y2=0
cc_526 N_VPWR_M1016_d N_A_437_309#_c_813_n 0.00450015f $X=5.755 $Y=1.545 $X2=0
+ $Y2=0
cc_527 N_VPWR_c_650_n N_A_437_309#_c_813_n 0.00312887f $X=5.685 $Y=2.72 $X2=0
+ $Y2=0
cc_528 N_VPWR_c_656_n N_A_437_309#_c_813_n 0.00305754f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_529 N_VPWR_c_646_n N_A_437_309#_c_813_n 0.0127308f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_530 N_VPWR_c_661_n N_A_437_309#_c_813_n 0.0235907f $X=5.9 $Y=2.36 $X2=0 $Y2=0
cc_531 N_VPWR_c_646_n N_Z_M1008_s 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_c_646_n N_Z_M1017_s 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_533 N_VPWR_c_646_n N_Z_M1028_s 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_534 N_VPWR_c_646_n N_Z_M1031_s 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_535 N_VPWR_M1000_d N_Z_c_900_n 0.00244559f $X=2.635 $Y=1.545 $X2=0 $Y2=0
cc_536 N_VPWR_M1002_d N_Z_c_900_n 0.00244559f $X=3.675 $Y=1.545 $X2=0 $Y2=0
cc_537 N_VPWR_M1006_d N_Z_c_900_n 0.00244559f $X=4.715 $Y=1.545 $X2=0 $Y2=0
cc_538 N_VPWR_M1016_d N_Z_c_900_n 0.00244559f $X=5.755 $Y=1.545 $X2=0 $Y2=0
cc_539 N_A_437_309#_c_791_n N_Z_M1008_s 0.00349548f $X=10.73 $Y=2.02 $X2=0 $Y2=0
cc_540 N_A_437_309#_c_791_n N_Z_M1017_s 0.00349548f $X=10.73 $Y=2.02 $X2=0 $Y2=0
cc_541 N_A_437_309#_c_791_n N_Z_M1028_s 0.00349548f $X=10.73 $Y=2.02 $X2=0 $Y2=0
cc_542 N_A_437_309#_c_791_n N_Z_M1031_s 0.00349548f $X=10.73 $Y=2.02 $X2=0 $Y2=0
cc_543 N_A_437_309#_M1035_d Z 0.00367994f $X=10.585 $Y=1.485 $X2=0 $Y2=0
cc_544 N_A_437_309#_c_791_n Z 0.0222273f $X=10.73 $Y=2.02 $X2=0 $Y2=0
cc_545 N_A_437_309#_M1000_s N_Z_c_900_n 0.00263554f $X=2.185 $Y=1.545 $X2=0
+ $Y2=0
cc_546 N_A_437_309#_M1001_s N_Z_c_900_n 0.00240864f $X=3.155 $Y=1.545 $X2=0
+ $Y2=0
cc_547 N_A_437_309#_M1003_s N_Z_c_900_n 0.00240864f $X=4.195 $Y=1.545 $X2=0
+ $Y2=0
cc_548 N_A_437_309#_M1012_s N_Z_c_900_n 0.00240864f $X=5.235 $Y=1.545 $X2=0
+ $Y2=0
cc_549 N_A_437_309#_M1021_s N_Z_c_900_n 0.0141146f $X=6.275 $Y=1.545 $X2=0 $Y2=0
cc_550 N_A_437_309#_M1015_d N_Z_c_900_n 0.00190453f $X=7.765 $Y=1.485 $X2=0
+ $Y2=0
cc_551 N_A_437_309#_M1020_d N_Z_c_900_n 0.00190453f $X=8.705 $Y=1.485 $X2=0
+ $Y2=0
cc_552 N_A_437_309#_M1030_d N_Z_c_900_n 0.00190453f $X=9.645 $Y=1.485 $X2=0
+ $Y2=0
cc_553 N_A_437_309#_M1035_d N_Z_c_900_n 3.46278e-19 $X=10.585 $Y=1.485 $X2=0
+ $Y2=0
cc_554 N_A_437_309#_c_793_n N_Z_c_900_n 0.0426593f $X=3.215 $Y=1.98 $X2=0 $Y2=0
cc_555 N_A_437_309#_c_790_n N_Z_c_900_n 0.0208868f $X=2.395 $Y=1.98 $X2=0 $Y2=0
cc_556 N_A_437_309#_c_799_n N_Z_c_900_n 0.0465044f $X=4.255 $Y=1.98 $X2=0 $Y2=0
cc_557 N_A_437_309#_c_804_n N_Z_c_900_n 0.0465044f $X=5.295 $Y=1.98 $X2=0 $Y2=0
cc_558 N_A_437_309#_c_810_n N_Z_c_900_n 0.0141171f $X=3.3 $Y=1.98 $X2=0 $Y2=0
cc_559 N_A_437_309#_c_811_n N_Z_c_900_n 0.0141171f $X=4.34 $Y=1.98 $X2=0 $Y2=0
cc_560 N_A_437_309#_c_812_n N_Z_c_900_n 0.0141171f $X=5.38 $Y=1.98 $X2=0 $Y2=0
cc_561 N_A_437_309#_c_813_n N_Z_c_900_n 0.321565f $X=6.335 $Y=2.18 $X2=0 $Y2=0
cc_562 N_Z_M1004_s N_VGND_c_1013_n 0.00256987f $X=7.255 $Y=0.235 $X2=0 $Y2=0
cc_563 N_Z_M1023_s N_VGND_c_1013_n 0.00256987f $X=8.195 $Y=0.235 $X2=0 $Y2=0
cc_564 N_Z_M1025_s N_VGND_c_1013_n 0.00256987f $X=9.135 $Y=0.235 $X2=0 $Y2=0
cc_565 N_Z_M1029_s N_VGND_c_1013_n 0.00297142f $X=10.075 $Y=0.235 $X2=0 $Y2=0
cc_566 N_Z_c_930_n N_A_485_47#_M1011_d 0.003954f $X=10.675 $Y=0.735 $X2=0 $Y2=0
cc_567 N_Z_c_930_n N_A_485_47#_M1024_d 0.00402091f $X=10.675 $Y=0.735 $X2=0
+ $Y2=0
cc_568 N_Z_c_930_n N_A_485_47#_M1027_d 0.00402091f $X=10.675 $Y=0.735 $X2=0
+ $Y2=0
cc_569 N_Z_c_930_n N_A_485_47#_M1037_d 6.34286e-19 $X=10.675 $Y=0.735 $X2=0
+ $Y2=0
cc_570 Z N_A_485_47#_M1037_d 4.96845e-19 $X=10.69 $Y=0.765 $X2=0 $Y2=0
cc_571 N_Z_c_897_n N_A_485_47#_M1037_d 0.00345418f $X=10.8 $Y=0.855 $X2=0 $Y2=0
cc_572 N_Z_M1004_s N_A_485_47#_c_1134_n 0.00400887f $X=7.255 $Y=0.235 $X2=0
+ $Y2=0
cc_573 N_Z_M1023_s N_A_485_47#_c_1134_n 0.00400887f $X=8.195 $Y=0.235 $X2=0
+ $Y2=0
cc_574 N_Z_M1025_s N_A_485_47#_c_1134_n 0.00400887f $X=9.135 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_Z_M1029_s N_A_485_47#_c_1134_n 0.00507048f $X=10.075 $Y=0.235 $X2=0
+ $Y2=0
cc_576 N_Z_c_930_n N_A_485_47#_c_1134_n 0.178251f $X=10.675 $Y=0.735 $X2=0 $Y2=0
cc_577 N_Z_c_897_n N_A_485_47#_c_1134_n 0.0194298f $X=10.8 $Y=0.855 $X2=0 $Y2=0
cc_578 N_Z_c_900_n N_A_485_47#_c_1168_n 0.00246104f $X=10.675 $Y=1.585 $X2=0
+ $Y2=0
cc_579 N_VGND_c_1013_n N_A_485_47#_M1009_d 0.00269999f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_580 N_VGND_c_1013_n N_A_485_47#_M1010_d 0.00355249f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_c_1013_n N_A_485_47#_M1019_d 0.00354571f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_582 N_VGND_c_1013_n N_A_485_47#_M1032_d 0.00355249f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_1013_n N_A_485_47#_M1036_d 0.00507211f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_c_1013_n N_A_485_47#_M1011_d 0.00255381f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_1013_n N_A_485_47#_M1024_d 0.00255381f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_1013_n N_A_485_47#_M1027_d 0.00255381f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_1013_n N_A_485_47#_M1037_d 0.00225742f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_1010_n N_A_485_47#_c_1132_n 0.0262933f $X=2.855 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_1013_n N_A_485_47#_c_1132_n 0.0145099f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_M1009_s N_A_485_47#_c_1137_n 0.00478863f $X=2.885 $Y=0.235 $X2=0
+ $Y2=0
cc_591 N_VGND_c_1006_n N_A_485_47#_c_1137_n 0.00313809f $X=3.895 $Y=0 $X2=0
+ $Y2=0
cc_592 N_VGND_c_1010_n N_A_485_47#_c_1137_n 0.00235235f $X=2.855 $Y=0 $X2=0
+ $Y2=0
cc_593 N_VGND_c_1013_n N_A_485_47#_c_1137_n 0.0116203f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_1014_n N_A_485_47#_c_1137_n 0.023992f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_1006_n N_A_485_47#_c_1144_n 0.0132487f $X=3.895 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_1013_n N_A_485_47#_c_1144_n 0.00827808f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_597 N_VGND_c_1014_n N_A_485_47#_c_1144_n 0.0132273f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_598 N_VGND_M1018_s N_A_485_47#_c_1145_n 0.00478863f $X=3.925 $Y=0.235 $X2=0
+ $Y2=0
cc_599 N_VGND_c_1006_n N_A_485_47#_c_1145_n 0.00235235f $X=3.895 $Y=0 $X2=0
+ $Y2=0
cc_600 N_VGND_c_1008_n N_A_485_47#_c_1145_n 0.00313809f $X=4.935 $Y=0 $X2=0
+ $Y2=0
cc_601 N_VGND_c_1013_n N_A_485_47#_c_1145_n 0.0116203f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_602 N_VGND_c_1015_n N_A_485_47#_c_1145_n 0.023992f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_603 N_VGND_c_1008_n N_A_485_47#_c_1150_n 0.014985f $X=4.935 $Y=0 $X2=0 $Y2=0
cc_604 N_VGND_c_1013_n N_A_485_47#_c_1150_n 0.00836816f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_605 N_VGND_c_1015_n N_A_485_47#_c_1150_n 0.014487f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_606 N_VGND_M1022_s N_A_485_47#_c_1151_n 0.00478863f $X=4.965 $Y=0.235 $X2=0
+ $Y2=0
cc_607 N_VGND_c_1007_n N_A_485_47#_c_1151_n 0.023992f $X=5.15 $Y=0 $X2=0 $Y2=0
cc_608 N_VGND_c_1008_n N_A_485_47#_c_1151_n 0.00235235f $X=4.935 $Y=0 $X2=0
+ $Y2=0
cc_609 N_VGND_c_1011_n N_A_485_47#_c_1151_n 0.00313809f $X=5.975 $Y=0 $X2=0
+ $Y2=0
cc_610 N_VGND_c_1013_n N_A_485_47#_c_1151_n 0.0116203f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_611 N_VGND_c_1007_n N_A_485_47#_c_1156_n 0.0132273f $X=5.15 $Y=0 $X2=0 $Y2=0
cc_612 N_VGND_c_1011_n N_A_485_47#_c_1156_n 0.0132487f $X=5.975 $Y=0 $X2=0 $Y2=0
cc_613 N_VGND_c_1013_n N_A_485_47#_c_1156_n 0.00827808f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_614 N_VGND_M1034_s N_A_485_47#_c_1157_n 0.00482866f $X=6.005 $Y=0.235 $X2=0
+ $Y2=0
cc_615 N_VGND_c_1011_n N_A_485_47#_c_1157_n 0.00235235f $X=5.975 $Y=0 $X2=0
+ $Y2=0
cc_616 N_VGND_c_1012_n N_A_485_47#_c_1157_n 0.00315225f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_617 N_VGND_c_1013_n N_A_485_47#_c_1157_n 0.0116364f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_618 N_VGND_c_1016_n N_A_485_47#_c_1157_n 0.023992f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_619 N_VGND_c_1012_n N_A_485_47#_c_1134_n 0.21887f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_620 N_VGND_c_1013_n N_A_485_47#_c_1134_n 0.13853f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_621 N_VGND_c_1012_n N_A_485_47#_c_1168_n 0.0296178f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_622 N_VGND_c_1013_n N_A_485_47#_c_1168_n 0.0164292f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_623 N_VGND_c_1016_n N_A_485_47#_c_1168_n 0.015242f $X=6.21 $Y=0 $X2=0 $Y2=0
