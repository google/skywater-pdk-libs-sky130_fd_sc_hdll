* File: sky130_fd_sc_hdll__o22a_4.pxi.spice
* Created: Wed Sep  2 08:45:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22A_4%A_96_21# N_A_96_21#_M1009_s N_A_96_21#_M1016_d
+ N_A_96_21#_M1003_s N_A_96_21#_M1017_s N_A_96_21#_c_104_n N_A_96_21#_M1007_g
+ N_A_96_21#_c_117_n N_A_96_21#_M1001_g N_A_96_21#_c_105_n N_A_96_21#_M1008_g
+ N_A_96_21#_c_118_n N_A_96_21#_M1005_g N_A_96_21#_c_106_n N_A_96_21#_M1014_g
+ N_A_96_21#_c_119_n N_A_96_21#_M1018_g N_A_96_21#_c_120_n N_A_96_21#_M1022_g
+ N_A_96_21#_c_107_n N_A_96_21#_M1015_g N_A_96_21#_c_108_n N_A_96_21#_c_109_n
+ N_A_96_21#_c_110_n N_A_96_21#_c_111_n N_A_96_21#_c_125_p N_A_96_21#_c_156_p
+ N_A_96_21#_c_112_n N_A_96_21#_c_113_n N_A_96_21#_c_131_p N_A_96_21#_c_114_n
+ N_A_96_21#_c_115_n N_A_96_21#_c_135_p N_A_96_21#_c_151_p N_A_96_21#_c_116_n
+ PM_SKY130_FD_SC_HDLL__O22A_4%A_96_21#
x_PM_SKY130_FD_SC_HDLL__O22A_4%B1 N_B1_c_250_n N_B1_M1013_g N_B1_c_251_n
+ N_B1_M1009_g N_B1_c_252_n N_B1_M1023_g N_B1_c_253_n N_B1_M1019_g N_B1_c_258_n
+ N_B1_c_254_n B1 B1 N_B1_c_255_n PM_SKY130_FD_SC_HDLL__O22A_4%B1
x_PM_SKY130_FD_SC_HDLL__O22A_4%B2 N_B2_c_327_n N_B2_M1010_g N_B2_c_331_n
+ N_B2_M1003_g N_B2_c_332_n N_B2_M1006_g N_B2_c_328_n N_B2_M1016_g B2
+ N_B2_c_330_n B2 PM_SKY130_FD_SC_HDLL__O22A_4%B2
x_PM_SKY130_FD_SC_HDLL__O22A_4%A1 N_A1_c_370_n N_A1_M1002_g N_A1_c_371_n
+ N_A1_M1000_g N_A1_c_372_n N_A1_M1011_g N_A1_c_373_n N_A1_M1004_g N_A1_c_380_n
+ N_A1_c_374_n N_A1_c_375_n A1 A1 PM_SKY130_FD_SC_HDLL__O22A_4%A1
x_PM_SKY130_FD_SC_HDLL__O22A_4%A2 N_A2_c_445_n N_A2_M1012_g N_A2_c_448_n
+ N_A2_M1017_g N_A2_c_449_n N_A2_M1021_g N_A2_c_446_n N_A2_M1020_g A2
+ N_A2_c_447_n A2 PM_SKY130_FD_SC_HDLL__O22A_4%A2
x_PM_SKY130_FD_SC_HDLL__O22A_4%VPWR N_VPWR_M1001_s N_VPWR_M1005_s N_VPWR_M1022_s
+ N_VPWR_M1023_s N_VPWR_M1011_s N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n
+ N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n
+ N_VPWR_c_500_n N_VPWR_c_501_n VPWR N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_491_n PM_SKY130_FD_SC_HDLL__O22A_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O22A_4%X N_X_M1007_d N_X_M1014_d N_X_M1001_d N_X_M1018_d
+ N_X_c_581_n N_X_c_582_n N_X_c_586_n N_X_c_587_n N_X_c_596_n N_X_c_628_n
+ N_X_c_588_n N_X_c_583_n N_X_c_611_n N_X_c_632_n N_X_c_584_n N_X_c_589_n X
+ PM_SKY130_FD_SC_HDLL__O22A_4%X
x_PM_SKY130_FD_SC_HDLL__O22A_4%A_614_297# N_A_614_297#_M1013_d
+ N_A_614_297#_M1006_d N_A_614_297#_c_656_n N_A_614_297#_c_660_n
+ N_A_614_297#_c_661_n PM_SKY130_FD_SC_HDLL__O22A_4%A_614_297#
x_PM_SKY130_FD_SC_HDLL__O22A_4%A_1006_297# N_A_1006_297#_M1002_d
+ N_A_1006_297#_M1021_d N_A_1006_297#_c_676_n N_A_1006_297#_c_683_n
+ N_A_1006_297#_c_679_n PM_SKY130_FD_SC_HDLL__O22A_4%A_1006_297#
x_PM_SKY130_FD_SC_HDLL__O22A_4%VGND N_VGND_M1007_s N_VGND_M1008_s N_VGND_M1015_s
+ N_VGND_M1000_d N_VGND_M1020_d N_VGND_c_692_n N_VGND_c_693_n N_VGND_c_694_n
+ N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n N_VGND_c_698_n N_VGND_c_699_n
+ N_VGND_c_700_n N_VGND_c_701_n N_VGND_c_702_n N_VGND_c_703_n N_VGND_c_704_n
+ VGND N_VGND_c_705_n N_VGND_c_706_n N_VGND_c_707_n
+ PM_SKY130_FD_SC_HDLL__O22A_4%VGND
x_PM_SKY130_FD_SC_HDLL__O22A_4%A_524_47# N_A_524_47#_M1009_d N_A_524_47#_M1010_s
+ N_A_524_47#_M1019_d N_A_524_47#_M1012_s N_A_524_47#_M1004_s
+ N_A_524_47#_c_794_n N_A_524_47#_c_846_n N_A_524_47#_c_795_n
+ N_A_524_47#_c_796_n N_A_524_47#_c_822_n N_A_524_47#_c_797_n
+ N_A_524_47#_c_798_n N_A_524_47#_c_799_n PM_SKY130_FD_SC_HDLL__O22A_4%A_524_47#
cc_1 VNB N_A_96_21#_c_104_n 0.0196598f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_2 VNB N_A_96_21#_c_105_n 0.0167602f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_3 VNB N_A_96_21#_c_106_n 0.0171978f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.995
cc_4 VNB N_A_96_21#_c_107_n 0.0200816f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.995
cc_5 VNB N_A_96_21#_c_108_n 6.30857e-19 $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=1.175
cc_6 VNB N_A_96_21#_c_109_n 6.59354e-19 $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.785
cc_7 VNB N_A_96_21#_c_110_n 0.00481211f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=1.075
cc_8 VNB N_A_96_21#_c_111_n 0.00193007f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=0.82
cc_9 VNB N_A_96_21#_c_112_n 0.002867f $X=-0.19 $Y=-0.24 $X2=2.745 $Y2=0.775
cc_10 VNB N_A_96_21#_c_113_n 0.0110516f $X=-0.19 $Y=-0.24 $X2=4.155 $Y2=0.73
cc_11 VNB N_A_96_21#_c_114_n 0.0042345f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.175
cc_12 VNB N_A_96_21#_c_115_n 0.00991332f $X=-0.19 $Y=-0.24 $X2=2.615 $Y2=0.775
cc_13 VNB N_A_96_21#_c_116_n 0.0801793f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.202
cc_14 VNB N_B1_c_250_n 0.0270532f $X=-0.19 $Y=-0.24 $X2=3.08 $Y2=0.235
cc_15 VNB N_B1_c_251_n 0.0199816f $X=-0.19 $Y=-0.24 $X2=5.5 $Y2=1.485
cc_16 VNB N_B1_c_252_n 0.0241936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_253_n 0.0180397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_c_254_n 0.00180472f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_19 VNB N_B1_c_255_n 0.00571858f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.41
cc_20 VNB N_B2_c_327_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=3.08 $Y2=0.235
cc_21 VNB N_B2_c_328_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB B2 0.00265411f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_23 VNB N_B2_c_330_n 0.0343022f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_24 VNB N_A1_c_370_n 0.0222035f $X=-0.19 $Y=-0.24 $X2=3.08 $Y2=0.235
cc_25 VNB N_A1_c_371_n 0.017338f $X=-0.19 $Y=-0.24 $X2=5.5 $Y2=1.485
cc_26 VNB N_A1_c_372_n 0.0295756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A1_c_373_n 0.0221445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A1_c_374_n 0.00395641f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.41
cc_29 VNB N_A1_c_375_n 2.74006e-19 $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_30 VNB A1 0.0022559f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.41
cc_31 VNB A1 0.0190447f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.985
cc_32 VNB N_A2_c_445_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=3.08 $Y2=0.235
cc_33 VNB N_A2_c_446_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A2_c_447_n 0.0369683f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_35 VNB N_VPWR_c_491_n 0.288713f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=1.202
cc_36 VNB N_X_c_581_n 0.0014432f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_37 VNB N_X_c_582_n 0.00986769f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.56
cc_38 VNB N_X_c_583_n 0.0052859f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.985
cc_39 VNB N_X_c_584_n 0.0025225f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.16
cc_40 VNB X 0.0213373f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.275
cc_41 VNB N_VGND_c_692_n 0.00471611f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.985
cc_42 VNB N_VGND_c_693_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.05 $Y2=1.41
cc_43 VNB N_VGND_c_694_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.56
cc_44 VNB N_VGND_c_695_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.52 $Y2=1.985
cc_45 VNB N_VGND_c_696_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.995
cc_46 VNB N_VGND_c_697_n 0.0194857f $X=-0.19 $Y=-0.24 $X2=2.1 $Y2=1.175
cc_47 VNB N_VGND_c_698_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.175
cc_48 VNB N_VGND_c_699_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_49 VNB N_VGND_c_700_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_701_n 0.064553f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.16
cc_51 VNB N_VGND_c_702_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.875 $Y2=1.16
cc_52 VNB N_VGND_c_703_n 0.0193035f $X=-0.19 $Y=-0.24 $X2=2.265 $Y2=1.785
cc_53 VNB N_VGND_c_704_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=2.285 $Y2=0.905
cc_54 VNB N_VGND_c_705_n 0.0130399f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=0.82
cc_55 VNB N_VGND_c_706_n 0.0200798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_707_n 0.339745f $X=-0.19 $Y=-0.24 $X2=5.645 $Y2=1.87
cc_57 VNB N_A_524_47#_c_794_n 0.00289463f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.41
cc_58 VNB N_A_524_47#_c_795_n 0.00343671f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.56
cc_59 VNB N_A_524_47#_c_796_n 0.00798888f $X=-0.19 $Y=-0.24 $X2=1.495 $Y2=0.56
cc_60 VNB N_A_524_47#_c_797_n 0.0135168f $X=-0.19 $Y=-0.24 $X2=1.99 $Y2=1.985
cc_61 VNB N_A_524_47#_c_798_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=2.015 $Y2=0.56
cc_62 VNB N_A_524_47#_c_799_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_63 VPB N_A_96_21#_c_117_n 0.019183f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_64 VPB N_A_96_21#_c_118_n 0.0158725f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.41
cc_65 VPB N_A_96_21#_c_119_n 0.0158895f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.41
cc_66 VPB N_A_96_21#_c_120_n 0.0191195f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.41
cc_67 VPB N_A_96_21#_c_109_n 0.00417399f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.785
cc_68 VPB N_A_96_21#_c_116_n 0.0467169f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.202
cc_69 VPB N_B1_c_250_n 0.030133f $X=-0.19 $Y=1.305 $X2=3.08 $Y2=0.235
cc_70 VPB N_B1_c_252_n 0.0257547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_B1_c_258_n 0.00726053f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_72 VPB N_B1_c_254_n 0.00224085f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_73 VPB N_B1_c_255_n 0.00307501f $X=-0.19 $Y=1.305 $X2=1.99 $Y2=1.41
cc_74 VPB N_B2_c_331_n 0.0159583f $X=-0.19 $Y=1.305 $X2=5.5 $Y2=1.485
cc_75 VPB N_B2_c_332_n 0.0159586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B2_c_330_n 0.0192444f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_77 VPB N_A1_c_370_n 0.0256643f $X=-0.19 $Y=1.305 $X2=3.08 $Y2=0.235
cc_78 VPB N_A1_c_372_n 0.0345571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A1_c_380_n 0.00607994f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_80 VPB N_A1_c_374_n 0.00272547f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_81 VPB N_A1_c_375_n 0.00131476f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_82 VPB N_A2_c_448_n 0.0159777f $X=-0.19 $Y=1.305 $X2=5.5 $Y2=1.485
cc_83 VPB N_A2_c_449_n 0.015974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A2_c_447_n 0.0192635f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=0.56
cc_85 VPB N_VPWR_c_492_n 0.0140014f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_86 VPB N_VPWR_c_493_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.985
cc_87 VPB N_VPWR_c_494_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.41
cc_88 VPB N_VPWR_c_495_n 0.00561515f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.56
cc_89 VPB N_VPWR_c_496_n 0.0121789f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.41
cc_90 VPB N_VPWR_c_497_n 0.00835273f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.985
cc_91 VPB N_VPWR_c_498_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.015 $Y2=0.56
cc_92 VPB N_VPWR_c_499_n 0.0047828f $X=-0.19 $Y=1.305 $X2=2.015 $Y2=0.56
cc_93 VPB N_VPWR_c_500_n 0.0403375f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.175
cc_94 VPB N_VPWR_c_501_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_95 VPB N_VPWR_c_502_n 0.0417635f $X=-0.19 $Y=1.305 $X2=4.155 $Y2=0.73
cc_96 VPB N_VPWR_c_503_n 0.0195604f $X=-0.19 $Y=1.305 $X2=5.645 $Y2=1.96
cc_97 VPB N_VPWR_c_504_n 0.0228965f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.202
cc_98 VPB N_VPWR_c_491_n 0.0507901f $X=-0.19 $Y=1.305 $X2=1.025 $Y2=1.202
cc_99 VPB N_X_c_586_n 0.00163065f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.56
cc_100 VPB N_X_c_587_n 0.0124524f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_101 VPB N_X_c_588_n 0.0037826f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=0.56
cc_102 VPB N_X_c_589_n 0.00150464f $X=-0.19 $Y=1.305 $X2=1.875 $Y2=1.16
cc_103 VPB X 0.00761414f $X=-0.19 $Y=1.305 $X2=2.265 $Y2=1.275
cc_104 N_A_96_21#_c_109_n N_B1_c_250_n 0.00617793f $X=2.265 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_96_21#_c_110_n N_B1_c_250_n 0.00249961f $X=2.285 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_106 N_A_96_21#_c_125_p N_B1_c_250_n 0.0156745f $X=3.56 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_96_21#_c_113_n N_B1_c_250_n 0.00441892f $X=4.155 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_108 N_A_96_21#_c_114_n N_B1_c_250_n 9.99723e-19 $X=2.265 $Y=1.175 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_96_21#_c_110_n N_B1_c_251_n 0.00229864f $X=2.285 $Y=1.075 $X2=0 $Y2=0
cc_110 N_A_96_21#_c_113_n N_B1_c_251_n 0.013855f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_111 N_A_96_21#_c_113_n N_B1_c_252_n 0.00233856f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_112 N_A_96_21#_c_131_p N_B1_c_252_n 0.0142943f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_113 N_A_96_21#_M1003_s N_B1_c_258_n 0.00187091f $X=3.54 $Y=1.485 $X2=0 $Y2=0
cc_114 N_A_96_21#_c_113_n N_B1_c_258_n 0.0118424f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_115 N_A_96_21#_c_131_p N_B1_c_258_n 0.0389168f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_116 N_A_96_21#_c_135_p N_B1_c_258_n 0.0135474f $X=3.685 $Y=1.87 $X2=0 $Y2=0
cc_117 N_A_96_21#_c_113_n N_B1_c_254_n 0.00976394f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_118 N_A_96_21#_c_109_n N_B1_c_255_n 0.0270316f $X=2.265 $Y=1.785 $X2=0 $Y2=0
cc_119 N_A_96_21#_c_125_p N_B1_c_255_n 0.0555873f $X=3.56 $Y=1.87 $X2=0 $Y2=0
cc_120 N_A_96_21#_c_112_n N_B1_c_255_n 0.0455576f $X=2.745 $Y=0.775 $X2=0 $Y2=0
cc_121 N_A_96_21#_c_114_n N_B1_c_255_n 0.0169778f $X=2.265 $Y=1.175 $X2=0 $Y2=0
cc_122 N_A_96_21#_c_116_n N_B1_c_255_n 9.87003e-19 $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_123 N_A_96_21#_c_113_n N_B2_c_327_n 0.0118103f $X=4.155 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_124 N_A_96_21#_c_125_p N_B2_c_331_n 0.0108425f $X=3.56 $Y=1.87 $X2=0 $Y2=0
cc_125 N_A_96_21#_c_131_p N_B2_c_332_n 0.0108425f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_126 N_A_96_21#_c_113_n N_B2_c_328_n 0.0118103f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_127 N_A_96_21#_c_113_n B2 0.0497757f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_128 N_A_96_21#_c_113_n N_B2_c_330_n 0.0047334f $X=4.155 $Y=0.73 $X2=0 $Y2=0
cc_129 N_A_96_21#_c_131_p N_A1_c_370_n 0.0140422f $X=5.52 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_96_21#_M1017_s N_A1_c_380_n 0.00187091f $X=5.5 $Y=1.485 $X2=0 $Y2=0
cc_131 N_A_96_21#_c_131_p N_A1_c_380_n 0.0218268f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_132 N_A_96_21#_c_151_p N_A1_c_380_n 0.0135474f $X=5.645 $Y=1.87 $X2=0 $Y2=0
cc_133 N_A_96_21#_c_131_p N_A1_c_374_n 0.0233516f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_134 N_A_96_21#_c_131_p N_A2_c_448_n 0.0108425f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_135 N_A_96_21#_c_109_n N_VPWR_M1022_s 0.00885389f $X=2.265 $Y=1.785 $X2=0
+ $Y2=0
cc_136 N_A_96_21#_c_125_p N_VPWR_M1022_s 0.0162575f $X=3.56 $Y=1.87 $X2=0 $Y2=0
cc_137 N_A_96_21#_c_156_p N_VPWR_M1022_s 0.00593207f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_138 N_A_96_21#_c_131_p N_VPWR_M1023_s 0.00987581f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_139 N_A_96_21#_c_117_n N_VPWR_c_493_n 0.00479105f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_96_21#_c_118_n N_VPWR_c_494_n 0.00300743f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_96_21#_c_119_n N_VPWR_c_494_n 0.00300743f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_96_21#_c_131_p N_VPWR_c_495_n 0.020234f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_143 N_A_96_21#_c_117_n N_VPWR_c_498_n 0.00702461f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_96_21#_c_118_n N_VPWR_c_498_n 0.00702461f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_96_21#_c_119_n N_VPWR_c_503_n 0.00702461f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_96_21#_c_120_n N_VPWR_c_503_n 0.00702461f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_96_21#_c_120_n N_VPWR_c_504_n 0.00514457f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_96_21#_c_125_p N_VPWR_c_504_n 0.0316562f $X=3.56 $Y=1.87 $X2=0 $Y2=0
cc_149 N_A_96_21#_c_156_p N_VPWR_c_504_n 0.0254138f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_150 N_A_96_21#_M1003_s N_VPWR_c_491_n 0.00231289f $X=3.54 $Y=1.485 $X2=0
+ $Y2=0
cc_151 N_A_96_21#_M1017_s N_VPWR_c_491_n 0.00232092f $X=5.5 $Y=1.485 $X2=0 $Y2=0
cc_152 N_A_96_21#_c_117_n N_VPWR_c_491_n 0.0133906f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_96_21#_c_118_n N_VPWR_c_491_n 0.0124092f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_96_21#_c_119_n N_VPWR_c_491_n 0.0124092f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_96_21#_c_120_n N_VPWR_c_491_n 0.0136891f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_96_21#_c_125_p N_VPWR_c_491_n 0.00923942f $X=3.56 $Y=1.87 $X2=0 $Y2=0
cc_157 N_A_96_21#_c_156_p N_VPWR_c_491_n 0.00133688f $X=2.43 $Y=1.87 $X2=0 $Y2=0
cc_158 N_A_96_21#_c_131_p N_VPWR_c_491_n 0.0165728f $X=5.52 $Y=1.87 $X2=0 $Y2=0
cc_159 N_A_96_21#_c_104_n N_X_c_581_n 0.0111251f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_96_21#_c_108_n N_X_c_581_n 0.00410208f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_161 N_A_96_21#_c_117_n N_X_c_586_n 0.0178749f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_96_21#_c_108_n N_X_c_586_n 0.0103328f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_163 N_A_96_21#_c_116_n N_X_c_586_n 9.44081e-19 $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_164 N_A_96_21#_c_104_n N_X_c_596_n 0.0109499f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_96_21#_c_105_n N_X_c_596_n 0.00676224f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_96_21#_c_106_n N_X_c_596_n 5.42233e-19 $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_96_21#_c_118_n N_X_c_588_n 0.0157513f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_96_21#_c_119_n N_X_c_588_n 0.015669f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_96_21#_c_120_n N_X_c_588_n 4.00176e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_96_21#_c_108_n N_X_c_588_n 0.0689039f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_171 N_A_96_21#_c_109_n N_X_c_588_n 0.00287394f $X=2.265 $Y=1.785 $X2=0 $Y2=0
cc_172 N_A_96_21#_c_116_n N_X_c_588_n 0.0151889f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_173 N_A_96_21#_c_105_n N_X_c_583_n 0.00901745f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_96_21#_c_106_n N_X_c_583_n 0.010179f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_96_21#_c_107_n N_X_c_583_n 2.14781e-19 $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_96_21#_c_108_n N_X_c_583_n 0.0704813f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_177 N_A_96_21#_c_111_n N_X_c_583_n 0.00148154f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_178 N_A_96_21#_c_116_n N_X_c_583_n 0.00831812f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_179 N_A_96_21#_c_105_n N_X_c_611_n 5.24597e-19 $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_96_21#_c_106_n N_X_c_611_n 0.00651696f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_96_21#_c_104_n N_X_c_584_n 0.00116607f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_96_21#_c_105_n N_X_c_584_n 0.00116607f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_96_21#_c_108_n N_X_c_584_n 0.0305614f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_184 N_A_96_21#_c_116_n N_X_c_584_n 0.00358132f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_185 N_A_96_21#_c_108_n N_X_c_589_n 0.020385f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_186 N_A_96_21#_c_116_n N_X_c_589_n 0.00664519f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_187 N_A_96_21#_c_104_n X 0.0186818f $X=0.555 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_96_21#_c_117_n X 0.00133332f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_96_21#_c_108_n X 0.0164324f $X=2.1 $Y=1.175 $X2=0 $Y2=0
cc_190 N_A_96_21#_c_125_p N_A_614_297#_M1013_d 0.00369247f $X=3.56 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_191 N_A_96_21#_c_131_p N_A_614_297#_M1006_d 0.00369141f $X=5.52 $Y=1.87 $X2=0
+ $Y2=0
cc_192 N_A_96_21#_M1003_s N_A_614_297#_c_656_n 0.00352392f $X=3.54 $Y=1.485
+ $X2=0 $Y2=0
cc_193 N_A_96_21#_c_125_p N_A_614_297#_c_656_n 0.00608347f $X=3.56 $Y=1.87 $X2=0
+ $Y2=0
cc_194 N_A_96_21#_c_131_p N_A_614_297#_c_656_n 0.00608347f $X=5.52 $Y=1.87 $X2=0
+ $Y2=0
cc_195 N_A_96_21#_c_135_p N_A_614_297#_c_656_n 0.0127274f $X=3.685 $Y=1.87 $X2=0
+ $Y2=0
cc_196 N_A_96_21#_c_125_p N_A_614_297#_c_660_n 0.0131392f $X=3.56 $Y=1.87 $X2=0
+ $Y2=0
cc_197 N_A_96_21#_c_131_p N_A_614_297#_c_661_n 0.0131392f $X=5.52 $Y=1.87 $X2=0
+ $Y2=0
cc_198 N_A_96_21#_c_131_p N_A_1006_297#_M1002_d 0.00367036f $X=5.52 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_199 N_A_96_21#_M1017_s N_A_1006_297#_c_676_n 0.00352392f $X=5.5 $Y=1.485
+ $X2=0 $Y2=0
cc_200 N_A_96_21#_c_131_p N_A_1006_297#_c_676_n 0.00608347f $X=5.52 $Y=1.87
+ $X2=0 $Y2=0
cc_201 N_A_96_21#_c_151_p N_A_1006_297#_c_676_n 0.0127274f $X=5.645 $Y=1.87
+ $X2=0 $Y2=0
cc_202 N_A_96_21#_c_131_p N_A_1006_297#_c_679_n 0.0130645f $X=5.52 $Y=1.87 $X2=0
+ $Y2=0
cc_203 N_A_96_21#_c_111_n N_VGND_M1015_s 0.00429247f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_204 N_A_96_21#_c_104_n N_VGND_c_692_n 0.00438629f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_96_21#_c_105_n N_VGND_c_693_n 0.00394736f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_96_21#_c_106_n N_VGND_c_693_n 0.00276126f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_96_21#_c_107_n N_VGND_c_694_n 0.00438629f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_96_21#_c_111_n N_VGND_c_694_n 0.0133599f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_209 N_A_96_21#_c_104_n N_VGND_c_697_n 0.00423737f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_96_21#_c_105_n N_VGND_c_697_n 0.00423737f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_96_21#_c_106_n N_VGND_c_699_n 0.00423334f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_212 N_A_96_21#_c_107_n N_VGND_c_699_n 0.00585385f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_96_21#_c_111_n N_VGND_c_701_n 0.00195943f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_214 N_A_96_21#_c_115_n N_VGND_c_701_n 0.00223545f $X=2.615 $Y=0.775 $X2=0
+ $Y2=0
cc_215 N_A_96_21#_M1009_s N_VGND_c_707_n 0.00216833f $X=3.08 $Y=0.235 $X2=0
+ $Y2=0
cc_216 N_A_96_21#_M1016_d N_VGND_c_707_n 0.00256987f $X=4.02 $Y=0.235 $X2=0
+ $Y2=0
cc_217 N_A_96_21#_c_104_n N_VGND_c_707_n 0.00687004f $X=0.555 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_96_21#_c_105_n N_VGND_c_707_n 0.0060934f $X=1.025 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_96_21#_c_106_n N_VGND_c_707_n 0.00608558f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_220 N_A_96_21#_c_107_n N_VGND_c_707_n 0.0121055f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_96_21#_c_111_n N_VGND_c_707_n 0.00413086f $X=2.43 $Y=0.82 $X2=0 $Y2=0
cc_222 N_A_96_21#_c_115_n N_VGND_c_707_n 0.004011f $X=2.615 $Y=0.775 $X2=0 $Y2=0
cc_223 N_A_96_21#_c_112_n N_A_524_47#_M1009_d 0.00295421f $X=2.745 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_224 N_A_96_21#_c_113_n N_A_524_47#_M1009_d 0.00137434f $X=4.155 $Y=0.73
+ $X2=-0.19 $Y2=-0.24
cc_225 N_A_96_21#_c_113_n N_A_524_47#_M1010_s 0.00279596f $X=4.155 $Y=0.73 $X2=0
+ $Y2=0
cc_226 N_A_96_21#_M1009_s N_A_524_47#_c_794_n 0.00312026f $X=3.08 $Y=0.235 $X2=0
+ $Y2=0
cc_227 N_A_96_21#_M1016_d N_A_524_47#_c_794_n 0.0041027f $X=4.02 $Y=0.235 $X2=0
+ $Y2=0
cc_228 N_A_96_21#_c_112_n N_A_524_47#_c_794_n 0.0939413f $X=2.745 $Y=0.775 $X2=0
+ $Y2=0
cc_229 N_A_96_21#_c_115_n N_A_524_47#_c_794_n 0.0018027f $X=2.615 $Y=0.775 $X2=0
+ $Y2=0
cc_230 N_A_96_21#_c_113_n N_A_524_47#_c_796_n 0.00140356f $X=4.155 $Y=0.73 $X2=0
+ $Y2=0
cc_231 N_B1_c_251_n N_B2_c_327_n 0.0270078f $X=3.005 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_232 N_B1_c_250_n N_B2_c_331_n 0.0378435f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B1_c_258_n N_B2_c_331_n 0.011867f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_234 N_B1_c_255_n N_B2_c_331_n 9.10997e-19 $X=3.18 $Y=1.345 $X2=0 $Y2=0
cc_235 N_B1_c_252_n N_B2_c_332_n 0.0378464f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B1_c_258_n N_B2_c_332_n 0.011867f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_237 N_B1_c_254_n N_B2_c_332_n 7.94204e-19 $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_238 N_B1_c_253_n N_B2_c_328_n 0.0219899f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B1_c_250_n B2 2.26386e-19 $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B1_c_252_n B2 6.9147e-19 $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B1_c_258_n B2 0.047909f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B1_c_254_n B2 0.0175463f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B1_c_255_n B2 0.0173858f $X=3.18 $Y=1.345 $X2=0 $Y2=0
cc_244 N_B1_c_250_n N_B2_c_330_n 0.0262945f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B1_c_252_n N_B2_c_330_n 0.0263033f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B1_c_258_n N_B2_c_330_n 0.00798993f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_247 N_B1_c_254_n N_B2_c_330_n 0.00383981f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_248 N_B1_c_255_n N_B2_c_330_n 0.0042972f $X=3.18 $Y=1.345 $X2=0 $Y2=0
cc_249 N_B1_c_252_n N_A1_c_370_n 0.0562911f $X=4.39 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_250 N_B1_c_258_n N_A1_c_370_n 5.2512e-19 $X=4.2 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_251 N_B1_c_254_n N_A1_c_370_n 5.96767e-19 $X=4.365 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_252 N_B1_c_253_n N_A1_c_371_n 0.0154445f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B1_c_252_n N_A1_c_374_n 0.00252166f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B1_c_258_n N_A1_c_374_n 0.0148627f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_255 N_B1_c_254_n N_A1_c_374_n 0.0303702f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_255_n N_VPWR_M1022_s 0.00421583f $X=3.18 $Y=1.345 $X2=0 $Y2=0
cc_257 N_B1_c_258_n N_VPWR_M1023_s 0.00118581f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_258 N_B1_c_252_n N_VPWR_c_495_n 0.00322023f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B1_c_250_n N_VPWR_c_500_n 0.00702461f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B1_c_252_n N_VPWR_c_500_n 0.00702461f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B1_c_250_n N_VPWR_c_504_n 0.00514457f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B1_c_250_n N_VPWR_c_491_n 0.00823967f $X=2.98 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B1_c_252_n N_VPWR_c_491_n 0.00716301f $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B1_c_258_n N_A_614_297#_M1013_d 0.00130005f $X=4.2 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_265 N_B1_c_255_n N_A_614_297#_M1013_d 5.85197e-19 $X=3.18 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_266 N_B1_c_258_n N_A_614_297#_M1006_d 0.00186927f $X=4.2 $Y=1.53 $X2=0 $Y2=0
cc_267 N_B1_c_251_n N_VGND_c_694_n 0.00179926f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B1_c_251_n N_VGND_c_701_n 0.00357877f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B1_c_253_n N_VGND_c_701_n 0.00357877f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B1_c_251_n N_VGND_c_707_n 0.00657948f $X=3.005 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B1_c_253_n N_VGND_c_707_n 0.00568976f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B1_c_251_n N_A_524_47#_c_794_n 0.00886996f $X=3.005 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_B1_c_252_n N_A_524_47#_c_794_n 3.99938e-19 $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_253_n N_A_524_47#_c_794_n 0.0112894f $X=4.415 $Y=0.995 $X2=0 $Y2=0
cc_275 N_B1_c_254_n N_A_524_47#_c_794_n 0.004983f $X=4.365 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B1_c_252_n N_A_524_47#_c_796_n 4.78733e-19 $X=4.39 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_253_n N_A_524_47#_c_796_n 2.31743e-19 $X=4.415 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_B2_c_331_n N_VPWR_c_500_n 0.00429453f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B2_c_332_n N_VPWR_c_500_n 0.00429453f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_280 N_B2_c_331_n N_VPWR_c_491_n 0.00609021f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B2_c_332_n N_VPWR_c_491_n 0.00609021f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B2_c_331_n N_A_614_297#_c_656_n 0.0099733f $X=3.45 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B2_c_332_n N_A_614_297#_c_656_n 0.0099733f $X=3.92 $Y=1.41 $X2=0 $Y2=0
cc_284 N_B2_c_327_n N_VGND_c_701_n 0.00357877f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B2_c_328_n N_VGND_c_701_n 0.00357877f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B2_c_327_n N_VGND_c_707_n 0.00549573f $X=3.425 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_328_n N_VGND_c_707_n 0.00561849f $X=3.945 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_327_n N_A_524_47#_c_794_n 0.00886996f $X=3.425 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_B2_c_328_n N_A_524_47#_c_794_n 0.00923997f $X=3.945 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A1_c_371_n N_A2_c_445_n 0.0258911f $X=4.965 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_291 N_A1_c_370_n N_A2_c_448_n 0.0378352f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A1_c_380_n N_A2_c_448_n 0.0116479f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_293 N_A1_c_374_n N_A2_c_448_n 0.00103157f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A1_c_372_n N_A2_c_449_n 0.0219395f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A1_c_380_n N_A2_c_449_n 0.0181096f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_296 N_A1_c_375_n N_A2_c_449_n 8.03195e-19 $X=6.18 $Y=1.445 $X2=0 $Y2=0
cc_297 N_A1_c_373_n N_A2_c_446_n 0.0213001f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A1_c_370_n A2 2.20437e-19 $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A1_c_380_n A2 0.0391785f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_300 N_A1_c_374_n A2 0.013729f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_301 A1 A2 0.0173958f $X=6.24 $Y=1.105 $X2=0 $Y2=0
cc_302 N_A1_c_370_n N_A2_c_447_n 0.0264727f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A1_c_372_n N_A2_c_447_n 0.0262388f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A1_c_380_n N_A2_c_447_n 0.00808788f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_305 N_A1_c_374_n N_A2_c_447_n 0.00472925f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A1_c_375_n N_A2_c_447_n 0.00319804f $X=6.18 $Y=1.445 $X2=0 $Y2=0
cc_307 A1 N_A2_c_447_n 0.00159526f $X=6.24 $Y=1.105 $X2=0 $Y2=0
cc_308 N_A1_c_374_n N_VPWR_M1023_s 0.00204417f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A1_c_370_n N_VPWR_c_495_n 0.00537492f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A1_c_372_n N_VPWR_c_497_n 0.0122183f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A1_c_380_n N_VPWR_c_497_n 0.0104762f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_312 A1 N_VPWR_c_497_n 0.0166332f $X=6.335 $Y=1.19 $X2=0 $Y2=0
cc_313 N_A1_c_370_n N_VPWR_c_502_n 0.00702461f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A1_c_372_n N_VPWR_c_502_n 0.00702461f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A1_c_370_n N_VPWR_c_491_n 0.00721773f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A1_c_372_n N_VPWR_c_491_n 0.013506f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A1_c_380_n N_A_1006_297#_M1002_d 0.00172342f $X=6.075 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_318 N_A1_c_374_n N_A_1006_297#_M1002_d 7.76441e-19 $X=4.915 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_319 N_A1_c_380_n N_A_1006_297#_M1021_d 0.00190617f $X=6.075 $Y=1.53 $X2=0
+ $Y2=0
cc_320 N_A1_c_380_n N_A_1006_297#_c_683_n 0.0152155f $X=6.075 $Y=1.53 $X2=0
+ $Y2=0
cc_321 N_A1_c_371_n N_VGND_c_695_n 0.00268723f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A1_c_373_n N_VGND_c_696_n 0.00359159f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A1_c_371_n N_VGND_c_701_n 0.00439206f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A1_c_373_n N_VGND_c_706_n 0.00396605f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A1_c_371_n N_VGND_c_707_n 0.00630876f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A1_c_373_n N_VGND_c_707_n 0.00670929f $X=6.375 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A1_c_370_n N_A_524_47#_c_795_n 0.00205406f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A1_c_371_n N_A_524_47#_c_795_n 0.0124528f $X=4.965 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A1_c_380_n N_A_524_47#_c_795_n 0.00717126f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_330 N_A1_c_374_n N_A_524_47#_c_795_n 0.0198504f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A1_c_370_n N_A_524_47#_c_796_n 0.00239959f $X=4.94 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A1_c_374_n N_A_524_47#_c_796_n 0.0141964f $X=4.915 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A1_c_371_n N_A_524_47#_c_822_n 5.32212e-19 $X=4.965 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A1_c_372_n N_A_524_47#_c_797_n 0.00443298f $X=6.35 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A1_c_373_n N_A_524_47#_c_797_n 0.00903373f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_336 N_A1_c_380_n N_A_524_47#_c_797_n 0.00522345f $X=6.075 $Y=1.53 $X2=0 $Y2=0
cc_337 A1 N_A_524_47#_c_797_n 0.0170528f $X=6.24 $Y=1.105 $X2=0 $Y2=0
cc_338 A1 N_A_524_47#_c_797_n 0.0372828f $X=6.335 $Y=1.19 $X2=0 $Y2=0
cc_339 N_A1_c_373_n N_A_524_47#_c_798_n 0.00850899f $X=6.375 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A2_c_448_n N_VPWR_c_502_n 0.00429453f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A2_c_449_n N_VPWR_c_502_n 0.00429453f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A2_c_448_n N_VPWR_c_491_n 0.00609021f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A2_c_449_n N_VPWR_c_491_n 0.00609021f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A2_c_448_n N_A_1006_297#_c_676_n 0.0100164f $X=5.41 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A2_c_449_n N_A_1006_297#_c_676_n 0.0143148f $X=5.88 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A2_c_445_n N_VGND_c_695_n 0.00268723f $X=5.385 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A2_c_446_n N_VGND_c_696_n 0.00276126f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A2_c_445_n N_VGND_c_703_n 0.00424416f $X=5.385 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A2_c_446_n N_VGND_c_703_n 0.00437852f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A2_c_445_n N_VGND_c_707_n 0.00600559f $X=5.385 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A2_c_446_n N_VGND_c_707_n 0.00627444f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A2_c_445_n N_A_524_47#_c_795_n 0.00891961f $X=5.385 $Y=0.995 $X2=0
+ $Y2=0
cc_353 A2 N_A_524_47#_c_795_n 0.00545718f $X=5.725 $Y=1.105 $X2=0 $Y2=0
cc_354 N_A2_c_445_n N_A_524_47#_c_822_n 0.00644736f $X=5.385 $Y=0.995 $X2=0
+ $Y2=0
cc_355 N_A2_c_446_n N_A_524_47#_c_797_n 0.0118054f $X=5.905 $Y=0.995 $X2=0 $Y2=0
cc_356 A2 N_A_524_47#_c_797_n 0.00658691f $X=5.725 $Y=1.105 $X2=0 $Y2=0
cc_357 N_A2_c_446_n N_A_524_47#_c_798_n 5.82315e-19 $X=5.905 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A2_c_445_n N_A_524_47#_c_799_n 0.00135102f $X=5.385 $Y=0.995 $X2=0
+ $Y2=0
cc_359 A2 N_A_524_47#_c_799_n 0.0307352f $X=5.725 $Y=1.105 $X2=0 $Y2=0
cc_360 N_A2_c_447_n N_A_524_47#_c_799_n 0.00486271f $X=5.88 $Y=1.202 $X2=0 $Y2=0
cc_361 N_VPWR_c_491_n N_X_M1001_d 0.00370124f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_362 N_VPWR_c_491_n N_X_M1018_d 0.00370124f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_363 N_VPWR_M1001_s N_X_c_586_n 7.22239e-19 $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_364 N_VPWR_c_493_n N_X_c_586_n 0.00434858f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_365 N_VPWR_M1001_s N_X_c_587_n 0.00354732f $X=0.2 $Y=1.485 $X2=0 $Y2=0
cc_366 N_VPWR_c_493_n N_X_c_587_n 0.011469f $X=0.345 $Y=1.99 $X2=0 $Y2=0
cc_367 N_VPWR_c_498_n N_X_c_628_n 0.0149311f $X=1.16 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_491_n N_X_c_628_n 0.00955092f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_M1005_s N_X_c_588_n 0.00191634f $X=1.14 $Y=1.485 $X2=0 $Y2=0
cc_370 N_VPWR_c_494_n N_X_c_588_n 0.0137198f $X=1.285 $Y=1.99 $X2=0 $Y2=0
cc_371 N_VPWR_c_503_n N_X_c_632_n 0.0149311f $X=2.1 $Y=2.465 $X2=0 $Y2=0
cc_372 N_VPWR_c_491_n N_X_c_632_n 0.00955092f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_c_491_n N_A_614_297#_M1013_d 0.00241598f $X=6.67 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_374 N_VPWR_c_491_n N_A_614_297#_M1006_d 0.00241598f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_500_n N_A_614_297#_c_656_n 0.0386815f $X=4.5 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_491_n N_A_614_297#_c_656_n 0.0239224f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_500_n N_A_614_297#_c_660_n 0.014332f $X=4.5 $Y=2.72 $X2=0 $Y2=0
cc_378 N_VPWR_c_491_n N_A_614_297#_c_660_n 0.00938745f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_500_n N_A_614_297#_c_661_n 0.014332f $X=4.5 $Y=2.72 $X2=0 $Y2=0
cc_380 N_VPWR_c_491_n N_A_614_297#_c_661_n 0.00938745f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_491_n N_A_1006_297#_M1002_d 0.00241598f $X=6.67 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_382 N_VPWR_c_491_n N_A_1006_297#_M1021_d 0.00297222f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_502_n N_A_1006_297#_c_676_n 0.0536835f $X=6.505 $Y=2.72 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_491_n N_A_1006_297#_c_676_n 0.0335464f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_502_n N_A_1006_297#_c_679_n 0.0143006f $X=6.505 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_491_n N_A_1006_297#_c_679_n 0.00938288f $X=6.67 $Y=2.72 $X2=0
+ $Y2=0
cc_387 N_X_c_581_n N_VGND_M1007_s 5.40298e-19 $X=0.6 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_388 N_X_c_582_n N_VGND_M1007_s 0.00329182f $X=0.37 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_389 N_X_c_583_n N_VGND_M1008_s 0.00251047f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_390 N_X_c_581_n N_VGND_c_692_n 0.00402428f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_391 N_X_c_582_n N_VGND_c_692_n 0.00920832f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_392 N_X_c_596_n N_VGND_c_693_n 0.0177507f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_393 N_X_c_583_n N_VGND_c_693_n 0.0127273f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_394 N_X_c_596_n N_VGND_c_697_n 0.0210053f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_395 N_X_c_583_n N_VGND_c_697_n 0.00266636f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_396 N_X_c_583_n N_VGND_c_699_n 0.00198695f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_397 N_X_c_611_n N_VGND_c_699_n 0.0231806f $X=1.755 $Y=0.39 $X2=0 $Y2=0
cc_398 N_X_c_581_n N_VGND_c_705_n 0.0019947f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_399 N_X_c_582_n N_VGND_c_705_n 0.00293744f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_400 N_X_M1007_d N_VGND_c_707_n 0.00255747f $X=0.63 $Y=0.235 $X2=0 $Y2=0
cc_401 N_X_M1014_d N_VGND_c_707_n 0.00364931f $X=1.57 $Y=0.235 $X2=0 $Y2=0
cc_402 N_X_c_581_n N_VGND_c_707_n 0.00407016f $X=0.6 $Y=0.815 $X2=0 $Y2=0
cc_403 N_X_c_582_n N_VGND_c_707_n 0.00542613f $X=0.37 $Y=0.815 $X2=0 $Y2=0
cc_404 N_X_c_596_n N_VGND_c_707_n 0.0140539f $X=0.815 $Y=0.39 $X2=0 $Y2=0
cc_405 N_X_c_583_n N_VGND_c_707_n 0.00972452f $X=1.54 $Y=0.815 $X2=0 $Y2=0
cc_406 N_X_c_611_n N_VGND_c_707_n 0.0143352f $X=1.755 $Y=0.39 $X2=0 $Y2=0
cc_407 N_VGND_c_707_n N_A_524_47#_M1009_d 0.00250339f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_408 N_VGND_c_707_n N_A_524_47#_M1010_s 0.00295535f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_707_n N_A_524_47#_M1019_d 0.00330638f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_c_707_n N_A_524_47#_M1012_s 0.00304143f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_411 N_VGND_c_707_n N_A_524_47#_M1004_s 0.00209319f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_412 N_VGND_c_694_n N_A_524_47#_c_794_n 0.0130084f $X=2.225 $Y=0.39 $X2=0
+ $Y2=0
cc_413 N_VGND_c_701_n N_A_524_47#_c_794_n 0.112077f $X=5.09 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_707_n N_A_524_47#_c_794_n 0.0703895f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_701_n N_A_524_47#_c_846_n 0.0216064f $X=5.09 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_707_n N_A_524_47#_c_846_n 0.0126938f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_417 N_VGND_M1000_d N_A_524_47#_c_795_n 0.00165819f $X=5.04 $Y=0.235 $X2=0
+ $Y2=0
cc_418 N_VGND_c_695_n N_A_524_47#_c_795_n 0.0116528f $X=5.175 $Y=0.39 $X2=0
+ $Y2=0
cc_419 N_VGND_c_701_n N_A_524_47#_c_795_n 0.00248756f $X=5.09 $Y=0 $X2=0 $Y2=0
cc_420 N_VGND_c_703_n N_A_524_47#_c_795_n 0.00193763f $X=6.03 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_707_n N_A_524_47#_c_795_n 0.00943347f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_703_n N_A_524_47#_c_822_n 0.0231806f $X=6.03 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_707_n N_A_524_47#_c_822_n 0.0143352f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_M1020_d N_A_524_47#_c_797_n 0.00251047f $X=5.98 $Y=0.235 $X2=0
+ $Y2=0
cc_425 N_VGND_c_696_n N_A_524_47#_c_797_n 0.0127273f $X=6.115 $Y=0.39 $X2=0
+ $Y2=0
cc_426 N_VGND_c_703_n N_A_524_47#_c_797_n 0.00254521f $X=6.03 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_706_n N_A_524_47#_c_797_n 0.00199443f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_707_n N_A_524_47#_c_797_n 0.00977515f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_429 N_VGND_c_696_n N_A_524_47#_c_798_n 0.0223967f $X=6.115 $Y=0.39 $X2=0
+ $Y2=0
cc_430 N_VGND_c_706_n N_A_524_47#_c_798_n 0.024373f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_707_n N_A_524_47#_c_798_n 0.0141066f $X=6.67 $Y=0 $X2=0 $Y2=0
