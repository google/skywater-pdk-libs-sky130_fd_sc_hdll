* File: sky130_fd_sc_hdll__o22a_2.pxi.spice
* Created: Thu Aug 27 19:21:07 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22A_2%A_83_21# N_A_83_21#_M1011_d N_A_83_21#_M1007_d
+ N_A_83_21#_c_58_n N_A_83_21#_M1006_g N_A_83_21#_c_65_n N_A_83_21#_M1001_g
+ N_A_83_21#_c_59_n N_A_83_21#_M1009_g N_A_83_21#_c_66_n N_A_83_21#_M1010_g
+ N_A_83_21#_c_60_n N_A_83_21#_c_61_n N_A_83_21#_c_68_n N_A_83_21#_c_98_p
+ N_A_83_21#_c_75_p N_A_83_21#_c_62_n N_A_83_21#_c_69_n N_A_83_21#_c_73_p
+ N_A_83_21#_c_63_n N_A_83_21#_c_64_n PM_SKY130_FD_SC_HDLL__O22A_2%A_83_21#
x_PM_SKY130_FD_SC_HDLL__O22A_2%B1 N_B1_c_145_n N_B1_M1005_g N_B1_c_142_n
+ N_B1_M1011_g B1 N_B1_c_144_n PM_SKY130_FD_SC_HDLL__O22A_2%B1
x_PM_SKY130_FD_SC_HDLL__O22A_2%B2 N_B2_c_173_n N_B2_M1007_g N_B2_c_174_n
+ N_B2_M1000_g B2 B2 PM_SKY130_FD_SC_HDLL__O22A_2%B2
x_PM_SKY130_FD_SC_HDLL__O22A_2%A2 N_A2_c_206_n N_A2_M1002_g N_A2_c_207_n
+ N_A2_M1008_g N_A2_c_208_n A2 PM_SKY130_FD_SC_HDLL__O22A_2%A2
x_PM_SKY130_FD_SC_HDLL__O22A_2%A1 N_A1_c_242_n N_A1_M1003_g N_A1_c_243_n
+ N_A1_M1004_g A1 A1 N_A1_c_244_n PM_SKY130_FD_SC_HDLL__O22A_2%A1
x_PM_SKY130_FD_SC_HDLL__O22A_2%VPWR N_VPWR_M1001_s N_VPWR_M1010_s N_VPWR_M1003_d
+ N_VPWR_c_266_n N_VPWR_c_267_n N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n
+ VPWR N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_265_n VPWR
+ PM_SKY130_FD_SC_HDLL__O22A_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O22A_2%X N_X_M1006_d N_X_M1001_d X N_X_c_311_n
+ PM_SKY130_FD_SC_HDLL__O22A_2%X
x_PM_SKY130_FD_SC_HDLL__O22A_2%VGND N_VGND_M1006_s N_VGND_M1009_s N_VGND_M1008_d
+ N_VGND_c_331_n N_VGND_c_332_n N_VGND_c_333_n N_VGND_c_334_n N_VGND_c_335_n
+ N_VGND_c_336_n N_VGND_c_337_n VGND N_VGND_c_338_n N_VGND_c_339_n
+ N_VGND_c_340_n VGND PM_SKY130_FD_SC_HDLL__O22A_2%VGND
x_PM_SKY130_FD_SC_HDLL__O22A_2%A_321_47# N_A_321_47#_M1011_s N_A_321_47#_M1000_d
+ N_A_321_47#_M1004_d N_A_321_47#_c_387_n N_A_321_47#_c_402_n
+ N_A_321_47#_c_394_n N_A_321_47#_c_388_n N_A_321_47#_c_389_n
+ PM_SKY130_FD_SC_HDLL__O22A_2%A_321_47#
cc_1 VNB N_A_83_21#_c_58_n 0.0223286f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_83_21#_c_59_n 0.0195121f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_3 VNB N_A_83_21#_c_60_n 0.00205011f $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.16
cc_4 VNB N_A_83_21#_c_61_n 4.23622e-19 $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=0.805
cc_5 VNB N_A_83_21#_c_62_n 0.00237603f $X=-0.19 $Y=-0.24 $X2=2.2 $Y2=0.73
cc_6 VNB N_A_83_21#_c_63_n 0.00931156f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.77
cc_7 VNB N_A_83_21#_c_64_n 0.0687335f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_8 VNB N_B1_c_142_n 0.0201528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB B1 0.00241597f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_10 VNB N_B1_c_144_n 0.0325403f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_11 VNB N_B2_c_173_n 0.0231649f $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=0.235
cc_12 VNB N_B2_c_174_n 0.018309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB B2 0.0061543f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.56
cc_14 VNB N_A2_c_206_n 0.023292f $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=0.235
cc_15 VNB N_A2_c_207_n 0.018564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A2_c_208_n 0.00314359f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_17 VNB N_A1_c_242_n 0.0384064f $X=-0.19 $Y=-0.24 $X2=2.065 $Y2=0.235
cc_18 VNB N_A1_c_243_n 0.0224126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_244_n 0.00151051f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.995
cc_20 VNB N_VPWR_c_265_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_311_n 0.0017201f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_22 VNB N_VGND_c_331_n 0.0113721f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_23 VNB N_VGND_c_332_n 0.00739463f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_24 VNB N_VGND_c_333_n 0.0223721f $X=-0.19 $Y=-0.24 $X2=0.95 $Y2=0.56
cc_25 VNB N_VGND_c_334_n 0.00479834f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.985
cc_26 VNB N_VGND_c_335_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.16
cc_27 VNB N_VGND_c_336_n 0.0461994f $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=0.805
cc_28 VNB N_VGND_c_337_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=2.34 $Y2=1.58
cc_29 VNB N_VGND_c_338_n 0.023064f $X=-0.19 $Y=-0.24 $X2=2.517 $Y2=1.58
cc_30 VNB N_VGND_c_339_n 0.230662f $X=-0.19 $Y=-0.24 $X2=2.61 $Y2=1.62
cc_31 VNB N_VGND_c_340_n 0.00343497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_321_47#_c_387_n 0.00248799f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_33 VNB N_A_321_47#_c_388_n 0.0089661f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_34 VNB N_A_321_47#_c_389_n 0.0164654f $X=-0.19 $Y=-0.24 $X2=1.215 $Y2=1.455
cc_35 VPB N_A_83_21#_c_65_n 0.0199934f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_36 VPB N_A_83_21#_c_66_n 0.0192904f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_37 VPB N_A_83_21#_c_60_n 0.00205805f $X=-0.19 $Y=1.305 $X2=1.235 $Y2=1.16
cc_38 VPB N_A_83_21#_c_68_n 0.00702546f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.58
cc_39 VPB N_A_83_21#_c_69_n 0.00248213f $X=-0.19 $Y=1.305 $X2=2.517 $Y2=1.705
cc_40 VPB N_A_83_21#_c_64_n 0.034369f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_41 VPB N_B1_c_145_n 0.0182539f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=0.235
cc_42 VPB N_B1_c_144_n 0.0143797f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_43 VPB N_B2_c_173_n 0.0271036f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=0.235
cc_44 VPB N_A2_c_206_n 0.028919f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=0.235
cc_45 VPB A2 0.00296899f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=0.995
cc_46 VPB N_A1_c_242_n 0.0320558f $X=-0.19 $Y=1.305 $X2=2.065 $Y2=0.235
cc_47 VPB N_A1_c_244_n 0.00713408f $X=-0.19 $Y=1.305 $X2=0.95 $Y2=0.995
cc_48 VPB N_VPWR_c_266_n 0.0106521f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_49 VPB N_VPWR_c_267_n 0.0497821f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_50 VPB N_VPWR_c_268_n 0.0208523f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_51 VPB N_VPWR_c_269_n 0.0163048f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_52 VPB N_VPWR_c_270_n 0.0346482f $X=-0.19 $Y=1.305 $X2=1.215 $Y2=1.455
cc_53 VPB N_VPWR_c_271_n 0.0464935f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.805
cc_54 VPB N_VPWR_c_272_n 0.0197075f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.77
cc_55 VPB N_VPWR_c_265_n 0.050548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_X_c_311_n 0.00158459f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_57 N_A_83_21#_c_60_n N_B1_c_145_n 0.00113072f $X=1.235 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_58 N_A_83_21#_c_68_n N_B1_c_145_n 0.0247424f $X=2.34 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_59 N_A_83_21#_c_73_p N_B1_c_145_n 0.00293076f $X=2.61 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_83_21#_c_60_n N_B1_c_142_n 0.0023965f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_83_21#_c_75_p N_B1_c_142_n 0.0100879f $X=2.075 $Y=0.77 $X2=0 $Y2=0
cc_62 N_A_83_21#_c_63_n N_B1_c_142_n 0.00628506f $X=1.95 $Y=0.77 $X2=0 $Y2=0
cc_63 N_A_83_21#_c_60_n B1 0.0156875f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_83_21#_c_68_n B1 0.026296f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_83_21#_c_63_n B1 0.0256743f $X=1.95 $Y=0.77 $X2=0 $Y2=0
cc_66 N_A_83_21#_c_64_n B1 0.00131724f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_67 N_A_83_21#_c_60_n N_B1_c_144_n 0.00337986f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_83_21#_c_68_n N_B1_c_144_n 0.00720194f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_69 N_A_83_21#_c_63_n N_B1_c_144_n 0.00826414f $X=1.95 $Y=0.77 $X2=0 $Y2=0
cc_70 N_A_83_21#_c_64_n N_B1_c_144_n 0.0216846f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_71 N_A_83_21#_c_68_n N_B2_c_173_n 0.00718525f $X=2.34 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_83_21#_c_62_n N_B2_c_173_n 0.00170855f $X=2.2 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_83_21#_c_69_n N_B2_c_173_n 0.00848516f $X=2.517 $Y=1.705 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_83_21#_c_73_p N_B2_c_173_n 0.0191259f $X=2.61 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_83_21#_c_62_n N_B2_c_174_n 0.00424953f $X=2.2 $Y=0.73 $X2=0 $Y2=0
cc_76 N_A_83_21#_c_68_n B2 0.0168386f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_83_21#_c_62_n B2 0.0187599f $X=2.2 $Y=0.73 $X2=0 $Y2=0
cc_78 N_A_83_21#_c_69_n B2 0.0218106f $X=2.517 $Y=1.705 $X2=0 $Y2=0
cc_79 N_A_83_21#_c_69_n N_A2_c_206_n 0.00106163f $X=2.517 $Y=1.705 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_83_21#_c_73_p N_A2_c_206_n 0.00405045f $X=2.61 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_83_21#_c_62_n N_A2_c_207_n 2.53164e-19 $X=2.2 $Y=0.73 $X2=0 $Y2=0
cc_82 N_A_83_21#_c_69_n A2 0.0106557f $X=2.517 $Y=1.705 $X2=0 $Y2=0
cc_83 N_A_83_21#_c_68_n N_VPWR_M1010_s 0.00888207f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_83_21#_c_98_p N_VPWR_M1010_s 0.00431066f $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_83_21#_c_65_n N_VPWR_c_267_n 0.00981714f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_83_21#_c_65_n N_VPWR_c_268_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_83_21#_c_66_n N_VPWR_c_268_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_83_21#_c_73_p N_VPWR_c_271_n 0.0225392f $X=2.61 $Y=2.3 $X2=0 $Y2=0
cc_89 N_A_83_21#_c_66_n N_VPWR_c_272_n 0.00513552f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_83_21#_c_68_n N_VPWR_c_272_n 0.0400793f $X=2.34 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_83_21#_c_98_p N_VPWR_c_272_n 0.0201061f $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_92 N_A_83_21#_c_73_p N_VPWR_c_272_n 0.021613f $X=2.61 $Y=2.3 $X2=0 $Y2=0
cc_93 N_A_83_21#_c_64_n N_VPWR_c_272_n 9.14481e-19 $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_94 N_A_83_21#_M1007_d N_VPWR_c_265_n 0.0113163f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_95 N_A_83_21#_c_65_n N_VPWR_c_265_n 0.0134391f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_83_21#_c_66_n N_VPWR_c_265_n 0.0136916f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_83_21#_c_73_p N_VPWR_c_265_n 0.0129551f $X=2.61 $Y=2.3 $X2=0 $Y2=0
cc_98 N_A_83_21#_c_58_n N_X_c_311_n 0.00351484f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_83_21#_c_65_n N_X_c_311_n 0.00135141f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_83_21#_c_59_n N_X_c_311_n 0.0016326f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_83_21#_c_66_n N_X_c_311_n 6.37934e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_83_21#_c_60_n N_X_c_311_n 0.0345116f $X=1.235 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_83_21#_c_61_n N_X_c_311_n 6.5033e-19 $X=1.355 $Y=0.805 $X2=0 $Y2=0
cc_104 N_A_83_21#_c_98_p N_X_c_311_n 0.00952835f $X=1.355 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A_83_21#_c_64_n N_X_c_311_n 0.0406344f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_106 N_A_83_21#_c_68_n A_411_297# 0.00463738f $X=2.34 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_107 N_A_83_21#_c_61_n N_VGND_M1009_s 0.00477615f $X=1.355 $Y=0.805 $X2=0
+ $Y2=0
cc_108 N_A_83_21#_c_58_n N_VGND_c_332_n 0.00882727f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_83_21#_c_58_n N_VGND_c_333_n 0.00585385f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_83_21#_c_59_n N_VGND_c_333_n 0.00585385f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_83_21#_c_61_n N_VGND_c_333_n 7.52196e-19 $X=1.355 $Y=0.805 $X2=0
+ $Y2=0
cc_112 N_A_83_21#_c_59_n N_VGND_c_334_n 0.00714755f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_83_21#_c_61_n N_VGND_c_334_n 0.0153534f $X=1.355 $Y=0.805 $X2=0 $Y2=0
cc_114 N_A_83_21#_c_64_n N_VGND_c_334_n 7.54704e-19 $X=0.985 $Y=1.202 $X2=0
+ $Y2=0
cc_115 N_A_83_21#_c_61_n N_VGND_c_336_n 8.30317e-19 $X=1.355 $Y=0.805 $X2=0
+ $Y2=0
cc_116 N_A_83_21#_c_63_n N_VGND_c_336_n 0.00326925f $X=1.95 $Y=0.77 $X2=0 $Y2=0
cc_117 N_A_83_21#_M1011_d N_VGND_c_339_n 0.00219239f $X=2.065 $Y=0.235 $X2=0
+ $Y2=0
cc_118 N_A_83_21#_c_58_n N_VGND_c_339_n 0.0117174f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_83_21#_c_59_n N_VGND_c_339_n 0.0121683f $X=0.95 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_83_21#_c_61_n N_VGND_c_339_n 0.00370573f $X=1.355 $Y=0.805 $X2=0
+ $Y2=0
cc_121 N_A_83_21#_c_63_n N_VGND_c_339_n 0.00649634f $X=1.95 $Y=0.77 $X2=0 $Y2=0
cc_122 N_A_83_21#_c_63_n N_A_321_47#_M1011_s 0.00426421f $X=1.95 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_123 N_A_83_21#_M1011_d N_A_321_47#_c_387_n 0.00323205f $X=2.065 $Y=0.235
+ $X2=0 $Y2=0
cc_124 N_A_83_21#_c_75_p N_A_321_47#_c_387_n 0.0207168f $X=2.075 $Y=0.77 $X2=0
+ $Y2=0
cc_125 N_A_83_21#_c_63_n N_A_321_47#_c_387_n 0.0170223f $X=1.95 $Y=0.77 $X2=0
+ $Y2=0
cc_126 N_A_83_21#_c_62_n N_A_321_47#_c_394_n 0.015009f $X=2.2 $Y=0.73 $X2=0
+ $Y2=0
cc_127 N_A_83_21#_c_69_n N_A_321_47#_c_394_n 0.00257981f $X=2.517 $Y=1.705 $X2=0
+ $Y2=0
cc_128 N_B1_c_145_n N_B2_c_173_n 0.0668085f $X=1.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_129 N_B1_c_144_n N_B2_c_173_n 0.0284609f $X=1.965 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_130 N_B1_c_142_n N_B2_c_174_n 0.0270391f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_131 B1 B2 0.0135933f $X=1.62 $Y=1.105 $X2=0 $Y2=0
cc_132 N_B1_c_144_n B2 0.00176813f $X=1.965 $Y=1.202 $X2=0 $Y2=0
cc_133 N_B1_c_145_n N_VPWR_c_271_n 0.0062441f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B1_c_145_n N_VPWR_c_272_n 0.0164221f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B1_c_145_n N_VPWR_c_265_n 0.0103479f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_136 N_B1_c_142_n N_VGND_c_334_n 0.00228359f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_142_n N_VGND_c_336_n 0.00366111f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_142_n N_VGND_c_339_n 0.0065944f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_142_n N_A_321_47#_c_387_n 0.00819977f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B2_c_173_n N_A2_c_206_n 0.0389782f $X=2.375 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_141 B2 N_A2_c_206_n 6.8902e-19 $X=2.355 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_142 N_B2_c_174_n N_A2_c_207_n 0.0173647f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B2_c_173_n N_A2_c_208_n 6.19643e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_144 B2 N_A2_c_208_n 0.0173093f $X=2.355 $Y=1.19 $X2=0 $Y2=0
cc_145 N_B2_c_173_n A2 0.00270205f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B2_c_173_n N_VPWR_c_271_n 0.00514216f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_147 N_B2_c_173_n N_VPWR_c_272_n 0.00272235f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_148 N_B2_c_173_n N_VPWR_c_265_n 0.00843094f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B2_c_174_n N_VGND_c_336_n 0.00366111f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B2_c_174_n N_VGND_c_339_n 0.00583513f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B2_c_173_n N_A_321_47#_c_387_n 0.00164267f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B2_c_174_n N_A_321_47#_c_387_n 0.0127348f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_153 B2 N_A_321_47#_c_387_n 0.00487113f $X=2.355 $Y=1.19 $X2=0 $Y2=0
cc_154 N_B2_c_174_n N_A_321_47#_c_394_n 0.007118f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_155 B2 N_A_321_47#_c_394_n 0.00245662f $X=2.355 $Y=1.19 $X2=0 $Y2=0
cc_156 N_A2_c_206_n N_A1_c_242_n 0.0943384f $X=3.045 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_157 N_A2_c_208_n N_A1_c_242_n 0.00107607f $X=2.96 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_158 A2 N_A1_c_242_n 3.27034e-19 $X=2.93 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_159 N_A2_c_207_n N_A1_c_243_n 0.025512f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_206_n N_A1_c_244_n 0.00136551f $X=3.045 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A2_c_208_n N_A1_c_244_n 0.034149f $X=2.96 $Y=1.16 $X2=0 $Y2=0
cc_162 N_A2_c_206_n N_VPWR_c_271_n 0.00443901f $X=3.045 $Y=1.41 $X2=0 $Y2=0
cc_163 A2 N_VPWR_c_271_n 0.0110916f $X=2.93 $Y=1.785 $X2=0 $Y2=0
cc_164 N_A2_c_206_n N_VPWR_c_265_n 0.00645065f $X=3.045 $Y=1.41 $X2=0 $Y2=0
cc_165 A2 N_VPWR_c_265_n 0.00915489f $X=2.93 $Y=1.785 $X2=0 $Y2=0
cc_166 N_A2_c_207_n N_VGND_c_335_n 0.00271724f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A2_c_207_n N_VGND_c_336_n 0.00433717f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A2_c_207_n N_VGND_c_339_n 0.00646074f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A2_c_207_n N_A_321_47#_c_402_n 0.00224788f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A2_c_206_n N_A_321_47#_c_394_n 0.00311655f $X=3.045 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A2_c_207_n N_A_321_47#_c_394_n 0.00336464f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_208_n N_A_321_47#_c_394_n 0.00917875f $X=2.96 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A2_c_206_n N_A_321_47#_c_388_n 0.00156902f $X=3.045 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_207_n N_A_321_47#_c_388_n 0.0130731f $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_c_208_n N_A_321_47#_c_388_n 0.0133344f $X=2.96 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A2_c_207_n N_A_321_47#_c_389_n 5.35028e-19 $X=3.07 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A1_c_244_n N_VPWR_M1003_d 0.00657895f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A1_c_242_n N_VPWR_c_270_n 0.00666012f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A1_c_244_n N_VPWR_c_270_n 0.00866122f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A1_c_242_n N_VPWR_c_271_n 0.00702461f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A1_c_242_n N_VPWR_c_265_n 0.0134147f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_c_243_n N_VGND_c_335_n 0.00416635f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_243_n N_VGND_c_338_n 0.00421028f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A1_c_243_n N_VGND_c_339_n 0.00686073f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A1_c_242_n N_A_321_47#_c_388_n 0.00666272f $X=3.455 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A1_c_243_n N_A_321_47#_c_388_n 0.00955327f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_244_n N_A_321_47#_c_388_n 0.0201063f $X=3.54 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A1_c_243_n N_A_321_47#_c_389_n 0.00621202f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_189 N_VPWR_c_265_n N_X_M1001_d 0.00370124f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_267_n N_X_c_311_n 0.0624127f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_191 N_VPWR_c_268_n N_X_c_311_n 0.0149311f $X=1.095 $Y=2.72 $X2=0 $Y2=0
cc_192 N_VPWR_c_265_n N_X_c_311_n 0.00955092f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_193 N_VPWR_c_265_n A_411_297# 0.00983149f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_194 N_VPWR_c_265_n A_627_297# 0.00848405f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_195 N_VPWR_c_267_n N_VGND_c_332_n 0.00652169f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_196 N_X_c_311_n N_VGND_c_333_n 0.00915701f $X=0.74 $Y=0.595 $X2=0 $Y2=0
cc_197 N_X_M1006_d N_VGND_c_339_n 0.00475625f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_198 N_X_c_311_n N_VGND_c_339_n 0.00899302f $X=0.74 $Y=0.595 $X2=0 $Y2=0
cc_199 N_VGND_c_339_n N_A_321_47#_M1011_s 0.00253093f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_200 N_VGND_c_339_n N_A_321_47#_M1000_d 0.00445357f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_201 N_VGND_c_339_n N_A_321_47#_M1004_d 0.00210425f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_334_n N_A_321_47#_c_387_n 0.0109506f $X=1.21 $Y=0.38 $X2=0 $Y2=0
cc_203 N_VGND_c_336_n N_A_321_47#_c_387_n 0.0464573f $X=3.195 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_339_n N_A_321_47#_c_387_n 0.0358315f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_205 N_VGND_c_336_n N_A_321_47#_c_402_n 0.0187671f $X=3.195 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_339_n N_A_321_47#_c_402_n 0.0127684f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_M1008_d N_A_321_47#_c_388_n 0.00772066f $X=3.145 $Y=0.235 $X2=0
+ $Y2=0
cc_208 N_VGND_c_335_n N_A_321_47#_c_388_n 0.0125799f $X=3.28 $Y=0.36 $X2=0 $Y2=0
cc_209 N_VGND_c_336_n N_A_321_47#_c_388_n 0.00314714f $X=3.195 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_338_n N_A_321_47#_c_388_n 0.00237788f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_339_n N_A_321_47#_c_388_n 0.0115771f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_212 N_VGND_c_335_n N_A_321_47#_c_389_n 0.0166203f $X=3.28 $Y=0.36 $X2=0 $Y2=0
cc_213 N_VGND_c_338_n N_A_321_47#_c_389_n 0.0182739f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_214 N_VGND_c_339_n N_A_321_47#_c_389_n 0.0124095f $X=3.91 $Y=0 $X2=0 $Y2=0
