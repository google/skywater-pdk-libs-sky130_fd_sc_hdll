* File: sky130_fd_sc_hdll__nor4b_4.pxi.spice
* Created: Wed Sep  2 08:41:48 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%A N_A_c_132_n N_A_M1008_g N_A_c_138_n
+ N_A_M1002_g N_A_c_133_n N_A_M1010_g N_A_c_139_n N_A_M1016_g N_A_c_134_n
+ N_A_M1025_g N_A_c_140_n N_A_M1022_g N_A_c_141_n N_A_M1030_g N_A_c_135_n
+ N_A_M1032_g A N_A_c_136_n N_A_c_137_n A PM_SKY130_FD_SC_HDLL__NOR4B_4%A
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%B N_B_c_207_n N_B_M1011_g N_B_c_213_n
+ N_B_M1000_g N_B_c_208_n N_B_M1019_g N_B_c_214_n N_B_M1006_g N_B_c_209_n
+ N_B_M1028_g N_B_c_215_n N_B_M1009_g N_B_c_216_n N_B_M1017_g N_B_c_210_n
+ N_B_M1029_g B N_B_c_211_n N_B_c_212_n B PM_SKY130_FD_SC_HDLL__NOR4B_4%B
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%C N_C_c_284_n N_C_M1005_g N_C_c_290_n
+ N_C_M1004_g N_C_c_285_n N_C_M1015_g N_C_c_291_n N_C_M1007_g N_C_c_286_n
+ N_C_M1024_g N_C_c_292_n N_C_M1020_g N_C_c_293_n N_C_M1031_g N_C_c_287_n
+ N_C_M1033_g C N_C_c_288_n N_C_c_289_n C PM_SKY130_FD_SC_HDLL__NOR4B_4%C
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%A_1311_21# N_A_1311_21#_M1027_s
+ N_A_1311_21#_M1013_s N_A_1311_21#_c_362_n N_A_1311_21#_M1001_g
+ N_A_1311_21#_c_371_n N_A_1311_21#_M1012_g N_A_1311_21#_c_363_n
+ N_A_1311_21#_M1003_g N_A_1311_21#_c_372_n N_A_1311_21#_M1018_g
+ N_A_1311_21#_c_364_n N_A_1311_21#_M1014_g N_A_1311_21#_c_373_n
+ N_A_1311_21#_M1023_g N_A_1311_21#_c_365_n N_A_1311_21#_M1021_g
+ N_A_1311_21#_c_374_n N_A_1311_21#_M1026_g N_A_1311_21#_c_419_p
+ N_A_1311_21#_c_366_n N_A_1311_21#_c_375_n N_A_1311_21#_c_376_n
+ N_A_1311_21#_c_377_n N_A_1311_21#_c_367_n N_A_1311_21#_c_368_n
+ N_A_1311_21#_c_378_n N_A_1311_21#_c_392_p N_A_1311_21#_c_369_n
+ N_A_1311_21#_c_370_n PM_SKY130_FD_SC_HDLL__NOR4B_4%A_1311_21#
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%D_N N_D_N_c_480_n N_D_N_M1027_g N_D_N_c_481_n
+ N_D_N_M1013_g D_N D_N PM_SKY130_FD_SC_HDLL__NOR4B_4%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%A_27_297# N_A_27_297#_M1002_d
+ N_A_27_297#_M1016_d N_A_27_297#_M1030_d N_A_27_297#_M1006_d
+ N_A_27_297#_M1017_d N_A_27_297#_c_507_n N_A_27_297#_c_508_n
+ N_A_27_297#_c_509_n N_A_27_297#_c_538_p N_A_27_297#_c_510_n
+ N_A_27_297#_c_511_n N_A_27_297#_c_540_p N_A_27_297#_c_530_n
+ N_A_27_297#_c_560_p N_A_27_297#_c_512_n N_A_27_297#_c_564_p
+ N_A_27_297#_c_513_n N_A_27_297#_c_543_p
+ PM_SKY130_FD_SC_HDLL__NOR4B_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%VPWR N_VPWR_M1002_s N_VPWR_M1022_s
+ N_VPWR_M1013_d N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n
+ N_VPWR_c_578_n VPWR N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n
+ N_VPWR_c_573_n PM_SKY130_FD_SC_HDLL__NOR4B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%A_493_297# N_A_493_297#_M1000_s
+ N_A_493_297#_M1009_s N_A_493_297#_M1004_d N_A_493_297#_M1020_d
+ N_A_493_297#_c_677_n N_A_493_297#_c_678_n N_A_493_297#_c_679_n
+ N_A_493_297#_c_680_n N_A_493_297#_c_681_n N_A_493_297#_c_682_n
+ N_A_493_297#_c_683_n PM_SKY130_FD_SC_HDLL__NOR4B_4%A_493_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%A_883_297# N_A_883_297#_M1004_s
+ N_A_883_297#_M1007_s N_A_883_297#_M1031_s N_A_883_297#_M1018_s
+ N_A_883_297#_M1026_s N_A_883_297#_c_757_n N_A_883_297#_c_740_n
+ N_A_883_297#_c_737_n N_A_883_297#_c_787_n N_A_883_297#_c_742_n
+ N_A_883_297#_c_738_n N_A_883_297#_c_747_n N_A_883_297#_c_749_n
+ N_A_883_297#_c_739_n N_A_883_297#_c_753_n N_A_883_297#_c_774_n
+ N_A_883_297#_c_776_n N_A_883_297#_c_778_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_4%A_883_297#
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%Y N_Y_M1008_d N_Y_M1025_d N_Y_M1011_s
+ N_Y_M1028_s N_Y_M1005_s N_Y_M1024_s N_Y_M1001_s N_Y_M1014_s N_Y_M1012_d
+ N_Y_M1023_d N_Y_c_820_n N_Y_c_802_n N_Y_c_803_n N_Y_c_831_n N_Y_c_804_n
+ N_Y_c_835_n N_Y_c_805_n N_Y_c_848_n N_Y_c_806_n N_Y_c_861_n N_Y_c_807_n
+ N_Y_c_868_n N_Y_c_808_n N_Y_c_872_n N_Y_c_809_n N_Y_c_810_n N_Y_c_818_n
+ N_Y_c_903_n N_Y_c_811_n N_Y_c_812_n N_Y_c_813_n N_Y_c_814_n N_Y_c_815_n
+ N_Y_c_816_n N_Y_c_909_n N_Y_c_819_n Y PM_SKY130_FD_SC_HDLL__NOR4B_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR4B_4%VGND N_VGND_M1008_s N_VGND_M1010_s
+ N_VGND_M1032_s N_VGND_M1019_d N_VGND_M1029_d N_VGND_M1015_d N_VGND_M1033_d
+ N_VGND_M1003_d N_VGND_M1021_d N_VGND_M1027_d N_VGND_c_998_n N_VGND_c_999_n
+ N_VGND_c_1000_n N_VGND_c_1001_n N_VGND_c_1002_n N_VGND_c_1003_n
+ N_VGND_c_1004_n N_VGND_c_1005_n N_VGND_c_1006_n N_VGND_c_1007_n
+ N_VGND_c_1008_n N_VGND_c_1009_n N_VGND_c_1010_n N_VGND_c_1011_n
+ N_VGND_c_1012_n N_VGND_c_1013_n N_VGND_c_1014_n N_VGND_c_1015_n
+ N_VGND_c_1016_n N_VGND_c_1017_n N_VGND_c_1018_n N_VGND_c_1019_n
+ N_VGND_c_1020_n VGND N_VGND_c_1021_n N_VGND_c_1022_n N_VGND_c_1023_n
+ N_VGND_c_1024_n N_VGND_c_1025_n N_VGND_c_1026_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_4%VGND
cc_1 VNB N_A_c_132_n 0.0221045f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_133_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_c_134_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_A_c_135_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A_c_136_n 0.0100386f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_6 VNB N_A_c_137_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_7 VNB N_B_c_207_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_8 VNB N_B_c_208_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_9 VNB N_B_c_209_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_10 VNB N_B_c_210_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_11 VNB N_B_c_211_n 0.00882304f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_12 VNB N_B_c_212_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_13 VNB N_C_c_284_n 0.021971f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_C_c_285_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_15 VNB N_C_c_286_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_16 VNB N_C_c_287_n 0.0169154f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_17 VNB N_C_c_288_n 0.0098547f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_18 VNB N_C_c_289_n 0.0801646f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_19 VNB N_A_1311_21#_c_362_n 0.0164576f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_20 VNB N_A_1311_21#_c_363_n 0.015981f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_21 VNB N_A_1311_21#_c_364_n 0.0167056f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_22 VNB N_A_1311_21#_c_365_n 0.0196183f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.105
cc_23 VNB N_A_1311_21#_c_366_n 0.0025053f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.16
cc_24 VNB N_A_1311_21#_c_367_n 0.0104937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_1311_21#_c_368_n 0.00685504f $X=-0.19 $Y=-0.24 $X2=1.135 $Y2=1.19
cc_26 VNB N_A_1311_21#_c_369_n 0.0303949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_1311_21#_c_370_n 0.0722793f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_D_N_c_480_n 0.0253661f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_29 VNB N_D_N_c_481_n 0.0427565f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_30 VNB D_N 0.0208841f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_31 VNB N_VPWR_c_573_n 0.402575f $X=-0.19 $Y=-0.24 $X2=1.235 $Y2=1.18
cc_32 VNB N_Y_c_802_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_33 VNB N_Y_c_803_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.202
cc_34 VNB N_Y_c_804_n 0.00447396f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.18
cc_35 VNB N_Y_c_805_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=1.18
cc_36 VNB N_Y_c_806_n 0.00915678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_807_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_808_n 0.00470652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_809_n 0.00194903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_810_n 0.00469873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_811_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_Y_c_812_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_813_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_814_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_815_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_816_n 0.00243026f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_998_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_48 VNB N_VGND_c_999_n 0.00779204f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_49 VNB N_VGND_c_1000_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_50 VNB N_VGND_c_1001_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_51 VNB N_VGND_c_1002_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.18
cc_52 VNB N_VGND_c_1003_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_1004_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_1005_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1006_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_1007_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_1008_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_1009_n 0.0138021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1010_n 0.00745006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_1011_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_1012_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1013_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1014_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1015_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1016_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1017_n 0.0191731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1018_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1019_n 0.0200006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1020_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1021_n 0.0215605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1022_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1023_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1024_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1025_n 0.0208752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1026_n 0.456715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VPB N_A_c_138_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_77 VPB N_A_c_139_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_78 VPB N_A_c_140_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_79 VPB N_A_c_141_n 0.0161064f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_80 VPB N_A_c_137_n 0.048391f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_81 VPB N_B_c_213_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_82 VPB N_B_c_214_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_83 VPB N_B_c_215_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_84 VPB N_B_c_216_n 0.0203443f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_85 VPB N_B_c_212_n 0.0492916f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_86 VPB N_C_c_290_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_87 VPB N_C_c_291_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_88 VPB N_C_c_292_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_89 VPB N_C_c_293_n 0.0164209f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_90 VPB N_C_c_289_n 0.0492868f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_91 VPB N_A_1311_21#_c_371_n 0.0164077f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_92 VPB N_A_1311_21#_c_372_n 0.0155712f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_93 VPB N_A_1311_21#_c_373_n 0.0159298f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_94 VPB N_A_1311_21#_c_374_n 0.0191625f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_95 VPB N_A_1311_21#_c_375_n 0.00287727f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_96 VPB N_A_1311_21#_c_376_n 0.0145923f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.202
cc_97 VPB N_A_1311_21#_c_377_n 8.55739e-19 $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.18
cc_98 VPB N_A_1311_21#_c_378_n 0.00932478f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_1311_21#_c_369_n 0.0113164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_1311_21#_c_370_n 0.0473565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_D_N_c_481_n 0.0428394f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_102 VPB N_A_27_297#_c_507_n 0.0327625f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_103 VPB N_A_27_297#_c_508_n 0.0018222f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_104 VPB N_A_27_297#_c_509_n 0.01536f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_105 VPB N_A_27_297#_c_510_n 0.00201678f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_106 VPB N_A_27_297#_c_511_n 0.00416269f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_107 VPB N_A_27_297#_c_512_n 0.0014688f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_108 VPB N_A_27_297#_c_513_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_574_n 0.00495424f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.56
cc_110 VPB N_VPWR_c_575_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_111 VPB N_VPWR_c_576_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_112 VPB N_VPWR_c_577_n 0.0137762f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_113 VPB N_VPWR_c_578_n 0.0079748f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_114 VPB N_VPWR_c_579_n 0.173083f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_115 VPB N_VPWR_c_580_n 0.0234703f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_116 VPB N_VPWR_c_581_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_573_n 0.0713217f $X=-0.19 $Y=1.305 $X2=1.235 $Y2=1.18
cc_118 VPB N_A_493_297#_c_677_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=0.56
cc_119 VPB N_A_493_297#_c_678_n 0.0201481f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_120 VPB N_A_493_297#_c_679_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_121 VPB N_A_493_297#_c_680_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_122 VPB N_A_493_297#_c_681_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_123 VPB N_A_493_297#_c_682_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=1.202
cc_124 VPB N_A_493_297#_c_683_n 0.00175152f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.202
cc_125 VPB N_A_883_297#_c_737_n 0.0014688f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_126 VPB N_A_883_297#_c_738_n 0.00445834f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_127 VPB N_A_883_297#_c_739_n 0.00139236f $X=-0.19 $Y=1.305 $X2=1.73 $Y2=1.16
cc_128 VPB N_Y_c_809_n 0.0028187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Y_c_818_n 0.00195526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Y_c_819_n 0.00177663f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 N_A_c_135_n N_B_c_207_n 0.0243397f $X=1.93 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_132 N_A_c_141_n N_B_c_213_n 0.00971598f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_136_n N_B_c_211_n 0.0121231f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_137_n N_B_c_211_n 2.62535e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_135 N_A_c_136_n N_B_c_212_n 2.62535e-19 $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_137_n N_B_c_212_n 0.0243397f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_c_138_n N_A_27_297#_c_507_n 0.0113204f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_139_n N_A_27_297#_c_507_n 6.54703e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_138_n N_A_27_297#_c_508_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_139_n N_A_27_297#_c_508_n 0.0156273f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_136_n N_A_27_297#_c_508_n 0.0458726f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_142 N_A_c_137_n N_A_27_297#_c_508_n 0.00807006f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_143 N_A_c_138_n N_A_27_297#_c_509_n 0.001185f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_136_n N_A_27_297#_c_509_n 0.00236396f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_137_n N_A_27_297#_c_509_n 3.16729e-19 $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_146 N_A_c_140_n N_A_27_297#_c_510_n 0.0156273f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_141_n N_A_27_297#_c_510_n 0.0155666f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_136_n N_A_27_297#_c_510_n 0.0480109f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_c_137_n N_A_27_297#_c_510_n 0.00816971f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_150 N_A_c_136_n N_A_27_297#_c_513_n 0.0204509f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_c_137_n N_A_27_297#_c_513_n 0.00656533f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_152 N_A_c_138_n N_VPWR_c_574_n 0.00553644f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_139_n N_VPWR_c_574_n 0.00295479f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_139_n N_VPWR_c_575_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_140_n N_VPWR_c_575_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_140_n N_VPWR_c_576_n 0.00300743f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_141_n N_VPWR_c_576_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_141_n N_VPWR_c_579_n 0.00702461f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_138_n N_VPWR_c_580_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_138_n N_VPWR_c_573_n 0.0127552f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_139_n N_VPWR_c_573_n 0.0124092f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_140_n N_VPWR_c_573_n 0.0124092f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_141_n N_VPWR_c_573_n 0.0124344f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_132_n N_Y_c_820_n 0.00539651f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_133_n N_Y_c_820_n 0.00686626f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_134_n N_Y_c_820_n 5.45498e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_133_n N_Y_c_802_n 0.00901745f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_134_n N_Y_c_802_n 0.00901745f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_136_n N_Y_c_802_n 0.0398926f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_c_137_n N_Y_c_802_n 0.00345541f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_c_132_n N_Y_c_803_n 0.00302596f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_133_n N_Y_c_803_n 0.00116636f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_136_n N_Y_c_803_n 0.0307014f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_137_n N_Y_c_803_n 0.00358305f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_c_133_n N_Y_c_831_n 5.24597e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_134_n N_Y_c_831_n 0.00651696f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_135_n N_Y_c_804_n 0.0106151f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_136_n N_Y_c_804_n 0.0118017f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_c_135_n N_Y_c_835_n 5.32212e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_134_n N_Y_c_811_n 0.00119564f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_136_n N_Y_c_811_n 0.030835f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_c_137_n N_Y_c_811_n 0.00486271f $X=1.905 $Y=1.202 $X2=0 $Y2=0
cc_183 N_A_c_132_n N_VGND_c_999_n 0.00460404f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_c_132_n N_VGND_c_1000_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_133_n N_VGND_c_1000_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_133_n N_VGND_c_1001_n 0.00379224f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_134_n N_VGND_c_1001_n 0.00276126f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_134_n N_VGND_c_1002_n 0.00423334f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_c_135_n N_VGND_c_1002_n 0.00437852f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_c_135_n N_VGND_c_1003_n 0.00268723f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_132_n N_VGND_c_1026_n 0.0105827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_c_133_n N_VGND_c_1026_n 0.006093f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_134_n N_VGND_c_1026_n 0.00608558f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_135_n N_VGND_c_1026_n 0.00615622f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B_c_211_n N_C_c_288_n 0.0155079f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_196 N_B_c_212_n N_C_c_288_n 9.30294e-19 $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_197 N_B_c_211_n N_C_c_289_n 8.91304e-19 $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_c_213_n N_A_27_297#_c_511_n 2.98195e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_213_n N_A_27_297#_c_530_n 0.0143578f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_214_n N_A_27_297#_c_530_n 0.01161f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_215_n N_A_27_297#_c_512_n 0.01161f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_216_n N_A_27_297#_c_512_n 0.01161f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_213_n N_VPWR_c_579_n 0.00429453f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_214_n N_VPWR_c_579_n 0.00429453f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_c_215_n N_VPWR_c_579_n 0.00429453f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_216_n N_VPWR_c_579_n 0.00429453f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_213_n N_VPWR_c_573_n 0.00609021f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_214_n N_VPWR_c_573_n 0.00606499f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_215_n N_VPWR_c_573_n 0.00606499f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_216_n N_VPWR_c_573_n 0.00734734f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_214_n N_A_493_297#_c_677_n 0.0128188f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_c_215_n N_A_493_297#_c_677_n 0.0128795f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B_c_211_n N_A_493_297#_c_677_n 0.0486996f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B_c_212_n N_A_493_297#_c_677_n 0.00864922f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_215 N_B_c_216_n N_A_493_297#_c_678_n 0.0148794f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B_c_211_n N_A_493_297#_c_678_n 0.0348238f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_217 N_B_c_212_n N_A_493_297#_c_678_n 8.84531e-19 $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_218 N_B_c_213_n N_A_493_297#_c_680_n 2.98195e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_211_n N_A_493_297#_c_680_n 0.0204252f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B_c_212_n N_A_493_297#_c_680_n 0.00655199f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_221 N_B_c_211_n N_A_493_297#_c_681_n 0.0204252f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_222 N_B_c_212_n N_A_493_297#_c_681_n 0.00634604f $X=3.785 $Y=1.202 $X2=0
+ $Y2=0
cc_223 N_B_c_207_n N_Y_c_804_n 0.00865686f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_211_n N_Y_c_804_n 0.00826974f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_225 N_B_c_207_n N_Y_c_835_n 0.00644736f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_208_n N_Y_c_835_n 0.00686626f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_227 N_B_c_209_n N_Y_c_835_n 5.45498e-19 $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B_c_208_n N_Y_c_805_n 0.00901745f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_209_n N_Y_c_805_n 0.00901745f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_211_n N_Y_c_805_n 0.0398926f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_231 N_B_c_212_n N_Y_c_805_n 0.00345541f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_232 N_B_c_208_n N_Y_c_848_n 5.24597e-19 $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_209_n N_Y_c_848_n 0.00651696f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_210_n N_Y_c_806_n 0.01289f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B_c_211_n N_Y_c_806_n 0.0321692f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_236 N_B_c_207_n N_Y_c_812_n 0.00116636f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_208_n N_Y_c_812_n 0.00116636f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_211_n N_Y_c_812_n 0.0307014f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_239 N_B_c_212_n N_Y_c_812_n 0.00358305f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_240 N_B_c_209_n N_Y_c_813_n 0.00119564f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_211_n N_Y_c_813_n 0.030835f $X=3.61 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B_c_212_n N_Y_c_813_n 0.00486271f $X=3.785 $Y=1.202 $X2=0 $Y2=0
cc_243 N_B_c_207_n N_VGND_c_1003_n 0.00268723f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B_c_208_n N_VGND_c_1004_n 0.00379224f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_245 N_B_c_209_n N_VGND_c_1004_n 0.00276126f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B_c_207_n N_VGND_c_1011_n 0.00423334f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B_c_208_n N_VGND_c_1011_n 0.00423334f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B_c_209_n N_VGND_c_1024_n 0.00423334f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B_c_210_n N_VGND_c_1024_n 0.00437852f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B_c_210_n N_VGND_c_1025_n 0.00481673f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B_c_207_n N_VGND_c_1026_n 0.00587047f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B_c_208_n N_VGND_c_1026_n 0.006093f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B_c_209_n N_VGND_c_1026_n 0.00608558f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B_c_210_n N_VGND_c_1026_n 0.00745263f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_255 N_C_c_287_n N_A_1311_21#_c_362_n 0.0237457f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_256 N_C_c_293_n N_A_1311_21#_c_371_n 0.00937092f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_257 N_C_c_288_n N_A_1311_21#_c_370_n 0.00101333f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_258 N_C_c_289_n N_A_1311_21#_c_370_n 0.0237457f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_259 N_C_c_290_n N_VPWR_c_579_n 0.00429453f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_260 N_C_c_291_n N_VPWR_c_579_n 0.00429453f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_261 N_C_c_292_n N_VPWR_c_579_n 0.00429453f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_262 N_C_c_293_n N_VPWR_c_579_n 0.00429453f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_263 N_C_c_290_n N_VPWR_c_573_n 0.00734734f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_264 N_C_c_291_n N_VPWR_c_573_n 0.00606499f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_265 N_C_c_292_n N_VPWR_c_573_n 0.00606499f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_266 N_C_c_293_n N_VPWR_c_573_n 0.00609021f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_267 N_C_c_290_n N_A_493_297#_c_678_n 0.0148794f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_268 N_C_c_288_n N_A_493_297#_c_678_n 0.036737f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_269 N_C_c_289_n N_A_493_297#_c_678_n 8.84531e-19 $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_270 N_C_c_291_n N_A_493_297#_c_679_n 0.0128795f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_271 N_C_c_292_n N_A_493_297#_c_679_n 0.0128188f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_272 N_C_c_288_n N_A_493_297#_c_679_n 0.0486996f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_273 N_C_c_289_n N_A_493_297#_c_679_n 0.00864922f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_274 N_C_c_288_n N_A_493_297#_c_682_n 0.0204252f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_275 N_C_c_289_n N_A_493_297#_c_682_n 0.00655199f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_276 N_C_c_293_n N_A_493_297#_c_683_n 2.98817e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_277 N_C_c_288_n N_A_493_297#_c_683_n 0.0204252f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_278 N_C_c_289_n N_A_493_297#_c_683_n 0.00634604f $X=6.185 $Y=1.202 $X2=0
+ $Y2=0
cc_279 N_C_c_290_n N_A_883_297#_c_740_n 0.01161f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_280 N_C_c_291_n N_A_883_297#_c_740_n 0.01161f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_281 N_C_c_292_n N_A_883_297#_c_742_n 0.01161f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_282 N_C_c_293_n N_A_883_297#_c_742_n 0.0143578f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_283 N_C_c_293_n N_A_883_297#_c_738_n 2.65342e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_284 N_C_c_284_n N_Y_c_806_n 0.0109318f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_285 N_C_c_288_n N_Y_c_806_n 0.0305587f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_286 N_C_c_284_n N_Y_c_861_n 0.0110728f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_287 N_C_c_285_n N_Y_c_861_n 0.00686626f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_288 N_C_c_286_n N_Y_c_861_n 5.45498e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_289 N_C_c_285_n N_Y_c_807_n 0.00901745f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_290 N_C_c_286_n N_Y_c_807_n 0.00901745f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_291 N_C_c_288_n N_Y_c_807_n 0.0398926f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_292 N_C_c_289_n N_Y_c_807_n 0.00345541f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_293 N_C_c_285_n N_Y_c_868_n 5.24597e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C_c_286_n N_Y_c_868_n 0.00651696f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_c_287_n N_Y_c_808_n 0.0106151f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_296 N_C_c_288_n N_Y_c_808_n 0.0118017f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_297 N_C_c_287_n N_Y_c_872_n 5.32212e-19 $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_c_288_n N_Y_c_809_n 0.00731834f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_299 N_C_c_289_n N_Y_c_809_n 8.00432e-19 $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_300 N_C_c_284_n N_Y_c_814_n 0.00116636f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_285_n N_Y_c_814_n 0.00116636f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_302 N_C_c_288_n N_Y_c_814_n 0.0307014f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_c_289_n N_Y_c_814_n 0.00358305f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_304 N_C_c_286_n N_Y_c_815_n 0.00119564f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_305 N_C_c_288_n N_Y_c_815_n 0.030835f $X=6.01 $Y=1.16 $X2=0 $Y2=0
cc_306 N_C_c_289_n N_Y_c_815_n 0.00486271f $X=6.185 $Y=1.202 $X2=0 $Y2=0
cc_307 N_C_c_285_n N_VGND_c_1005_n 0.00379224f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_308 N_C_c_286_n N_VGND_c_1005_n 0.00276126f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_309 N_C_c_287_n N_VGND_c_1006_n 0.00268723f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_310 N_C_c_284_n N_VGND_c_1013_n 0.00423334f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_311 N_C_c_285_n N_VGND_c_1013_n 0.00423334f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_312 N_C_c_286_n N_VGND_c_1015_n 0.00423334f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_313 N_C_c_287_n N_VGND_c_1015_n 0.00437852f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_314 N_C_c_284_n N_VGND_c_1025_n 0.00481673f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_315 N_C_c_284_n N_VGND_c_1026_n 0.00716687f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_316 N_C_c_285_n N_VGND_c_1026_n 0.006093f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_317 N_C_c_286_n N_VGND_c_1026_n 0.00608558f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_318 N_C_c_287_n N_VGND_c_1026_n 0.00615622f $X=6.21 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_1311_21#_c_366_n N_D_N_c_480_n 0.00213537f $X=8.355 $Y=1.075
+ $X2=-0.19 $Y2=-0.24
cc_320 N_A_1311_21#_c_367_n N_D_N_c_480_n 0.00307527f $X=8.797 $Y=0.735
+ $X2=-0.19 $Y2=-0.24
cc_321 N_A_1311_21#_c_368_n N_D_N_c_480_n 0.00625705f $X=8.82 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_322 N_A_1311_21#_c_366_n N_D_N_c_481_n 4.5229e-19 $X=8.355 $Y=1.075 $X2=0
+ $Y2=0
cc_323 N_A_1311_21#_c_375_n N_D_N_c_481_n 0.0033817f $X=8.355 $Y=1.455 $X2=0
+ $Y2=0
cc_324 N_A_1311_21#_c_376_n N_D_N_c_481_n 0.00340445f $X=8.65 $Y=1.54 $X2=0
+ $Y2=0
cc_325 N_A_1311_21#_c_378_n N_D_N_c_481_n 0.0105084f $X=8.82 $Y=1.63 $X2=0 $Y2=0
cc_326 N_A_1311_21#_c_392_p N_D_N_c_481_n 2.01987e-19 $X=8.355 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_1311_21#_c_369_n N_D_N_c_481_n 0.00963129f $X=8.355 $Y=1.16 $X2=0
+ $Y2=0
cc_328 N_A_1311_21#_c_376_n D_N 0.0109334f $X=8.65 $Y=1.54 $X2=0 $Y2=0
cc_329 N_A_1311_21#_c_367_n D_N 0.00971996f $X=8.797 $Y=0.735 $X2=0 $Y2=0
cc_330 N_A_1311_21#_c_392_p D_N 0.00950329f $X=8.355 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_1311_21#_c_369_n D_N 0.00210458f $X=8.355 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_1311_21#_c_376_n N_VPWR_c_578_n 0.0112654f $X=8.65 $Y=1.54 $X2=0
+ $Y2=0
cc_333 N_A_1311_21#_c_378_n N_VPWR_c_578_n 0.0520518f $X=8.82 $Y=1.63 $X2=0
+ $Y2=0
cc_334 N_A_1311_21#_c_371_n N_VPWR_c_579_n 0.00429453f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_335 N_A_1311_21#_c_372_n N_VPWR_c_579_n 0.00429453f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_336 N_A_1311_21#_c_373_n N_VPWR_c_579_n 0.00429453f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_337 N_A_1311_21#_c_374_n N_VPWR_c_579_n 0.00429453f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_338 N_A_1311_21#_c_378_n N_VPWR_c_579_n 0.021418f $X=8.82 $Y=1.63 $X2=0 $Y2=0
cc_339 N_A_1311_21#_M1013_s N_VPWR_c_573_n 0.00217517f $X=8.695 $Y=1.485 $X2=0
+ $Y2=0
cc_340 N_A_1311_21#_c_371_n N_VPWR_c_573_n 0.00609021f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A_1311_21#_c_372_n N_VPWR_c_573_n 0.00606499f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_342 N_A_1311_21#_c_373_n N_VPWR_c_573_n 0.00606499f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A_1311_21#_c_374_n N_VPWR_c_573_n 0.00734734f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_344 N_A_1311_21#_c_378_n N_VPWR_c_573_n 0.0126651f $X=8.82 $Y=1.63 $X2=0
+ $Y2=0
cc_345 N_A_1311_21#_c_377_n N_A_883_297#_M1026_s 0.00426111f $X=8.44 $Y=1.54
+ $X2=0 $Y2=0
cc_346 N_A_1311_21#_c_371_n N_A_883_297#_c_738_n 2.65342e-19 $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_347 N_A_1311_21#_c_371_n N_A_883_297#_c_747_n 0.0143578f $X=6.655 $Y=1.41
+ $X2=0 $Y2=0
cc_348 N_A_1311_21#_c_372_n N_A_883_297#_c_747_n 0.0116061f $X=7.125 $Y=1.41
+ $X2=0 $Y2=0
cc_349 N_A_1311_21#_c_370_n N_A_883_297#_c_749_n 3.19626e-19 $X=8.165 $Y=1.16
+ $X2=0 $Y2=0
cc_350 N_A_1311_21#_c_373_n N_A_883_297#_c_739_n 0.01161f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_351 N_A_1311_21#_c_374_n N_A_883_297#_c_739_n 0.0143578f $X=8.065 $Y=1.41
+ $X2=0 $Y2=0
cc_352 N_A_1311_21#_c_378_n N_A_883_297#_c_739_n 0.0120455f $X=8.82 $Y=1.63
+ $X2=0 $Y2=0
cc_353 N_A_1311_21#_c_419_p N_A_883_297#_c_753_n 0.0024768f $X=8.27 $Y=1.18
+ $X2=0 $Y2=0
cc_354 N_A_1311_21#_c_377_n N_A_883_297#_c_753_n 0.0139284f $X=8.44 $Y=1.54
+ $X2=0 $Y2=0
cc_355 N_A_1311_21#_c_378_n N_A_883_297#_c_753_n 0.0327603f $X=8.82 $Y=1.63
+ $X2=0 $Y2=0
cc_356 N_A_1311_21#_c_369_n N_A_883_297#_c_753_n 0.00230337f $X=8.355 $Y=1.16
+ $X2=0 $Y2=0
cc_357 N_A_1311_21#_c_362_n N_Y_c_808_n 0.0122977f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A_1311_21#_c_362_n N_Y_c_872_n 0.00644736f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A_1311_21#_c_363_n N_Y_c_872_n 0.00686626f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A_1311_21#_c_364_n N_Y_c_872_n 5.45498e-19 $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A_1311_21#_c_362_n N_Y_c_809_n 0.00263038f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A_1311_21#_c_371_n N_Y_c_809_n 0.00135799f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_1311_21#_c_363_n N_Y_c_809_n 0.00272547f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_1311_21#_c_372_n N_Y_c_809_n 0.00134741f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_1311_21#_c_364_n N_Y_c_809_n 0.00210171f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A_1311_21#_c_373_n N_Y_c_809_n 0.00102052f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_1311_21#_c_419_p N_Y_c_809_n 0.0170792f $X=8.27 $Y=1.18 $X2=0 $Y2=0
cc_368 N_A_1311_21#_c_370_n N_Y_c_809_n 0.0477562f $X=8.165 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A_1311_21#_c_364_n N_Y_c_810_n 0.0101705f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_370 N_A_1311_21#_c_365_n N_Y_c_810_n 0.00320625f $X=8.04 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_1311_21#_c_419_p N_Y_c_810_n 0.0444453f $X=8.27 $Y=1.18 $X2=0 $Y2=0
cc_372 N_A_1311_21#_c_367_n N_Y_c_810_n 0.010195f $X=8.797 $Y=0.735 $X2=0 $Y2=0
cc_373 N_A_1311_21#_c_368_n N_Y_c_810_n 3.17939e-19 $X=8.82 $Y=0.39 $X2=0 $Y2=0
cc_374 N_A_1311_21#_c_370_n N_Y_c_810_n 0.00768007f $X=8.165 $Y=1.16 $X2=0 $Y2=0
cc_375 N_A_1311_21#_c_373_n N_Y_c_818_n 0.0128188f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_1311_21#_c_419_p N_Y_c_818_n 0.0199914f $X=8.27 $Y=1.18 $X2=0 $Y2=0
cc_377 N_A_1311_21#_c_370_n N_Y_c_818_n 0.00778251f $X=8.165 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_1311_21#_c_363_n N_Y_c_903_n 5.24597e-19 $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A_1311_21#_c_364_n N_Y_c_903_n 0.00651696f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_1311_21#_c_365_n N_Y_c_903_n 0.00758151f $X=8.04 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_1311_21#_c_368_n N_Y_c_903_n 0.00517465f $X=8.82 $Y=0.39 $X2=0 $Y2=0
cc_382 N_A_1311_21#_c_362_n N_Y_c_816_n 0.00224457f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A_1311_21#_c_363_n N_Y_c_816_n 0.0082196f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A_1311_21#_c_371_n N_Y_c_909_n 2.98817e-19 $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A_1311_21#_c_372_n N_Y_c_909_n 0.0107664f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A_1311_21#_c_374_n N_Y_c_819_n 3.54824e-19 $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A_1311_21#_c_419_p N_Y_c_819_n 0.0204252f $X=8.27 $Y=1.18 $X2=0 $Y2=0
cc_388 N_A_1311_21#_c_377_n N_Y_c_819_n 0.00581892f $X=8.44 $Y=1.54 $X2=0 $Y2=0
cc_389 N_A_1311_21#_c_370_n N_Y_c_819_n 0.00655199f $X=8.165 $Y=1.16 $X2=0 $Y2=0
cc_390 N_A_1311_21#_c_367_n N_VGND_M1021_d 0.00423552f $X=8.797 $Y=0.735 $X2=0
+ $Y2=0
cc_391 N_A_1311_21#_c_362_n N_VGND_c_1006_n 0.00268723f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_392 N_A_1311_21#_c_363_n N_VGND_c_1007_n 0.00379224f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_393 N_A_1311_21#_c_364_n N_VGND_c_1007_n 0.00276126f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_394 N_A_1311_21#_c_365_n N_VGND_c_1008_n 0.00530265f $X=8.04 $Y=0.995 $X2=0
+ $Y2=0
cc_395 N_A_1311_21#_c_419_p N_VGND_c_1008_n 0.00178945f $X=8.27 $Y=1.18 $X2=0
+ $Y2=0
cc_396 N_A_1311_21#_c_367_n N_VGND_c_1008_n 0.00851553f $X=8.797 $Y=0.735 $X2=0
+ $Y2=0
cc_397 N_A_1311_21#_c_368_n N_VGND_c_1008_n 0.0193253f $X=8.82 $Y=0.39 $X2=0
+ $Y2=0
cc_398 N_A_1311_21#_c_369_n N_VGND_c_1008_n 0.00110459f $X=8.355 $Y=1.16 $X2=0
+ $Y2=0
cc_399 N_A_1311_21#_c_367_n N_VGND_c_1010_n 0.0111174f $X=8.797 $Y=0.735 $X2=0
+ $Y2=0
cc_400 N_A_1311_21#_c_368_n N_VGND_c_1010_n 0.0300175f $X=8.82 $Y=0.39 $X2=0
+ $Y2=0
cc_401 N_A_1311_21#_c_362_n N_VGND_c_1017_n 0.00423334f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_A_1311_21#_c_363_n N_VGND_c_1017_n 0.00423225f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_403 N_A_1311_21#_c_364_n N_VGND_c_1019_n 0.00423334f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_404 N_A_1311_21#_c_365_n N_VGND_c_1019_n 0.00541359f $X=8.04 $Y=0.995 $X2=0
+ $Y2=0
cc_405 N_A_1311_21#_c_367_n N_VGND_c_1021_n 0.00335436f $X=8.797 $Y=0.735 $X2=0
+ $Y2=0
cc_406 N_A_1311_21#_c_368_n N_VGND_c_1021_n 0.0237059f $X=8.82 $Y=0.39 $X2=0
+ $Y2=0
cc_407 N_A_1311_21#_M1027_s N_VGND_c_1026_n 0.00209319f $X=8.695 $Y=0.235 $X2=0
+ $Y2=0
cc_408 N_A_1311_21#_c_362_n N_VGND_c_1026_n 0.00587047f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_409 N_A_1311_21#_c_363_n N_VGND_c_1026_n 0.00609103f $X=7.1 $Y=0.995 $X2=0
+ $Y2=0
cc_410 N_A_1311_21#_c_364_n N_VGND_c_1026_n 0.00597024f $X=7.57 $Y=0.995 $X2=0
+ $Y2=0
cc_411 N_A_1311_21#_c_365_n N_VGND_c_1026_n 0.0110773f $X=8.04 $Y=0.995 $X2=0
+ $Y2=0
cc_412 N_A_1311_21#_c_367_n N_VGND_c_1026_n 0.00642555f $X=8.797 $Y=0.735 $X2=0
+ $Y2=0
cc_413 N_A_1311_21#_c_368_n N_VGND_c_1026_n 0.0140329f $X=8.82 $Y=0.39 $X2=0
+ $Y2=0
cc_414 N_D_N_c_481_n N_VPWR_c_578_n 0.0141495f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_415 D_N N_VPWR_c_578_n 0.0187446f $X=9.28 $Y=1.105 $X2=0 $Y2=0
cc_416 N_D_N_c_481_n N_VPWR_c_579_n 0.00673617f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_417 N_D_N_c_481_n N_VPWR_c_573_n 0.0141249f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_418 N_D_N_c_480_n N_VGND_c_1008_n 0.00194637f $X=9.03 $Y=0.995 $X2=0 $Y2=0
cc_419 N_D_N_c_480_n N_VGND_c_1010_n 0.00706728f $X=9.03 $Y=0.995 $X2=0 $Y2=0
cc_420 N_D_N_c_481_n N_VGND_c_1010_n 0.00523789f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_421 D_N N_VGND_c_1010_n 0.0187437f $X=9.28 $Y=1.105 $X2=0 $Y2=0
cc_422 N_D_N_c_480_n N_VGND_c_1021_n 0.00540385f $X=9.03 $Y=0.995 $X2=0 $Y2=0
cc_423 N_D_N_c_480_n N_VGND_c_1026_n 0.0119805f $X=9.03 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A_27_297#_c_508_n N_VPWR_M1002_s 0.00182839f $X=1.075 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_425 N_A_27_297#_c_510_n N_VPWR_M1022_s 0.00187091f $X=2.015 $Y=1.54 $X2=0
+ $Y2=0
cc_426 N_A_27_297#_c_507_n N_VPWR_c_574_n 0.0412102f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_427 N_A_27_297#_c_508_n N_VPWR_c_574_n 0.0139937f $X=1.075 $Y=1.54 $X2=0
+ $Y2=0
cc_428 N_A_27_297#_c_538_p N_VPWR_c_575_n 0.0149311f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_429 N_A_27_297#_c_510_n N_VPWR_c_576_n 0.0143191f $X=2.015 $Y=1.54 $X2=0
+ $Y2=0
cc_430 N_A_27_297#_c_540_p N_VPWR_c_579_n 0.015002f $X=2.14 $Y=2.295 $X2=0 $Y2=0
cc_431 N_A_27_297#_c_530_n N_VPWR_c_579_n 0.0386815f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_432 N_A_27_297#_c_512_n N_VPWR_c_579_n 0.0549564f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_433 N_A_27_297#_c_543_p N_VPWR_c_579_n 0.0149886f $X=3.08 $Y=2.38 $X2=0 $Y2=0
cc_434 N_A_27_297#_c_507_n N_VPWR_c_580_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_435 N_A_27_297#_M1002_d N_VPWR_c_573_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_436 N_A_27_297#_M1016_d N_VPWR_c_573_n 0.00370124f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_437 N_A_27_297#_M1030_d N_VPWR_c_573_n 0.00297222f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_438 N_A_27_297#_M1006_d N_VPWR_c_573_n 0.00231264f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_439 N_A_27_297#_M1017_d N_VPWR_c_573_n 0.00217519f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_440 N_A_27_297#_c_507_n N_VPWR_c_573_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_441 N_A_27_297#_c_538_p N_VPWR_c_573_n 0.00955092f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_442 N_A_27_297#_c_540_p N_VPWR_c_573_n 0.00962794f $X=2.14 $Y=2.295 $X2=0
+ $Y2=0
cc_443 N_A_27_297#_c_530_n N_VPWR_c_573_n 0.0239144f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_444 N_A_27_297#_c_512_n N_VPWR_c_573_n 0.0335386f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_445 N_A_27_297#_c_543_p N_VPWR_c_573_n 0.00962421f $X=3.08 $Y=2.38 $X2=0
+ $Y2=0
cc_446 N_A_27_297#_c_530_n N_A_493_297#_M1000_s 0.00352392f $X=2.955 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_447 N_A_27_297#_c_512_n N_A_493_297#_M1009_s 0.00352392f $X=3.895 $Y=2.38
+ $X2=0 $Y2=0
cc_448 N_A_27_297#_M1006_d N_A_493_297#_c_677_n 0.00187091f $X=2.935 $Y=1.485
+ $X2=0 $Y2=0
cc_449 N_A_27_297#_c_530_n N_A_493_297#_c_677_n 0.00385532f $X=2.955 $Y=2.38
+ $X2=0 $Y2=0
cc_450 N_A_27_297#_c_560_p N_A_493_297#_c_677_n 0.0143018f $X=3.08 $Y=1.96 $X2=0
+ $Y2=0
cc_451 N_A_27_297#_c_512_n N_A_493_297#_c_677_n 0.00385532f $X=3.895 $Y=2.38
+ $X2=0 $Y2=0
cc_452 N_A_27_297#_M1017_d N_A_493_297#_c_678_n 0.00294603f $X=3.875 $Y=1.485
+ $X2=0 $Y2=0
cc_453 N_A_27_297#_c_512_n N_A_493_297#_c_678_n 0.00385532f $X=3.895 $Y=2.38
+ $X2=0 $Y2=0
cc_454 N_A_27_297#_c_564_p N_A_493_297#_c_678_n 0.0172271f $X=4.02 $Y=1.96 $X2=0
+ $Y2=0
cc_455 N_A_27_297#_c_511_n N_A_493_297#_c_680_n 0.00226124f $X=2.14 $Y=1.625
+ $X2=0 $Y2=0
cc_456 N_A_27_297#_c_530_n N_A_493_297#_c_680_n 0.013395f $X=2.955 $Y=2.38 $X2=0
+ $Y2=0
cc_457 N_A_27_297#_c_512_n N_A_493_297#_c_681_n 0.013395f $X=3.895 $Y=2.38 $X2=0
+ $Y2=0
cc_458 N_A_27_297#_c_564_p N_A_883_297#_c_757_n 0.027317f $X=4.02 $Y=1.96 $X2=0
+ $Y2=0
cc_459 N_A_27_297#_c_512_n N_A_883_297#_c_737_n 0.0108671f $X=3.895 $Y=2.38
+ $X2=0 $Y2=0
cc_460 N_A_27_297#_c_510_n N_Y_c_804_n 3.18413e-19 $X=2.015 $Y=1.54 $X2=0 $Y2=0
cc_461 N_A_27_297#_c_511_n N_Y_c_804_n 0.00936521f $X=2.14 $Y=1.625 $X2=0 $Y2=0
cc_462 N_A_27_297#_c_509_n N_VGND_c_999_n 0.00684525f $X=0.425 $Y=1.54 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_573_n N_A_493_297#_M1000_s 0.00232895f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_464 N_VPWR_c_573_n N_A_493_297#_M1009_s 0.00232895f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_573_n N_A_493_297#_M1004_d 0.00232895f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_573_n N_A_493_297#_M1020_d 0.00232895f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_573_n N_A_883_297#_M1004_s 0.00217519f $X=9.43 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_468 N_VPWR_c_573_n N_A_883_297#_M1007_s 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_573_n N_A_883_297#_M1031_s 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_573_n N_A_883_297#_M1018_s 0.00231264f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_573_n N_A_883_297#_M1026_s 0.00217519f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_579_n N_A_883_297#_c_740_n 0.0386815f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_573_n N_A_883_297#_c_740_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_579_n N_A_883_297#_c_737_n 0.0162749f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_573_n N_A_883_297#_c_737_n 0.00962421f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_579_n N_A_883_297#_c_742_n 0.0386815f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_573_n N_A_883_297#_c_742_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_579_n N_A_883_297#_c_747_n 0.0386815f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_573_n N_A_883_297#_c_747_n 0.0239144f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_579_n N_A_883_297#_c_739_n 0.0549564f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_573_n N_A_883_297#_c_739_n 0.0335386f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_579_n N_A_883_297#_c_774_n 0.0149886f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_573_n N_A_883_297#_c_774_n 0.00962421f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_579_n N_A_883_297#_c_776_n 0.015002f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_573_n N_A_883_297#_c_776_n 0.00961749f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_579_n N_A_883_297#_c_778_n 0.0149886f $X=9.205 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_573_n N_A_883_297#_c_778_n 0.00962421f $X=9.43 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_573_n N_Y_M1012_d 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_489 N_VPWR_c_573_n N_Y_M1023_d 0.00232895f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_490 N_A_493_297#_c_678_n N_A_883_297#_M1004_s 0.00294603f $X=4.885 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_491 N_A_493_297#_c_679_n N_A_883_297#_M1007_s 0.00187091f $X=5.825 $Y=1.54
+ $X2=0 $Y2=0
cc_492 N_A_493_297#_c_678_n N_A_883_297#_c_757_n 0.0172271f $X=4.885 $Y=1.54
+ $X2=0 $Y2=0
cc_493 N_A_493_297#_M1004_d N_A_883_297#_c_740_n 0.00352392f $X=4.865 $Y=1.485
+ $X2=0 $Y2=0
cc_494 N_A_493_297#_c_678_n N_A_883_297#_c_740_n 0.00385532f $X=4.885 $Y=1.54
+ $X2=0 $Y2=0
cc_495 N_A_493_297#_c_679_n N_A_883_297#_c_740_n 0.00385532f $X=5.825 $Y=1.54
+ $X2=0 $Y2=0
cc_496 N_A_493_297#_c_682_n N_A_883_297#_c_740_n 0.013395f $X=5.01 $Y=1.62 $X2=0
+ $Y2=0
cc_497 N_A_493_297#_c_679_n N_A_883_297#_c_787_n 0.0143018f $X=5.825 $Y=1.54
+ $X2=0 $Y2=0
cc_498 N_A_493_297#_M1020_d N_A_883_297#_c_742_n 0.00352392f $X=5.805 $Y=1.485
+ $X2=0 $Y2=0
cc_499 N_A_493_297#_c_679_n N_A_883_297#_c_742_n 0.00385532f $X=5.825 $Y=1.54
+ $X2=0 $Y2=0
cc_500 N_A_493_297#_c_683_n N_A_883_297#_c_742_n 0.013395f $X=5.95 $Y=1.62 $X2=0
+ $Y2=0
cc_501 N_A_493_297#_c_683_n N_A_883_297#_c_738_n 0.00209545f $X=5.95 $Y=1.62
+ $X2=0 $Y2=0
cc_502 N_A_493_297#_c_678_n N_Y_c_806_n 0.00787473f $X=4.885 $Y=1.54 $X2=0 $Y2=0
cc_503 N_A_883_297#_c_747_n N_Y_M1012_d 0.00352392f $X=7.235 $Y=2.38 $X2=0 $Y2=0
cc_504 N_A_883_297#_c_739_n N_Y_M1023_d 0.00352392f $X=8.175 $Y=2.38 $X2=0 $Y2=0
cc_505 N_A_883_297#_c_738_n N_Y_c_808_n 0.00929029f $X=6.42 $Y=1.62 $X2=0 $Y2=0
cc_506 N_A_883_297#_M1018_s N_Y_c_818_n 0.00187091f $X=7.215 $Y=1.485 $X2=0
+ $Y2=0
cc_507 N_A_883_297#_c_749_n N_Y_c_818_n 0.0143018f $X=7.36 $Y=1.96 $X2=0 $Y2=0
cc_508 N_A_883_297#_c_739_n N_Y_c_818_n 0.00385532f $X=8.175 $Y=2.38 $X2=0 $Y2=0
cc_509 N_A_883_297#_c_738_n N_Y_c_909_n 0.00209545f $X=6.42 $Y=1.62 $X2=0 $Y2=0
cc_510 N_A_883_297#_c_747_n N_Y_c_909_n 0.00431849f $X=7.235 $Y=2.38 $X2=0 $Y2=0
cc_511 N_A_883_297#_c_739_n N_Y_c_819_n 0.013395f $X=8.175 $Y=2.38 $X2=0 $Y2=0
cc_512 N_A_883_297#_c_747_n Y 0.0134104f $X=7.235 $Y=2.38 $X2=0 $Y2=0
cc_513 N_Y_c_802_n N_VGND_M1010_s 0.00251047f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_514 N_Y_c_804_n N_VGND_M1032_s 0.00162089f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_515 N_Y_c_805_n N_VGND_M1019_d 0.00251047f $X=3.335 $Y=0.815 $X2=0 $Y2=0
cc_516 N_Y_c_806_n N_VGND_M1029_d 0.0108248f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_517 N_Y_c_807_n N_VGND_M1015_d 0.00251047f $X=5.735 $Y=0.815 $X2=0 $Y2=0
cc_518 N_Y_c_808_n N_VGND_M1033_d 0.00162089f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_519 N_Y_c_810_n N_VGND_M1003_d 0.00214495f $X=7.615 $Y=0.815 $X2=0 $Y2=0
cc_520 N_Y_c_816_n N_VGND_M1003_d 3.6276e-19 $X=6.962 $Y=0.815 $X2=0 $Y2=0
cc_521 N_Y_c_803_n N_VGND_c_999_n 0.00750114f $X=0.895 $Y=0.815 $X2=0 $Y2=0
cc_522 N_Y_c_820_n N_VGND_c_1000_n 0.0223596f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_523 N_Y_c_802_n N_VGND_c_1000_n 0.00266636f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_524 N_Y_c_820_n N_VGND_c_1001_n 0.0183628f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_525 N_Y_c_802_n N_VGND_c_1001_n 0.0127273f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_526 N_Y_c_802_n N_VGND_c_1002_n 0.00198695f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_527 N_Y_c_831_n N_VGND_c_1002_n 0.0231806f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_528 N_Y_c_804_n N_VGND_c_1002_n 0.00254521f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_529 N_Y_c_804_n N_VGND_c_1003_n 0.0122559f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_530 N_Y_c_835_n N_VGND_c_1004_n 0.0183628f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_531 N_Y_c_805_n N_VGND_c_1004_n 0.0127273f $X=3.335 $Y=0.815 $X2=0 $Y2=0
cc_532 N_Y_c_861_n N_VGND_c_1005_n 0.0183628f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_533 N_Y_c_807_n N_VGND_c_1005_n 0.0127273f $X=5.735 $Y=0.815 $X2=0 $Y2=0
cc_534 N_Y_c_808_n N_VGND_c_1006_n 0.0122559f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_535 N_Y_c_872_n N_VGND_c_1007_n 0.0183628f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_536 N_Y_c_810_n N_VGND_c_1007_n 0.0127273f $X=7.615 $Y=0.815 $X2=0 $Y2=0
cc_537 N_Y_c_903_n N_VGND_c_1008_n 0.0183628f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_538 N_Y_c_804_n N_VGND_c_1011_n 0.00198695f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_539 N_Y_c_835_n N_VGND_c_1011_n 0.0223596f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_540 N_Y_c_805_n N_VGND_c_1011_n 0.00266636f $X=3.335 $Y=0.815 $X2=0 $Y2=0
cc_541 N_Y_c_806_n N_VGND_c_1013_n 0.00198695f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_542 N_Y_c_861_n N_VGND_c_1013_n 0.0223596f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_543 N_Y_c_807_n N_VGND_c_1013_n 0.00266636f $X=5.735 $Y=0.815 $X2=0 $Y2=0
cc_544 N_Y_c_807_n N_VGND_c_1015_n 0.00198695f $X=5.735 $Y=0.815 $X2=0 $Y2=0
cc_545 N_Y_c_868_n N_VGND_c_1015_n 0.0231806f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_546 N_Y_c_808_n N_VGND_c_1015_n 0.00254521f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_547 N_Y_c_808_n N_VGND_c_1017_n 0.00198695f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_548 N_Y_c_872_n N_VGND_c_1017_n 0.022413f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_549 N_Y_c_810_n N_VGND_c_1017_n 3.48906e-19 $X=7.615 $Y=0.815 $X2=0 $Y2=0
cc_550 N_Y_c_816_n N_VGND_c_1017_n 0.00250291f $X=6.962 $Y=0.815 $X2=0 $Y2=0
cc_551 N_Y_c_810_n N_VGND_c_1019_n 0.00198695f $X=7.615 $Y=0.815 $X2=0 $Y2=0
cc_552 N_Y_c_903_n N_VGND_c_1019_n 0.0223596f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_553 N_Y_c_805_n N_VGND_c_1024_n 0.00198695f $X=3.335 $Y=0.815 $X2=0 $Y2=0
cc_554 N_Y_c_848_n N_VGND_c_1024_n 0.0231806f $X=3.55 $Y=0.39 $X2=0 $Y2=0
cc_555 N_Y_c_806_n N_VGND_c_1024_n 0.00254521f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_556 N_Y_c_806_n N_VGND_c_1025_n 0.0528344f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_557 N_Y_M1008_d N_VGND_c_1026_n 0.0025535f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_558 N_Y_M1025_d N_VGND_c_1026_n 0.00304143f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_559 N_Y_M1011_s N_VGND_c_1026_n 0.0025535f $X=2.425 $Y=0.235 $X2=0 $Y2=0
cc_560 N_Y_M1028_s N_VGND_c_1026_n 0.00304143f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_561 N_Y_M1005_s N_VGND_c_1026_n 0.0025535f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_562 N_Y_M1024_s N_VGND_c_1026_n 0.00304143f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_563 N_Y_M1001_s N_VGND_c_1026_n 0.0025535f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_564 N_Y_M1014_s N_VGND_c_1026_n 0.0025535f $X=7.645 $Y=0.235 $X2=0 $Y2=0
cc_565 N_Y_c_820_n N_VGND_c_1026_n 0.0141302f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_566 N_Y_c_802_n N_VGND_c_1026_n 0.00972452f $X=1.455 $Y=0.815 $X2=0 $Y2=0
cc_567 N_Y_c_831_n N_VGND_c_1026_n 0.0143352f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_568 N_Y_c_804_n N_VGND_c_1026_n 0.0094839f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_569 N_Y_c_835_n N_VGND_c_1026_n 0.0141302f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_570 N_Y_c_805_n N_VGND_c_1026_n 0.00972452f $X=3.335 $Y=0.815 $X2=0 $Y2=0
cc_571 N_Y_c_848_n N_VGND_c_1026_n 0.0143352f $X=3.55 $Y=0.39 $X2=0 $Y2=0
cc_572 N_Y_c_806_n N_VGND_c_1026_n 0.0114512f $X=4.795 $Y=0.815 $X2=0 $Y2=0
cc_573 N_Y_c_861_n N_VGND_c_1026_n 0.0141302f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_574 N_Y_c_807_n N_VGND_c_1026_n 0.00972452f $X=5.735 $Y=0.815 $X2=0 $Y2=0
cc_575 N_Y_c_868_n N_VGND_c_1026_n 0.0143352f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_576 N_Y_c_808_n N_VGND_c_1026_n 0.0094839f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_577 N_Y_c_872_n N_VGND_c_1026_n 0.0141433f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_578 N_Y_c_810_n N_VGND_c_1026_n 0.0051951f $X=7.615 $Y=0.815 $X2=0 $Y2=0
cc_579 N_Y_c_903_n N_VGND_c_1026_n 0.0141302f $X=7.83 $Y=0.39 $X2=0 $Y2=0
cc_580 N_Y_c_816_n N_VGND_c_1026_n 0.00483502f $X=6.962 $Y=0.815 $X2=0 $Y2=0
