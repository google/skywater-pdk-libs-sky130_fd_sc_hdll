* File: sky130_fd_sc_hdll__nand3b_1.pex.spice
* Created: Wed Sep  2 08:37:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%A_N 1 3 4 6 7
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.16 $X2=0.51 $Y2=1.16
r27 7 11 6.28605 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=0.69 $Y=1.16 $X2=0.51
+ $Y2=1.16
r28 4 10 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=0.65 $Y=0.995
+ $X2=0.535 $Y2=1.16
r29 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.65 $Y=0.995 $X2=0.65
+ $Y2=0.675
r30 1 10 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=0.625 $Y=1.41
+ $X2=0.535 $Y2=1.16
r31 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.625 $Y=1.41
+ $X2=0.625 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%C 1 3 4 6 7 14
r27 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.1
+ $Y=1.16 $X2=1.1 $Y2=1.16
r28 7 14 3.5621 $w=3.28e-07 $l=1.02e-07 $layer=LI1_cond $X=1.202 $Y=1.16 $X2=1.1
+ $Y2=1.16
r29 4 10 38.5562 $w=2.99e-07 $l=2.04316e-07 $layer=POLY_cond $X=1.185 $Y=0.995
+ $X2=1.097 $Y2=1.16
r30 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.185 $Y=0.995
+ $X2=1.185 $Y2=0.56
r31 1 10 47.8775 $w=2.99e-07 $l=2.79732e-07 $layer=POLY_cond $X=1.16 $Y=1.41
+ $X2=1.097 $Y2=1.16
r32 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.16 $Y=1.41 $X2=1.16
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%B 1 3 4 6 7 14
r31 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.16 $X2=1.605 $Y2=1.16
r32 7 14 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=1.71 $Y=1.16
+ $X2=1.605 $Y2=1.16
r33 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.665 $Y=0.995
+ $X2=1.605 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.665 $Y=0.995
+ $X2=1.665 $Y2=0.56
r35 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.64 $Y=1.41
+ $X2=1.605 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.64 $Y=1.41 $X2=1.64
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%A_53_93# 1 2 7 9 10 12 14 15 19 26 30
c61 19 0 1.78374e-19 $X=2.085 $Y=1.16
r62 27 30 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=0.17 $Y=1.76
+ $X2=0.39 $Y2=1.76
r63 25 26 7.20646 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=0.39 $Y=0.635
+ $X2=0.51 $Y2=0.635
r64 22 25 6.67204 $w=3.78e-07 $l=2.2e-07 $layer=LI1_cond $X=0.17 $Y=0.635
+ $X2=0.39 $Y2=0.635
r65 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.085
+ $Y=1.16 $X2=2.085 $Y2=1.16
r66 17 19 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=2.11 $Y=0.825
+ $X2=2.11 $Y2=1.16
r67 15 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2 $Y=0.74
+ $X2=2.11 $Y2=0.825
r68 15 26 97.2086 $w=1.68e-07 $l=1.49e-06 $layer=LI1_cond $X=2 $Y=0.74 $X2=0.51
+ $Y2=0.74
r69 14 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.17 $Y=1.595
+ $X2=0.17 $Y2=1.76
r70 13 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.635
r71 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.595
r72 10 20 39.2931 $w=2.55e-07 $l=1.90526e-07 $layer=POLY_cond $X=2.14 $Y=0.995
+ $X2=2.085 $Y2=1.16
r73 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.14 $Y=0.995
+ $X2=2.14 $Y2=0.56
r74 7 20 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.12 $Y=1.41
+ $X2=2.085 $Y2=1.16
r75 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.12 $Y=1.41 $X2=2.12
+ $Y2=1.985
r76 2 30 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=0.265
+ $Y=1.485 $X2=0.39 $Y2=1.76
r77 1 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.265
+ $Y=0.465 $X2=0.39 $Y2=0.61
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%VPWR 1 2 9 15 18 19 21 22 23 33 34
r37 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 27 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r41 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 23 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 21 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.79 $Y=2.72
+ $X2=1.61 $Y2=2.72
r44 21 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=2.72
+ $X2=1.875 $Y2=2.72
r45 20 33 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 20 22 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.96 $Y=2.72
+ $X2=1.875 $Y2=2.72
r47 18 26 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.76 $Y=2.72 $X2=0.69
+ $Y2=2.72
r48 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.76 $Y=2.72
+ $X2=0.885 $Y2=2.72
r49 17 30 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.01 $Y=2.72 $X2=1.61
+ $Y2=2.72
r50 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.01 $Y=2.72
+ $X2=0.885 $Y2=2.72
r51 13 22 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=2.635
+ $X2=1.875 $Y2=2.72
r52 13 15 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.875 $Y=2.635
+ $X2=1.875 $Y2=2
r53 9 12 15.6732 $w=2.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.885 $Y=1.66
+ $X2=0.885 $Y2=2
r54 7 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.885 $Y=2.635
+ $X2=0.885 $Y2=2.72
r55 7 12 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=0.885 $Y=2.635
+ $X2=0.885 $Y2=2
r56 2 15 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.73
+ $Y=1.485 $X2=1.875 $Y2=2
r57 1 12 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=0.715
+ $Y=1.485 $X2=0.925 $Y2=2
r58 1 9 600 $w=1.7e-07 $l=2.84341e-07 $layer=licon1_PDIFF $count=1 $X=0.715
+ $Y=1.485 $X2=0.925 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%Y 1 2 3 10 12 14 16 22 23 24 25 26 27 36
+ 39
r45 36 39 1.08721 $w=2.63e-07 $l=2.5e-08 $layer=LI1_cond $X=2.542 $Y=0.485
+ $X2=2.542 $Y2=0.51
r46 27 52 2.7433 $w=5.43e-07 $l=1.25e-07 $layer=LI1_cond $X=2.402 $Y=2.21
+ $X2=2.402 $Y2=2.335
r47 26 27 7.46177 $w=5.43e-07 $l=3.4e-07 $layer=LI1_cond $X=2.402 $Y=1.87
+ $X2=2.402 $Y2=2.21
r48 26 46 4.49901 $w=5.43e-07 $l=2.05e-07 $layer=LI1_cond $X=2.402 $Y=1.87
+ $X2=2.402 $Y2=1.665
r49 25 37 2.39067 $w=4.05e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.402 $Y=1.58
+ $X2=2.542 $Y2=1.495
r50 25 46 2.39067 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=2.402 $Y=1.58
+ $X2=2.402 $Y2=1.665
r51 25 37 1.08721 $w=2.63e-07 $l=2.5e-08 $layer=LI1_cond $X=2.542 $Y=1.47
+ $X2=2.542 $Y2=1.495
r52 24 25 12.1768 $w=2.63e-07 $l=2.8e-07 $layer=LI1_cond $X=2.542 $Y=1.19
+ $X2=2.542 $Y2=1.47
r53 23 24 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.542 $Y=0.85
+ $X2=2.542 $Y2=1.19
r54 22 36 3.19435 $w=2.65e-07 $l=1.15e-07 $layer=LI1_cond $X=2.542 $Y=0.37
+ $X2=2.542 $Y2=0.485
r55 22 23 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=2.542 $Y=0.54
+ $X2=2.542 $Y2=0.85
r56 22 39 1.30465 $w=2.63e-07 $l=3e-08 $layer=LI1_cond $X=2.542 $Y=0.54
+ $X2=2.542 $Y2=0.51
r57 16 22 3.66656 $w=2.3e-07 $l=1.32e-07 $layer=LI1_cond $X=2.41 $Y=0.37
+ $X2=2.542 $Y2=0.37
r58 16 18 2.75584 $w=2.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.41 $Y=0.37
+ $X2=2.355 $Y2=0.37
r59 15 21 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.56 $Y=1.58 $X2=1.37
+ $Y2=1.58
r60 14 25 4.59089 $w=1.7e-07 $l=2.72e-07 $layer=LI1_cond $X=2.13 $Y=1.58
+ $X2=2.402 $Y2=1.58
r61 14 15 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.13 $Y=1.58
+ $X2=1.56 $Y2=1.58
r62 10 21 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=1.665
+ $X2=1.37 $Y2=1.58
r63 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.37 $Y=1.665
+ $X2=1.37 $Y2=2.34
r64 3 25 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.485 $X2=2.355 $Y2=1.655
r65 3 52 400 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=2.21
+ $Y=1.485 $X2=2.355 $Y2=2.335
r66 2 21 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.485 $X2=1.395 $Y2=1.66
r67 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.25
+ $Y=1.485 $X2=1.395 $Y2=2.34
r68 1 18 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.235 $X2=2.355 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_1%VGND 1 6 9 10 11 21 22
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r31 19 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r32 18 21 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r33 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r34 15 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r35 14 15 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r36 11 15 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r37 9 14 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.69
+ $Y2=0
r38 9 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.76 $Y=0 $X2=0.925
+ $Y2=0
r39 8 18 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.15
+ $Y2=0
r40 8 10 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.925
+ $Y2=0
r41 4 10 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0
r42 4 6 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.925 $Y=0.085
+ $X2=0.925 $Y2=0.38
r43 1 6 182 $w=1.7e-07 $l=2.38747e-07 $layer=licon1_NDIFF $count=1 $X=0.725
+ $Y=0.465 $X2=0.925 $Y2=0.38
.ends

