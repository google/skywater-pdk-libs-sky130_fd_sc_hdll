* File: sky130_fd_sc_hdll__o211ai_2.pex.spice
* Created: Wed Sep  2 08:42:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%C1 1 3 4 6 7 9 10 12 13 17 20
c41 10 0 3.94966e-20 $X=1.025 $Y=0.995
r42 20 21 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=1 $Y=1.202
+ $X2=1.025 $Y2=1.202
r43 19 20 60.25 $w=3.64e-07 $l=4.55e-07 $layer=POLY_cond $X=0.545 $Y=1.202 $X2=1
+ $Y2=1.202
r44 18 19 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.545 $Y2=1.202
r45 16 18 37.0769 $w=3.64e-07 $l=2.8e-07 $layer=POLY_cond $X=0.24 $Y=1.202
+ $X2=0.52 $Y2=1.202
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r47 13 17 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=1.53
+ $X2=0.23 $Y2=1.16
r48 10 21 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.56
r50 7 20 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.985
r52 4 19 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=1.202
r53 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.545 $Y=0.995
+ $X2=0.545 $Y2=0.56
r54 1 18 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.202
r55 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41 $X2=0.52
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%B1 1 3 4 6 7 9 10 12 13 22 23 29
r49 23 24 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=1.96 $Y=1.202
+ $X2=1.985 $Y2=1.202
r50 22 29 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.835 $Y=1.22
+ $X2=1.61 $Y2=1.22
r51 21 23 16.0667 $w=3.75e-07 $l=1.25e-07 $layer=POLY_cond $X=1.835 $Y=1.202
+ $X2=1.96 $Y2=1.202
r52 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.835
+ $Y=1.16 $X2=1.835 $Y2=1.16
r53 19 21 42.416 $w=3.75e-07 $l=3.3e-07 $layer=POLY_cond $X=1.505 $Y=1.202
+ $X2=1.835 $Y2=1.202
r54 18 19 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=1.48 $Y=1.202
+ $X2=1.505 $Y2=1.202
r55 16 18 4.49867 $w=3.75e-07 $l=3.5e-08 $layer=POLY_cond $X=1.445 $Y=1.202
+ $X2=1.48 $Y2=1.202
r56 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.445
+ $Y=1.16 $X2=1.445 $Y2=1.16
r57 13 29 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=1.595 $Y=1.22
+ $X2=1.61 $Y2=1.22
r58 13 17 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=1.595 $Y=1.22
+ $X2=1.445 $Y2=1.22
r59 10 24 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=1.202
r60 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=0.56
r61 7 23 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.202
r62 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.96 $Y=1.41 $X2=1.96
+ $Y2=1.985
r63 4 19 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.505 $Y=0.995
+ $X2=1.505 $Y2=1.202
r64 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.505 $Y=0.995
+ $X2=1.505 $Y2=0.56
r65 1 18 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.48 $Y=1.41
+ $X2=1.48 $Y2=1.202
r66 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.48 $Y=1.41 $X2=1.48
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%A2 1 3 4 6 7 9 10 12 13 19 20 23
r43 20 21 6.39257 $w=3.77e-07 $l=5e-08 $layer=POLY_cond $X=3.48 $Y=1.202
+ $X2=3.53 $Y2=1.202
r44 18 20 7.67109 $w=3.77e-07 $l=6e-08 $layer=POLY_cond $X=3.42 $Y=1.202
+ $X2=3.48 $Y2=1.202
r45 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.42
+ $Y=1.16 $X2=3.42 $Y2=1.16
r46 16 18 50.5013 $w=3.77e-07 $l=3.95e-07 $layer=POLY_cond $X=3.025 $Y=1.202
+ $X2=3.42 $Y2=1.202
r47 15 16 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=3 $Y=1.202
+ $X2=3.025 $Y2=1.202
r48 13 19 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.99 $Y=1.215
+ $X2=3.42 $Y2=1.215
r49 13 23 0.823174 $w=2.78e-07 $l=2e-08 $layer=LI1_cond $X=2.99 $Y=1.215
+ $X2=2.97 $Y2=1.215
r50 10 21 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=1.202
r51 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.53 $Y=0.995
+ $X2=3.53 $Y2=0.56
r52 7 20 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.48 $Y2=1.202
r53 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.48 $Y=1.41 $X2=3.48
+ $Y2=1.985
r54 4 16 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=1.202
r55 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=0.56
r56 1 15 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3 $Y=1.41 $X2=3
+ $Y2=1.202
r57 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3 $Y=1.41 $X2=3
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%A1 1 3 4 6 7 9 10 12 13 18 23
c42 1 0 8.33369e-20 $X=3.96 $Y=1.41
r43 23 24 3.83554 $w=3.77e-07 $l=3e-08 $layer=POLY_cond $X=4.44 $Y=1.202
+ $X2=4.47 $Y2=1.202
r44 20 21 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=3.96 $Y=1.202
+ $X2=3.985 $Y2=1.202
r45 18 28 8.90414 $w=4.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.69 $Y=0.85
+ $X2=4.69 $Y2=1.185
r46 16 23 10.2281 $w=3.77e-07 $l=8e-08 $layer=POLY_cond $X=4.36 $Y=1.202
+ $X2=4.44 $Y2=1.202
r47 16 21 47.9443 $w=3.77e-07 $l=3.75e-07 $layer=POLY_cond $X=4.36 $Y=1.202
+ $X2=3.985 $Y2=1.202
r48 15 16 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.36
+ $Y=1.16 $X2=4.36 $Y2=1.16
r49 13 28 4.9351 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=4.465 $Y=1.185
+ $X2=4.69 $Y2=1.185
r50 13 15 5.5003 $w=2.18e-07 $l=1.05e-07 $layer=LI1_cond $X=4.465 $Y=1.185
+ $X2=4.36 $Y2=1.185
r51 10 24 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=1.202
r52 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.47 $Y=0.995
+ $X2=4.47 $Y2=0.56
r53 7 23 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.44 $Y=1.41
+ $X2=4.44 $Y2=1.202
r54 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.44 $Y=1.41 $X2=4.44
+ $Y2=1.985
r55 4 21 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.985 $Y2=1.202
r56 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.985 $Y2=0.56
r57 1 20 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.96 $Y=1.41
+ $X2=3.96 $Y2=1.202
r58 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.96 $Y=1.41 $X2=3.96
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%VPWR 1 2 3 4 13 15 19 23 27 30 31 32 34
+ 39 52 53 59 62
r69 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r70 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r72 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r73 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 47 50 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 47 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r76 46 49 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r77 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 44 62 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.175 $Y2=2.72
r79 44 46 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.365 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 43 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r81 43 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r82 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r83 40 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.405 $Y=2.72
+ $X2=1.215 $Y2=2.72
r84 40 42 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=1.405 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 39 62 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.985 $Y=2.72
+ $X2=2.175 $Y2=2.72
r86 39 42 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.985 $Y=2.72
+ $X2=1.61 $Y2=2.72
r87 38 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r89 35 56 4.09637 $w=1.7e-07 $l=1.88e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.187 $Y2=2.72
r90 35 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.375 $Y=2.72
+ $X2=0.69 $Y2=2.72
r91 34 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=1.215 $Y2=2.72
r92 34 37 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=0.69 $Y2=2.72
r93 32 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 32 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 30 49 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 30 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=4.175 $Y2=2.72
r97 29 52 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.365 $Y=2.72
+ $X2=4.83 $Y2=2.72
r98 29 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.365 $Y=2.72
+ $X2=4.175 $Y2=2.72
r99 25 31 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=2.635
+ $X2=4.175 $Y2=2.72
r100 25 27 20.7743 $w=3.78e-07 $l=6.85e-07 $layer=LI1_cond $X=4.175 $Y=2.635
+ $X2=4.175 $Y2=1.95
r101 21 62 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.175 $Y=2.635
+ $X2=2.175 $Y2=2.72
r102 21 23 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.175 $Y=2.635
+ $X2=2.175 $Y2=2
r103 17 59 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=2.72
r104 17 19 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=2
r105 13 56 3.11585 $w=2.6e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.187 $Y2=2.72
r106 13 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2.34
r107 4 27 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=4.05
+ $Y=1.485 $X2=4.2 $Y2=1.95
r108 3 23 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.485 $X2=2.2 $Y2=2
r109 2 19 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.24 $Y2=2
r110 1 15 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.155
+ $Y=1.485 $X2=0.28 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%Y 1 2 3 4 15 17 21 23 28 29 31 32 35
c50 31 0 8.33369e-20 $X=3.24 $Y=1.7
r51 32 35 2.72947 $w=3.78e-07 $l=9e-08 $layer=LI1_cond $X=0.735 $Y=0.85
+ $X2=0.735 $Y2=0.76
r52 27 32 20.9259 $w=3.78e-07 $l=6.9e-07 $layer=LI1_cond $X=0.735 $Y=1.54
+ $X2=0.735 $Y2=0.85
r53 27 28 2.7724 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.54
+ $X2=0.735 $Y2=1.625
r54 24 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.815 $Y=1.625
+ $X2=1.72 $Y2=1.625
r55 23 31 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.025 $Y=1.625
+ $X2=3.215 $Y2=1.625
r56 23 24 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.025 $Y=1.625
+ $X2=1.815 $Y2=1.625
r57 19 29 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=1.71
+ $X2=1.72 $Y2=1.625
r58 19 21 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.72 $Y=1.71
+ $X2=1.72 $Y2=1.845
r59 18 28 3.97867 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.925 $Y=1.625
+ $X2=0.735 $Y2=1.625
r60 17 29 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.625 $Y=1.625
+ $X2=1.72 $Y2=1.625
r61 17 18 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.625 $Y=1.625
+ $X2=0.925 $Y2=1.625
r62 13 28 2.7724 $w=3.45e-07 $l=1.00995e-07 $layer=LI1_cond $X=0.7 $Y=1.71
+ $X2=0.735 $Y2=1.625
r63 13 15 4.08931 $w=3.08e-07 $l=1.1e-07 $layer=LI1_cond $X=0.7 $Y=1.71 $X2=0.7
+ $Y2=1.82
r64 4 31 300 $w=1.7e-07 $l=2.80134e-07 $layer=licon1_PDIFF $count=2 $X=3.09
+ $Y=1.485 $X2=3.24 $Y2=1.7
r65 3 21 300 $w=1.7e-07 $l=4.28486e-07 $layer=licon1_PDIFF $count=2 $X=1.57
+ $Y=1.485 $X2=1.72 $Y2=1.845
r66 2 15 300 $w=1.7e-07 $l=4.03082e-07 $layer=licon1_PDIFF $count=2 $X=0.61
+ $Y=1.485 $X2=0.76 $Y2=1.82
r67 1 35 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.62
+ $Y=0.235 $X2=0.76 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%A_527_297# 1 2 3 10 16 17 20 23
r29 23 25 3.54598 $w=2.58e-07 $l=8e-08 $layer=LI1_cond $X=2.725 $Y=2.3 $X2=2.725
+ $Y2=2.38
r30 18 20 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=4.715 $Y=1.695
+ $X2=4.715 $Y2=1.96
r31 16 18 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.585 $Y=1.61
+ $X2=4.715 $Y2=1.695
r32 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.585 $Y=1.61
+ $X2=3.815 $Y2=1.61
r33 13 15 27.4354 $w=1.88e-07 $l=4.7e-07 $layer=LI1_cond $X=3.72 $Y=2.295
+ $X2=3.72 $Y2=1.825
r34 12 17 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.72 $Y=1.695
+ $X2=3.815 $Y2=1.61
r35 12 15 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=3.72 $Y=1.695
+ $X2=3.72 $Y2=1.825
r36 11 25 3.22376 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.855 $Y=2.38
+ $X2=2.725 $Y2=2.38
r37 10 13 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=3.625 $Y=2.38
+ $X2=3.72 $Y2=2.295
r38 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.625 $Y=2.38
+ $X2=2.855 $Y2=2.38
r39 3 20 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=4.53
+ $Y=1.485 $X2=4.68 $Y2=1.96
r40 2 15 300 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=2 $X=3.57
+ $Y=1.485 $X2=3.72 $Y2=1.825
r41 1 23 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.485 $X2=2.76 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%A_27_47# 1 2 3 10 16 20 23
c32 16 0 3.94966e-20 $X=1.24 $Y=0.705
r33 18 23 4.9491 $w=2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.335 $Y=0.36 $X2=1.24
+ $Y2=0.36
r34 18 20 45.684 $w=2.08e-07 $l=8.65e-07 $layer=LI1_cond $X=1.335 $Y=0.36
+ $X2=2.2 $Y2=0.36
r35 14 23 1.5279 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=1.24 $Y=0.465
+ $X2=1.24 $Y2=0.36
r36 14 16 14.0096 $w=1.88e-07 $l=2.4e-07 $layer=LI1_cond $X=1.24 $Y=0.465
+ $X2=1.24 $Y2=0.705
r37 10 23 4.9491 $w=2e-07 $l=9.98749e-08 $layer=LI1_cond $X=1.145 $Y=0.35
+ $X2=1.24 $Y2=0.36
r38 10 12 50.4928 $w=1.88e-07 $l=8.65e-07 $layer=LI1_cond $X=1.145 $Y=0.35
+ $X2=0.28 $Y2=0.35
r39 3 20 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.235 $X2=2.2 $Y2=0.36
r40 2 23 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.24 $Y2=0.36
r41 2 16 182 $w=1.7e-07 $l=5.35444e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.24 $Y2=0.705
r42 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%A_316_47# 1 2 3 10 17
r32 17 19 3.50239 $w=1.88e-07 $l=6e-08 $layer=LI1_cond $X=4.2 $Y=0.68 $X2=4.2
+ $Y2=0.74
r33 12 15 80.2771 $w=2.08e-07 $l=1.52e-06 $layer=LI1_cond $X=1.72 $Y=0.74
+ $X2=3.24 $Y2=0.74
r34 10 19 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=4.105 $Y=0.74
+ $X2=4.2 $Y2=0.74
r35 10 15 45.684 $w=2.08e-07 $l=8.65e-07 $layer=LI1_cond $X=4.105 $Y=0.74
+ $X2=3.24 $Y2=0.74
r36 3 17 182 $w=1.7e-07 $l=5.10221e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.2 $Y2=0.68
r37 2 15 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.235 $X2=3.24 $Y2=0.74
r38 1 12 182 $w=1.7e-07 $l=5.70723e-07 $layer=licon1_NDIFF $count=1 $X=1.58
+ $Y=0.235 $X2=1.72 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_2%VGND 1 2 3 12 15 16 17 18 24 36 41 42
r58 41 44 9.44516 $w=4.65e-07 $l=3.6e-07 $layer=LI1_cond $X=4.762 $Y=0 $X2=4.762
+ $Y2=0.36
r59 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r60 39 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r61 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r62 36 41 6.7035 $w=1.7e-07 $l=2.97e-07 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.762
+ $Y2=0
r63 36 38 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.465 $Y=0 $X2=4.37
+ $Y2=0
r64 35 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r65 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r66 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r67 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r68 27 31 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r69 24 32 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r70 24 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r71 20 38 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.905 $Y=0 $X2=4.37
+ $Y2=0
r72 18 34 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.525 $Y=0 $X2=3.45
+ $Y2=0
r73 17 22 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.715
+ $Y2=0.36
r74 17 20 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.905
+ $Y2=0
r75 17 18 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.715 $Y=0 $X2=3.525
+ $Y2=0
r76 15 31 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.53
+ $Y2=0
r77 15 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.595 $Y=0 $X2=2.76
+ $Y2=0
r78 14 34 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.45
+ $Y2=0
r79 14 16 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.76
+ $Y2=0
r80 10 16 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0
r81 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.76 $Y=0.085
+ $X2=2.76 $Y2=0.36
r82 3 44 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=4.545
+ $Y=0.235 $X2=4.705 $Y2=0.36
r83 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.605
+ $Y=0.235 $X2=3.74 $Y2=0.36
r84 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.76 $Y2=0.36
.ends

