* File: sky130_fd_sc_hdll__o2bb2a_1.pxi.spice
* Created: Wed Sep  2 08:45:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_76_199# N_A_76_199#_M1010_s
+ N_A_76_199#_M1011_d N_A_76_199#_c_80_n N_A_76_199#_M1002_g N_A_76_199#_c_81_n
+ N_A_76_199#_M1009_g N_A_76_199#_c_82_n N_A_76_199#_c_89_n N_A_76_199#_c_99_p
+ N_A_76_199#_c_142_p N_A_76_199#_c_83_n N_A_76_199#_c_91_n N_A_76_199#_c_84_n
+ N_A_76_199#_c_85_n N_A_76_199#_c_86_n N_A_76_199#_c_92_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_76_199#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%A1_N N_A1_N_c_181_n N_A1_N_c_182_n
+ N_A1_N_M1006_g N_A1_N_M1001_g A1_N N_A1_N_c_179_n A1_N
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%A2_N N_A2_N_M1004_g N_A2_N_c_223_n
+ N_A2_N_c_230_n N_A2_N_M1000_g N_A2_N_c_224_n N_A2_N_c_225_n N_A2_N_c_226_n
+ A2_N N_A2_N_c_228_n PM_SKY130_FD_SC_HDLL__O2BB2A_1%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_224_369# N_A_224_369#_M1004_d
+ N_A_224_369#_M1006_d N_A_224_369#_c_279_n N_A_224_369#_M1011_g
+ N_A_224_369#_M1010_g N_A_224_369#_c_281_n N_A_224_369#_c_282_n
+ N_A_224_369#_c_283_n N_A_224_369#_c_277_n N_A_224_369#_c_284_n
+ N_A_224_369#_c_278_n PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_224_369#
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%B2 N_B2_M1003_g N_B2_c_349_n N_B2_c_350_n
+ N_B2_M1005_g N_B2_c_347_n N_B2_c_348_n B2 N_B2_c_353_n B2
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%B1 N_B1_M1008_g N_B1_c_397_n N_B1_c_398_n
+ N_B1_M1007_g B1 B1 N_B1_c_396_n PM_SKY130_FD_SC_HDLL__O2BB2A_1%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%X N_X_M1009_s N_X_M1002_s N_X_c_423_n
+ N_X_c_424_n N_X_c_426_n N_X_c_425_n X N_X_c_428_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%X
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%VPWR N_VPWR_M1002_d N_VPWR_M1000_d
+ N_VPWR_M1007_d N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n VPWR
+ N_VPWR_c_448_n N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n
+ N_VPWR_c_444_n PM_SKY130_FD_SC_HDLL__O2BB2A_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%VGND N_VGND_M1009_d N_VGND_M1003_d
+ N_VGND_c_498_n N_VGND_c_499_n N_VGND_c_500_n N_VGND_c_501_n VGND
+ N_VGND_c_502_n N_VGND_c_503_n N_VGND_c_504_n VGND
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_529_47# N_A_529_47#_M1010_d
+ N_A_529_47#_M1008_d N_A_529_47#_c_552_n N_A_529_47#_c_553_n
+ N_A_529_47#_c_554_n N_A_529_47#_c_555_n
+ PM_SKY130_FD_SC_HDLL__O2BB2A_1%A_529_47#
cc_1 VNB N_A_76_199#_c_80_n 0.02825f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_76_199#_c_81_n 0.0204983f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A_76_199#_c_82_n 0.00263372f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_4 VNB N_A_76_199#_c_83_n 5.22012e-19 $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=1.495
cc_5 VNB N_A_76_199#_c_84_n 0.00208406f $X=-0.19 $Y=-0.24 $X2=2.31 $Y2=0.485
cc_6 VNB N_A_76_199#_c_85_n 0.00751946f $X=-0.19 $Y=-0.24 $X2=2.402 $Y2=1.075
cc_7 VNB N_A_76_199#_c_86_n 0.002487f $X=-0.19 $Y=-0.24 $X2=2.402 $Y2=1.245
cc_8 VNB N_A1_N_M1001_g 0.0299214f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_9 VNB N_A1_N_c_179_n 0.0250453f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.445
cc_10 VNB A1_N 0.00852564f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.97
cc_11 VNB N_A2_N_c_223_n 0.0130279f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A2_N_c_224_n 0.00597738f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_13 VNB N_A2_N_c_225_n 0.00126844f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB N_A2_N_c_226_n 0.0369002f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_15 VNB A2_N 7.41212e-19 $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.615
cc_16 VNB N_A2_N_c_228_n 0.0203621f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.97
cc_17 VNB N_A_224_369#_M1010_g 0.0537332f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_18 VNB N_A_224_369#_c_277_n 0.00359901f $X=-0.19 $Y=-0.24 $X2=2.33 $Y2=1.97
cc_19 VNB N_A_224_369#_c_278_n 0.0141663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_M1003_g 0.0301413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B2_c_347_n 0.0088251f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_22 VNB N_B2_c_348_n 0.023929f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.445
cc_23 VNB N_B1_M1008_g 0.0379047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB B1 0.00881129f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_25 VNB N_B1_c_396_n 0.042002f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.615
cc_26 VNB N_X_c_423_n 0.0160045f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_27 VNB N_X_c_424_n 0.00666696f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.445
cc_28 VNB N_X_c_425_n 0.0220799f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_29 VNB N_VPWR_c_444_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_498_n 0.0047376f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_31 VNB N_VGND_c_499_n 0.00574137f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_32 VNB N_VGND_c_500_n 0.0615553f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.615
cc_33 VNB N_VGND_c_501_n 0.0067041f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=1.885
cc_34 VNB N_VGND_c_502_n 0.0190948f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.485
cc_35 VNB N_VGND_c_503_n 0.22578f $X=-0.19 $Y=-0.24 $X2=2.31 $Y2=0.485
cc_36 VNB N_VGND_c_504_n 0.0235541f $X=-0.19 $Y=-0.24 $X2=2.402 $Y2=1.075
cc_37 VNB N_A_529_47#_c_552_n 0.00129968f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_38 VNB N_A_529_47#_c_553_n 0.0196434f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_39 VNB N_A_529_47#_c_554_n 0.00390584f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_40 VNB N_A_529_47#_c_555_n 0.0168304f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_41 VPB N_A_76_199#_c_80_n 0.0313058f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_A_76_199#_c_82_n 0.0014802f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_43 VPB N_A_76_199#_c_89_n 0.00185155f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.885
cc_44 VPB N_A_76_199#_c_83_n 4.42383e-19 $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.495
cc_45 VPB N_A_76_199#_c_91_n 0.00657038f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.53
cc_46 VPB N_A_76_199#_c_92_n 0.0139764f $X=-0.19 $Y=1.305 $X2=2.632 $Y2=1.97
cc_47 VPB N_A1_N_c_181_n 0.0215714f $X=-0.19 $Y=1.305 $X2=2.635 $Y2=1.845
cc_48 VPB N_A1_N_c_182_n 0.024986f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A1_N_c_179_n 0.00447281f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.445
cc_50 VPB N_A2_N_c_223_n 0.0203767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A2_N_c_230_n 0.0263053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_224_369#_c_279_n 0.0177168f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_53 VPB N_A_224_369#_M1010_g 0.00309964f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_54 VPB N_A_224_369#_c_281_n 0.0508903f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_55 VPB N_A_224_369#_c_282_n 0.0200887f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_56 VPB N_A_224_369#_c_283_n 0.00878984f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_57 VPB N_A_224_369#_c_284_n 0.00849787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_224_369#_c_278_n 8.66278e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B2_c_349_n 0.0220397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_B2_c_350_n 0.0253638f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_61 VPB N_B2_c_347_n 0.00734023f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_62 VPB N_B2_c_348_n 0.00520446f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.445
cc_63 VPB N_B2_c_353_n 0.0175474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_B1_c_397_n 0.0251152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_B1_c_398_n 0.0300241f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_66 VPB B1 0.0163181f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_67 VPB N_B1_c_396_n 0.0103535f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.615
cc_68 VPB N_X_c_426_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_69 VPB N_X_c_425_n 0.0195719f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_70 VPB N_X_c_428_n 0.0208429f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=1.885
cc_71 VPB N_VPWR_c_445_n 0.0077704f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_72 VPB N_VPWR_c_446_n 0.0116186f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_73 VPB N_VPWR_c_447_n 0.0368842f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_74 VPB N_VPWR_c_448_n 0.0150576f $X=-0.19 $Y=1.305 $X2=2.33 $Y2=1.97
cc_75 VPB N_VPWR_c_449_n 0.0267798f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.495
cc_76 VPB N_VPWR_c_450_n 0.0402951f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=0.485
cc_77 VPB N_VPWR_c_451_n 0.005797f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_78 VPB N_VPWR_c_452_n 0.0153178f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_444_n 0.0785117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 N_A_76_199#_c_80_n N_A1_N_c_181_n 0.0132797f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_76_199#_c_82_n N_A1_N_c_181_n 0.00237013f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A_76_199#_c_89_n N_A1_N_c_181_n 0.00220402f $X=0.79 $Y=1.885 $X2=0 $Y2=0
cc_83 N_A_76_199#_c_91_n N_A1_N_c_181_n 0.00254159f $X=0.79 $Y=1.53 $X2=0 $Y2=0
cc_84 N_A_76_199#_c_80_n N_A1_N_c_182_n 0.0144107f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_76_199#_c_89_n N_A1_N_c_182_n 0.00281836f $X=0.79 $Y=1.885 $X2=0 $Y2=0
cc_86 N_A_76_199#_c_99_p N_A1_N_c_182_n 0.0151259f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_87 N_A_76_199#_c_81_n N_A1_N_M1001_g 0.0200796f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_76_199#_c_80_n N_A1_N_c_179_n 0.0212212f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_76_199#_c_82_n N_A1_N_c_179_n 0.00102926f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_76_199#_c_80_n A1_N 0.00128482f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_76_199#_c_82_n A1_N 0.0158298f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_76_199#_c_99_p A1_N 0.00351608f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_93 N_A_76_199#_c_91_n A1_N 0.00419335f $X=0.79 $Y=1.53 $X2=0 $Y2=0
cc_94 N_A_76_199#_c_99_p N_A2_N_c_230_n 0.0159089f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_95 N_A_76_199#_c_92_n N_A2_N_c_230_n 0.00399922f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_96 N_A_76_199#_c_81_n N_A2_N_c_225_n 7.04993e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_76_199#_c_99_p N_A_224_369#_M1006_d 0.00927633f $X=2.33 $Y=1.97 $X2=0
+ $Y2=0
cc_98 N_A_76_199#_c_92_n N_A_224_369#_c_279_n 0.0252753f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_99 N_A_76_199#_c_83_n N_A_224_369#_M1010_g 0.00314477f $X=2.415 $Y=1.495
+ $X2=0 $Y2=0
cc_100 N_A_76_199#_c_84_n N_A_224_369#_M1010_g 0.00961943f $X=2.31 $Y=0.485
+ $X2=0 $Y2=0
cc_101 N_A_76_199#_c_86_n N_A_224_369#_M1010_g 0.00466522f $X=2.402 $Y=1.245
+ $X2=0 $Y2=0
cc_102 N_A_76_199#_c_99_p N_A_224_369#_c_281_n 0.00738394f $X=2.33 $Y=1.97 $X2=0
+ $Y2=0
cc_103 N_A_76_199#_c_83_n N_A_224_369#_c_281_n 0.00610077f $X=2.415 $Y=1.495
+ $X2=0 $Y2=0
cc_104 N_A_76_199#_c_84_n N_A_224_369#_c_281_n 0.00194568f $X=2.31 $Y=0.485
+ $X2=0 $Y2=0
cc_105 N_A_76_199#_c_86_n N_A_224_369#_c_281_n 7.75851e-19 $X=2.402 $Y=1.245
+ $X2=0 $Y2=0
cc_106 N_A_76_199#_c_92_n N_A_224_369#_c_281_n 0.0070843f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_107 N_A_76_199#_c_83_n N_A_224_369#_c_282_n 0.00407164f $X=2.415 $Y=1.495
+ $X2=0 $Y2=0
cc_108 N_A_76_199#_c_92_n N_A_224_369#_c_282_n 0.017313f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_109 N_A_76_199#_c_89_n N_A_224_369#_c_283_n 0.00786855f $X=0.79 $Y=1.885
+ $X2=0 $Y2=0
cc_110 N_A_76_199#_c_99_p N_A_224_369#_c_283_n 0.0551054f $X=2.33 $Y=1.97 $X2=0
+ $Y2=0
cc_111 N_A_76_199#_c_91_n N_A_224_369#_c_283_n 0.0101776f $X=0.79 $Y=1.53 $X2=0
+ $Y2=0
cc_112 N_A_76_199#_c_84_n N_A_224_369#_c_277_n 0.0141351f $X=2.31 $Y=0.485 $X2=0
+ $Y2=0
cc_113 N_A_76_199#_c_99_p N_A_224_369#_c_284_n 0.0222516f $X=2.33 $Y=1.97 $X2=0
+ $Y2=0
cc_114 N_A_76_199#_c_83_n N_A_224_369#_c_284_n 0.00981918f $X=2.415 $Y=1.495
+ $X2=0 $Y2=0
cc_115 N_A_76_199#_c_92_n N_A_224_369#_c_284_n 0.0174234f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_116 N_A_76_199#_c_83_n N_A_224_369#_c_278_n 0.00587569f $X=2.415 $Y=1.495
+ $X2=0 $Y2=0
cc_117 N_A_76_199#_c_84_n N_A_224_369#_c_278_n 0.0095286f $X=2.31 $Y=0.485 $X2=0
+ $Y2=0
cc_118 N_A_76_199#_c_85_n N_A_224_369#_c_278_n 0.0319889f $X=2.402 $Y=1.075
+ $X2=0 $Y2=0
cc_119 N_A_76_199#_c_83_n N_B2_c_349_n 8.08053e-19 $X=2.415 $Y=1.495 $X2=0 $Y2=0
cc_120 N_A_76_199#_c_92_n N_B2_c_349_n 0.00370502f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_121 N_A_76_199#_c_92_n N_B2_c_350_n 0.0014571f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_122 N_A_76_199#_c_86_n N_B2_c_347_n 0.0165753f $X=2.402 $Y=1.245 $X2=0 $Y2=0
cc_123 N_A_76_199#_c_92_n N_B2_c_347_n 0.018331f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_124 N_A_76_199#_c_86_n N_B2_c_348_n 2.00411e-19 $X=2.402 $Y=1.245 $X2=0 $Y2=0
cc_125 N_A_76_199#_c_92_n N_B2_c_348_n 0.00186365f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_126 N_A_76_199#_c_92_n N_B2_c_353_n 0.0256721f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_127 N_A_76_199#_c_80_n N_X_c_424_n 0.00116024f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_76_199#_c_89_n N_X_c_426_n 0.00386336f $X=0.79 $Y=1.885 $X2=0 $Y2=0
cc_129 N_A_76_199#_c_142_p N_X_c_426_n 0.00815002f $X=0.875 $Y=1.97 $X2=0 $Y2=0
cc_130 N_A_76_199#_c_80_n N_X_c_425_n 0.0174815f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_76_199#_c_81_n N_X_c_425_n 0.0047149f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_76_199#_c_82_n N_X_c_425_n 0.0328403f $X=0.515 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_76_199#_c_89_n N_X_c_425_n 0.00640837f $X=0.79 $Y=1.885 $X2=0 $Y2=0
cc_134 N_A_76_199#_c_91_n N_X_c_425_n 0.0128407f $X=0.79 $Y=1.53 $X2=0 $Y2=0
cc_135 N_A_76_199#_c_89_n N_VPWR_M1002_d 0.00480398f $X=0.79 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_76_199#_c_99_p N_VPWR_M1002_d 2.1423e-19 $X=2.33 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_137 N_A_76_199#_c_142_p N_VPWR_M1002_d 0.00432679f $X=0.875 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_76_199#_c_91_n N_VPWR_M1002_d 0.00226067f $X=0.79 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_139 N_A_76_199#_c_99_p N_VPWR_M1000_d 0.0160105f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_140 N_A_76_199#_c_92_n N_VPWR_M1000_d 0.00207403f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_141 N_A_76_199#_c_80_n N_VPWR_c_445_n 0.013365f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_76_199#_c_99_p N_VPWR_c_445_n 5.54398e-19 $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_143 N_A_76_199#_c_142_p N_VPWR_c_445_n 0.0132919f $X=0.875 $Y=1.97 $X2=0
+ $Y2=0
cc_144 N_A_76_199#_c_91_n N_VPWR_c_445_n 0.00369081f $X=0.79 $Y=1.53 $X2=0 $Y2=0
cc_145 N_A_76_199#_c_80_n N_VPWR_c_448_n 0.00427505f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_76_199#_c_99_p N_VPWR_c_449_n 0.0139061f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_147 N_A_76_199#_c_99_p N_VPWR_c_450_n 0.00105858f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_148 N_A_76_199#_c_92_n N_VPWR_c_450_n 0.0160361f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_149 N_A_76_199#_c_99_p N_VPWR_c_452_n 0.0291396f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_150 N_A_76_199#_c_92_n N_VPWR_c_452_n 0.00291694f $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_151 N_A_76_199#_c_80_n N_VPWR_c_444_n 0.0082412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_76_199#_c_99_p N_VPWR_c_444_n 0.0301679f $X=2.33 $Y=1.97 $X2=0 $Y2=0
cc_153 N_A_76_199#_c_142_p N_VPWR_c_444_n 7.98136e-19 $X=0.875 $Y=1.97 $X2=0
+ $Y2=0
cc_154 N_A_76_199#_c_92_n N_VPWR_c_444_n 0.0196265f $X=2.632 $Y=1.97 $X2=0 $Y2=0
cc_155 N_A_76_199#_c_80_n N_VGND_c_498_n 0.00118907f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_76_199#_c_81_n N_VGND_c_498_n 0.00553486f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_76_199#_c_84_n N_VGND_c_500_n 0.0112593f $X=2.31 $Y=0.485 $X2=0 $Y2=0
cc_158 N_A_76_199#_M1010_s N_VGND_c_503_n 0.0047105f $X=2.185 $Y=0.235 $X2=0
+ $Y2=0
cc_159 N_A_76_199#_c_81_n N_VGND_c_503_n 0.0119587f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_76_199#_c_84_n N_VGND_c_503_n 0.00918075f $X=2.31 $Y=0.485 $X2=0
+ $Y2=0
cc_161 N_A_76_199#_c_81_n N_VGND_c_504_n 0.00585385f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_76_199#_c_84_n N_A_529_47#_c_552_n 0.00446296f $X=2.31 $Y=0.485 $X2=0
+ $Y2=0
cc_163 N_A_76_199#_c_85_n N_A_529_47#_c_554_n 0.0126647f $X=2.402 $Y=1.075 $X2=0
+ $Y2=0
cc_164 N_A_76_199#_c_92_n N_A_529_47#_c_554_n 9.70378e-19 $X=2.632 $Y=1.97 $X2=0
+ $Y2=0
cc_165 N_A1_N_c_181_n N_A2_N_c_223_n 0.0071273f $X=1.03 $Y=1.67 $X2=0 $Y2=0
cc_166 N_A1_N_c_179_n N_A2_N_c_223_n 0.00907223f $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_167 A1_N N_A2_N_c_223_n 0.0019023f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_168 N_A1_N_c_182_n N_A2_N_c_230_n 0.0267183f $X=1.03 $Y=1.77 $X2=0 $Y2=0
cc_169 N_A1_N_M1001_g N_A2_N_c_224_n 5.97299e-19 $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_170 N_A1_N_c_179_n N_A2_N_c_224_n 5.37172e-19 $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_171 A1_N N_A2_N_c_224_n 0.0034089f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_172 N_A1_N_M1001_g N_A2_N_c_225_n 0.00796716f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_173 N_A1_N_c_179_n N_A2_N_c_225_n 0.00269131f $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_174 A1_N N_A2_N_c_225_n 0.0225271f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_175 N_A1_N_c_179_n N_A2_N_c_226_n 0.00701716f $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_176 N_A1_N_M1001_g A2_N 0.0103229f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_177 N_A1_N_M1001_g N_A2_N_c_228_n 0.0344453f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_178 N_A1_N_c_181_n N_A_224_369#_c_283_n 0.00671979f $X=1.03 $Y=1.67 $X2=0
+ $Y2=0
cc_179 N_A1_N_c_182_n N_A_224_369#_c_283_n 0.0024725f $X=1.03 $Y=1.77 $X2=0
+ $Y2=0
cc_180 N_A1_N_c_179_n N_A_224_369#_c_283_n 0.00231747f $X=1.045 $Y=1.16 $X2=0
+ $Y2=0
cc_181 A1_N N_A_224_369#_c_283_n 0.0166076f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_182 A1_N N_A_224_369#_c_278_n 0.00614761f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_183 N_A1_N_c_182_n N_VPWR_c_445_n 0.00396483f $X=1.03 $Y=1.77 $X2=0 $Y2=0
cc_184 N_A1_N_c_182_n N_VPWR_c_449_n 0.00479146f $X=1.03 $Y=1.77 $X2=0 $Y2=0
cc_185 N_A1_N_c_182_n N_VPWR_c_444_n 0.00619141f $X=1.03 $Y=1.77 $X2=0 $Y2=0
cc_186 N_A1_N_M1001_g N_VGND_c_498_n 0.00827125f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_187 A1_N N_VGND_c_498_n 9.9771e-19 $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_188 N_A1_N_M1001_g N_VGND_c_500_n 0.00437915f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A1_N_M1001_g N_VGND_c_503_n 0.00727435f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A2_N_c_226_n N_A_224_369#_M1010_g 0.00277126f $X=1.575 $Y=0.935 $X2=0
+ $Y2=0
cc_191 N_A2_N_c_223_n N_A_224_369#_c_281_n 0.020771f $X=1.63 $Y=1.67 $X2=0 $Y2=0
cc_192 N_A2_N_c_230_n N_A_224_369#_c_282_n 8.59035e-19 $X=1.63 $Y=1.77 $X2=0
+ $Y2=0
cc_193 N_A2_N_c_223_n N_A_224_369#_c_283_n 0.0116706f $X=1.63 $Y=1.67 $X2=0
+ $Y2=0
cc_194 N_A2_N_c_230_n N_A_224_369#_c_283_n 0.00462887f $X=1.63 $Y=1.77 $X2=0
+ $Y2=0
cc_195 N_A2_N_c_224_n N_A_224_369#_c_283_n 0.0135699f $X=1.49 $Y=0.82 $X2=0
+ $Y2=0
cc_196 N_A2_N_c_226_n N_A_224_369#_c_283_n 0.00297086f $X=1.575 $Y=0.935 $X2=0
+ $Y2=0
cc_197 N_A2_N_c_224_n N_A_224_369#_c_277_n 0.00939206f $X=1.49 $Y=0.82 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_226_n N_A_224_369#_c_277_n 0.00311395f $X=1.575 $Y=0.935 $X2=0
+ $Y2=0
cc_199 A2_N N_A_224_369#_c_277_n 0.00962703f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_200 N_A2_N_c_228_n N_A_224_369#_c_277_n 0.00294085f $X=1.61 $Y=0.77 $X2=0
+ $Y2=0
cc_201 N_A2_N_c_223_n N_A_224_369#_c_284_n 2.19802e-19 $X=1.63 $Y=1.67 $X2=0
+ $Y2=0
cc_202 N_A2_N_c_223_n N_A_224_369#_c_278_n 0.0103574f $X=1.63 $Y=1.67 $X2=0
+ $Y2=0
cc_203 N_A2_N_c_224_n N_A_224_369#_c_278_n 0.0267861f $X=1.49 $Y=0.82 $X2=0
+ $Y2=0
cc_204 N_A2_N_c_226_n N_A_224_369#_c_278_n 0.00408182f $X=1.575 $Y=0.935 $X2=0
+ $Y2=0
cc_205 A2_N N_A_224_369#_c_278_n 0.00529005f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_206 N_A2_N_c_228_n N_A_224_369#_c_278_n 0.0022268f $X=1.61 $Y=0.77 $X2=0
+ $Y2=0
cc_207 N_A2_N_c_230_n N_VPWR_c_449_n 0.00479146f $X=1.63 $Y=1.77 $X2=0 $Y2=0
cc_208 N_A2_N_c_230_n N_VPWR_c_452_n 0.00636594f $X=1.63 $Y=1.77 $X2=0 $Y2=0
cc_209 N_A2_N_c_230_n N_VPWR_c_444_n 0.00619141f $X=1.63 $Y=1.77 $X2=0 $Y2=0
cc_210 N_A2_N_c_225_n N_VGND_c_498_n 0.00112201f $X=1.3 $Y=0.82 $X2=0 $Y2=0
cc_211 A2_N N_VGND_c_498_n 0.0253059f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_212 N_A2_N_c_224_n N_VGND_c_500_n 0.0036955f $X=1.49 $Y=0.82 $X2=0 $Y2=0
cc_213 A2_N N_VGND_c_500_n 0.00958867f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_214 N_A2_N_c_228_n N_VGND_c_500_n 0.0042936f $X=1.61 $Y=0.77 $X2=0 $Y2=0
cc_215 N_A2_N_c_224_n N_VGND_c_503_n 0.00653356f $X=1.49 $Y=0.82 $X2=0 $Y2=0
cc_216 A2_N N_VGND_c_503_n 0.00954404f $X=1.07 $Y=0.425 $X2=0 $Y2=0
cc_217 N_A2_N_c_228_n N_VGND_c_503_n 0.00747565f $X=1.61 $Y=0.77 $X2=0 $Y2=0
cc_218 A2_N A_225_47# 0.00459468f $X=1.07 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_219 N_A_224_369#_M1010_g N_B2_M1003_g 0.0194674f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_220 N_A_224_369#_M1010_g N_B2_c_349_n 0.0078775f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_221 N_A_224_369#_c_279_n N_B2_c_350_n 0.00831609f $X=2.545 $Y=1.77 $X2=0
+ $Y2=0
cc_222 N_A_224_369#_c_282_n N_B2_c_350_n 0.0078775f $X=2.545 $Y=1.562 $X2=0
+ $Y2=0
cc_223 N_A_224_369#_M1010_g N_B2_c_347_n 0.00193645f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_224_369#_M1010_g N_B2_c_348_n 0.0198675f $X=2.57 $Y=0.445 $X2=0 $Y2=0
cc_225 N_A_224_369#_c_279_n N_VPWR_c_450_n 0.0046716f $X=2.545 $Y=1.77 $X2=0
+ $Y2=0
cc_226 N_A_224_369#_c_279_n N_VPWR_c_452_n 0.00515589f $X=2.545 $Y=1.77 $X2=0
+ $Y2=0
cc_227 N_A_224_369#_c_279_n N_VPWR_c_444_n 0.00619141f $X=2.545 $Y=1.77 $X2=0
+ $Y2=0
cc_228 N_A_224_369#_M1010_g N_VGND_c_500_n 0.00585385f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_229 N_A_224_369#_c_277_n N_VGND_c_500_n 0.0164014f $X=1.885 $Y=0.48 $X2=0
+ $Y2=0
cc_230 N_A_224_369#_M1004_d N_VGND_c_503_n 0.00273077f $X=1.59 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_A_224_369#_M1010_g N_VGND_c_503_n 0.0123397f $X=2.57 $Y=0.445 $X2=0
+ $Y2=0
cc_232 N_A_224_369#_c_277_n N_VGND_c_503_n 0.0169233f $X=1.885 $Y=0.48 $X2=0
+ $Y2=0
cc_233 N_A_224_369#_M1010_g N_A_529_47#_c_552_n 5.98067e-19 $X=2.57 $Y=0.445
+ $X2=0 $Y2=0
cc_234 N_A_224_369#_M1010_g N_A_529_47#_c_554_n 0.00174989f $X=2.57 $Y=0.445
+ $X2=0 $Y2=0
cc_235 N_B2_M1003_g N_B1_M1008_g 0.0216135f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_236 N_B2_c_349_n N_B1_c_397_n 0.00729364f $X=3.075 $Y=1.67 $X2=0 $Y2=0
cc_237 N_B2_c_353_n N_B1_c_397_n 0.00647259f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_238 N_B2_c_350_n N_B1_c_398_n 0.0212288f $X=3.075 $Y=1.77 $X2=0 $Y2=0
cc_239 N_B2_c_353_n N_B1_c_398_n 0.00535582f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_240 N_B2_c_347_n B1 0.021165f $X=3.335 $Y=1.2 $X2=0 $Y2=0
cc_241 N_B2_c_348_n B1 2.23297e-19 $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_242 N_B2_c_353_n B1 0.0243797f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_243 N_B2_c_347_n N_B1_c_396_n 0.00299034f $X=3.335 $Y=1.2 $X2=0 $Y2=0
cc_244 N_B2_c_348_n N_B1_c_396_n 0.00729364f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B2_c_353_n N_VPWR_c_447_n 0.0304709f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_246 N_B2_c_350_n N_VPWR_c_450_n 0.00620597f $X=3.075 $Y=1.77 $X2=0 $Y2=0
cc_247 N_B2_c_353_n N_VPWR_c_450_n 0.0113264f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_248 N_B2_c_350_n N_VPWR_c_444_n 0.00619141f $X=3.075 $Y=1.77 $X2=0 $Y2=0
cc_249 N_B2_c_353_n N_VPWR_c_444_n 0.00747463f $X=3.435 $Y=1.325 $X2=0 $Y2=0
cc_250 N_B2_c_353_n A_633_369# 0.00880371f $X=3.435 $Y=1.325 $X2=-0.19 $Y2=-0.24
cc_251 N_B2_M1003_g N_VGND_c_499_n 0.0053916f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_252 N_B2_M1003_g N_VGND_c_500_n 0.00437852f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_253 N_B2_M1003_g N_VGND_c_503_n 0.00643597f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_254 N_B2_M1003_g N_A_529_47#_c_552_n 0.0018743f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_255 N_B2_M1003_g N_A_529_47#_c_553_n 0.0131548f $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_256 N_B2_c_347_n N_A_529_47#_c_553_n 0.0457798f $X=3.335 $Y=1.2 $X2=0 $Y2=0
cc_257 N_B2_c_348_n N_A_529_47#_c_553_n 0.00222979f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B2_c_347_n N_A_529_47#_c_554_n 0.0189241f $X=3.335 $Y=1.2 $X2=0 $Y2=0
cc_259 N_B2_c_348_n N_A_529_47#_c_554_n 0.00229607f $X=2.99 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B2_M1003_g N_A_529_47#_c_555_n 8.23015e-19 $X=3.04 $Y=0.445 $X2=0 $Y2=0
cc_261 N_B1_c_398_n N_VPWR_c_447_n 0.011855f $X=3.645 $Y=1.77 $X2=0 $Y2=0
cc_262 B1 N_VPWR_c_447_n 0.0318759f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_263 N_B1_c_396_n N_VPWR_c_447_n 0.00115968f $X=3.875 $Y=1.16 $X2=0 $Y2=0
cc_264 N_B1_c_398_n N_VPWR_c_450_n 0.00515958f $X=3.645 $Y=1.77 $X2=0 $Y2=0
cc_265 N_B1_c_398_n N_VPWR_c_444_n 0.00519391f $X=3.645 $Y=1.77 $X2=0 $Y2=0
cc_266 N_B1_M1008_g N_VGND_c_499_n 0.00768374f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_267 N_B1_M1008_g N_VGND_c_502_n 0.00425893f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_268 N_B1_M1008_g N_VGND_c_503_n 0.00724352f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_269 N_B1_M1008_g N_A_529_47#_c_553_n 0.0189313f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_270 B1 N_A_529_47#_c_553_n 0.0303523f $X=3.825 $Y=1.105 $X2=0 $Y2=0
cc_271 N_B1_c_396_n N_A_529_47#_c_553_n 0.00912169f $X=3.875 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B1_M1008_g N_A_529_47#_c_555_n 0.00845291f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_273 N_X_c_428_n N_VPWR_c_445_n 0.0177194f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_274 N_X_c_428_n N_VPWR_c_448_n 0.0182037f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_275 N_X_M1002_s N_VPWR_c_444_n 0.00425811f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_276 N_X_c_428_n N_VPWR_c_444_n 0.00993477f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_277 N_X_M1009_s N_VGND_c_503_n 0.0031974f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_278 N_X_c_423_n N_VGND_c_503_n 0.0129881f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_279 N_X_c_423_n N_VGND_c_504_n 0.0224663f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_280 N_VGND_c_503_n A_225_47# 0.00333848f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_281 N_VGND_c_503_n N_A_529_47#_M1010_d 0.00447847f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_282 N_VGND_c_503_n N_A_529_47#_M1008_d 0.00256165f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_283 N_VGND_c_500_n N_A_529_47#_c_552_n 0.0111709f $X=3.135 $Y=0 $X2=0 $Y2=0
cc_284 N_VGND_c_503_n N_A_529_47#_c_552_n 0.00919097f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_285 N_VGND_c_499_n N_A_529_47#_c_553_n 0.0261732f $X=3.315 $Y=0.39 $X2=0
+ $Y2=0
cc_286 N_VGND_c_500_n N_A_529_47#_c_553_n 0.00261274f $X=3.135 $Y=0 $X2=0 $Y2=0
cc_287 N_VGND_c_502_n N_A_529_47#_c_553_n 0.00251757f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_288 N_VGND_c_503_n N_A_529_47#_c_553_n 0.00980822f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_289 N_VGND_c_499_n N_A_529_47#_c_555_n 0.0177522f $X=3.315 $Y=0.39 $X2=0
+ $Y2=0
cc_290 N_VGND_c_502_n N_A_529_47#_c_555_n 0.0176634f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_291 N_VGND_c_503_n N_A_529_47#_c_555_n 0.0141724f $X=3.91 $Y=0 $X2=0 $Y2=0
