* File: sky130_fd_sc_hdll__nand4b_2.spice
* Created: Wed Sep  2 08:38:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4b_2.pex.spice"
.subckt sky130_fd_sc_hdll__nand4b_2  VNB VPB A_N B C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_A_N_M1011_g N_A_27_47#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_A_225_47#_M1004_d N_A_27_47#_M1004_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1014 N_A_225_47#_M1014_d N_A_27_47#_M1014_g N_Y_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1008 N_A_225_47#_M1014_d N_B_M1008_g N_A_495_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_A_225_47#_M1010_d N_B_M1010_g N_A_495_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_A_705_47#_M1005_d N_C_M1005_g N_A_495_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1015 N_A_705_47#_M1015_d N_C_M1015_g N_A_495_47#_M1005_s VNB NSHORT L=0.15
+ W=0.65 AD=0.13325 AS=0.104 PD=1.06 PS=0.97 NRD=7.38 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_705_47#_M1015_d N_D_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13325 AS=0.104 PD=1.06 PS=0.97 NRD=16.608 NRS=0 M=1 R=4.33333 SA=75001.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_705_47#_M1007_d N_D_M1007_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_47#_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_47#_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_27_47#_M1016_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1016_d N_B_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90003.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.38
+ AS=0.145 PD=1.76 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1006_d N_C_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.38
+ AS=0.145 PD=1.76 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90001.8 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_C_M1017_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.19
+ AS=0.145 PD=1.38 PS=1.29 NRD=7.8603 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1017_d N_D_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.19
+ AS=0.145 PD=1.38 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90003.6
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_D_M1013_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.41
+ AS=0.145 PD=2.82 PS=1.29 NRD=16.7253 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX18_noxref VNB VPB NWDIODE A=10.2078 P=15.93
*
.include "sky130_fd_sc_hdll__nand4b_2.pxi.spice"
*
.ends
*
*
