* File: sky130_fd_sc_hdll__nand3_2.pxi.spice
* Created: Thu Aug 27 19:13:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3_2%A N_A_c_56_n N_A_M1000_g N_A_c_52_n N_A_M1001_g
+ N_A_c_57_n N_A_M1005_g N_A_c_53_n N_A_M1008_g A N_A_c_55_n
+ PM_SKY130_FD_SC_HDLL__NAND3_2%A
x_PM_SKY130_FD_SC_HDLL__NAND3_2%B N_B_c_100_n N_B_M1007_g N_B_M1009_g
+ N_B_c_101_n N_B_M1010_g N_B_M1011_g B B B N_B_c_98_n B B B
+ PM_SKY130_FD_SC_HDLL__NAND3_2%B
x_PM_SKY130_FD_SC_HDLL__NAND3_2%C N_C_M1004_g N_C_c_149_n N_C_M1002_g
+ N_C_c_146_n N_C_M1006_g N_C_c_150_n N_C_M1003_g C C C N_C_c_148_n C C
+ PM_SKY130_FD_SC_HDLL__NAND3_2%C
x_PM_SKY130_FD_SC_HDLL__NAND3_2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d
+ N_VPWR_M1010_d N_VPWR_M1002_d N_VPWR_M1003_d N_VPWR_c_187_n N_VPWR_c_188_n
+ N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n N_VPWR_c_192_n N_VPWR_c_193_n
+ N_VPWR_c_194_n VPWR N_VPWR_c_195_n N_VPWR_c_196_n N_VPWR_c_197_n
+ N_VPWR_c_186_n PM_SKY130_FD_SC_HDLL__NAND3_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3_2%Y N_Y_M1001_s N_Y_M1000_s N_Y_M1007_s
+ N_Y_M1002_s N_Y_c_248_n N_Y_c_244_n N_Y_c_252_n N_Y_c_245_n N_Y_c_246_n
+ N_Y_c_283_n N_Y_c_247_n Y Y Y N_Y_c_243_n PM_SKY130_FD_SC_HDLL__NAND3_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND3_2%A_27_47# N_A_27_47#_M1001_d N_A_27_47#_M1008_d
+ N_A_27_47#_M1011_d N_A_27_47#_c_313_n N_A_27_47#_c_314_n N_A_27_47#_c_315_n
+ PM_SKY130_FD_SC_HDLL__NAND3_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND3_2%A_307_47# N_A_307_47#_M1009_s
+ N_A_307_47#_M1004_s N_A_307_47#_c_340_n
+ PM_SKY130_FD_SC_HDLL__NAND3_2%A_307_47#
x_PM_SKY130_FD_SC_HDLL__NAND3_2%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_c_363_n N_VGND_c_364_n N_VGND_c_365_n VGND N_VGND_c_366_n
+ N_VGND_c_367_n N_VGND_c_368_n N_VGND_c_369_n
+ PM_SKY130_FD_SC_HDLL__NAND3_2%VGND
cc_1 VNB N_A_c_52_n 0.0219834f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_c_53_n 0.0171408f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB A 0.0134856f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_c_55_n 0.059491f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_B_M1009_g 0.0181911f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_6 VNB N_B_M1011_g 0.023617f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_7 VNB N_B_c_98_n 0.0498353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB B 0.0150192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_C_M1004_g 0.0225343f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_10 VNB N_C_c_146_n 0.0235983f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_11 VNB C 0.0231427f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_12 VNB N_C_c_148_n 0.0562975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_186_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_243_n 0.00106845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_313_n 0.0123949f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_16 VNB N_A_27_47#_c_314_n 0.00754845f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB N_A_27_47#_c_315_n 0.00218948f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_18 VNB N_A_307_47#_c_340_n 0.0185818f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_19 VNB N_VGND_c_363_n 0.00560444f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_20 VNB N_VGND_c_364_n 0.0173253f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_21 VNB N_VGND_c_365_n 0.0365407f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_22 VNB N_VGND_c_366_n 0.0614619f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_23 VNB N_VGND_c_367_n 0.018763f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_368_n 0.00507168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_369_n 0.22719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_c_56_n 0.0207437f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_27 VPB N_A_c_57_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_28 VPB A 0.00291996f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_29 VPB N_A_c_55_n 0.032798f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_30 VPB N_B_c_100_n 0.0159796f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_31 VPB N_B_c_101_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_32 VPB N_B_c_98_n 0.0283568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_C_c_149_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_34 VPB N_C_c_150_n 0.0198539f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_35 VPB N_C_c_148_n 0.0319527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_187_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_37 VPB N_VPWR_c_188_n 0.0427361f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_38 VPB N_VPWR_c_189_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_190_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_191_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_192_n 0.0166326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_193_n 0.0172994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_194_n 0.0534625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_195_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_196_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_197_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_186_n 0.0491407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_Y_c_244_n 0.00520112f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_49 VPB N_Y_c_245_n 0.0126876f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_246_n 0.00175503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_Y_c_247_n 0.00175503f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_A_c_57_n N_B_c_100_n 0.0229911f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_53 N_A_c_53_n N_B_M1009_g 0.0221472f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_c_55_n N_B_c_98_n 0.025615f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_55 N_A_c_55_n B 0.00189651f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_56 N_A_c_56_n N_VPWR_c_188_n 0.00777002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 A N_VPWR_c_188_n 0.0199082f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_55_n N_VPWR_c_188_n 0.00239995f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_59 N_A_c_56_n N_VPWR_c_189_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_57_n N_VPWR_c_189_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_57_n N_VPWR_c_190_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_c_56_n N_VPWR_c_186_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A_c_57_n N_VPWR_c_186_n 0.011869f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_56_n N_Y_c_248_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_Y_c_248_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_57_n N_Y_c_244_n 0.020382f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_c_55_n N_Y_c_244_n 4.93319e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_68 N_A_c_57_n N_Y_c_252_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_56_n Y 0.00551099f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_c_57_n Y 8.77306e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_c_56_n N_Y_c_243_n 0.00199531f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_52_n N_Y_c_243_n 0.0146242f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_57_n N_Y_c_243_n 0.00103355f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_53_n N_Y_c_243_n 0.00296985f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_75 A N_Y_c_243_n 0.0228434f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_55_n N_Y_c_243_n 0.0390452f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_77 N_A_c_52_n N_A_27_47#_c_313_n 0.00534663f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_313_n 0.016487f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_55_n N_A_27_47#_c_313_n 0.00223477f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_80 N_A_c_52_n N_A_27_47#_c_315_n 0.010732f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_53_n N_A_27_47#_c_315_n 0.0127383f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_55_n N_A_27_47#_c_315_n 0.00246449f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_83 N_A_c_53_n N_A_307_47#_c_340_n 8.96673e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A_c_52_n N_VGND_c_366_n 0.00366111f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_c_53_n N_VGND_c_366_n 0.00366111f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_c_52_n N_VGND_c_369_n 0.00644821f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_c_53_n N_VGND_c_369_n 0.00551736f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B_c_98_n C 3.83125e-19 $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_89 B C 0.0185484f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_90 N_B_c_98_n N_C_c_148_n 0.00552895f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_91 B N_C_c_148_n 9.3524e-19 $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_92 N_B_c_100_n N_VPWR_c_190_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_100_n N_VPWR_c_191_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_101_n N_VPWR_c_191_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_101_n N_VPWR_c_192_n 0.00825342f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_100_n N_VPWR_c_186_n 0.0100198f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_101_n N_VPWR_c_186_n 0.0131262f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B_c_100_n N_Y_c_248_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_100_n N_Y_c_244_n 0.0113403f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_98_n N_Y_c_244_n 0.00164063f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_101 B N_Y_c_244_n 0.0210009f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_102 N_B_c_100_n N_Y_c_252_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B_c_101_n N_Y_c_252_n 0.0153658f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_101_n N_Y_c_245_n 0.0179883f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B_c_98_n N_Y_c_245_n 0.00440776f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_106 B N_Y_c_245_n 0.0586349f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_107 N_B_c_100_n N_Y_c_247_n 0.00292783f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B_c_101_n N_Y_c_247_n 0.00116723f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B_c_98_n N_Y_c_247_n 0.00760751f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_110 B N_Y_c_247_n 0.0305804f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_111 N_B_c_98_n N_Y_c_243_n 0.00113945f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_112 B N_Y_c_243_n 0.0117738f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_113 N_B_M1009_g N_A_27_47#_c_315_n 0.00914262f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_114 N_B_M1011_g N_A_27_47#_c_315_n 0.00818766f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_115 N_B_c_98_n N_A_27_47#_c_315_n 0.00176769f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_116 B N_A_27_47#_c_315_n 0.00685365f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_117 N_B_M1009_g N_A_307_47#_c_340_n 0.0083047f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_118 N_B_M1011_g N_A_307_47#_c_340_n 0.0146104f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_119 N_B_c_98_n N_A_307_47#_c_340_n 0.00758944f $X=1.93 $Y=1.212 $X2=0 $Y2=0
cc_120 B N_A_307_47#_c_340_n 0.0878841f $X=2.505 $Y=1.19 $X2=0 $Y2=0
cc_121 N_B_M1011_g N_VGND_c_363_n 0.00294182f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_122 N_B_M1009_g N_VGND_c_366_n 0.00366111f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_123 N_B_M1011_g N_VGND_c_366_n 0.00366111f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_124 N_B_M1009_g N_VGND_c_369_n 0.00551736f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_125 N_B_M1011_g N_VGND_c_369_n 0.00669801f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_126 N_C_c_149_n N_VPWR_c_192_n 0.00762417f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_127 N_C_c_150_n N_VPWR_c_194_n 0.0100482f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_128 C N_VPWR_c_194_n 0.0317849f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_129 N_C_c_148_n N_VPWR_c_194_n 0.00310533f $X=3.365 $Y=1.21 $X2=0 $Y2=0
cc_130 N_C_c_149_n N_VPWR_c_195_n 0.00597712f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C_c_150_n N_VPWR_c_195_n 0.00673617f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C_c_149_n N_VPWR_c_186_n 0.0112769f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_133 N_C_c_150_n N_VPWR_c_186_n 0.0129313f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_134 N_C_c_149_n N_Y_c_245_n 0.0139912f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_135 C N_Y_c_245_n 0.00918194f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_136 N_C_c_148_n N_Y_c_245_n 3.10838e-19 $X=3.365 $Y=1.21 $X2=0 $Y2=0
cc_137 N_C_c_149_n N_Y_c_246_n 0.00292783f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_138 N_C_c_150_n N_Y_c_246_n 0.00349846f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_139 C N_Y_c_246_n 0.0305804f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_140 N_C_c_148_n N_Y_c_246_n 0.00760751f $X=3.365 $Y=1.21 $X2=0 $Y2=0
cc_141 N_C_c_149_n N_Y_c_283_n 0.0178402f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_142 N_C_c_150_n N_Y_c_283_n 0.0100147f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_143 N_C_M1004_g N_A_307_47#_c_340_n 0.0156754f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_144 N_C_c_146_n N_A_307_47#_c_340_n 0.00529891f $X=3.34 $Y=1.01 $X2=0 $Y2=0
cc_145 C N_A_307_47#_c_340_n 0.0376347f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_146 N_C_c_148_n N_A_307_47#_c_340_n 0.00332038f $X=3.365 $Y=1.21 $X2=0 $Y2=0
cc_147 N_C_M1004_g N_VGND_c_363_n 0.0108095f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_148 N_C_c_146_n N_VGND_c_363_n 0.00208456f $X=3.34 $Y=1.01 $X2=0 $Y2=0
cc_149 N_C_c_146_n N_VGND_c_365_n 0.0259861f $X=3.34 $Y=1.01 $X2=0 $Y2=0
cc_150 C N_VGND_c_365_n 0.0288662f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_151 N_C_c_148_n N_VGND_c_365_n 0.00317081f $X=3.365 $Y=1.21 $X2=0 $Y2=0
cc_152 N_C_M1004_g N_VGND_c_367_n 0.00339367f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_153 N_C_c_146_n N_VGND_c_367_n 0.00553327f $X=3.34 $Y=1.01 $X2=0 $Y2=0
cc_154 N_C_M1004_g N_VGND_c_369_n 0.00411889f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_155 N_C_c_146_n N_VGND_c_369_n 0.0113336f $X=3.34 $Y=1.01 $X2=0 $Y2=0
cc_156 N_VPWR_c_186_n N_Y_M1000_s 0.00231261f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_186_n N_Y_M1007_s 0.00231261f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_186_n N_Y_M1002_s 0.00231261f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_c_188_n N_Y_c_248_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_160 N_VPWR_c_189_n N_Y_c_248_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_190_n N_Y_c_248_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_162 N_VPWR_c_186_n N_Y_c_248_n 0.0140101f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_M1005_d N_Y_c_244_n 0.00180012f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_164 N_VPWR_c_190_n N_Y_c_244_n 0.0139097f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_165 N_VPWR_c_190_n N_Y_c_252_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_166 N_VPWR_c_191_n N_Y_c_252_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_192_n N_Y_c_252_n 0.0429581f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_168 N_VPWR_c_186_n N_Y_c_252_n 0.0140101f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_169 N_VPWR_M1010_d N_Y_c_245_n 0.00313113f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_170 N_VPWR_M1002_d N_Y_c_245_n 0.00313113f $X=2.535 $Y=1.485 $X2=0 $Y2=0
cc_171 N_VPWR_c_192_n N_Y_c_245_n 0.0578207f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_172 N_VPWR_c_194_n N_Y_c_246_n 0.0150684f $X=3.63 $Y=1.66 $X2=0 $Y2=0
cc_173 N_VPWR_c_192_n N_Y_c_283_n 0.0523533f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_174 N_VPWR_c_194_n N_Y_c_283_n 0.0520038f $X=3.63 $Y=1.66 $X2=0 $Y2=0
cc_175 N_VPWR_c_195_n N_Y_c_283_n 0.0223557f $X=3.515 $Y=2.72 $X2=0 $Y2=0
cc_176 N_VPWR_c_186_n N_Y_c_283_n 0.0140101f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_177 N_VPWR_c_188_n Y 0.0137498f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_178 N_Y_c_243_n N_A_27_47#_c_313_n 0.0115394f $X=0.73 $Y=0.72 $X2=0 $Y2=0
cc_179 N_Y_M1001_s N_A_27_47#_c_315_n 0.00414409f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_180 N_Y_c_243_n N_A_27_47#_c_315_n 0.0214701f $X=0.73 $Y=0.72 $X2=0 $Y2=0
cc_181 N_Y_c_245_n N_A_307_47#_c_340_n 0.00607047f $X=2.915 $Y=1.555 $X2=0 $Y2=0
cc_182 N_Y_c_243_n N_A_307_47#_c_340_n 0.00455089f $X=0.73 $Y=0.72 $X2=0 $Y2=0
cc_183 N_Y_M1001_s N_VGND_c_369_n 0.00259839f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_315_n N_A_307_47#_M1009_s 0.00415666f $X=2.14 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_185 N_A_27_47#_M1011_d N_A_307_47#_c_340_n 0.00321334f $X=2.005 $Y=0.235
+ $X2=0 $Y2=0
cc_186 N_A_27_47#_c_315_n N_A_307_47#_c_340_n 0.0473162f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_315_n N_VGND_c_363_n 0.0137364f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_314_n N_VGND_c_366_n 0.0139838f $X=0.345 $Y=0.38 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_315_n N_VGND_c_366_n 0.0880312f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_190 N_A_27_47#_M1001_d N_VGND_c_369_n 0.00253833f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1008_d N_VGND_c_369_n 0.00258215f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1011_d N_VGND_c_369_n 0.00211652f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_314_n N_VGND_c_369_n 0.00953535f $X=0.345 $Y=0.38 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_315_n N_VGND_c_369_n 0.0682273f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_195 N_A_307_47#_c_340_n N_VGND_M1004_d 0.00320842f $X=3.13 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A_307_47#_c_340_n N_VGND_c_363_n 0.0212463f $X=3.13 $Y=0.72 $X2=0 $Y2=0
cc_197 N_A_307_47#_c_340_n N_VGND_c_365_n 0.0169814f $X=3.13 $Y=0.72 $X2=0 $Y2=0
cc_198 N_A_307_47#_c_340_n N_VGND_c_366_n 0.00358f $X=3.13 $Y=0.72 $X2=0 $Y2=0
cc_199 N_A_307_47#_c_340_n N_VGND_c_367_n 0.00733853f $X=3.13 $Y=0.72 $X2=0
+ $Y2=0
cc_200 N_A_307_47#_M1009_s N_VGND_c_369_n 0.00259839f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_A_307_47#_M1004_s N_VGND_c_369_n 0.003737f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_202 N_A_307_47#_c_340_n N_VGND_c_369_n 0.0215685f $X=3.13 $Y=0.72 $X2=0 $Y2=0
