* File: sky130_fd_sc_hdll__einvn_2.pex.spice
* Created: Wed Sep  2 08:31:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%TE_B 1 2 3 5 8 10 12 14 15 17 19 20 21
c49 17 0 1.829e-19 $X=1.49 $Y=1.47
c50 15 0 9.48564e-20 $X=1.4 $Y=1.395
r51 21 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r52 17 19 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.49 $Y=1.47
+ $X2=1.49 $Y2=2.015
r53 16 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.11 $Y=1.395 $X2=1.02
+ $Y2=1.395
r54 15 17 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.4 $Y=1.395
+ $X2=1.49 $Y2=1.47
r55 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.4 $Y=1.395
+ $X2=1.11 $Y2=1.395
r56 12 20 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.47 $X2=1.02
+ $Y2=1.395
r57 12 14 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.02 $Y=1.47
+ $X2=1.02 $Y2=2.015
r58 11 24 28.2469 $w=4.01e-07 $l=3.42929e-07 $layer=POLY_cond $X=0.595 $Y=1.395
+ $X2=0.35 $Y2=1.16
r59 10 20 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=0.93 $Y=1.395 $X2=1.02
+ $Y2=1.395
r60 10 11 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.93 $Y=1.395
+ $X2=0.595 $Y2=1.395
r61 6 24 39.605 $w=4.01e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.35 $Y2=1.16
r62 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r63 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r64 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r65 1 11 21.1201 $w=4.01e-07 $l=1.32288e-07 $layer=POLY_cond $X=0.495 $Y=1.47
+ $X2=0.595 $Y2=1.395
r66 1 2 66.3154 $w=2e-07 $l=2e-07 $layer=POLY_cond $X=0.495 $Y=1.47 $X2=0.495
+ $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%A_27_47# 1 2 7 9 10 11 12 14 17 21 24 25
+ 27 36
c68 24 0 1.829e-19 $X=0.72 $Y=1.555
r69 28 36 22.4813 $w=2.68e-07 $l=1.25e-07 $layer=POLY_cond $X=1.935 $Y=1.16
+ $X2=1.935 $Y2=1.035
r70 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.16 $X2=1.935 $Y2=1.16
r71 25 27 40.7471 $w=2.78e-07 $l=9.9e-07 $layer=LI1_cond $X=0.945 $Y=1.135
+ $X2=1.935 $Y2=1.135
r72 23 25 8.0722 $w=3.83e-07 $l=2.98119e-07 $layer=LI1_cond $X=0.72 $Y=0.965
+ $X2=0.945 $Y2=1.135
r73 23 24 7.44227 $w=4.48e-07 $l=2.8e-07 $layer=LI1_cond $X=0.72 $Y=1.275
+ $X2=0.72 $Y2=1.555
r74 19 24 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=0.215 $Y=1.64
+ $X2=0.72 $Y2=1.64
r75 19 21 19.5029 $w=2.58e-07 $l=4.4e-07 $layer=LI1_cond $X=0.215 $Y=1.725
+ $X2=0.215 $Y2=2.165
r76 15 23 16.0862 $w=3.83e-07 $l=6.41541e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.72 $Y2=0.965
r77 15 17 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r78 12 36 22.7584 $w=2.68e-07 $l=9.28709e-08 $layer=POLY_cond $X=1.975 $Y=0.96
+ $X2=1.935 $Y2=1.035
r79 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.975 $Y=0.96
+ $X2=1.975 $Y2=0.56
r80 10 36 16.3317 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.8 $Y=1.035
+ $X2=1.935 $Y2=1.035
r81 10 11 87.1702 $w=1.5e-07 $l=1.7e-07 $layer=POLY_cond $X=1.8 $Y=1.035
+ $X2=1.63 $Y2=1.035
r82 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.555 $Y=0.96
+ $X2=1.63 $Y2=1.035
r83 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.555 $Y=0.96 $X2=1.555
+ $Y2=0.56
r84 2 21 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r85 1 17 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%A 3 5 7 8 10 11 13 14 19 27
r47 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.15
+ $Y=1.16 $X2=3.15 $Y2=1.16
r48 19 21 18.9157 $w=3.44e-07 $l=1.35e-07 $layer=POLY_cond $X=3.015 $Y=1.202
+ $X2=3.15 $Y2=1.202
r49 18 19 3.50291 $w=3.44e-07 $l=2.5e-08 $layer=POLY_cond $X=2.99 $Y=1.202
+ $X2=3.015 $Y2=1.202
r50 17 18 62.3517 $w=3.44e-07 $l=4.45e-07 $layer=POLY_cond $X=2.545 $Y=1.202
+ $X2=2.99 $Y2=1.202
r51 16 17 3.50291 $w=3.44e-07 $l=2.5e-08 $layer=POLY_cond $X=2.52 $Y=1.202
+ $X2=2.545 $Y2=1.202
r52 14 27 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.29 $Y=1.175
+ $X2=3.295 $Y2=1.175
r53 14 22 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=3.29 $Y=1.175
+ $X2=3.15 $Y2=1.175
r54 11 19 17.902 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.202
r55 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.985
r56 8 18 22.2144 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=1.202
r57 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.99 $Y=0.995
+ $X2=2.99 $Y2=0.56
r58 5 17 17.902 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.202
r59 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.985
r60 1 16 22.2144 $w=1.5e-07 $l=1.77e-07 $layer=POLY_cond $X=2.52 $Y=1.025
+ $X2=2.52 $Y2=1.202
r61 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.52 $Y=1.025
+ $X2=2.52 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%VPWR 1 2 9 11 15 17 18 19 21 37 38 41
r55 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 34 37 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r59 34 35 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r60 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 29 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r65 26 41 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.945 $Y=2.72
+ $X2=0.73 $Y2=2.72
r66 26 28 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.945 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 21 41 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.73 $Y2=2.72
r68 21 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 19 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 19 23 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 18 34 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 17 31 2.82709 $w=5.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.2 $Y=2.53 $X2=2.07
+ $Y2=2.53
r73 17 18 12.2241 $w=5.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.2 $Y=2.53
+ $X2=2.475 $Y2=2.53
r74 15 28 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 14 15 10.9193 $w=5.48e-07 $l=2.15e-07 $layer=LI1_cond $X=1.725 $Y=2.53
+ $X2=1.51 $Y2=2.53
r76 11 31 6.19786 $w=5.48e-07 $l=2.85e-07 $layer=LI1_cond $X=1.785 $Y=2.53
+ $X2=2.07 $Y2=2.53
r77 11 14 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=1.785 $Y=2.53
+ $X2=1.725 $Y2=2.53
r78 7 41 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r79 7 9 16.4826 $w=4.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.02
r80 2 14 600 $w=1.7e-07 $l=8.64465e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.545 $X2=1.725 $Y2=2.34
r81 1 9 300 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.845 $X2=0.755 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%A_222_309# 1 2 9 11 15 20
r43 18 20 18.0146 $w=6.38e-07 $l=6.7e-07 $layer=LI1_cond $X=1.255 $Y=1.765
+ $X2=1.925 $Y2=1.765
r44 13 15 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.78 $Y=2.085
+ $X2=2.78 $Y2=2.265
r45 11 13 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.695 $Y=1.975
+ $X2=2.78 $Y2=2.085
r46 11 20 40.3355 $w=2.18e-07 $l=7.7e-07 $layer=LI1_cond $X=2.695 $Y=1.975
+ $X2=1.925 $Y2=1.975
r47 7 18 8.73481 $w=1.7e-07 $l=3.2e-07 $layer=LI1_cond $X=1.255 $Y=2.085
+ $X2=1.255 $Y2=1.765
r48 7 9 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.255 $Y=2.085
+ $X2=1.255 $Y2=2.265
r49 2 15 600 $w=1.7e-07 $l=8.49412e-07 $layer=licon1_PDIFF $count=1 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=2.265
r50 1 18 600 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.545 $X2=1.255 $Y2=1.925
r51 1 9 600 $w=1.7e-07 $l=7.89177e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.545 $X2=1.255 $Y2=2.265
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%Z 1 2 3 10 11 12 13 14 15 16 24 28 32 47
+ 50
c41 24 0 9.48564e-20 $X=2.445 $Y=1.57
r42 38 50 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=3.285 $Y=1.57
+ $X2=3.26 $Y2=1.57
r43 30 47 5.9927 $w=2.48e-07 $l=1.3e-07 $layer=LI1_cond $X=2.63 $Y=1.57 $X2=2.76
+ $Y2=1.57
r44 24 30 8.52808 $w=2.48e-07 $l=1.85e-07 $layer=LI1_cond $X=2.445 $Y=1.57
+ $X2=2.63 $Y2=1.57
r45 24 28 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=2.445 $Y=1.57
+ $X2=2.3 $Y2=1.57
r46 15 16 9.44902 $w=4.98e-07 $l=3.95e-07 $layer=LI1_cond $X=3.285 $Y=1.815
+ $X2=3.285 $Y2=2.21
r47 15 38 2.87059 $w=4.98e-07 $l=1.2e-07 $layer=LI1_cond $X=3.285 $Y=1.815
+ $X2=3.285 $Y2=1.695
r48 14 38 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.29 $Y=1.57
+ $X2=3.285 $Y2=1.57
r49 13 50 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=2.78 $Y=1.57
+ $X2=3.26 $Y2=1.57
r50 13 47 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=2.78 $Y=1.57 $X2=2.76
+ $Y2=1.57
r51 12 32 2.80324 $w=3.68e-07 $l=9e-08 $layer=LI1_cond $X=2.63 $Y=0.85 $X2=2.63
+ $Y2=0.76
r52 11 30 7.94251 $w=3.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.63 $Y=1.19
+ $X2=2.63 $Y2=1.445
r53 11 12 10.59 $w=3.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.63 $Y=1.19 $X2=2.63
+ $Y2=0.85
r54 10 28 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=2.27 $Y=1.57 $X2=2.3
+ $Y2=1.57
r55 3 15 300 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.485 $X2=3.25 $Y2=1.815
r56 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.485 $X2=2.31 $Y2=1.61
r57 1 32 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.73 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%VGND 1 2 9 11 15 17 19 29 30 33 36
r48 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r50 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 27 30 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r53 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r54 26 29 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r55 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r56 24 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.765
+ $Y2=0
r57 24 26 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.07
+ $Y2=0
r58 19 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r59 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r60 17 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r62 13 36 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=0.085
+ $X2=1.765 $Y2=0
r63 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.765 $Y=0.085
+ $X2=1.765 $Y2=0.36
r64 12 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r65 11 36 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.765
+ $Y2=0
r66 11 12 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.6 $Y=0 $X2=0.895
+ $Y2=0
r67 7 33 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r68 7 9 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.38
r69 2 15 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.63
+ $Y=0.235 $X2=1.765 $Y2=0.36
r70 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_2%A_234_47# 1 2 3 12 17 18 19 22 25
r42 20 22 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.3 $Y=0.425
+ $X2=3.3 $Y2=0.56
r43 18 20 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.165 $Y=0.34
+ $X2=3.3 $Y2=0.425
r44 18 19 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=3.165 $Y=0.34
+ $X2=2.27 $Y2=0.34
r45 15 17 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.185 $Y=0.655
+ $X2=2.185 $Y2=0.56
r46 14 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.185 $Y=0.425
+ $X2=2.27 $Y2=0.34
r47 14 17 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.185 $Y=0.425
+ $X2=2.185 $Y2=0.56
r48 13 25 4.96789 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=1.38 $Y=0.74
+ $X2=1.222 $Y2=0.74
r49 12 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.1 $Y=0.74
+ $X2=2.185 $Y2=0.655
r50 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=2.1 $Y=0.74 $X2=1.38
+ $Y2=0.74
r51 3 22 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.25 $Y2=0.56
r52 2 17 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.05
+ $Y=0.235 $X2=2.185 $Y2=0.56
r53 1 25 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=1.17
+ $Y=0.235 $X2=1.295 $Y2=0.74
.ends

