* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o221a_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 a_38_47# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_38_47# C1 a_151_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VGND a_38_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_38_47# A2 a_535_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_535_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND A2 a_245_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_245_47# B2 a_151_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR B1 a_255_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 X a_38_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 X a_38_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_151_47# B1 a_245_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_255_297# B2 a_38_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR a_38_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_245_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
