* File: sky130_fd_sc_hdll__or3b_1.pxi.spice
* Created: Wed Sep  2 08:48:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3B_1%C_N N_C_N_c_70_n N_C_N_M1003_g N_C_N_c_67_n
+ N_C_N_M1006_g C_N N_C_N_c_69_n C_N PM_SKY130_FD_SC_HDLL__OR3B_1%C_N
x_PM_SKY130_FD_SC_HDLL__OR3B_1%A_117_297# N_A_117_297#_M1006_d
+ N_A_117_297#_M1003_d N_A_117_297#_c_94_n N_A_117_297#_M1007_g
+ N_A_117_297#_M1002_g N_A_117_297#_c_91_n N_A_117_297#_c_92_n
+ N_A_117_297#_c_93_n N_A_117_297#_c_98_n
+ PM_SKY130_FD_SC_HDLL__OR3B_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__OR3B_1%B N_B_c_132_n N_B_c_133_n N_B_c_135_n N_B_c_136_n
+ N_B_M1005_g N_B_M1000_g N_B_c_134_n B B B N_B_c_138_n B B B
+ PM_SKY130_FD_SC_HDLL__OR3B_1%B
x_PM_SKY130_FD_SC_HDLL__OR3B_1%A N_A_c_172_n N_A_M1004_g N_A_M1001_g A A A
+ N_A_c_174_n N_A_c_175_n A PM_SKY130_FD_SC_HDLL__OR3B_1%A
x_PM_SKY130_FD_SC_HDLL__OR3B_1%A_225_53# N_A_225_53#_M1002_s N_A_225_53#_M1000_d
+ N_A_225_53#_M1007_s N_A_225_53#_c_221_n N_A_225_53#_M1008_g
+ N_A_225_53#_c_222_n N_A_225_53#_M1009_g N_A_225_53#_c_223_n
+ N_A_225_53#_c_231_n N_A_225_53#_c_224_n N_A_225_53#_c_225_n
+ N_A_225_53#_c_232_n N_A_225_53#_c_233_n N_A_225_53#_c_300_p
+ N_A_225_53#_c_226_n N_A_225_53#_c_269_n N_A_225_53#_c_234_n
+ N_A_225_53#_c_227_n N_A_225_53#_c_235_n N_A_225_53#_c_228_n
+ N_A_225_53#_c_229_n PM_SKY130_FD_SC_HDLL__OR3B_1%A_225_53#
x_PM_SKY130_FD_SC_HDLL__OR3B_1%VPWR N_VPWR_M1003_s N_VPWR_M1004_d N_VPWR_c_315_n
+ N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n N_VPWR_c_319_n VPWR
+ N_VPWR_c_320_n N_VPWR_c_314_n PM_SKY130_FD_SC_HDLL__OR3B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3B_1%X N_X_M1009_d N_X_M1008_d N_X_c_351_n N_X_c_353_n
+ N_X_c_352_n X PM_SKY130_FD_SC_HDLL__OR3B_1%X
x_PM_SKY130_FD_SC_HDLL__OR3B_1%VGND N_VGND_M1006_s N_VGND_M1002_d N_VGND_M1001_d
+ N_VGND_c_369_n N_VGND_c_370_n N_VGND_c_371_n VGND N_VGND_c_372_n
+ N_VGND_c_373_n N_VGND_c_374_n N_VGND_c_375_n N_VGND_c_376_n
+ PM_SKY130_FD_SC_HDLL__OR3B_1%VGND
cc_1 VNB N_C_N_c_67_n 0.0214087f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB C_N 0.00874107f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_69_n 0.0453644f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_117_297#_M1002_g 0.0311171f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_5 VNB N_A_117_297#_c_91_n 0.0259433f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_6 VNB N_A_117_297#_c_92_n 0.0111748f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_A_117_297#_c_93_n 0.0220809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B_c_132_n 0.00670441f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_B_c_133_n 0.0216074f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_10 VNB N_B_c_134_n 0.0142901f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_11 VNB N_A_c_172_n 0.0214548f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_A_M1001_g 0.0284569f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.675
cc_13 VNB N_A_c_174_n 0.0026363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_c_175_n 0.00172512f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_15 VNB N_A_225_53#_c_221_n 0.0242891f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_16 VNB N_A_225_53#_c_222_n 0.0209442f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_17 VNB N_A_225_53#_c_223_n 0.0088433f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_53#_c_224_n 0.00387737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_225_53#_c_225_n 0.00393129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_53#_c_226_n 0.00177504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_225_53#_c_227_n 0.00150105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_225_53#_c_228_n 0.00290988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_225_53#_c_229_n 0.0018431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_314_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_351_n 0.0177099f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_26 VNB N_X_c_352_n 0.0290836f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_27 VNB N_VGND_c_369_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_VGND_c_370_n 0.0388559f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_29 VNB N_VGND_c_371_n 0.0010436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_372_n 0.0305624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_373_n 0.023165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_374_n 0.0249567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_375_n 0.22599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_376_n 0.00544933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_C_N_c_70_n 0.0235164f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB C_N 8.94523e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_37 VPB N_C_N_c_69_n 0.0191905f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_38 VPB N_A_117_297#_c_94_n 0.0187575f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_39 VPB N_A_117_297#_c_91_n 0.0103639f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_40 VPB N_A_117_297#_c_92_n 0.00650162f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_41 VPB N_A_117_297#_c_93_n 0.0120926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_117_297#_c_98_n 0.00461033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B_c_135_n 0.00617305f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_44 VPB N_B_c_136_n 0.0488187f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_45 VPB N_B_M1005_g 0.0111419f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.675
cc_46 VPB N_B_c_138_n 0.0511848f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_c_172_n 0.0273426f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB A 0.00149589f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_49 VPB N_A_c_174_n 0.00354214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_225_53#_c_221_n 0.0323221f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_51 VPB N_A_225_53#_c_231_n 0.00319925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_225_53#_c_232_n 0.0039877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_225_53#_c_233_n 0.00462889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_225_53#_c_234_n 0.00156472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_225_53#_c_235_n 0.00139614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_315_n 0.00983572f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_57 VPB N_VPWR_c_316_n 0.0568304f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_58 VPB N_VPWR_c_317_n 0.0113669f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_59 VPB N_VPWR_c_318_n 0.0549492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_319_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_61 VPB N_VPWR_c_320_n 0.0245761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_314_n 0.0742847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_X_c_353_n 0.0097098f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_64 VPB N_X_c_352_n 0.010412f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_65 VPB X 0.0361203f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_66 N_C_N_c_69_n N_A_117_297#_c_91_n 0.00706646f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_67 N_C_N_c_67_n N_A_117_297#_c_93_n 0.0224674f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_68 C_N N_A_117_297#_c_93_n 0.0171994f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_69 N_C_N_c_70_n N_A_117_297#_c_98_n 0.00610416f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 N_C_N_c_69_n N_A_117_297#_c_98_n 0.00340849f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_71 N_C_N_c_67_n N_A_225_53#_c_223_n 0.00428704f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_72 N_C_N_c_70_n N_A_225_53#_c_233_n 0.00234292f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C_N_c_70_n N_VPWR_c_316_n 0.00877297f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 C_N N_VPWR_c_316_n 0.020735f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 N_C_N_c_69_n N_VPWR_c_316_n 0.00545118f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_76 N_C_N_c_70_n N_VPWR_c_318_n 0.00393512f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_77 N_C_N_c_70_n N_VPWR_c_314_n 0.00500987f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_78 N_C_N_c_67_n N_VGND_c_370_n 0.0082712f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_79 C_N N_VGND_c_370_n 0.0210991f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_80 N_C_N_c_69_n N_VGND_c_370_n 0.00600816f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_81 N_C_N_c_67_n N_VGND_c_372_n 0.00439675f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_82 N_C_N_c_67_n N_VGND_c_375_n 0.00512902f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_117_297#_M1002_g N_B_c_132_n 0.0199102f $X=1.51 $Y=0.475 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_117_297#_c_92_n N_B_c_133_n 0.0199102f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_85 N_A_117_297#_c_94_n N_B_M1005_g 0.0332289f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_117_297#_M1002_g N_B_c_134_n 0.0137274f $X=1.51 $Y=0.475 $X2=0 $Y2=0
cc_87 N_A_117_297#_c_94_n N_B_c_138_n 0.00528678f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_117_297#_c_98_n N_B_c_138_n 0.0106665f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_89 N_A_117_297#_c_94_n A 0.00761075f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_117_297#_c_92_n A 0.00457154f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_91 N_A_117_297#_c_92_n N_A_c_175_n 0.0118108f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_92 N_A_117_297#_c_93_n N_A_c_175_n 0.020012f $X=0.73 $Y=1.325 $X2=0 $Y2=0
cc_93 N_A_117_297#_M1002_g N_A_225_53#_c_223_n 0.00504015f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_94 N_A_117_297#_c_93_n N_A_225_53#_c_223_n 0.0135221f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_95 N_A_117_297#_c_91_n N_A_225_53#_c_231_n 0.00334724f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_117_297#_c_93_n N_A_225_53#_c_231_n 0.0156876f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_97 N_A_117_297#_c_98_n N_A_225_53#_c_231_n 0.0163366f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_98 N_A_117_297#_M1002_g N_A_225_53#_c_224_n 0.0151676f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_99 N_A_117_297#_c_91_n N_A_225_53#_c_224_n 0.00388751f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_117_297#_c_91_n N_A_225_53#_c_225_n 0.00345493f $X=1.385 $Y=1.16
+ $X2=0 $Y2=0
cc_101 N_A_117_297#_c_93_n N_A_225_53#_c_225_n 0.0309385f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_102 N_A_117_297#_c_94_n N_A_225_53#_c_232_n 0.0137869f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_A_117_297#_c_98_n N_A_225_53#_c_233_n 0.00612897f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_104 N_A_117_297#_c_98_n N_VPWR_c_316_n 0.0192564f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_105 N_A_117_297#_c_93_n N_VGND_c_370_n 0.032547f $X=0.73 $Y=1.325 $X2=0 $Y2=0
cc_106 N_A_117_297#_M1002_g N_VGND_c_371_n 0.0107839f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_107 N_A_117_297#_M1002_g N_VGND_c_372_n 0.00187556f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_108 N_A_117_297#_c_93_n N_VGND_c_372_n 0.00967825f $X=0.73 $Y=1.325 $X2=0
+ $Y2=0
cc_109 N_A_117_297#_M1002_g N_VGND_c_375_n 0.00356717f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_110 N_A_117_297#_c_93_n N_VGND_c_375_n 0.012569f $X=0.73 $Y=1.325 $X2=0 $Y2=0
cc_111 N_B_c_133_n N_A_c_172_n 0.0180488f $X=1.905 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_112 N_B_c_135_n N_A_c_172_n 0.00367285f $X=1.905 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_113 N_B_M1005_g N_A_c_172_n 0.0219568f $X=1.905 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_114 N_B_c_138_n N_A_c_172_n 6.06139e-19 $X=1.94 $Y=2.31 $X2=-0.19 $Y2=-0.24
cc_115 N_B_c_134_n N_A_M1001_g 0.0169001f $X=1.905 $Y=0.76 $X2=0 $Y2=0
cc_116 N_B_c_135_n A 0.00215744f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B_M1005_g A 0.00239676f $X=1.905 $Y=1.695 $X2=0 $Y2=0
cc_118 N_B_c_133_n N_A_c_174_n 0.0147857f $X=1.905 $Y=1.31 $X2=0 $Y2=0
cc_119 N_B_c_135_n N_A_c_174_n 0.00522181f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B_c_132_n N_A_225_53#_c_224_n 0.00628546f $X=1.905 $Y=0.86 $X2=0 $Y2=0
cc_121 N_B_c_134_n N_A_225_53#_c_224_n 0.00712359f $X=1.905 $Y=0.76 $X2=0 $Y2=0
cc_122 N_B_c_136_n N_A_225_53#_c_232_n 7.17844e-19 $X=1.905 $Y=2.035 $X2=0 $Y2=0
cc_123 N_B_M1005_g N_A_225_53#_c_232_n 0.0128616f $X=1.905 $Y=1.695 $X2=0 $Y2=0
cc_124 N_B_c_138_n N_A_225_53#_c_232_n 0.0628104f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_125 N_B_c_138_n N_A_225_53#_c_233_n 0.0215827f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_126 N_B_M1005_g N_A_225_53#_c_235_n 0.00481342f $X=1.905 $Y=1.695 $X2=0 $Y2=0
cc_127 N_B_c_138_n N_A_225_53#_c_235_n 0.0138656f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_128 N_B_c_138_n N_VPWR_c_316_n 0.0196594f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_129 N_B_c_136_n N_VPWR_c_317_n 0.00415023f $X=1.905 $Y=2.035 $X2=0 $Y2=0
cc_130 N_B_c_138_n N_VPWR_c_317_n 0.0239207f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_131 N_B_c_136_n N_VPWR_c_318_n 0.00676986f $X=1.905 $Y=2.035 $X2=0 $Y2=0
cc_132 N_B_c_138_n N_VPWR_c_318_n 0.108123f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_133 N_B_c_136_n N_VPWR_c_314_n 0.00939765f $X=1.905 $Y=2.035 $X2=0 $Y2=0
cc_134 N_B_c_138_n N_VPWR_c_314_n 0.0643141f $X=1.94 $Y=2.31 $X2=0 $Y2=0
cc_135 N_B_c_134_n N_VGND_c_371_n 0.00720054f $X=1.905 $Y=0.76 $X2=0 $Y2=0
cc_136 N_B_c_134_n N_VGND_c_373_n 0.00376964f $X=1.905 $Y=0.76 $X2=0 $Y2=0
cc_137 N_B_c_134_n N_VGND_c_375_n 0.0040746f $X=1.905 $Y=0.76 $X2=0 $Y2=0
cc_138 N_A_c_172_n N_A_225_53#_c_221_n 0.0340889f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_174_n N_A_225_53#_c_221_n 3.50713e-19 $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_A_225_53#_c_222_n 0.017558f $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_141 A N_A_225_53#_c_231_n 0.00821086f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_142 N_A_c_174_n N_A_225_53#_c_224_n 0.0249068f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_175_n N_A_225_53#_c_224_n 0.0200426f $X=1.647 $Y=1.325 $X2=0 $Y2=0
cc_144 N_A_c_172_n N_A_225_53#_c_232_n 2.14526e-19 $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_145 A N_A_225_53#_c_232_n 0.013878f $X=1.525 $Y=1.445 $X2=0 $Y2=0
cc_146 N_A_c_174_n N_A_225_53#_c_232_n 0.01267f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_c_172_n N_A_225_53#_c_226_n 0.00229621f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_M1001_g N_A_225_53#_c_226_n 0.0125258f $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_149 N_A_c_174_n N_A_225_53#_c_226_n 0.0138864f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_c_172_n N_A_225_53#_c_269_n 0.0147951f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_174_n N_A_225_53#_c_269_n 0.00821244f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_c_172_n N_A_225_53#_c_234_n 0.00173315f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_172_n N_A_225_53#_c_227_n 5.36764e-19 $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_174_n N_A_225_53#_c_227_n 0.0146459f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_c_172_n N_A_225_53#_c_235_n 0.0113409f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_174_n N_A_225_53#_c_235_n 0.0112473f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_c_172_n N_A_225_53#_c_228_n 0.00375514f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_174_n N_A_225_53#_c_228_n 0.020012f $X=2.38 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_M1001_g N_A_225_53#_c_229_n 0.00375514f $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_160 N_A_c_172_n N_VPWR_c_317_n 0.00330158f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_172_n N_VPWR_c_318_n 0.00351015f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_172_n N_VPWR_c_314_n 0.00445321f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_163 A A_315_297# 0.00139384f $X=1.525 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_164 N_A_M1001_g N_VGND_c_371_n 5.04903e-19 $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_165 N_A_M1001_g N_VGND_c_373_n 0.0118414f $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_166 N_A_M1001_g N_VGND_c_375_n 0.00282535f $X=2.445 $Y=0.475 $X2=0 $Y2=0
cc_167 N_A_225_53#_c_269_n N_VPWR_M1004_d 0.00563715f $X=2.72 $Y=1.58 $X2=0
+ $Y2=0
cc_168 N_A_225_53#_c_221_n N_VPWR_c_317_n 0.00505337f $X=2.96 $Y=1.41 $X2=0
+ $Y2=0
cc_169 N_A_225_53#_c_269_n N_VPWR_c_317_n 0.0204259f $X=2.72 $Y=1.58 $X2=0 $Y2=0
cc_170 N_A_225_53#_c_235_n N_VPWR_c_317_n 0.00726621f $X=2.265 $Y=1.58 $X2=0
+ $Y2=0
cc_171 N_A_225_53#_c_221_n N_VPWR_c_320_n 0.00702461f $X=2.96 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_225_53#_c_221_n N_VPWR_c_314_n 0.014874f $X=2.96 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_225_53#_c_232_n A_315_297# 0.0013394f $X=2.18 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_225_53#_c_232_n A_399_297# 0.00249728f $X=2.18 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_225_53#_c_235_n A_399_297# 0.00469227f $X=2.265 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_225_53#_c_221_n N_X_c_353_n 0.0127049f $X=2.96 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_225_53#_c_269_n N_X_c_353_n 0.0114924f $X=2.72 $Y=1.58 $X2=0 $Y2=0
cc_178 N_A_225_53#_c_221_n N_X_c_352_n 7.62883e-19 $X=2.96 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_225_53#_c_222_n N_X_c_352_n 0.0136361f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_225_53#_c_234_n N_X_c_352_n 0.00554781f $X=2.805 $Y=1.495 $X2=0 $Y2=0
cc_181 N_A_225_53#_c_228_n N_X_c_352_n 0.021207f $X=2.91 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_225_53#_c_229_n N_X_c_352_n 0.00697759f $X=2.857 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_225_53#_c_224_n N_VGND_M1002_d 0.00160115f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_184 N_A_225_53#_c_226_n N_VGND_M1001_d 0.00660803f $X=2.72 $Y=0.74 $X2=0
+ $Y2=0
cc_185 N_A_225_53#_c_229_n N_VGND_M1001_d 6.98847e-19 $X=2.857 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_225_53#_c_223_n N_VGND_c_371_n 0.0177338f $X=1.25 $Y=0.42 $X2=0 $Y2=0
cc_187 N_A_225_53#_c_224_n N_VGND_c_371_n 0.0196541f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_188 N_A_225_53#_c_300_p N_VGND_c_371_n 0.0110177f $X=2.19 $Y=0.47 $X2=0 $Y2=0
cc_189 N_A_225_53#_c_223_n N_VGND_c_372_n 0.0182527f $X=1.25 $Y=0.42 $X2=0 $Y2=0
cc_190 N_A_225_53#_c_224_n N_VGND_c_372_n 0.00232694f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_191 N_A_225_53#_c_221_n N_VGND_c_373_n 3.3049e-19 $X=2.96 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_225_53#_c_222_n N_VGND_c_373_n 0.00498441f $X=2.985 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_225_53#_c_224_n N_VGND_c_373_n 0.00310196f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_194 N_A_225_53#_c_300_p N_VGND_c_373_n 0.0223186f $X=2.19 $Y=0.47 $X2=0 $Y2=0
cc_195 N_A_225_53#_c_226_n N_VGND_c_373_n 0.0298237f $X=2.72 $Y=0.74 $X2=0 $Y2=0
cc_196 N_A_225_53#_c_222_n N_VGND_c_374_n 0.00585385f $X=2.985 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_225_53#_c_222_n N_VGND_c_375_n 0.0123608f $X=2.985 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_225_53#_c_223_n N_VGND_c_375_n 0.00989054f $X=1.25 $Y=0.42 $X2=0
+ $Y2=0
cc_199 N_A_225_53#_c_224_n N_VGND_c_375_n 0.0115556f $X=2.105 $Y=0.74 $X2=0
+ $Y2=0
cc_200 N_A_225_53#_c_300_p N_VGND_c_375_n 0.00625722f $X=2.19 $Y=0.47 $X2=0
+ $Y2=0
cc_201 N_A_225_53#_c_226_n N_VGND_c_375_n 0.00684962f $X=2.72 $Y=0.74 $X2=0
+ $Y2=0
cc_202 N_VPWR_c_314_n N_X_M1008_d 0.00442383f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_c_320_n X 0.0300192f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_204 N_VPWR_c_314_n X 0.0162905f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_205 N_X_c_351_n N_VGND_c_374_n 0.014483f $X=3.195 $Y=0.59 $X2=0 $Y2=0
cc_206 N_X_M1009_d N_VGND_c_375_n 0.00419212f $X=3.06 $Y=0.235 $X2=0 $Y2=0
cc_207 N_X_c_351_n N_VGND_c_375_n 0.0147712f $X=3.195 $Y=0.59 $X2=0 $Y2=0
