# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__mux2_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.40000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.105000 1.075000 9.455000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.075000 1.915000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.665000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.925000 1.075000 4.275000 1.325000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  3.724000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.585000 0.255000 10.915000 0.725000 ;
        RECT 10.585000 0.725000 17.495000 0.905000 ;
        RECT 10.585000 1.495000 17.495000 1.665000 ;
        RECT 10.585000 1.665000 10.915000 2.465000 ;
        RECT 11.525000 0.255000 11.855000 0.725000 ;
        RECT 11.525000 1.665000 11.855000 2.465000 ;
        RECT 12.465000 0.255000 12.795000 0.725000 ;
        RECT 12.465000 1.665000 12.795000 2.465000 ;
        RECT 13.405000 0.255000 13.735000 0.725000 ;
        RECT 13.405000 1.665000 13.735000 2.465000 ;
        RECT 14.345000 0.255000 14.675000 0.725000 ;
        RECT 14.345000 1.665000 14.675000 2.465000 ;
        RECT 15.285000 0.255000 15.615000 0.725000 ;
        RECT 15.285000 1.665000 15.615000 2.465000 ;
        RECT 16.225000 0.255000 16.555000 0.725000 ;
        RECT 16.225000 1.665000 16.555000 2.465000 ;
        RECT 17.085000 0.905000 17.495000 1.495000 ;
        RECT 17.165000 0.255000 17.495000 0.725000 ;
        RECT 17.165000 1.665000 17.495000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 18.400000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 18.400000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.400000 0.085000 ;
      RECT  0.000000  2.635000 18.400000 2.805000 ;
      RECT  0.095000  0.255000  2.305000 0.425000 ;
      RECT  0.095000  0.425000  0.395000 2.295000 ;
      RECT  0.095000  2.295000  2.305000 2.465000 ;
      RECT  0.565000  0.595000  0.895000 0.725000 ;
      RECT  0.565000  0.725000  4.235000 0.905000 ;
      RECT  0.565000  1.495000  1.835000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.125000 ;
      RECT  1.065000  0.425000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.295000 ;
      RECT  1.505000  0.595000  1.835000 0.725000 ;
      RECT  1.505000  1.665000  1.835000 2.125000 ;
      RECT  2.005000  0.425000  2.305000 0.550000 ;
      RECT  2.005000  1.495000  2.305000 2.295000 ;
      RECT  2.525000  0.085000  2.795000 0.550000 ;
      RECT  2.525000  1.495000  2.795000 2.635000 ;
      RECT  2.965000  0.255000  3.295000 0.725000 ;
      RECT  2.965000  1.495000  4.235000 1.665000 ;
      RECT  2.965000  1.665000  3.295000 2.465000 ;
      RECT  3.465000  0.085000  3.735000 0.545000 ;
      RECT  3.465000  1.835000  3.735000 2.635000 ;
      RECT  3.905000  0.255000  4.235000 0.725000 ;
      RECT  3.905000  1.665000  4.235000 2.465000 ;
      RECT  4.405000  0.085000  4.675000 0.905000 ;
      RECT  4.405000  1.495000  4.675000 2.635000 ;
      RECT  4.845000  0.255000  5.175000 1.075000 ;
      RECT  4.845000  1.075000  7.095000 1.325000 ;
      RECT  4.845000  1.325000  5.175000 2.465000 ;
      RECT  5.345000  0.085000  5.615000 0.905000 ;
      RECT  5.345000  1.495000  5.615000 2.635000 ;
      RECT  5.785000  0.255000  6.115000 0.725000 ;
      RECT  5.785000  0.725000  9.455000 0.905000 ;
      RECT  5.785000  1.495000  7.055000 1.665000 ;
      RECT  5.785000  1.665000  6.115000 2.465000 ;
      RECT  6.285000  0.085000  6.555000 0.545000 ;
      RECT  6.285000  1.835000  6.555000 2.635000 ;
      RECT  6.725000  0.255000  7.055000 0.725000 ;
      RECT  6.725000  1.665000  7.055000 2.465000 ;
      RECT  7.225000  0.085000  7.495000 0.550000 ;
      RECT  7.225000  1.495000  7.495000 2.635000 ;
      RECT  7.715000  0.255000  9.925000 0.425000 ;
      RECT  7.715000  0.425000  8.015000 0.550000 ;
      RECT  7.715000  1.495000  8.015000 2.295000 ;
      RECT  7.715000  2.295000  9.925000 2.465000 ;
      RECT  8.185000  0.595000  8.515000 0.725000 ;
      RECT  8.185000  1.495000  9.455000 1.665000 ;
      RECT  8.185000  1.665000  8.515000 2.125000 ;
      RECT  8.685000  0.425000  8.955000 0.545000 ;
      RECT  8.685000  1.835000  8.955000 2.295000 ;
      RECT  9.125000  0.595000  9.455000 0.725000 ;
      RECT  9.125000  1.665000  9.455000 2.125000 ;
      RECT  9.625000  0.425000  9.925000 1.075000 ;
      RECT  9.625000  1.075000 16.865000 1.325000 ;
      RECT  9.625000  1.325000  9.925000 2.295000 ;
      RECT 10.145000  0.085000 10.415000 0.905000 ;
      RECT 10.145000  1.495000 10.415000 2.635000 ;
      RECT 11.085000  0.085000 11.355000 0.545000 ;
      RECT 11.085000  1.835000 11.355000 2.635000 ;
      RECT 12.025000  0.085000 12.295000 0.545000 ;
      RECT 12.025000  1.835000 12.295000 2.635000 ;
      RECT 12.965000  0.085000 13.235000 0.545000 ;
      RECT 12.965000  1.835000 13.235000 2.635000 ;
      RECT 13.905000  0.085000 14.175000 0.550000 ;
      RECT 13.905000  1.835000 14.175000 2.635000 ;
      RECT 14.845000  0.085000 15.115000 0.545000 ;
      RECT 14.845000  1.835000 15.115000 2.635000 ;
      RECT 15.785000  0.085000 16.055000 0.545000 ;
      RECT 15.785000  1.835000 16.055000 2.635000 ;
      RECT 16.725000  0.085000 16.995000 0.545000 ;
      RECT 16.725000  1.835000 16.995000 2.635000 ;
      RECT 17.665000  0.085000 17.935000 0.905000 ;
      RECT 17.665000  1.495000 17.935000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.175000  0.425000  0.345000 0.595000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.645000  1.785000  0.815000 1.955000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.585000  1.785000  1.755000 1.955000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.045000  2.125000  3.215000 2.295000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.985000  2.125000  4.155000 2.295000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  5.865000  1.785000  6.035000 1.955000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  6.805000  1.785000  6.975000 1.955000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.265000  1.785000  8.435000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.205000  1.785000  9.375000 1.955000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.675000  0.425000  9.845000 0.595000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
    LAYER met1 ;
      RECT 0.115000 0.395000 0.405000 0.440000 ;
      RECT 0.115000 0.440000 9.905000 0.580000 ;
      RECT 0.115000 0.580000 0.405000 0.625000 ;
      RECT 0.585000 1.755000 0.875000 1.800000 ;
      RECT 0.585000 1.800000 7.035000 1.940000 ;
      RECT 0.585000 1.940000 0.875000 1.985000 ;
      RECT 1.525000 1.755000 1.815000 1.800000 ;
      RECT 1.525000 1.940000 1.815000 1.985000 ;
      RECT 2.985000 2.095000 3.275000 2.140000 ;
      RECT 2.985000 2.140000 7.660000 2.280000 ;
      RECT 2.985000 2.280000 3.275000 2.325000 ;
      RECT 3.925000 2.095000 4.215000 2.140000 ;
      RECT 3.925000 2.280000 4.215000 2.325000 ;
      RECT 5.805000 1.755000 6.095000 1.800000 ;
      RECT 5.805000 1.940000 6.095000 1.985000 ;
      RECT 6.745000 1.755000 7.035000 1.800000 ;
      RECT 6.745000 1.940000 7.035000 1.985000 ;
      RECT 7.520000 1.800000 9.435000 1.940000 ;
      RECT 7.520000 1.940000 7.660000 2.140000 ;
      RECT 8.205000 1.755000 8.495000 1.800000 ;
      RECT 8.205000 1.940000 8.495000 1.985000 ;
      RECT 9.145000 1.755000 9.435000 1.800000 ;
      RECT 9.145000 1.940000 9.435000 1.985000 ;
      RECT 9.615000 0.395000 9.905000 0.440000 ;
      RECT 9.615000 0.580000 9.905000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_16
END LIBRARY
