* File: sky130_fd_sc_hdll__a31o_4.pex.spice
* Created: Wed Sep  2 08:20:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31O_4%A3 1 3 4 6 7 9 10 12 13 16 21 22 27
c81 10 0 2.32895e-19 $X=2.905 $Y=1.41
c82 7 0 1.74322e-19 $X=2.88 $Y=0.995
r83 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r84 21 22 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=0.335 $Y=1.19
+ $X2=0.335 $Y2=1.53
r85 21 27 0.909823 $w=3.78e-07 $l=3e-08 $layer=LI1_cond $X=0.335 $Y=1.19
+ $X2=0.335 $Y2=1.16
r86 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=2.965 $Y=1.16
+ $X2=2.965 $Y2=1.53
r87 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.94
+ $Y=1.16 $X2=2.94 $Y2=1.16
r88 14 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=1.53
+ $X2=0.335 $Y2=1.53
r89 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.53
+ $X2=2.965 $Y2=1.53
r90 13 14 146.791 $w=1.68e-07 $l=2.25e-06 $layer=LI1_cond $X=2.775 $Y=1.53
+ $X2=0.525 $Y2=1.53
r91 10 17 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.965 $Y2=1.16
r92 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.905 $Y=1.41
+ $X2=2.905 $Y2=1.985
r93 7 17 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.88 $Y=0.995
+ $X2=2.965 $Y2=1.16
r94 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.88 $Y=0.995 $X2=2.88
+ $Y2=0.56
r95 4 26 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.41 $Y2=1.16
r96 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r97 1 26 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.41 $Y2=1.16
r98 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%A2 1 3 4 6 7 9 10 12 13 16 19 22 23 30
c75 13 0 1.74322e-19 $X=2.185 $Y=0.82
c76 7 0 1.92338e-19 $X=2.375 $Y=1.41
c77 1 0 1.63932e-19 $X=0.965 $Y=1.41
r78 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r79 23 28 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=1.015 $Y=1.19
+ $X2=1.015 $Y2=1.16
r80 22 28 7.72467 $w=4.78e-07 $l=3.1e-07 $layer=LI1_cond $X=1.015 $Y=0.85
+ $X2=1.015 $Y2=1.16
r81 22 30 0.747549 $w=4.78e-07 $l=3e-08 $layer=LI1_cond $X=1.015 $Y=0.85
+ $X2=1.015 $Y2=0.82
r82 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.35
+ $Y=1.16 $X2=2.35 $Y2=1.16
r83 16 19 1.21796 $w=1.85e-07 $l=1e-07 $layer=LI1_cond $X=2.277 $Y=1.075
+ $X2=2.277 $Y2=1.175
r84 15 16 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=2.277 $Y=0.905
+ $X2=2.277 $Y2=1.075
r85 14 30 6.90116 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=1.255 $Y=0.82
+ $X2=1.015 $Y2=0.82
r86 13 15 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=2.185 $Y=0.82
+ $X2=2.277 $Y2=0.905
r87 13 14 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.185 $Y=0.82
+ $X2=1.255 $Y2=0.82
r88 10 20 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.375 $Y2=1.16
r89 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995 $X2=2.4
+ $Y2=0.56
r90 7 20 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.16
r91 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r92 4 27 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.965 $Y2=1.16
r93 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r94 1 27 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r95 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%A1 3 5 7 8 10 13 15 22
c43 15 0 3.5627e-19 $X=1.61 $Y=1.19
r44 22 23 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r45 20 22 34.2249 $w=3.38e-07 $l=2.4e-07 $layer=POLY_cond $X=1.665 $Y=1.217
+ $X2=1.905 $Y2=1.217
r46 18 20 32.7988 $w=3.38e-07 $l=2.3e-07 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.665 $Y2=1.217
r47 17 18 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.217
+ $X2=1.435 $Y2=1.217
r48 15 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.665
+ $Y=1.16 $X2=1.665 $Y2=1.16
r49 11 23 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r50 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r51 8 22 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r52 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r53 5 18 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r54 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r55 1 17 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.217
r56 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%B1 1 3 4 6 7 9 10 12 13 18 21 23 24 29
r66 24 29 3.19945 $w=2.4e-07 $l=1.05e-07 $layer=LI1_cond $X=4.335 $Y=1.18
+ $X2=4.335 $Y2=1.075
r67 23 29 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=4.335 $Y=0.85
+ $X2=4.335 $Y2=1.075
r68 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.16 $X2=4.14 $Y2=1.16
r69 18 24 3.65652 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=4.215 $Y=1.18
+ $X2=4.335 $Y2=1.18
r70 18 20 3.96104 $w=2.08e-07 $l=7.5e-08 $layer=LI1_cond $X=4.215 $Y=1.18
+ $X2=4.14 $Y2=1.18
r71 16 17 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=3.88 $Y=1.202
+ $X2=3.905 $Y2=1.202
r72 15 16 56.7434 $w=3.78e-07 $l=4.45e-07 $layer=POLY_cond $X=3.435 $Y=1.202
+ $X2=3.88 $Y2=1.202
r73 14 15 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=3.41 $Y=1.202
+ $X2=3.435 $Y2=1.202
r74 13 21 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=4.005 $Y=1.16
+ $X2=4.14 $Y2=1.16
r75 13 17 16.7575 $w=3.78e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.005 $Y=1.16
+ $X2=3.905 $Y2=1.202
r76 10 17 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.905 $Y=1.41
+ $X2=3.905 $Y2=1.202
r77 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.905 $Y=1.41
+ $X2=3.905 $Y2=1.985
r78 7 16 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=1.202
r79 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.88 $Y=0.995 $X2=3.88
+ $Y2=0.56
r80 4 15 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.202
r81 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.985
r82 1 14 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.202
r83 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995 $X2=3.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%A_297_47# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 38 42 45 48 50 52 57 60 64 65 78
c152 65 0 1.90952e-19 $X=3.645 $Y=1.54
r153 78 79 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=6.305 $Y=1.202
+ $X2=6.33 $Y2=1.202
r154 75 76 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=5.835 $Y=1.202
+ $X2=5.86 $Y2=1.202
r155 74 75 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=5.39 $Y=1.202
+ $X2=5.835 $Y2=1.202
r156 73 74 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=5.365 $Y=1.202
+ $X2=5.39 $Y2=1.202
r157 72 73 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=4.92 $Y=1.202
+ $X2=5.365 $Y2=1.202
r158 71 72 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.895 $Y=1.202
+ $X2=4.92 $Y2=1.202
r159 60 62 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.685 $Y=0.48
+ $X2=2.685 $Y2=0.785
r160 58 78 31.8302 $w=3.71e-07 $l=2.45e-07 $layer=POLY_cond $X=6.06 $Y=1.202
+ $X2=6.305 $Y2=1.202
r161 58 76 25.9838 $w=3.71e-07 $l=2e-07 $layer=POLY_cond $X=6.06 $Y=1.202
+ $X2=5.86 $Y2=1.202
r162 57 58 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.06
+ $Y=1.16 $X2=6.06 $Y2=1.16
r163 55 71 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=4.89 $Y=1.202
+ $X2=4.895 $Y2=1.202
r164 54 57 40.8593 $w=3.28e-07 $l=1.17e-06 $layer=LI1_cond $X=4.89 $Y=1.16
+ $X2=6.06 $Y2=1.16
r165 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.89
+ $Y=1.16 $X2=4.89 $Y2=1.16
r166 52 68 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=4.735 $Y=1.16
+ $X2=4.735 $Y2=1.54
r167 52 54 2.44458 $w=3.28e-07 $l=7e-08 $layer=LI1_cond $X=4.82 $Y=1.16 $X2=4.89
+ $Y2=1.16
r168 51 65 3.57226 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.835 $Y=1.54
+ $X2=3.645 $Y2=1.54
r169 50 68 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=1.54
+ $X2=4.735 $Y2=1.54
r170 50 51 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=4.65 $Y=1.54
+ $X2=3.835 $Y2=1.54
r171 46 65 3.05675 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=1.625
+ $X2=3.645 $Y2=1.54
r172 46 48 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=3.645 $Y=1.625
+ $X2=3.645 $Y2=1.63
r173 45 65 3.05675 $w=3.1e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.575 $Y=1.455
+ $X2=3.645 $Y2=1.54
r174 44 64 3.05675 $w=3.1e-07 $l=2.22036e-07 $layer=LI1_cond $X=3.575 $Y=0.87
+ $X2=3.455 $Y2=0.7
r175 44 45 28.0908 $w=2.38e-07 $l=5.85e-07 $layer=LI1_cond $X=3.575 $Y=0.87
+ $X2=3.575 $Y2=1.455
r176 40 64 3.05675 $w=3.1e-07 $l=1.9e-07 $layer=LI1_cond $X=3.645 $Y=0.7
+ $X2=3.455 $Y2=0.7
r177 40 42 9.70478 $w=3.78e-07 $l=3.2e-07 $layer=LI1_cond $X=3.645 $Y=0.7
+ $X2=3.645 $Y2=0.38
r178 39 62 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.77 $Y=0.785
+ $X2=2.685 $Y2=0.785
r179 38 64 3.57226 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.455 $Y=0.785
+ $X2=3.455 $Y2=0.7
r180 38 39 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.455 $Y=0.785
+ $X2=2.77 $Y2=0.785
r181 34 60 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=0.48
+ $X2=2.685 $Y2=0.48
r182 34 36 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=2.6 $Y=0.48
+ $X2=1.67 $Y2=0.48
r183 31 79 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.33 $Y=0.995
+ $X2=6.33 $Y2=1.202
r184 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.33 $Y=0.995
+ $X2=6.33 $Y2=0.56
r185 28 78 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.305 $Y=1.41
+ $X2=6.305 $Y2=1.202
r186 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.305 $Y=1.41
+ $X2=6.305 $Y2=1.985
r187 25 76 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.86 $Y=0.995
+ $X2=5.86 $Y2=1.202
r188 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.86 $Y=0.995
+ $X2=5.86 $Y2=0.56
r189 22 75 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.835 $Y=1.41
+ $X2=5.835 $Y2=1.202
r190 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.835 $Y=1.41
+ $X2=5.835 $Y2=1.985
r191 19 74 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.39 $Y=0.995
+ $X2=5.39 $Y2=1.202
r192 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.39 $Y=0.995
+ $X2=5.39 $Y2=0.56
r193 16 73 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.202
r194 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.985
r195 13 72 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.92 $Y=0.995
+ $X2=4.92 $Y2=1.202
r196 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.92 $Y=0.995
+ $X2=4.92 $Y2=0.56
r197 10 71 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.895 $Y=1.41
+ $X2=4.895 $Y2=1.202
r198 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.895 $Y=1.41
+ $X2=4.895 $Y2=1.985
r199 3 48 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.525
+ $Y=1.485 $X2=3.67 $Y2=1.63
r200 2 42 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.485
+ $Y=0.235 $X2=3.67 $Y2=0.38
r201 1 36 182 $w=1.7e-07 $l=3.24577e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.48
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%A_27_297# 1 2 3 4 5 18 22 26 28 29 30 31 34
+ 37 39 41
c65 28 0 4.1943e-20 $X=3.2 $Y=1.955
r66 32 34 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=4.14 $Y=2.295
+ $X2=4.14 $Y2=1.96
r67 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.055 $Y=2.38
+ $X2=4.14 $Y2=2.295
r68 30 31 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.055 $Y=2.38
+ $X2=3.285 $Y2=2.38
r69 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.2 $Y=2.295
+ $X2=3.285 $Y2=2.38
r70 28 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=1.955 $X2=3.2
+ $Y2=1.87
r71 28 29 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=3.2 $Y=1.955 $X2=3.2
+ $Y2=2.295
r72 27 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.87
+ $X2=2.14 $Y2=1.87
r73 26 43 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=1.87 $X2=3.2
+ $Y2=1.87
r74 26 27 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.115 $Y=1.87
+ $X2=2.225 $Y2=1.87
r75 23 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.87 $X2=1.2
+ $Y2=1.87
r76 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=1.87
+ $X2=2.14 $Y2=1.87
r77 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=1.87
+ $X2=1.285 $Y2=1.87
r78 19 37 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.26 $Y2=1.87
r79 18 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.87 $X2=1.2
+ $Y2=1.87
r80 18 19 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=1.87
+ $X2=0.345 $Y2=1.87
r81 5 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.995
+ $Y=1.485 $X2=4.14 $Y2=1.96
r82 4 43 300 $w=1.7e-07 $l=5.58167e-07 $layer=licon1_PDIFF $count=2 $X=2.995
+ $Y=1.485 $X2=3.2 $Y2=1.95
r83 3 41 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.95
r84 2 39 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.95
r85 1 37 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 44 45
+ 47 48 49 51 56 61 76 81 84 87 91
r120 90 91 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r124 79 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r125 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r126 76 90 5.01588 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=6.325 $Y=2.72
+ $X2=6.612 $Y2=2.72
r127 76 78 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.325 $Y=2.72
+ $X2=6.21 $Y2=2.72
r128 75 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r129 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r130 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r131 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 69 72 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 69 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 68 71 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r135 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r136 66 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.585 $Y2=2.72
r137 66 68 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r138 65 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r139 65 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r140 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 62 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r142 62 64 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 61 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.585 $Y2=2.72
r144 61 64 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 60 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r146 60 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 57 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r149 57 59 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r150 56 84 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r151 56 59 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r152 51 81 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r153 51 53 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r154 49 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 49 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r156 47 74 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.29 $Y2=2.72
r157 47 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.575 $Y2=2.72
r158 46 78 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=6.21 $Y2=2.72
r159 46 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.575 $Y2=2.72
r160 44 71 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.495 $Y=2.72
+ $X2=4.37 $Y2=2.72
r161 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.495 $Y=2.72
+ $X2=4.66 $Y2=2.72
r162 43 74 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=5.29 $Y2=2.72
r163 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.66 $Y2=2.72
r164 39 90 3.1808 $w=3.8e-07 $l=1.32868e-07 $layer=LI1_cond $X=6.515 $Y=2.635
+ $X2=6.612 $Y2=2.72
r165 39 41 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=6.515 $Y=2.635
+ $X2=6.515 $Y2=2.21
r166 35 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=2.635
+ $X2=5.575 $Y2=2.72
r167 35 37 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=5.575 $Y=2.635
+ $X2=5.575 $Y2=2.21
r168 31 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.66 $Y=2.635
+ $X2=4.66 $Y2=2.72
r169 31 33 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=4.66 $Y=2.635
+ $X2=4.66 $Y2=2.21
r170 27 87 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.72
r171 27 29 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=2.585 $Y=2.635
+ $X2=2.585 $Y2=2.21
r172 23 84 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.72
r173 23 25 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=1.645 $Y=2.635
+ $X2=1.645 $Y2=2.21
r174 19 81 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r175 19 21 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.21
r176 6 41 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=6.395
+ $Y=1.485 $X2=6.54 $Y2=2.21
r177 5 37 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=1.485 $X2=5.6 $Y2=2.21
r178 4 33 600 $w=1.7e-07 $l=7.85016e-07 $layer=licon1_PDIFF $count=1 $X=4.535
+ $Y=1.485 $X2=4.66 $Y2=2.21
r179 3 29 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.21
r180 2 25 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.21
r181 1 21 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%X 1 2 3 4 15 20 23 24 25 26 27 36 39
r57 48 51 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.13 $Y=0.74
+ $X2=6.07 $Y2=0.74
r58 36 39 1.42191 $w=1.93e-07 $l=2.5e-08 $layer=LI1_cond $X=6.682 $Y=0.825
+ $X2=6.682 $Y2=0.85
r59 26 27 10.5363 $w=3.63e-07 $l=2.55e-07 $layer=LI1_cond $X=6.682 $Y=1.53
+ $X2=6.682 $Y2=1.785
r60 25 26 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=6.682 $Y=1.19
+ $X2=6.682 $Y2=1.53
r61 24 36 3.20299 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=6.682 $Y=0.74
+ $X2=6.682 $Y2=0.825
r62 24 51 26.6124 $w=2.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.585 $Y=0.74
+ $X2=6.07 $Y2=0.74
r63 24 25 17.6317 $w=1.93e-07 $l=3.1e-07 $layer=LI1_cond $X=6.682 $Y=0.88
+ $X2=6.682 $Y2=1.19
r64 24 39 1.70629 $w=1.93e-07 $l=3e-08 $layer=LI1_cond $X=6.682 $Y=0.88
+ $X2=6.682 $Y2=0.85
r65 21 27 16.0146 $w=3.38e-07 $l=4.3e-07 $layer=LI1_cond $X=6.155 $Y=1.87
+ $X2=6.585 $Y2=1.87
r66 21 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=1.87
+ $X2=6.07 $Y2=1.87
r67 16 20 3.40825 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=5.215 $Y=1.87
+ $X2=5.075 $Y2=1.87
r68 15 23 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=1.87
+ $X2=6.07 $Y2=1.87
r69 15 16 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.985 $Y=1.87
+ $X2=5.215 $Y2=1.87
r70 4 23 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=5.925
+ $Y=1.485 $X2=6.07 $Y2=1.95
r71 3 20 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=4.985
+ $Y=1.485 $X2=5.13 $Y2=1.95
r72 2 51 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.235 $X2=6.07 $Y2=0.74
r73 1 48 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=4.995
+ $Y=0.235 $X2=5.13 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_4%VGND 1 2 3 4 5 16 18 22 26 28 30 33 34 35
+ 37 42 51 59 63 70
r94 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r95 63 66 9.02701 $w=5.28e-07 $l=4e-07 $layer=LI1_cond $X=4.4 $Y=0 $X2=4.4
+ $Y2=0.4
r96 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r97 59 60 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r98 54 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r99 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r100 51 69 5.01588 $w=1.7e-07 $l=2.87e-07 $layer=LI1_cond $X=6.325 $Y=0
+ $X2=6.612 $Y2=0
r101 51 53 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.325 $Y=0
+ $X2=6.21 $Y2=0
r102 50 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r103 50 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r104 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r105 47 63 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=4.665 $Y=0 $X2=4.4
+ $Y2=0
r106 47 49 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.665 $Y=0
+ $X2=5.29 $Y2=0
r107 46 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r108 46 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r109 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r110 43 59 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.117 $Y2=0
r111 43 45 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.91 $Y2=0
r112 42 63 7.52407 $w=1.7e-07 $l=2.65e-07 $layer=LI1_cond $X=4.135 $Y=0 $X2=4.4
+ $Y2=0
r113 42 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=4.135 $Y=0
+ $X2=3.91 $Y2=0
r114 41 60 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.99
+ $Y2=0
r115 40 41 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 38 56 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r117 38 40 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r118 37 59 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=3.117
+ $Y2=0
r119 37 40 147.444 $w=1.68e-07 $l=2.26e-06 $layer=LI1_cond $X=2.95 $Y=0 $X2=0.69
+ $Y2=0
r120 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r121 35 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r122 33 49 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.29
+ $Y2=0
r123 33 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.385 $Y=0 $X2=5.575
+ $Y2=0
r124 32 53 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=5.765 $Y=0
+ $X2=6.21 $Y2=0
r125 32 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.765 $Y=0 $X2=5.575
+ $Y2=0
r126 28 69 3.1808 $w=3.8e-07 $l=1.32868e-07 $layer=LI1_cond $X=6.515 $Y=0.085
+ $X2=6.612 $Y2=0
r127 28 30 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=6.515 $Y=0.085
+ $X2=6.515 $Y2=0.4
r128 24 34 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0
r129 24 26 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=5.575 $Y=0.085
+ $X2=5.575 $Y2=0.4
r130 20 59 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=3.117 $Y=0.085
+ $X2=3.117 $Y2=0
r131 20 22 9.63236 $w=3.33e-07 $l=2.8e-07 $layer=LI1_cond $X=3.117 $Y=0.085
+ $X2=3.117 $Y2=0.365
r132 16 56 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r133 16 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r134 5 30 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=6.405
+ $Y=0.235 $X2=6.54 $Y2=0.4
r135 4 26 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.235 $X2=5.6 $Y2=0.4
r136 3 66 91 $w=1.7e-07 $l=7.02673e-07 $layer=licon1_NDIFF $count=2 $X=3.955
+ $Y=0.235 $X2=4.58 $Y2=0.4
r137 2 22 182 $w=1.7e-07 $l=2.82622e-07 $layer=licon1_NDIFF $count=1 $X=2.955
+ $Y=0.235 $X2=3.18 $Y2=0.365
r138 1 18 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

