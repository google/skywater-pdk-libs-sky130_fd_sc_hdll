* File: sky130_fd_sc_hdll__a21oi_4.pex.spice
* Created: Thu Aug 27 18:53:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 30 31 40 43 46
c75 22 0 6.06305e-20 $X=1.965 $Y=0.995
c76 4 0 3.22468e-20 $X=0.5 $Y=1.41
r77 43 44 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.94 $Y=1.202
+ $X2=1.965 $Y2=1.202
r78 42 43 60.0849 $w=3.65e-07 $l=4.55e-07 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.94 $Y2=1.202
r79 41 42 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.485 $Y2=1.202
r80 39 41 12.5452 $w=3.65e-07 $l=9.5e-08 $layer=POLY_cond $X=1.365 $Y=1.202
+ $X2=1.46 $Y2=1.202
r81 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.365
+ $Y=1.16 $X2=1.365 $Y2=1.16
r82 37 39 47.5397 $w=3.65e-07 $l=3.6e-07 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.365 $Y2=1.202
r83 36 37 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.005 $Y2=1.202
r84 35 36 63.3863 $w=3.65e-07 $l=4.8e-07 $layer=POLY_cond $X=0.5 $Y=1.202
+ $X2=0.98 $Y2=1.202
r85 34 35 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.475 $Y=1.202
+ $X2=0.5 $Y2=1.202
r86 31 40 6.21713 $w=3.78e-07 $l=2.05e-07 $layer=LI1_cond $X=1.16 $Y=1.225
+ $X2=1.365 $Y2=1.225
r87 31 46 0.151637 $w=3.78e-07 $l=5e-09 $layer=LI1_cond $X=1.16 $Y=1.225
+ $X2=1.155 $Y2=1.225
r88 30 46 22.8972 $w=3.78e-07 $l=7.55e-07 $layer=LI1_cond $X=0.4 $Y=1.225
+ $X2=1.155 $Y2=1.225
r89 28 34 30.3726 $w=3.65e-07 $l=2.3e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.475 $Y2=1.202
r90 27 30 4.3816 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.245 $Y=1.205
+ $X2=0.4 $Y2=1.205
r91 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r92 22 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.965 $Y2=1.202
r93 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.965 $Y=0.995
+ $X2=1.965 $Y2=0.56
r94 19 43 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.202
r95 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.985
r96 16 42 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=1.202
r97 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=0.56
r98 13 41 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.202
r99 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.985
r100 10 37 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r101 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r102 7 36 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r104 4 35 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.202
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
r106 1 34 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r107 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 31 32 33 34 48 51 54
c128 31 0 3.14505e-20 $X=2.645 $Y=1.592
r129 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.855
+ $Y=1.16 $X2=5.855 $Y2=1.16
r130 48 50 4.57182 $w=3.69e-07 $l=3.5e-08 $layer=POLY_cond $X=5.82 $Y=1.202
+ $X2=5.855 $Y2=1.202
r131 47 48 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.795 $Y=1.202
+ $X2=5.82 $Y2=1.202
r132 46 54 3.22751 $w=6.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.465 $Y=1.39
+ $X2=5.295 $Y2=1.39
r133 45 47 43.1057 $w=3.69e-07 $l=3.3e-07 $layer=POLY_cond $X=5.465 $Y=1.202
+ $X2=5.795 $Y2=1.202
r134 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=1.16 $X2=5.465 $Y2=1.16
r135 43 45 16.3279 $w=3.69e-07 $l=1.25e-07 $layer=POLY_cond $X=5.34 $Y=1.202
+ $X2=5.465 $Y2=1.202
r136 42 43 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.315 $Y=1.202
+ $X2=5.34 $Y2=1.202
r137 41 54 3.22751 $w=6.28e-07 $l=1.7e-07 $layer=LI1_cond $X=5.125 $Y=1.39
+ $X2=5.295 $Y2=1.39
r138 40 42 24.8184 $w=3.69e-07 $l=1.9e-07 $layer=POLY_cond $X=5.125 $Y=1.202
+ $X2=5.315 $Y2=1.202
r139 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.125
+ $Y=1.16 $X2=5.125 $Y2=1.16
r140 38 40 34.6152 $w=3.69e-07 $l=2.65e-07 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=5.125 $Y2=1.202
r141 37 38 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.835 $Y=1.202
+ $X2=4.86 $Y2=1.202
r142 34 51 1.80361 $w=6.28e-07 $l=9.5e-08 $layer=LI1_cond $X=5.76 $Y=1.39
+ $X2=5.855 $Y2=1.39
r143 34 46 5.60068 $w=6.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.76 $Y=1.39
+ $X2=5.465 $Y2=1.39
r144 32 41 2.56303 $w=6.28e-07 $l=1.35e-07 $layer=LI1_cond $X=4.99 $Y=1.39
+ $X2=5.125 $Y2=1.39
r145 32 33 11.207 $w=6.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.99 $Y=1.39
+ $X2=4.675 $Y2=1.39
r146 31 33 103.976 $w=2.23e-07 $l=2.03e-06 $layer=LI1_cond $X=2.645 $Y=1.592
+ $X2=4.675 $Y2=1.592
r147 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.415
+ $Y=1.16 $X2=2.415 $Y2=1.16
r148 25 31 7.50513 $w=2.25e-07 $l=2.4775e-07 $layer=LI1_cond $X=2.447 $Y=1.48
+ $X2=2.645 $Y2=1.592
r149 25 27 9.33625 $w=3.93e-07 $l=3.2e-07 $layer=LI1_cond $X=2.447 $Y=1.48
+ $X2=2.447 $Y2=1.16
r150 22 48 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.202
r151 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.985
r152 19 47 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=1.202
r153 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=0.56
r154 16 43 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.202
r155 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.34 $Y=1.41
+ $X2=5.34 $Y2=1.985
r156 13 42 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.315 $Y=0.995
+ $X2=5.315 $Y2=1.202
r157 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.315 $Y=0.995
+ $X2=5.315 $Y2=0.56
r158 10 38 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.202
r159 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.985
r160 7 37 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=1.202
r161 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.835 $Y=0.995
+ $X2=4.835 $Y2=0.56
r162 4 28 45.964 $w=3.43e-07 $l=2.54951e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.44 $Y2=1.16
r163 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.45 $Y2=1.985
r164 1 28 38.7084 $w=3.43e-07 $l=1.67481e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.44 $Y2=1.16
r165 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.435 $Y=0.995
+ $X2=2.435 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 44 45 52
c71 22 0 9.39532e-20 $X=4.405 $Y=0.99
r72 45 46 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=4.38 $Y=1.2
+ $X2=4.405 $Y2=1.2
r73 43 45 22.0305 $w=3.61e-07 $l=1.65e-07 $layer=POLY_cond $X=4.215 $Y=1.2
+ $X2=4.38 $Y2=1.2
r74 43 44 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.215
+ $Y=1.16 $X2=4.215 $Y2=1.16
r75 41 43 42.0582 $w=3.61e-07 $l=3.15e-07 $layer=POLY_cond $X=3.9 $Y=1.2
+ $X2=4.215 $Y2=1.2
r76 40 41 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=3.875 $Y=1.2
+ $X2=3.9 $Y2=1.2
r77 39 52 4.23346 $w=2.43e-07 $l=9e-08 $layer=LI1_cond $X=3.825 $Y=1.187
+ $X2=3.915 $Y2=1.187
r78 38 40 6.6759 $w=3.61e-07 $l=5e-08 $layer=POLY_cond $X=3.825 $Y=1.2 $X2=3.875
+ $Y2=1.2
r79 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.825
+ $Y=1.16 $X2=3.825 $Y2=1.16
r80 36 39 18.345 $w=2.43e-07 $l=3.9e-07 $layer=LI1_cond $X=3.435 $Y=1.187
+ $X2=3.825 $Y2=1.187
r81 35 38 52.072 $w=3.61e-07 $l=3.9e-07 $layer=POLY_cond $X=3.435 $Y=1.2
+ $X2=3.825 $Y2=1.2
r82 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.435
+ $Y=1.16 $X2=3.435 $Y2=1.16
r83 33 35 2.00277 $w=3.61e-07 $l=1.5e-08 $layer=POLY_cond $X=3.42 $Y=1.2
+ $X2=3.435 $Y2=1.2
r84 32 33 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=3.395 $Y=1.2
+ $X2=3.42 $Y2=1.2
r85 31 36 18.345 $w=2.43e-07 $l=3.9e-07 $layer=LI1_cond $X=3.045 $Y=1.187
+ $X2=3.435 $Y2=1.187
r86 30 32 46.7313 $w=3.61e-07 $l=3.5e-07 $layer=POLY_cond $X=3.045 $Y=1.2
+ $X2=3.395 $Y2=1.2
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.045
+ $Y=1.16 $X2=3.045 $Y2=1.16
r88 28 30 14.0194 $w=3.61e-07 $l=1.05e-07 $layer=POLY_cond $X=2.94 $Y=1.2
+ $X2=3.045 $Y2=1.2
r89 27 28 3.33795 $w=3.61e-07 $l=2.5e-08 $layer=POLY_cond $X=2.915 $Y=1.2
+ $X2=2.94 $Y2=1.2
r90 25 44 13.6412 $w=2.43e-07 $l=2.9e-07 $layer=LI1_cond $X=3.925 $Y=1.187
+ $X2=4.215 $Y2=1.187
r91 25 52 0.470385 $w=2.43e-07 $l=1e-08 $layer=LI1_cond $X=3.925 $Y=1.187
+ $X2=3.915 $Y2=1.187
r92 22 46 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.405 $Y=0.99
+ $X2=4.405 $Y2=1.2
r93 22 24 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.405 $Y=0.99
+ $X2=4.405 $Y2=0.56
r94 19 45 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.38 $Y=1.41
+ $X2=4.38 $Y2=1.2
r95 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.38 $Y=1.41
+ $X2=4.38 $Y2=1.985
r96 16 41 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.9 $Y=1.41 $X2=3.9
+ $Y2=1.2
r97 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.9 $Y=1.41 $X2=3.9
+ $Y2=1.985
r98 13 40 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.875 $Y=0.99
+ $X2=3.875 $Y2=1.2
r99 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.875 $Y=0.99
+ $X2=3.875 $Y2=0.56
r100 10 33 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.2
r101 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.985
r102 7 32 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.395 $Y=0.99
+ $X2=3.395 $Y2=1.2
r103 7 9 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.395 $Y=0.99
+ $X2=3.395 $Y2=0.56
r104 4 28 19.0337 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.94 $Y2=1.2
r105 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.94 $Y2=1.985
r106 1 27 23.3725 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.915 $Y=0.99
+ $X2=2.915 $Y2=1.2
r107 1 3 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.915 $Y=0.99
+ $X2=2.915 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%A_28_297# 1 2 3 4 5 6 7 22 24 26 28 29 32
+ 34 38 40 44 46 48 50 59 61 62
c83 29 0 3.22468e-20 $X=2.315 $Y=1.99
r84 55 57 38.9613 $w=3.1e-07 $l=9.9e-07 $layer=LI1_cond $X=1.22 $Y=2.205
+ $X2=2.21 $Y2=2.205
r85 48 64 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=6.095 $Y=2.105
+ $X2=6.095 $Y2=1.99
r86 48 50 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=6.095 $Y=2.105
+ $X2=6.095 $Y2=2.3
r87 47 62 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.185 $Y=1.99 $X2=5.095
+ $Y2=1.99
r88 46 64 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=5.965 $Y=1.99
+ $X2=6.095 $Y2=1.99
r89 46 47 39.0829 $w=2.28e-07 $l=7.8e-07 $layer=LI1_cond $X=5.965 $Y=1.99
+ $X2=5.185 $Y2=1.99
r90 42 62 2.23839 $w=1.8e-07 $l=1.15e-07 $layer=LI1_cond $X=5.095 $Y=2.105
+ $X2=5.095 $Y2=1.99
r91 42 44 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=5.095 $Y=2.105
+ $X2=5.095 $Y2=2.3
r92 41 61 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.235 $Y=1.99
+ $X2=4.14 $Y2=1.99
r93 40 62 4.19361 $w=2.3e-07 $l=9e-08 $layer=LI1_cond $X=5.005 $Y=1.99 $X2=5.095
+ $Y2=1.99
r94 40 41 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=5.005 $Y=1.99
+ $X2=4.235 $Y2=1.99
r95 36 61 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=4.14 $Y=2.105
+ $X2=4.14 $Y2=1.99
r96 36 38 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=4.14 $Y=2.105
+ $X2=4.14 $Y2=2.3
r97 35 59 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.275 $Y=1.99
+ $X2=3.18 $Y2=1.99
r98 34 61 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=4.045 $Y=1.99
+ $X2=4.14 $Y2=1.99
r99 34 35 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=4.045 $Y=1.99
+ $X2=3.275 $Y2=1.99
r100 30 59 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.18 $Y=2.105
+ $X2=3.18 $Y2=1.99
r101 30 32 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.18 $Y=2.105
+ $X2=3.18 $Y2=2.3
r102 29 57 4.97025 $w=3.1e-07 $l=2.62298e-07 $layer=LI1_cond $X=2.315 $Y=1.99
+ $X2=2.21 $Y2=2.205
r103 28 59 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.085 $Y=1.99
+ $X2=3.18 $Y2=1.99
r104 28 29 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.085 $Y=1.99
+ $X2=2.315 $Y2=1.99
r105 27 53 3.05549 $w=2.5e-07 $l=9.8e-08 $layer=LI1_cond $X=0.375 $Y=2.34
+ $X2=0.277 $Y2=2.34
r106 26 55 8.95388 $w=3.1e-07 $l=2.74317e-07 $layer=LI1_cond $X=1.005 $Y=2.34
+ $X2=1.22 $Y2=2.205
r107 26 27 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=1.005 $Y=2.34
+ $X2=0.375 $Y2=2.34
r108 22 53 3.89731 $w=1.95e-07 $l=1.25e-07 $layer=LI1_cond $X=0.277 $Y=2.215
+ $X2=0.277 $Y2=2.34
r109 22 24 14.5035 $w=1.93e-07 $l=2.55e-07 $layer=LI1_cond $X=0.277 $Y=2.215
+ $X2=0.277 $Y2=1.96
r110 7 64 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.485 $X2=6.06 $Y2=1.96
r111 7 50 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.91
+ $Y=1.485 $X2=6.06 $Y2=2.3
r112 6 44 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=4.95
+ $Y=1.485 $X2=5.1 $Y2=2.3
r113 5 61 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.485 $X2=4.14 $Y2=1.96
r114 5 38 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=3.99
+ $Y=1.485 $X2=4.14 $Y2=2.3
r115 4 59 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.485 $X2=3.18 $Y2=1.96
r116 4 32 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.485 $X2=3.18 $Y2=2.3
r117 3 57 600 $w=1.7e-07 $l=9.00514e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.485 $X2=2.21 $Y2=2.3
r118 2 55 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.485 $X2=1.22 $Y2=2.36
r119 1 53 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.3
r120 1 24 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%Y 1 2 3 4 5 6 19 23 26 29 33 36 41 42 43
+ 44 50
c80 41 0 1.1531e-19 $X=1.7 $Y=0.76
c81 33 0 9.39532e-20 $X=4.14 $Y=0.76
c82 29 0 3.99762e-19 $X=2.585 $Y=0.785
r83 47 50 23.2571 $w=4.48e-07 $l=8.75e-07 $layer=LI1_cond $X=0.74 $Y=1.81
+ $X2=1.615 $Y2=1.81
r84 44 50 0.132898 $w=4.48e-07 $l=5e-09 $layer=LI1_cond $X=1.62 $Y=1.81
+ $X2=1.615 $Y2=1.81
r85 42 44 3.45534 $w=4.48e-07 $l=1.3e-07 $layer=LI1_cond $X=1.75 $Y=1.81
+ $X2=1.62 $Y2=1.81
r86 31 33 50.2884 $w=2.18e-07 $l=9.6e-07 $layer=LI1_cond $X=3.18 $Y=0.785
+ $X2=4.14 $Y2=0.785
r87 29 43 5.8804 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=2.585 $Y=0.785
+ $X2=2.475 $Y2=0.785
r88 29 31 31.1683 $w=2.18e-07 $l=5.95e-07 $layer=LI1_cond $X=2.585 $Y=0.785
+ $X2=3.18 $Y2=0.785
r89 28 41 3.50213 $w=2e-07 $l=5.57786e-07 $layer=LI1_cond $X=2.08 $Y=0.795
+ $X2=1.605 $Y2=0.615
r90 28 43 21.9045 $w=1.98e-07 $l=3.95e-07 $layer=LI1_cond $X=2.08 $Y=0.795
+ $X2=2.475 $Y2=0.795
r91 26 42 8.75241 $w=3.13e-07 $l=2.96226e-07 $layer=LI1_cond $X=1.915 $Y=1.585
+ $X2=1.75 $Y2=1.81
r92 25 41 2.62102 $w=3.3e-07 $l=4.27668e-07 $layer=LI1_cond $X=1.915 $Y=0.895
+ $X2=1.605 $Y2=0.615
r93 25 26 24.0965 $w=3.28e-07 $l=6.9e-07 $layer=LI1_cond $X=1.915 $Y=0.895
+ $X2=1.915 $Y2=1.585
r94 21 41 2.62102 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.7 $Y=0.615
+ $X2=1.605 $Y2=0.615
r95 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=1.7 $Y=0.615
+ $X2=1.7 $Y2=0.42
r96 20 36 11.9665 $w=1.88e-07 $l=2.05e-07 $layer=LI1_cond $X=0.74 $Y=0.74
+ $X2=0.74 $Y2=0.535
r97 19 41 3.50213 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.605 $Y=0.74
+ $X2=1.605 $Y2=0.615
r98 19 20 35.4952 $w=2.48e-07 $l=7.7e-07 $layer=LI1_cond $X=1.605 $Y=0.74
+ $X2=0.835 $Y2=0.74
r99 6 44 600 $w=1.7e-07 $l=4.74104e-07 $layer=licon1_PDIFF $count=1 $X=1.55
+ $Y=1.485 $X2=1.7 $Y2=1.89
r100 5 47 600 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.85
r101 4 33 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.14 $Y2=0.76
r102 3 31 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.235 $X2=3.18 $Y2=0.76
r103 2 41 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.76
r104 2 23 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.42
r105 1 36 182 $w=1.7e-07 $l=3.83406e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.74 $Y2=0.535
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%VPWR 1 2 3 4 13 16 19 23 26 29 31 44 45 48
+ 55
r100 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r101 55 58 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.635 $Y=2.36
+ $X2=3.635 $Y2=2.72
r102 52 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r103 51 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r104 48 51 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.675 $Y=2.36
+ $X2=2.675 $Y2=2.72
r105 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r106 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r107 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r108 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r109 39 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.45 $Y2=2.72
r110 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r111 36 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.635 $Y2=2.72
r112 36 38 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=4.37 $Y2=2.72
r113 31 51 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.675 $Y2=2.72
r114 31 33 147.118 $w=1.68e-07 $l=2.255e-06 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=0.23 $Y2=2.72
r115 29 52 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r116 29 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r117 27 44 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.745 $Y=2.72
+ $X2=6.21 $Y2=2.72
r118 26 41 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.365 $Y=2.72
+ $X2=5.29 $Y2=2.72
r119 25 27 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.555 $Y=2.72
+ $X2=5.745 $Y2=2.72
r120 25 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.555 $Y=2.72
+ $X2=5.365 $Y2=2.72
r121 23 25 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.555 $Y=2.36
+ $X2=5.555 $Y2=2.72
r122 20 41 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 19 38 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.37 $Y2=2.72
r124 18 20 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.785 $Y2=2.72
r125 18 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.595 $Y=2.72
+ $X2=4.405 $Y2=2.72
r126 16 18 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.595 $Y=2.36
+ $X2=4.595 $Y2=2.72
r127 14 51 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.675 $Y2=2.72
r128 13 58 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=3.635 $Y2=2.72
r129 13 14 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.445 $Y=2.72
+ $X2=2.865 $Y2=2.72
r130 4 23 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=5.43
+ $Y=1.485 $X2=5.58 $Y2=2.36
r131 3 16 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=4.47
+ $Y=1.485 $X2=4.62 $Y2=2.36
r132 2 55 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.485 $X2=3.66 $Y2=2.36
r133 1 48 600 $w=1.7e-07 $l=9.51643e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.485 $X2=2.7 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%VGND 1 2 3 4 5 16 18 22 26 28 30 33 34 35
+ 37 42 54 63 69 73
c97 33 0 1.51849e-19 $X=5.005 $Y=0
r98 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r99 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r100 63 66 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.195 $Y=0
+ $X2=1.195 $Y2=0.36
r101 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r102 57 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r103 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r104 54 72 3.98437 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=6.202 $Y2=0
r105 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.965 $Y=0
+ $X2=5.75 $Y2=0
r106 53 57 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r107 52 53 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r108 50 53 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r109 50 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r110 49 52 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r111 49 50 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r112 47 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.315 $Y=0 $X2=2.15
+ $Y2=0
r113 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.315 $Y=0
+ $X2=2.53 $Y2=0
r114 46 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r115 46 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r116 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r117 43 63 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.195
+ $Y2=0
r118 43 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.385 $Y=0
+ $X2=1.61 $Y2=0
r119 42 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.15
+ $Y2=0
r120 42 45 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.985 $Y=0
+ $X2=1.61 $Y2=0
r121 41 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r122 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 38 59 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r124 38 40 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r125 37 63 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.195
+ $Y2=0
r126 37 40 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=0
+ $X2=0.69 $Y2=0
r127 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r128 35 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r129 33 52 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.005 $Y=0
+ $X2=4.83 $Y2=0
r130 33 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.005 $Y=0 $X2=5.1
+ $Y2=0
r131 32 56 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.195 $Y=0
+ $X2=5.75 $Y2=0
r132 32 34 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=5.195 $Y=0 $X2=5.1
+ $Y2=0
r133 28 72 3.22785 $w=2.6e-07 $l=1.43332e-07 $layer=LI1_cond $X=6.095 $Y=0.085
+ $X2=6.202 $Y2=0
r134 28 30 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.095 $Y=0.085
+ $X2=6.095 $Y2=0.38
r135 24 34 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.1 $Y=0.085
+ $X2=5.1 $Y2=0
r136 24 26 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=5.1 $Y=0.085
+ $X2=5.1 $Y2=0.4
r137 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0
r138 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.15 $Y=0.085
+ $X2=2.15 $Y2=0.36
r139 16 59 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r140 16 18 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r141 5 30 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=5.87
+ $Y=0.235 $X2=6.06 $Y2=0.38
r142 4 26 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.235 $X2=5.1 $Y2=0.4
r143 3 22 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.22 $Y2=0.36
r144 2 66 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.36
r145 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_4%A_502_47# 1 2 3 4 13 19 22 23 24 27
c49 1 0 1.87282e-19 $X=2.51 $Y=0.235
r50 25 27 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=5.555 $Y=0.735
+ $X2=5.555 $Y2=0.395
r51 23 25 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.365 $Y=0.82
+ $X2=5.555 $Y2=0.735
r52 23 24 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=5.365 $Y=0.82
+ $X2=4.785 $Y2=0.82
r53 20 24 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.655 $Y=0.735
+ $X2=4.785 $Y2=0.82
r54 20 22 1.55137 $w=2.58e-07 $l=3.5e-08 $layer=LI1_cond $X=4.655 $Y=0.735
+ $X2=4.655 $Y2=0.7
r55 19 30 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=4.655 $Y=0.505
+ $X2=4.655 $Y2=0.38
r56 19 22 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=4.655 $Y=0.505
+ $X2=4.655 $Y2=0.7
r57 15 18 44.2538 $w=2.48e-07 $l=9.6e-07 $layer=LI1_cond $X=2.7 $Y=0.38 $X2=3.66
+ $Y2=0.38
r58 13 30 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=4.525 $Y=0.38
+ $X2=4.655 $Y2=0.38
r59 13 18 39.8745 $w=2.48e-07 $l=8.65e-07 $layer=LI1_cond $X=4.525 $Y=0.38
+ $X2=3.66 $Y2=0.38
r60 4 27 91 $w=1.7e-07 $l=2.57876e-07 $layer=licon1_NDIFF $count=2 $X=5.39
+ $Y=0.235 $X2=5.58 $Y2=0.395
r61 3 30 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.235 $X2=4.62 $Y2=0.36
r62 3 22 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=4.48
+ $Y=0.235 $X2=4.62 $Y2=0.7
r63 2 18 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.235 $X2=3.66 $Y2=0.42
r64 1 15 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.7 $Y2=0.42
.ends

