* File: sky130_fd_sc_hdll__xor3_2.spice
* Created: Thu Aug 27 19:30:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xor3_2.pex.spice"
.subckt sky130_fd_sc_hdll__xor3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 N_X_M1001_d N_A_81_21#_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.1755 PD=1 PS=1.84 NRD=12.912 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1016 N_X_M1001_d N_A_81_21#_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.175105 PD=1 PS=1.36075 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75000.7 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1008 N_A_335_93#_M1008_d N_C_M1008_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1974 AS=0.113145 PD=1.78 PS=0.879252 NRD=52.848 NRS=61.248 M=1 R=2.8
+ SA=75001.3 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_81_21#_M1002_d N_C_M1002_g N_A_483_49#_M1002_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1424 AS=0.208 PD=1.085 PS=1.93 NRD=0 NRS=9.372 M=1 R=4.26667
+ SA=75000.2 SB=75001 A=0.096 P=1.58 MULT=1
MM1019 N_A_465_325#_M1019_d N_A_335_93#_M1019_g N_A_81_21#_M1002_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3168 AS=0.1424 PD=2.27 PS=1.085 NRD=38.436 NRS=31.872 M=1
+ R=4.26667 SA=75000.8 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1018 N_A_934_297#_M1018_d N_B_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1978 AS=0.2275 PD=1.92 PS=2 NRD=8.304 NRS=8.304 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_A_483_49#_M1009_d N_B_M1009_g N_A_1050_365#_M1009_s VNB NSHORT L=0.15
+ W=0.64 AD=0.234445 AS=0.1948 PD=1.56981 PS=1.9 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75000.2 SB=75002.5 A=0.096 P=1.58 MULT=1
MM1011 N_A_1335_297#_M1011_d N_A_934_297#_M1011_g N_A_483_49#_M1009_d VNB NSHORT
+ L=0.15 W=0.42 AD=0.152666 AS=0.153855 PD=1.0183 PS=1.03019 NRD=88.14
+ NRS=109.992 M=1 R=2.8 SA=75001 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1005 N_A_465_325#_M1005_d N_B_M1005_g N_A_1335_297#_M1011_d VNB NSHORT L=0.15
+ W=0.64 AD=0.177368 AS=0.232634 PD=1.23871 PS=1.5517 NRD=10.308 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75001.8 A=0.096 P=1.58 MULT=1
MM1015 N_A_1050_365#_M1015_d N_A_934_297#_M1015_g N_A_465_325#_M1005_d VNB
+ NSHORT L=0.15 W=0.6 AD=0.121935 AS=0.166282 PD=1.00645 PS=1.16129 NRD=15
+ NRS=42.996 M=1 R=4 SA=75002.1 SB=75001.2 A=0.09 P=1.5 MULT=1
MM1006 N_VGND_M1006_d N_A_M1006_g N_A_1050_365#_M1015_d VNB NSHORT L=0.15 W=0.64
+ AD=0.1024 AS=0.130065 PD=0.96 PS=1.07355 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75002.5 SB=75000.7 A=0.096 P=1.58 MULT=1
MM1023 N_A_1335_297#_M1023_d N_A_1050_365#_M1023_g N_VGND_M1006_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1664 AS=0.1024 PD=1.8 PS=0.96 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75003 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1007 N_X_M1007_d N_A_81_21#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1022 N_X_M1007_d N_A_81_21#_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.267927 PD=1.29 PS=1.79268 NRD=0.9653 NRS=17.73 M=1 R=5.55556
+ SA=90000.6 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1012 N_A_335_93#_M1012_d N_C_M1012_g N_VPWR_M1022_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1856 AS=0.171473 PD=1.86 PS=1.14732 NRD=1.5366 NRS=65.5222 M=1 R=3.55556
+ SA=90001.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1013 N_A_81_21#_M1013_d N_C_M1013_g N_A_465_325#_M1013_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.168 AS=0.2772 PD=1.24 PS=2.34 NRD=11.7215 NRS=1.1623 M=1 R=4.66667
+ SA=90000.2 SB=90001 A=0.1512 P=2.04 MULT=1
MM1003 N_A_483_49#_M1003_d N_A_335_93#_M1003_g N_A_81_21#_M1013_d VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.4494 AS=0.168 PD=2.75 PS=1.24 NRD=59.7895 NRS=16.4101 M=1
+ R=4.66667 SA=90000.8 SB=90000.4 A=0.1512 P=2.04 MULT=1
MM1004 N_A_934_297#_M1004_d N_B_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.3126 AS=0.27 PD=2.64 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1021 N_A_465_325#_M1021_d N_B_M1021_g N_A_1050_365#_M1021_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.286735 AS=0.362 PD=1.66865 PS=2.55 NRD=49.2303 NRS=39.8531 M=1
+ R=4.66667 SA=90000.3 SB=90002.3 A=0.1512 P=2.04 MULT=1
MM1017 N_A_1335_297#_M1017_d N_A_934_297#_M1017_g N_A_465_325#_M1021_d VPB
+ PHIGHVT L=0.18 W=0.64 AD=0.2524 AS=0.218465 PD=1.545 PS=1.27135 NRD=141.584
+ NRS=43.0839 M=1 R=3.55556 SA=90001.1 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1014 N_A_483_49#_M1014_d N_B_M1014_g N_A_1335_297#_M1017_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.132497 AS=0.2524 PD=1.05946 PS=1.545 NRD=46.7875 NRS=0 M=1
+ R=3.55556 SA=90001.6 SB=90001.8 A=0.1152 P=1.64 MULT=1
MM1010 N_A_1050_365#_M1010_d N_A_934_297#_M1010_g N_A_483_49#_M1014_d VPB
+ PHIGHVT L=0.18 W=0.84 AD=0.164987 AS=0.173903 PD=1.25543 PS=1.39054
+ NRD=33.1551 NRS=0 M=1 R=4.66667 SA=90001.7 SB=90001.2 A=0.1512 P=2.04 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_A_1050_365#_M1010_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.196413 PD=1.29 PS=1.49457 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1020 N_A_1335_297#_M1020_d N_A_1050_365#_M1020_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.275 AS=0.145 PD=2.55 PS=1.29 NRD=1.9503 NRS=0.9653 M=1
+ R=5.55556 SA=90002.4 SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.1142 P=23.29
pX25_noxref noxref_16 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__xor3_2.pxi.spice"
*
.ends
*
*
