* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkinvlp_2 A VGND VNB VPB VPWR Y
M1000 Y A a_150_67# VNB nshort w=550000u l=150000u
+  ad=1.5675e+11p pd=1.67e+06u as=1.98e+11p ps=1.82e+06u
M1001 VPWR A Y VPB phighvt w=1e+06u l=250000u
+  ad=6.5e+11p pd=5.3e+06u as=2.8e+11p ps=2.56e+06u
M1002 a_150_67# A VGND VNB nshort w=550000u l=150000u
+  ad=0p pd=0u as=1.5675e+11p ps=1.67e+06u
M1003 Y A VPWR VPB phighvt w=1e+06u l=250000u
+  ad=0p pd=0u as=0p ps=0u
.ends
