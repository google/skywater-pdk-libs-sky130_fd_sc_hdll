* File: sky130_fd_sc_hdll__or4b_1.pex.spice
* Created: Thu Aug 27 19:25:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%D_N 1 3 6 8 9 15
c26 8 0 1.95301e-19 $X=0.265 $Y=0.85
r27 15 16 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r28 13 15 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r29 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r30 8 9 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.255 $Y=0.85
+ $X2=0.255 $Y2=1.16
r31 4 16 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r32 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r33 1 15 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r34 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%A_117_297# 1 2 7 9 12 16 20 26 30
c41 30 0 1.95301e-19 $X=1.485 $Y=1.202
r42 30 31 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r43 27 30 35.8512 $w=3.63e-07 $l=2.7e-07 $layer=POLY_cond $X=1.215 $Y=1.202
+ $X2=1.485 $Y2=1.202
r44 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r45 24 26 15.6453 $w=3.28e-07 $l=4.48e-07 $layer=LI1_cond $X=0.767 $Y=1.16
+ $X2=1.215 $Y2=1.16
r46 22 24 0.069845 $w=3.28e-07 $l=2e-09 $layer=LI1_cond $X=0.765 $Y=1.16
+ $X2=0.767 $Y2=1.16
r47 18 22 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.16
r48 18 20 18.9673 $w=2.38e-07 $l=3.95e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.72
r49 14 24 2.50173 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=0.767 $Y=0.995
+ $X2=0.767 $Y2=1.16
r50 14 16 23.2841 $w=2.43e-07 $l=4.95e-07 $layer=LI1_cond $X=0.767 $Y=0.995
+ $X2=0.767 $Y2=0.5
r51 10 31 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r52 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.475
r53 7 30 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r54 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.695
r55 2 20 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.72
r56 1 16 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=0.73 $Y2=0.5
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%C 1 3 6 8 10 22 26
r36 18 26 2.70082 $w=6.18e-07 $l=1.4e-07 $layer=LI1_cond $X=1.93 $Y=1.305
+ $X2=2.07 $Y2=1.305
r37 18 22 3.56894 $w=6.18e-07 $l=1.85e-07 $layer=LI1_cond $X=1.93 $Y=1.305
+ $X2=1.745 $Y2=1.305
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.16 $X2=1.93 $Y2=1.16
r39 10 26 2.89374 $w=6.18e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.305
+ $X2=2.07 $Y2=1.305
r40 8 22 0.675206 $w=6.18e-07 $l=3.5e-08 $layer=LI1_cond $X=1.71 $Y=1.305
+ $X2=1.745 $Y2=1.305
r41 4 17 38.8084 $w=2.75e-07 $l=1.98167e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=1.942 $Y2=1.16
r42 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.475
r43 1 17 49.5676 $w=2.75e-07 $l=2.72947e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.942 $Y2=1.16
r44 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.99 $Y=1.41 $X2=1.99
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%B 1 2 3 4 6 9 10 11 12 13 14 21 25 28 31 35
c42 2 0 8.49032e-20 $X=2.43 $Y=1.31
r43 25 28 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.27 $X2=1.15
+ $Y2=2.27
r44 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=2.31 $X2=2.47 $Y2=2.31
r45 14 21 9.93485 $w=2.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.22 $Y=2.27
+ $X2=2.47 $Y2=2.27
r46 14 35 5.96091 $w=2.88e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=2.27
+ $X2=2.07 $Y2=2.27
r47 13 35 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.71 $Y=2.27
+ $X2=2.07 $Y2=2.27
r48 13 31 3.97394 $w=2.88e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=2.27 $X2=1.61
+ $Y2=2.27
r49 12 31 16.2932 $w=2.88e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=2.27 $X2=1.61
+ $Y2=2.27
r50 12 28 1.98697 $w=2.88e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=2.27 $X2=1.15
+ $Y2=2.27
r51 11 25 4.96743 $w=2.88e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=2.27
+ $X2=0.87 $Y2=2.27
r52 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=2.455 $Y=0.475
+ $X2=2.455 $Y2=0.76
r53 4 20 56.0837 $w=2.56e-07 $l=2.92916e-07 $layer=POLY_cond $X=2.43 $Y=2.035
+ $X2=2.467 $Y2=2.31
r54 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=2.43 $Y=2.035 $X2=2.43
+ $Y2=1.695
r55 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.43 $Y=1.41 $X2=2.43
+ $Y2=1.695
r56 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.43 $Y=1.31 $X2=2.43
+ $Y2=1.41
r57 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.43 $Y=0.86 $X2=2.43
+ $Y2=0.76
r58 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=2.43 $Y=0.86 $X2=2.43
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%A 1 3 6 8 12 16
r38 12 16 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=2.89 $Y=1.16
+ $X2=2.765 $Y2=1.16
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=1.16 $X2=2.89 $Y2=1.16
r40 8 16 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.73 $Y=1.16
+ $X2=2.765 $Y2=1.16
r41 4 11 39.1718 $w=2.59e-07 $l=1.93959e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=2.892 $Y2=1.16
r42 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.955 $Y=0.995
+ $X2=2.955 $Y2=0.475
r43 1 11 51.0578 $w=2.59e-07 $l=2.68328e-07 $layer=POLY_cond $X=2.93 $Y=1.41
+ $X2=2.892 $Y2=1.16
r44 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.93 $Y=1.41 $X2=2.93
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%A_225_297# 1 2 3 10 12 13 15 16 20 22 23 26
+ 28 30 35 37 41 42 47 49
c94 47 0 1.17306e-19 $X=3.42 $Y=1.16
c95 35 0 1.08657e-19 $X=3.33 $Y=1.495
r96 47 50 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=1.16
+ $X2=3.375 $Y2=1.325
r97 47 49 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=1.16
+ $X2=3.375 $Y2=0.995
r98 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.16 $X2=3.42 $Y2=1.16
r99 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.775 $Y2=1.87
r100 37 39 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=1.24 $Y=1.685
+ $X2=1.24 $Y2=1.87
r101 35 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.33 $Y=1.495
+ $X2=3.33 $Y2=1.325
r102 32 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.33 $Y=0.825
+ $X2=3.33 $Y2=0.995
r103 31 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.86 $Y=1.58
+ $X2=2.775 $Y2=1.58
r104 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=1.58
+ $X2=3.33 $Y2=1.495
r105 30 31 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.245 $Y=1.58
+ $X2=2.86 $Y2=1.58
r106 29 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.78 $Y=0.74
+ $X2=2.695 $Y2=0.74
r107 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=0.74
+ $X2=3.33 $Y2=0.825
r108 28 29 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.245 $Y=0.74
+ $X2=2.78 $Y2=0.74
r109 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.655
+ $X2=2.695 $Y2=0.74
r110 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.695 $Y=0.655
+ $X2=2.695 $Y2=0.47
r111 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.74
+ $X2=2.695 $Y2=0.74
r112 22 23 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.61 $Y=0.74
+ $X2=1.835 $Y2=0.74
r113 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.75 $Y=0.655
+ $X2=1.835 $Y2=0.74
r114 18 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.75 $Y=0.655
+ $X2=1.75 $Y2=0.47
r115 17 39 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=1.4 $Y=1.87 $X2=1.24
+ $Y2=1.87
r116 16 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.69 $Y=1.87
+ $X2=2.775 $Y2=1.87
r117 16 17 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=2.69 $Y=1.87
+ $X2=1.4 $Y2=1.87
r118 13 48 38.9672 $w=2.67e-07 $l=1.96074e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.427 $Y2=1.16
r119 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.495 $Y2=0.56
r120 10 48 50.2707 $w=2.67e-07 $l=2.70647e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.427 $Y2=1.16
r121 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.985
r122 3 37 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.685
r123 2 26 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.265 $X2=2.695 $Y2=0.47
r124 1 20 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.265 $X2=1.75 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%VPWR 1 2 7 9 13 16 17 18 28 29
c35 2 0 1.08657e-19 $X=3.02 $Y=1.485
r36 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r37 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r38 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 23 26 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.99 $Y2=2.72
r40 22 25 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.99 $Y2=2.72
r41 22 23 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 20 32 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r43 20 22 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 16 25 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=3.08 $Y=2.72 $X2=2.99
+ $Y2=2.72
r47 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.08 $Y=2.72 $X2=3.22
+ $Y2=2.72
r48 15 28 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.36 $Y=2.72
+ $X2=3.91 $Y2=2.72
r49 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=3.36 $Y=2.72 $X2=3.22
+ $Y2=2.72
r50 11 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r51 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2
r52 7 32 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.212 $Y2=2.72
r53 7 9 31.0143 $w=3.38e-07 $l=9.15e-07 $layer=LI1_cond $X=0.255 $Y=2.635
+ $X2=0.255 $Y2=1.72
r54 2 13 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=3.02
+ $Y=1.485 $X2=3.23 $Y2=2
r55 1 9 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%X 1 2 10 13 14 15
r18 13 15 5.00929 $w=3.73e-07 $l=1.63e-07 $layer=LI1_cond $X=3.807 $Y=1.682
+ $X2=3.807 $Y2=1.845
r19 13 14 6.669 $w=3.73e-07 $l=1.87e-07 $layer=LI1_cond $X=3.807 $Y=1.682
+ $X2=3.807 $Y2=1.495
r20 12 14 31.3721 $w=2.68e-07 $l=7.35e-07 $layer=LI1_cond $X=3.86 $Y=0.76
+ $X2=3.86 $Y2=1.495
r21 10 12 6.14656 $w=3.73e-07 $l=1.7e-07 $layer=LI1_cond $X=3.807 $Y=0.59
+ $X2=3.807 $Y2=0.76
r22 2 15 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.485 $X2=3.705 $Y2=1.845
r23 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.705 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4B_1%VGND 1 2 3 4 13 15 17 21 23 27 29 31 35 36
+ 42 45 49
r63 49 52 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.165
+ $Y2=0.4
r64 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r65 46 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r66 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r67 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r68 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r69 36 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r70 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r71 33 49 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.165
+ $Y2=0
r72 33 35 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.91
+ $Y2=0
r73 31 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r74 31 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r75 30 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.2
+ $Y2=0
r76 29 49 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=3.165
+ $Y2=0
r77 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.95 $Y=0 $X2=2.39
+ $Y2=0
r78 25 45 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=0.085 $X2=2.2
+ $Y2=0
r79 25 27 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.2 $Y=0.085
+ $X2=2.2 $Y2=0.4
r80 24 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.415 $Y=0 $X2=1.25
+ $Y2=0
r81 23 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=2.2
+ $Y2=0
r82 23 24 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.01 $Y=0 $X2=1.415
+ $Y2=0
r83 19 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0
r84 19 21 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0.5
r85 18 39 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r86 17 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=1.25
+ $Y2=0
r87 17 18 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.085 $Y=0 $X2=0.425
+ $Y2=0
r88 13 39 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.212 $Y2=0
r89 13 15 14.0666 $w=3.38e-07 $l=4.15e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.5
r90 4 52 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.03
+ $Y=0.265 $X2=3.215 $Y2=0.4
r91 3 27 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.265 $X2=2.225 $Y2=0.4
r92 2 21 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.265 $X2=1.25 $Y2=0.5
r93 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends

