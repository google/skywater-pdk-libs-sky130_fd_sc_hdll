* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfxtp_4 CLK D SCD SCE VGND VNB VPB VPWR Q
M1000 VPWR a_1189_183# a_1121_413# VPB phighvt w=420000u l=180000u
+  ad=1.98115e+12p pd=1.754e+07u as=1.47e+11p ps=1.54e+06u
M1001 VPWR CLK a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1002 a_608_369# D a_517_47# VNB nshort w=420000u l=150000u
+  ad=2.604e+11p pd=2.88e+06u as=1.428e+11p ps=1.52e+06u
M1003 a_1474_413# a_27_47# a_1189_183# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.307e+11p ps=2.19e+06u
M1004 VPWR a_1667_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 VGND a_1667_315# a_1625_47# VNB nshort w=420000u l=150000u
+  ad=1.48085e+12p pd=1.433e+07u as=1.32e+11p ps=1.49e+06u
M1006 VGND a_1667_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.485e+11p ps=3.98e+06u
M1007 VGND a_1189_183# a_1127_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.584e+11p ps=1.62e+06u
M1008 a_504_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=2.176e+11p pd=1.96e+06u as=0p ps=0u
M1009 a_203_47# a_27_47# VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1010 VPWR a_1667_315# a_1568_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.121e+11p ps=1.85e+06u
M1011 VGND a_1667_315# Q VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR SCE a_319_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 a_1121_413# a_27_47# a_1011_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1014 a_1474_413# a_203_47# a_1189_183# VNB nshort w=360000u l=150000u
+  ad=1.854e+11p pd=1.75e+06u as=1.978e+11p ps=1.99e+06u
M1015 Q a_1667_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND SCE a_319_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1017 Q a_1667_315# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_1667_315# Q VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND a_1474_413# a_1667_315# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1020 a_517_47# a_319_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1127_47# a_203_47# a_1011_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.548e+11p ps=1.58e+06u
M1022 a_1189_183# a_1011_47# VPWR VPB phighvt w=750000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 Q a_1667_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_1011_47# a_203_47# a_608_369# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=3.2e+11p ps=3.34e+06u
M1025 Q a_1667_315# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_203_47# a_27_47# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1027 a_1625_47# a_27_47# a_1474_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 VPWR SCD a_702_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=2.144e+11p ps=1.95e+06u
M1029 VGND SCD a_721_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=9.66e+10p ps=1.3e+06u
M1030 VPWR a_1474_413# a_1667_315# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1031 a_702_369# a_319_47# a_608_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1032 a_1189_183# a_1011_47# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_1568_413# a_203_47# a_1474_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_1011_47# a_27_47# a_608_369# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 VGND CLK a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1036 a_721_47# SCE a_608_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_608_369# D a_504_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
