* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb4to1_1 D[3] D[2] D[1] D[0] S[3] S[2] S[1] S[0] VGND
+ VNB VPB VPWR Z
X0 VPWR S[1] a_533_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND D[2] a_937_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1012_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 a_1574_47# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1012_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_109_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X7 VPWR D[2] a_945_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR S[3] a_1361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_117_297# a_184_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X10 Z a_533_47# a_734_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_184_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X12 VGND S[3] a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X13 VGND S[1] a_533_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X14 a_1562_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_945_297# a_1012_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 VGND D[0] a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Z a_1361_47# a_1562_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X18 a_937_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X19 Z S[3] a_1574_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 Z S[1] a_746_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_734_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_184_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_746_47# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
