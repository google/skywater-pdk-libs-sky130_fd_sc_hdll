* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor3_4 A B C VGND VNB VPB VPWR X
M1000 X a_101_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.50095e+12p ps=1.307e+07u
M1001 a_1490_297# a_1207_297# VGND VNB nshort w=640000u l=150000u
+  ad=5.677e+11p pd=4.42e+06u as=1.0748e+12p ps=9.85e+06u
M1002 a_532_93# C VPWR VPB phighvt w=640000u l=180000u
+  ad=1.856e+11p pd=1.86e+06u as=0p ps=0u
M1003 VGND A a_1207_297# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=4.44e+11p ps=3.96e+06u
M1004 a_1089_297# B VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1005 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 a_657_325# B a_1207_297# VNB nshort w=640000u l=150000u
+  ad=5.835e+11p pd=4.49e+06u as=0p ps=0u
M1007 VGND a_101_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_681_49# B a_1207_297# VPB phighvt w=840000u l=180000u
+  ad=8.3175e+11p pd=5.4e+06u as=7.226e+11p ps=5.29e+06u
M1009 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_1207_297# a_1089_297# a_657_325# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=5.878e+11p ps=4.8e+06u
M1011 a_1490_297# a_1089_297# a_657_325# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_101_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_1490_297# a_1207_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.998e+11p pd=5.68e+06u as=0p ps=0u
M1014 a_681_49# B a_1490_297# VNB nshort w=640000u l=150000u
+  ad=5.4845e+11p pd=4.32e+06u as=0p ps=0u
M1015 a_1207_297# a_1089_297# a_681_49# VNB nshort w=600000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_657_325# B a_1490_297# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_101_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR A a_1207_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_101_21# C a_657_325# VPB phighvt w=840000u l=180000u
+  ad=3.227e+11p pd=2.67e+06u as=0p ps=0u
M1020 a_657_325# a_532_93# a_101_21# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=2.432e+11p ps=2.04e+06u
M1021 a_1490_297# a_1089_297# a_681_49# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_101_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_101_21# C a_681_49# VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VPWR a_101_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1025 a_681_49# a_532_93# a_101_21# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_532_93# C VGND VNB nshort w=420000u l=150000u
+  ad=1.995e+11p pd=1.79e+06u as=0p ps=0u
M1027 a_1089_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.2e+11p pd=2.64e+06u as=0p ps=0u
.ends
