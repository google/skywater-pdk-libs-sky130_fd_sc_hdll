* File: sky130_fd_sc_hdll__sdfbbp_1.pxi.spice
* Created: Wed Sep  2 08:50:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%CLK N_CLK_c_297_n N_CLK_c_298_n N_CLK_M1008_g
+ N_CLK_c_292_n N_CLK_M1033_g N_CLK_c_293_n CLK CLK N_CLK_c_295_n N_CLK_c_296_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%CLK
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_27_47# N_A_27_47#_M1033_s N_A_27_47#_M1008_s
+ N_A_27_47#_c_344_n N_A_27_47#_c_345_n N_A_27_47#_M1038_g N_A_27_47#_M1001_g
+ N_A_27_47#_c_334_n N_A_27_47#_M1027_g N_A_27_47#_c_346_n N_A_27_47#_M1006_g
+ N_A_27_47#_c_347_n N_A_27_47#_c_348_n N_A_27_47#_M1042_g N_A_27_47#_c_335_n
+ N_A_27_47#_c_336_n N_A_27_47#_M1046_g N_A_27_47#_c_576_p N_A_27_47#_c_338_n
+ N_A_27_47#_c_339_n N_A_27_47#_c_351_n N_A_27_47#_c_463_p N_A_27_47#_c_340_n
+ N_A_27_47#_c_341_n N_A_27_47#_c_342_n N_A_27_47#_c_354_n N_A_27_47#_c_355_n
+ N_A_27_47#_c_356_n N_A_27_47#_c_357_n N_A_27_47#_c_358_n N_A_27_47#_c_359_n
+ N_A_27_47#_c_343_n N_A_27_47#_c_361_n N_A_27_47#_c_362_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCD N_SCD_c_591_n N_SCD_M1018_g N_SCD_M1023_g
+ SCD SCD N_SCD_c_594_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCD
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_453_315# N_A_453_315#_M1003_s
+ N_A_453_315#_M1011_s N_A_453_315#_c_634_n N_A_453_315#_M1022_g
+ N_A_453_315#_c_635_n N_A_453_315#_c_636_n N_A_453_315#_c_628_n
+ N_A_453_315#_M1045_g N_A_453_315#_c_637_n N_A_453_315#_c_659_p
+ N_A_453_315#_c_638_n N_A_453_315#_c_629_n N_A_453_315#_c_630_n
+ N_A_453_315#_c_631_n N_A_453_315#_c_632_n N_A_453_315#_c_640_n
+ N_A_453_315#_c_633_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_453_315#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCE N_SCE_c_737_n N_SCE_M1024_g N_SCE_c_738_n
+ N_SCE_c_739_n N_SCE_c_747_n N_SCE_M1011_g N_SCE_c_740_n N_SCE_M1003_g
+ N_SCE_c_748_n N_SCE_c_749_n N_SCE_M1004_g N_SCE_c_741_n N_SCE_c_750_n
+ N_SCE_c_742_n N_SCE_c_757_n SCE SCE SCE N_SCE_c_745_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%SCE
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%D N_D_c_847_n N_D_c_848_n N_D_M1044_g
+ N_D_M1035_g D D N_D_c_850_n N_D_c_851_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%D
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_211_363# N_A_211_363#_M1001_d
+ N_A_211_363#_M1038_d N_A_211_363#_c_911_n N_A_211_363#_c_912_n
+ N_A_211_363#_M1020_g N_A_211_363#_c_893_n N_A_211_363#_c_894_n
+ N_A_211_363#_M1019_g N_A_211_363#_c_896_n N_A_211_363#_c_897_n
+ N_A_211_363#_M1010_g N_A_211_363#_c_915_n N_A_211_363#_M1032_g
+ N_A_211_363#_c_898_n N_A_211_363#_c_899_n N_A_211_363#_c_900_n
+ N_A_211_363#_c_916_n N_A_211_363#_c_901_n N_A_211_363#_c_902_n
+ N_A_211_363#_c_903_n N_A_211_363#_c_904_n N_A_211_363#_c_905_n
+ N_A_211_363#_c_906_n N_A_211_363#_c_907_n N_A_211_363#_c_908_n
+ N_A_211_363#_c_909_n N_A_211_363#_c_910_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_211_363#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1197_21# N_A_1197_21#_M1013_d
+ N_A_1197_21#_M1012_d N_A_1197_21#_M1025_g N_A_1197_21#_c_1131_n
+ N_A_1197_21#_M1015_g N_A_1197_21#_c_1132_n N_A_1197_21#_c_1133_n
+ N_A_1197_21#_M1041_g N_A_1197_21#_c_1124_n N_A_1197_21#_M1037_g
+ N_A_1197_21#_c_1134_n N_A_1197_21#_c_1181_p N_A_1197_21#_c_1146_n
+ N_A_1197_21#_c_1125_n N_A_1197_21#_c_1126_n N_A_1197_21#_c_1127_n
+ N_A_1197_21#_c_1136_n N_A_1197_21#_c_1148_n N_A_1197_21#_c_1128_n
+ N_A_1197_21#_c_1129_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1197_21#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%SET_B N_SET_B_c_1270_n N_SET_B_c_1282_n
+ N_SET_B_M1012_g N_SET_B_M1009_g N_SET_B_c_1272_n N_SET_B_c_1284_n
+ N_SET_B_M1002_g N_SET_B_M1000_g N_SET_B_c_1274_n N_SET_B_c_1275_n
+ N_SET_B_c_1276_n N_SET_B_c_1277_n SET_B N_SET_B_c_1278_n N_SET_B_c_1279_n
+ N_SET_B_c_1280_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%SET_B
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1003_47# N_A_1003_47#_M1027_d
+ N_A_1003_47#_M1020_d N_A_1003_47#_c_1400_n N_A_1003_47#_M1031_g
+ N_A_1003_47#_M1013_g N_A_1003_47#_c_1409_n N_A_1003_47#_c_1414_n
+ N_A_1003_47#_c_1406_n N_A_1003_47#_c_1402_n N_A_1003_47#_c_1403_n
+ N_A_1003_47#_c_1404_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1003_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1525_21# N_A_1525_21#_M1028_s
+ N_A_1525_21#_M1017_s N_A_1525_21#_M1021_g N_A_1525_21#_c_1516_n
+ N_A_1525_21#_M1026_g N_A_1525_21#_c_1517_n N_A_1525_21#_M1036_g
+ N_A_1525_21#_M1007_g N_A_1525_21#_c_1509_n N_A_1525_21#_c_1510_n
+ N_A_1525_21#_c_1518_n N_A_1525_21#_c_1519_n N_A_1525_21#_c_1511_n
+ N_A_1525_21#_c_1512_n N_A_1525_21#_c_1521_n N_A_1525_21#_c_1522_n
+ N_A_1525_21#_c_1523_n N_A_1525_21#_c_1524_n N_A_1525_21#_c_1513_n
+ N_A_1525_21#_c_1514_n N_A_1525_21#_c_1515_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1525_21#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2058_21# N_A_2058_21#_M1040_d
+ N_A_2058_21#_M1002_d N_A_2058_21#_M1014_g N_A_2058_21#_c_1674_n
+ N_A_2058_21#_M1029_g N_A_2058_21#_c_1663_n N_A_2058_21#_M1039_g
+ N_A_2058_21#_c_1664_n N_A_2058_21#_M1005_g N_A_2058_21#_c_1665_n
+ N_A_2058_21#_c_1666_n N_A_2058_21#_c_1667_n N_A_2058_21#_c_1677_n
+ N_A_2058_21#_M1030_g N_A_2058_21#_c_1668_n N_A_2058_21#_M1043_g
+ N_A_2058_21#_c_1669_n N_A_2058_21#_c_1670_n N_A_2058_21#_c_1678_n
+ N_A_2058_21#_c_1679_n N_A_2058_21#_c_1680_n N_A_2058_21#_c_1738_p
+ N_A_2058_21#_c_1698_n N_A_2058_21#_c_1707_n N_A_2058_21#_c_1671_n
+ N_A_2058_21#_c_1682_n N_A_2058_21#_c_1683_n N_A_2058_21#_c_1724_n
+ N_A_2058_21#_c_1700_n N_A_2058_21#_c_1726_n N_A_2058_21#_c_1672_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2058_21#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1864_47# N_A_1864_47#_M1010_d
+ N_A_1864_47#_M1042_d N_A_1864_47#_c_1845_n N_A_1864_47#_M1034_g
+ N_A_1864_47#_M1040_g N_A_1864_47#_c_1856_n N_A_1864_47#_c_1859_n
+ N_A_1864_47#_c_1847_n N_A_1864_47#_c_1852_n N_A_1864_47#_c_1848_n
+ N_A_1864_47#_c_1849_n N_A_1864_47#_c_1850_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1864_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%RESET_B N_RESET_B_c_1940_n N_RESET_B_M1017_g
+ N_RESET_B_M1028_g RESET_B N_RESET_B_c_1942_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%RESET_B
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2845_47# N_A_2845_47#_M1043_s
+ N_A_2845_47#_M1030_s N_A_2845_47#_c_1972_n N_A_2845_47#_M1016_g
+ N_A_2845_47#_c_1973_n N_A_2845_47#_M1047_g N_A_2845_47#_c_1978_n
+ N_A_2845_47#_c_1979_n N_A_2845_47#_c_1974_n N_A_2845_47#_c_1975_n
+ N_A_2845_47#_c_1981_n N_A_2845_47#_c_1976_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2845_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%VPWR N_VPWR_M1008_d N_VPWR_M1018_s
+ N_VPWR_M1011_d N_VPWR_M1015_d N_VPWR_M1026_d N_VPWR_M1029_d N_VPWR_M1036_d
+ N_VPWR_M1017_d N_VPWR_M1030_d N_VPWR_c_2028_n N_VPWR_c_2029_n N_VPWR_c_2030_n
+ N_VPWR_c_2031_n N_VPWR_c_2032_n N_VPWR_c_2033_n N_VPWR_c_2034_n
+ N_VPWR_c_2035_n N_VPWR_c_2036_n N_VPWR_c_2037_n N_VPWR_c_2038_n VPWR VPWR
+ N_VPWR_c_2039_n N_VPWR_c_2040_n N_VPWR_c_2041_n N_VPWR_c_2042_n
+ N_VPWR_c_2043_n N_VPWR_c_2044_n N_VPWR_c_2045_n N_VPWR_c_2027_n
+ N_VPWR_c_2047_n N_VPWR_c_2048_n N_VPWR_c_2049_n N_VPWR_c_2050_n
+ N_VPWR_c_2051_n N_VPWR_c_2052_n N_VPWR_c_2053_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_483_47# N_A_483_47#_M1024_d
+ N_A_483_47#_M1035_d N_A_483_47#_M1022_d N_A_483_47#_M1044_d
+ N_A_483_47#_c_2240_n N_A_483_47#_c_2248_n N_A_483_47#_c_2249_n
+ N_A_483_47#_c_2241_n N_A_483_47#_c_2242_n N_A_483_47#_c_2243_n
+ N_A_483_47#_c_2244_n N_A_483_47#_c_2245_n N_A_483_47#_c_2246_n
+ N_A_483_47#_c_2247_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_483_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q_N N_Q_N_M1005_d N_Q_N_M1039_d N_Q_N_c_2380_n
+ Q_N Q_N Q_N PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q_N
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q N_Q_M1047_d N_Q_M1016_d N_Q_c_2410_n
+ N_Q_c_2413_n N_Q_c_2411_n Q Q Q PM_SKY130_FD_SC_HDLL__SDFBBP_1%Q
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%VGND N_VGND_M1033_d N_VGND_M1023_s
+ N_VGND_M1003_d N_VGND_M1025_d N_VGND_M1037_s N_VGND_M1014_d N_VGND_M1028_d
+ N_VGND_M1043_d N_VGND_c_2427_n N_VGND_c_2428_n N_VGND_c_2429_n N_VGND_c_2430_n
+ N_VGND_c_2431_n N_VGND_c_2432_n N_VGND_c_2433_n N_VGND_c_2434_n
+ N_VGND_c_2435_n N_VGND_c_2436_n N_VGND_c_2437_n VGND VGND N_VGND_c_2438_n
+ N_VGND_c_2439_n N_VGND_c_2440_n N_VGND_c_2441_n N_VGND_c_2442_n
+ N_VGND_c_2443_n N_VGND_c_2444_n N_VGND_c_2445_n N_VGND_c_2446_n
+ N_VGND_c_2447_n N_VGND_c_2448_n N_VGND_c_2449_n
+ PM_SKY130_FD_SC_HDLL__SDFBBP_1%VGND
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1353_47# N_A_1353_47#_M1009_d
+ N_A_1353_47#_M1021_d N_A_1353_47#_c_2647_n N_A_1353_47#_c_2650_n
+ N_A_1353_47#_c_2657_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_1353_47#
x_PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2216_47# N_A_2216_47#_M1000_d
+ N_A_2216_47#_M1007_d N_A_2216_47#_c_2675_n N_A_2216_47#_c_2678_n
+ N_A_2216_47#_c_2687_n PM_SKY130_FD_SC_HDLL__SDFBBP_1%A_2216_47#
cc_1 VNB N_CLK_c_292_n 0.0173562f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_CLK_c_293_n 0.0274923f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB CLK 0.0190059f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_CLK_c_295_n 0.0200795f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_5 VNB N_CLK_c_296_n 0.012957f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_6 VNB N_A_27_47#_M1001_g 0.0399088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_334_n 0.0184212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_335_n 0.0140217f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_9 VNB N_A_27_47#_c_336_n 0.00421248f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_10 VNB N_A_27_47#_M1046_g 0.0485955f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_11 VNB N_A_27_47#_c_338_n 0.00306944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_339_n 0.00649157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_340_n 0.00697621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_341_n 0.00495758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_342_n 0.0354975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_343_n 0.0266073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_SCD_M1023_g 0.0515243f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_18 VNB SCD 0.00765024f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_19 VNB N_A_453_315#_c_628_n 0.0172836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_453_315#_c_629_n 0.00171575f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_21 VNB N_A_453_315#_c_630_n 7.51239e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_22 VNB N_A_453_315#_c_631_n 0.00739396f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.4
cc_23 VNB N_A_453_315#_c_632_n 0.0043798f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_24 VNB N_A_453_315#_c_633_n 0.0335168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_SCE_c_737_n 0.0175345f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_26 VNB N_SCE_c_738_n 0.0503975f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.59
cc_27 VNB N_SCE_c_739_n 0.0306073f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_28 VNB N_SCE_c_740_n 0.0186337f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_29 VNB N_SCE_c_741_n 0.00495818f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_30 VNB N_SCE_c_742_n 0.00165072f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_31 VNB SCE 9.00566e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB SCE 0.00350585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_SCE_c_745_n 0.0332322f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_D_M1035_g 0.0497285f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_35 VNB N_A_211_363#_c_893_n 0.0136597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_211_363#_c_894_n 0.00503487f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_37 VNB N_A_211_363#_M1019_g 0.0207598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_211_363#_c_896_n 0.00970036f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_39 VNB N_A_211_363#_c_897_n 0.0187478f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_40 VNB N_A_211_363#_c_898_n 0.00393559f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_41 VNB N_A_211_363#_c_899_n 0.0358981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_211_363#_c_900_n 0.00519746f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_43 VNB N_A_211_363#_c_901_n 0.0307224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_211_363#_c_902_n 0.00717892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_211_363#_c_903_n 0.0012696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_211_363#_c_904_n 0.0226005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_211_363#_c_905_n 0.00244668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_211_363#_c_906_n 0.00200585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_211_363#_c_907_n 0.00147534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_211_363#_c_908_n 0.0281305f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_211_363#_c_909_n 0.00544606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_211_363#_c_910_n 0.0144647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_1197_21#_M1025_g 0.0441094f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_54 VNB N_A_1197_21#_c_1124_n 0.0201729f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_55 VNB N_A_1197_21#_c_1125_n 0.00234062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1197_21#_c_1126_n 0.00458496f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_57 VNB N_A_1197_21#_c_1127_n 0.0106807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1197_21#_c_1128_n 0.00509217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1197_21#_c_1129_n 0.0403718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_SET_B_c_1270_n 0.00806415f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=1.07
cc_61 VNB N_SET_B_M1009_g 0.0219221f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_62 VNB N_SET_B_c_1272_n 0.00905407f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.805
cc_63 VNB N_SET_B_M1000_g 0.0219371f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_64 VNB N_SET_B_c_1274_n 0.0178189f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_65 VNB N_SET_B_c_1275_n 0.00236707f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_66 VNB N_SET_B_c_1276_n 0.00377633f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_SET_B_c_1277_n 0.00499724f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_68 VNB N_SET_B_c_1278_n 0.0343481f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_69 VNB N_SET_B_c_1279_n 0.0363063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_SET_B_c_1280_n 0.00766748f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1003_47#_c_1400_n 0.0164642f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_72 VNB N_A_1003_47#_M1013_g 0.0270526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1003_47#_c_1402_n 0.00436764f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_74 VNB N_A_1003_47#_c_1403_n 0.00920304f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_75 VNB N_A_1003_47#_c_1404_n 0.00397751f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.53
cc_76 VNB N_A_1525_21#_M1021_g 0.0290482f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_77 VNB N_A_1525_21#_M1007_g 0.0302025f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_78 VNB N_A_1525_21#_c_1509_n 0.0128915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1525_21#_c_1510_n 9.06558e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1525_21#_c_1511_n 0.00275664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1525_21#_c_1512_n 9.08783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1525_21#_c_1513_n 0.0229813f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1525_21#_c_1514_n 0.0216754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1525_21#_c_1515_n 0.00430752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_2058_21#_M1014_g 0.047147f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_86 VNB N_A_2058_21#_c_1663_n 0.0185038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_2058_21#_c_1664_n 0.0205943f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.665
cc_88 VNB N_A_2058_21#_c_1665_n 0.0695137f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_89 VNB N_A_2058_21#_c_1666_n 0.00922379f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_90 VNB N_A_2058_21#_c_1667_n 5.47963e-19 $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_91 VNB N_A_2058_21#_c_1668_n 0.0182233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2058_21#_c_1669_n 0.022776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_2058_21#_c_1670_n 0.00868848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_2058_21#_c_1671_n 0.00768762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2058_21#_c_1672_n 0.00274082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_1864_47#_c_1845_n 0.0207574f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_97 VNB N_A_1864_47#_M1040_g 0.0230717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_1864_47#_c_1847_n 0.0121665f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_99 VNB N_A_1864_47#_c_1848_n 0.0121507f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_100 VNB N_A_1864_47#_c_1849_n 5.15456e-19 $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.19
cc_101 VNB N_A_1864_47#_c_1850_n 0.00278937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_RESET_B_c_1940_n 0.0330627f $X=-0.19 $Y=-0.24 $X2=0.3 $Y2=0.88
cc_103 VNB N_RESET_B_M1028_g 0.036034f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.135
cc_104 VNB N_RESET_B_c_1942_n 0.00445413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_A_2845_47#_c_1972_n 0.0296875f $X=-0.19 $Y=-0.24 $X2=0.495
+ $Y2=2.135
cc_106 VNB N_A_2845_47#_c_1973_n 0.0209122f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_107 VNB N_A_2845_47#_c_1974_n 0.0055399f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_108 VNB N_A_2845_47#_c_1975_n 0.00577182f $X=-0.19 $Y=-0.24 $X2=0.24
+ $Y2=1.235
cc_109 VNB N_A_2845_47#_c_1976_n 3.97688e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VPWR_c_2027_n 0.649277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_A_483_47#_c_2240_n 0.00646091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_A_483_47#_c_2241_n 0.00649828f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_113 VNB N_A_483_47#_c_2242_n 0.00691332f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.07
cc_114 VNB N_A_483_47#_c_2243_n 0.0105956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_A_483_47#_c_2244_n 0.00216713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_A_483_47#_c_2245_n 0.00650741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_A_483_47#_c_2246_n 0.00342916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_A_483_47#_c_2247_n 0.0141494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB Q_N 0.00724219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB Q_N 0.00435453f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_121 VNB N_Q_c_2410_n 0.00558658f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_122 VNB N_Q_c_2411_n 0.0239385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB Q 0.0173379f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_124 VNB N_VGND_c_2427_n 0.0193693f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.235
cc_125 VNB N_VGND_c_2428_n 0.00902838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2429_n 0.00561552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2430_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2431_n 0.00270706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2432_n 0.0084514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2433_n 0.00540497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2434_n 0.0652777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2435_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_VGND_c_2436_n 0.0456676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2437_n 0.00469069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2438_n 0.0153731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2439_n 0.0485686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2440_n 0.0583156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2441_n 0.0589514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2442_n 0.0362874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2443_n 0.0185741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2444_n 0.717564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2445_n 0.00803343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2446_n 0.00478425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2447_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2448_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2449_n 0.00554993f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VPB N_CLK_c_297_n 0.0103472f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.59
cc_148 VPB N_CLK_c_298_n 0.0469586f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.74
cc_149 VPB CLK 0.0180386f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_150 VPB N_CLK_c_295_n 0.0102811f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_151 VPB N_A_27_47#_c_344_n 0.0182013f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_152 VPB N_A_27_47#_c_345_n 0.0249569f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_153 VPB N_A_27_47#_c_346_n 0.0535589f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_154 VPB N_A_27_47#_c_347_n 0.0136389f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_155 VPB N_A_27_47#_c_348_n 0.0560417f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_156 VPB N_A_27_47#_c_335_n 0.0188976f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.4
cc_157 VPB N_A_27_47#_c_336_n 0.00462609f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_158 VPB N_A_27_47#_c_351_n 0.00118717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_27_47#_c_340_n 0.00383268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_27_47#_c_341_n 0.00305141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_27_47#_c_354_n 0.00363921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_27_47#_c_355_n 0.0348058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_27_47#_c_356_n 0.00241915f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_27_47#_c_357_n 0.00875464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_27_47#_c_358_n 0.00166538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_27_47#_c_359_n 0.00352609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_27_47#_c_343_n 0.0123596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_27_47#_c_361_n 0.0062255f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_27_47#_c_362_n 0.00243614f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_SCD_c_591_n 0.0186886f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.88
cc_171 VPB N_SCD_M1023_g 0.00126351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_172 VPB SCD 0.00536826f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_173 VPB N_SCD_c_594_n 0.0583117f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_174 VPB N_A_453_315#_c_634_n 0.0190875f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_175 VPB N_A_453_315#_c_635_n 0.0629439f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_176 VPB N_A_453_315#_c_636_n 0.0125601f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_177 VPB N_A_453_315#_c_637_n 0.00301632f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.665
cc_178 VPB N_A_453_315#_c_638_n 0.00860618f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_179 VPB N_A_453_315#_c_632_n 0.00586331f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_180 VPB N_A_453_315#_c_640_n 0.00654809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_SCE_c_739_n 0.0361068f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_182 VPB N_SCE_c_747_n 0.0187356f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_183 VPB N_SCE_c_748_n 0.0326077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_SCE_c_749_n 0.0162468f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_SCE_c_750_n 0.00721158f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_186 VPB SCE 0.00666805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_D_c_847_n 0.01732f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.07
cc_188 VPB N_D_c_848_n 0.0225192f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_189 VPB N_D_M1035_g 0.00318633f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_190 VPB N_D_c_850_n 0.00784376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_D_c_851_n 0.042205f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_192 VPB N_A_211_363#_c_911_n 0.029172f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_193 VPB N_A_211_363#_c_912_n 0.0231835f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_194 VPB N_A_211_363#_c_893_n 0.0196492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_211_363#_c_894_n 0.00386093f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_196 VPB N_A_211_363#_c_915_n 0.0561794f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_197 VPB N_A_211_363#_c_916_n 0.00430496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_211_363#_c_907_n 2.53141e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_211_363#_c_910_n 0.0128307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1197_21#_M1025_g 0.0154962f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_201 VPB N_A_1197_21#_c_1131_n 0.0581122f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_202 VPB N_A_1197_21#_c_1132_n 0.00987662f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_203 VPB N_A_1197_21#_c_1133_n 0.0259332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_A_1197_21#_c_1134_n 0.00575753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_A_1197_21#_c_1126_n 0.00666344f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_206 VPB N_A_1197_21#_c_1136_n 0.00635064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_A_1197_21#_c_1129_n 0.00787197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_1270_n 0.0340648f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.07
cc_209 VPB N_SET_B_c_1282_n 0.0235956f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.4
cc_210 VPB N_SET_B_c_1272_n 0.0334405f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_211 VPB N_SET_B_c_1284_n 0.0229713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1003_47#_c_1400_n 0.04097f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.135
cc_213 VPB N_A_1003_47#_c_1406_n 0.0123514f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_214 VPB N_A_1003_47#_c_1403_n 0.00805778f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_215 VPB N_A_1003_47#_c_1404_n 0.00302582f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.53
cc_216 VPB N_A_1525_21#_c_1516_n 0.0177579f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_217 VPB N_A_1525_21#_c_1517_n 0.0174941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1525_21#_c_1518_n 0.00109772f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_219 VPB N_A_1525_21#_c_1519_n 0.00655658f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_220 VPB N_A_1525_21#_c_1512_n 0.00163792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1525_21#_c_1521_n 0.0348043f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_1525_21#_c_1522_n 0.00261931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1525_21#_c_1523_n 0.00860559f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1525_21#_c_1524_n 0.00357303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1525_21#_c_1513_n 0.0286231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1525_21#_c_1514_n 0.0356097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1525_21#_c_1515_n 0.00149955f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_2058_21#_M1014_g 0.016378f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_229 VPB N_A_2058_21#_c_1674_n 0.0597226f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_230 VPB N_A_2058_21#_c_1663_n 0.0309364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_2058_21#_c_1667_n 0.0147366f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_232 VPB N_A_2058_21#_c_1677_n 0.0203315f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_233 VPB N_A_2058_21#_c_1678_n 0.0222659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_2058_21#_c_1679_n 0.0044592f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_2058_21#_c_1680_n 0.00304218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_2058_21#_c_1671_n 0.00355641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_2058_21#_c_1682_n 0.00738916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_2058_21#_c_1683_n 0.00169275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_2058_21#_c_1672_n 2.41561e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_1864_47#_c_1845_n 0.0349234f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.135
cc_241 VPB N_A_1864_47#_c_1852_n 0.0119786f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.235
cc_242 VPB N_A_1864_47#_c_1848_n 0.00624517f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_243 VPB N_A_1864_47#_c_1849_n 7.65226e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_244 VPB N_A_1864_47#_c_1850_n 0.00126723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_RESET_B_c_1940_n 0.0372403f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.88
cc_246 VPB N_RESET_B_c_1942_n 0.0016954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_A_2845_47#_c_1972_n 0.0333263f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.135
cc_248 VPB N_A_2845_47#_c_1978_n 0.00101005f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.805
cc_249 VPB N_A_2845_47#_c_1979_n 0.00191687f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=1.665
cc_250 VPB N_A_2845_47#_c_1975_n 0.00574119f $X=-0.19 $Y=1.305 $X2=0.24
+ $Y2=1.235
cc_251 VPB N_A_2845_47#_c_1981_n 0.00668049f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.19
cc_252 VPB N_VPWR_c_2028_n 0.00108335f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_2029_n 0.0181798f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_2030_n 0.00852905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_2031_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_2032_n 0.00319272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_2033_n 0.00562899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_2034_n 0.00366828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_2035_n 0.0451296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_2036_n 0.00502902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_2037_n 0.0335239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_2038_n 0.00476476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_2039_n 0.0154511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_2040_n 0.0603463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_2041_n 0.0336449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_2042_n 0.0660042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_2043_n 0.00419147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_2044_n 0.035015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_2045_n 0.0175273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_2027_n 0.0780946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_2047_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_2048_n 0.00535993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_2049_n 0.00615406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_2050_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_2051_n 0.00939565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_2052_n 0.0257275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_2053_n 0.00446479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_A_483_47#_c_2248_n 0.00569182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_A_483_47#_c_2249_n 0.00673857f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_280 VPB N_A_483_47#_c_2242_n 0.00237862f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.07
cc_281 VPB N_A_483_47#_c_2244_n 3.39779e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_A_483_47#_c_2245_n 0.0033882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_A_483_47#_c_2246_n 0.00134466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_A_483_47#_c_2247_n 0.0126288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_Q_N_c_2380_n 0.015633f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_286 VPB Q_N 9.76594e-19 $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_287 VPB N_Q_c_2413_n 0.00558658f $X=-0.19 $Y=1.305 $X2=0.3 $Y2=0.805
cc_288 VPB N_Q_c_2411_n 0.0142359f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB Q 0.0287471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 N_CLK_c_298_n N_A_27_47#_c_344_n 0.00668884f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_291 CLK N_A_27_47#_c_344_n 7.96209e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_292 N_CLK_c_295_n N_A_27_47#_c_344_n 0.00257439f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_293 N_CLK_c_298_n N_A_27_47#_c_345_n 0.0193438f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_294 N_CLK_c_292_n N_A_27_47#_M1001_g 0.0154215f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_295 N_CLK_c_296_n N_A_27_47#_M1001_g 0.00188341f $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_296 N_CLK_c_292_n N_A_27_47#_c_338_n 0.0064334f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_297 N_CLK_c_293_n N_A_27_47#_c_338_n 0.0110008f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_298 CLK N_A_27_47#_c_338_n 0.00698378f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_299 N_CLK_c_293_n N_A_27_47#_c_339_n 0.00621081f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_300 CLK N_A_27_47#_c_339_n 0.0148236f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_301 N_CLK_c_295_n N_A_27_47#_c_339_n 3.2891e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_302 N_CLK_c_298_n N_A_27_47#_c_351_n 0.0172023f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_303 CLK N_A_27_47#_c_351_n 0.00693999f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_304 N_CLK_c_298_n N_A_27_47#_c_340_n 0.00449089f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_305 N_CLK_c_293_n N_A_27_47#_c_340_n 0.00198234f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_306 CLK N_A_27_47#_c_340_n 0.0429447f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_307 N_CLK_c_295_n N_A_27_47#_c_340_n 7.54672e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_308 N_CLK_c_296_n N_A_27_47#_c_340_n 5.50669e-19 $X=0.24 $Y=1.07 $X2=0 $Y2=0
cc_309 N_CLK_c_298_n N_A_27_47#_c_354_n 0.00818228f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_310 CLK N_A_27_47#_c_354_n 0.0157801f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_311 N_CLK_c_295_n N_A_27_47#_c_354_n 2.59784e-19 $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_312 N_CLK_c_298_n N_A_27_47#_c_356_n 0.00104874f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_313 CLK N_A_27_47#_c_343_n 0.00184694f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_314 N_CLK_c_295_n N_A_27_47#_c_343_n 0.0131315f $X=0.24 $Y=1.235 $X2=0 $Y2=0
cc_315 N_CLK_c_298_n N_VPWR_c_2028_n 0.0125197f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_316 N_CLK_c_298_n N_VPWR_c_2039_n 0.00304525f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_317 N_CLK_c_298_n N_VPWR_c_2027_n 0.00454898f $X=0.495 $Y=1.74 $X2=0 $Y2=0
cc_318 N_CLK_c_292_n N_VGND_c_2438_n 0.00198377f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_319 N_CLK_c_293_n N_VGND_c_2438_n 6.54873e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_320 N_CLK_c_292_n N_VGND_c_2444_n 0.00367064f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_321 N_CLK_c_292_n N_VGND_c_2445_n 0.0142867f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_322 N_A_27_47#_c_355_n N_SCD_c_591_n 0.00771316f $X=5.085 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_323 N_A_27_47#_c_355_n SCD 0.00953786f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_355_n N_SCD_c_594_n 0.00279472f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_325 N_A_27_47#_c_343_n N_SCD_c_594_n 0.00611744f $X=0.99 $Y=1.235 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_355_n N_A_453_315#_c_634_n 0.00930383f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_355_n N_A_453_315#_c_635_n 0.00802107f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_355_n N_A_453_315#_c_636_n 4.59039e-19 $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_355_n N_A_453_315#_c_637_n 0.00712494f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_355_n N_A_453_315#_c_638_n 0.0154757f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_355_n N_A_453_315#_c_640_n 0.0162289f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_355_n N_SCE_c_739_n 0.00274302f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_355_n N_SCE_c_748_n 0.0114282f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_355_n N_SCE_c_750_n 0.00455867f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_355_n SCE 0.0170101f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_336 N_A_27_47#_c_355_n N_D_c_847_n 0.00157584f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_355_n N_D_c_848_n 0.00122534f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_334_n N_D_M1035_g 0.0258618f $X=4.94 $Y=0.705 $X2=0 $Y2=0
cc_339 N_A_27_47#_c_355_n N_D_c_850_n 0.0281754f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_340 N_A_27_47#_c_355_n N_D_c_851_n 0.00132861f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_341 N_A_27_47#_c_355_n N_A_211_363#_M1038_d 9.36802e-19 $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_346_n N_A_211_363#_c_911_n 0.0230152f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_341_n N_A_211_363#_c_911_n 0.0062194f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_355_n N_A_211_363#_c_911_n 0.00493484f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_361_n N_A_211_363#_c_911_n 0.00800436f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_346_n N_A_211_363#_c_912_n 0.0127701f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_347 N_A_27_47#_c_355_n N_A_211_363#_c_912_n 0.00228218f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_358_n N_A_211_363#_c_912_n 5.32023e-19 $X=5.375 $Y=1.87
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_361_n N_A_211_363#_c_912_n 0.00321127f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_350 N_A_27_47#_c_346_n N_A_211_363#_c_893_n 0.0245098f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_351 N_A_27_47#_c_341_n N_A_211_363#_c_893_n 0.0105477f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_352 N_A_27_47#_c_357_n N_A_211_363#_c_893_n 3.79612e-19 $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_361_n N_A_211_363#_c_893_n 0.00709305f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_354 N_A_27_47#_c_341_n N_A_211_363#_c_894_n 0.00300385f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_355 N_A_27_47#_c_342_n N_A_211_363#_c_894_n 0.0266356f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_356 N_A_27_47#_c_334_n N_A_211_363#_M1019_g 0.0114115f $X=4.94 $Y=0.705 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_341_n N_A_211_363#_M1019_g 4.47076e-19 $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_358 N_A_27_47#_c_342_n N_A_211_363#_M1019_g 0.0215755f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_359 N_A_27_47#_M1046_g N_A_211_363#_c_897_n 0.015077f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_348_n N_A_211_363#_c_915_n 0.0363699f $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_361 N_A_27_47#_c_335_n N_A_211_363#_c_915_n 0.0245423f $X=9.81 $Y=1.32 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_359_n N_A_211_363#_c_915_n 0.00343993f $X=9.26 $Y=1.87 $X2=0
+ $Y2=0
cc_363 N_A_27_47#_c_362_n N_A_211_363#_c_915_n 0.00189925f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_364 N_A_27_47#_c_336_n N_A_211_363#_c_898_n 3.14726e-19 $X=9.38 $Y=1.32 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_M1046_g N_A_211_363#_c_898_n 0.00307895f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_c_336_n N_A_211_363#_c_899_n 0.0242058f $X=9.38 $Y=1.32 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_M1046_g N_A_211_363#_c_899_n 0.017261f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_c_335_n N_A_211_363#_c_900_n 0.0121244f $X=9.81 $Y=1.32 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_c_336_n N_A_211_363#_c_900_n 0.005116f $X=9.38 $Y=1.32 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1046_g N_A_211_363#_c_900_n 0.00646476f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_362_n N_A_211_363#_c_900_n 0.00677084f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_c_347_n N_A_211_363#_c_916_n 0.00545761f $X=9.28 $Y=1.575
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_c_348_n N_A_211_363#_c_916_n 9.69034e-19 $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_374 N_A_27_47#_c_335_n N_A_211_363#_c_916_n 0.00968845f $X=9.81 $Y=1.32 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_359_n N_A_211_363#_c_916_n 0.00468874f $X=9.26 $Y=1.87 $X2=0
+ $Y2=0
cc_376 N_A_27_47#_c_362_n N_A_211_363#_c_916_n 0.0132738f $X=9.195 $Y=1.74 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_341_n N_A_211_363#_c_901_n 0.018011f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_378 N_A_27_47#_c_342_n N_A_211_363#_c_901_n 0.00555754f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_M1001_g N_A_211_363#_c_902_n 0.00662116f $X=0.99 $Y=0.445
+ $X2=0 $Y2=0
cc_380 N_A_27_47#_c_338_n N_A_211_363#_c_902_n 0.00218461f $X=0.655 $Y=0.72
+ $X2=0 $Y2=0
cc_381 N_A_27_47#_c_340_n N_A_211_363#_c_902_n 0.0050932f $X=0.8 $Y=1.235 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_341_n N_A_211_363#_c_903_n 0.0090349f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_348_n N_A_211_363#_c_904_n 2.37019e-19 $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_357_n N_A_211_363#_c_905_n 0.124057f $X=9.115 $Y=1.87 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_341_n N_A_211_363#_c_906_n 4.33096e-19 $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_336_n N_A_211_363#_c_907_n 0.00131409f $X=9.38 $Y=1.32 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_362_n N_A_211_363#_c_907_n 0.00151402f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_388 N_A_27_47#_c_341_n N_A_211_363#_c_908_n 0.00709421f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_334_n N_A_211_363#_c_909_n 4.98615e-19 $X=4.94 $Y=0.705
+ $X2=0 $Y2=0
cc_390 N_A_27_47#_c_346_n N_A_211_363#_c_909_n 3.55508e-19 $X=5.435 $Y=1.99
+ $X2=0 $Y2=0
cc_391 N_A_27_47#_c_341_n N_A_211_363#_c_909_n 0.0213902f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_342_n N_A_211_363#_c_909_n 0.00158268f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_361_n N_A_211_363#_c_909_n 0.00503336f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_345_n N_A_211_363#_c_910_n 0.00704502f $X=0.965 $Y=1.74
+ $X2=0 $Y2=0
cc_395 N_A_27_47#_M1001_g N_A_211_363#_c_910_n 0.0222495f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_338_n N_A_211_363#_c_910_n 0.00926283f $X=0.655 $Y=0.72
+ $X2=0 $Y2=0
cc_397 N_A_27_47#_c_463_p N_A_211_363#_c_910_n 0.00824887f $X=0.77 $Y=1.795
+ $X2=0 $Y2=0
cc_398 N_A_27_47#_c_340_n N_A_211_363#_c_910_n 0.0569443f $X=0.8 $Y=1.235 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_355_n N_A_211_363#_c_910_n 0.0249106f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_356_n N_A_211_363#_c_910_n 0.00203677f $X=0.885 $Y=1.87
+ $X2=0 $Y2=0
cc_401 N_A_27_47#_c_346_n N_A_1197_21#_c_1131_n 0.025095f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_402 N_A_27_47#_c_357_n N_A_1197_21#_c_1131_n 0.00386067f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_336_n N_A_1197_21#_c_1132_n 0.00250207f $X=9.38 $Y=1.32
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_c_347_n N_A_1197_21#_c_1133_n 0.00256251f $X=9.28 $Y=1.575
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_c_348_n N_A_1197_21#_c_1133_n 0.0234456f $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_406 N_A_27_47#_c_357_n N_A_1197_21#_c_1133_n 0.00860239f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_c_362_n N_A_1197_21#_c_1133_n 0.00251036f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_c_357_n N_A_1197_21#_c_1134_n 0.0264788f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_357_n N_A_1197_21#_c_1146_n 0.0305977f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_357_n N_A_1197_21#_c_1136_n 0.0168828f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_357_n N_A_1197_21#_c_1148_n 0.00959465f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_412 N_A_27_47#_c_336_n N_A_1197_21#_c_1129_n 0.00276634f $X=9.38 $Y=1.32
+ $X2=0 $Y2=0
cc_413 N_A_27_47#_M1046_g N_SET_B_c_1274_n 0.00588147f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_c_346_n N_A_1003_47#_c_1409_n 0.0125372f $X=5.435 $Y=1.99
+ $X2=0 $Y2=0
cc_415 N_A_27_47#_c_355_n N_A_1003_47#_c_1409_n 2.16481e-19 $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_416 N_A_27_47#_c_357_n N_A_1003_47#_c_1409_n 0.00528022f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_417 N_A_27_47#_c_358_n N_A_1003_47#_c_1409_n 0.00304252f $X=5.375 $Y=1.87
+ $X2=0 $Y2=0
cc_418 N_A_27_47#_c_361_n N_A_1003_47#_c_1409_n 0.0168604f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_c_334_n N_A_1003_47#_c_1414_n 0.00310961f $X=4.94 $Y=0.705
+ $X2=0 $Y2=0
cc_420 N_A_27_47#_c_341_n N_A_1003_47#_c_1414_n 0.0070258f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_342_n N_A_1003_47#_c_1414_n 9.58359e-19 $X=5.07 $Y=0.87
+ $X2=0 $Y2=0
cc_422 N_A_27_47#_c_346_n N_A_1003_47#_c_1406_n 0.00861559f $X=5.435 $Y=1.99
+ $X2=0 $Y2=0
cc_423 N_A_27_47#_c_341_n N_A_1003_47#_c_1406_n 0.00627038f $X=5.07 $Y=0.87
+ $X2=0 $Y2=0
cc_424 N_A_27_47#_c_357_n N_A_1003_47#_c_1406_n 0.013911f $X=9.115 $Y=1.87 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_c_358_n N_A_1003_47#_c_1406_n 0.00140757f $X=5.375 $Y=1.87
+ $X2=0 $Y2=0
cc_426 N_A_27_47#_c_361_n N_A_1003_47#_c_1406_n 0.028593f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_357_n N_A_1003_47#_c_1403_n 0.0037128f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_428 N_A_27_47#_c_341_n N_A_1003_47#_c_1404_n 0.00673762f $X=5.07 $Y=0.87
+ $X2=0 $Y2=0
cc_429 N_A_27_47#_c_357_n N_A_1003_47#_c_1404_n 0.0047069f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_430 N_A_27_47#_c_357_n N_A_1525_21#_c_1516_n 0.00714084f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_431 N_A_27_47#_c_357_n N_A_1525_21#_c_1512_n 0.00482524f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_432 N_A_27_47#_c_347_n N_A_1525_21#_c_1521_n 0.00403803f $X=9.28 $Y=1.575
+ $X2=0 $Y2=0
cc_433 N_A_27_47#_c_348_n N_A_1525_21#_c_1521_n 0.00251754f $X=9.28 $Y=1.99
+ $X2=0 $Y2=0
cc_434 N_A_27_47#_c_335_n N_A_1525_21#_c_1521_n 0.00399632f $X=9.81 $Y=1.32
+ $X2=0 $Y2=0
cc_435 N_A_27_47#_c_357_n N_A_1525_21#_c_1521_n 0.0139809f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_436 N_A_27_47#_c_359_n N_A_1525_21#_c_1521_n 0.0254967f $X=9.26 $Y=1.87 $X2=0
+ $Y2=0
cc_437 N_A_27_47#_c_362_n N_A_1525_21#_c_1521_n 0.00664405f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_438 N_A_27_47#_c_347_n N_A_1525_21#_c_1522_n 7.54777e-19 $X=9.28 $Y=1.575
+ $X2=0 $Y2=0
cc_439 N_A_27_47#_c_348_n N_A_1525_21#_c_1522_n 8.27492e-19 $X=9.28 $Y=1.99
+ $X2=0 $Y2=0
cc_440 N_A_27_47#_c_357_n N_A_1525_21#_c_1522_n 0.0264578f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_441 N_A_27_47#_c_362_n N_A_1525_21#_c_1522_n 0.00130051f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_442 N_A_27_47#_c_347_n N_A_1525_21#_c_1523_n 0.00291473f $X=9.28 $Y=1.575
+ $X2=0 $Y2=0
cc_443 N_A_27_47#_c_348_n N_A_1525_21#_c_1523_n 7.11393e-19 $X=9.28 $Y=1.99
+ $X2=0 $Y2=0
cc_444 N_A_27_47#_c_357_n N_A_1525_21#_c_1523_n 0.0232209f $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_445 N_A_27_47#_c_362_n N_A_1525_21#_c_1523_n 0.00461714f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_446 N_A_27_47#_c_357_n N_A_1525_21#_c_1513_n 2.01181e-19 $X=9.115 $Y=1.87
+ $X2=0 $Y2=0
cc_447 N_A_27_47#_M1046_g N_A_2058_21#_M1014_g 0.0419655f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_448 N_A_27_47#_c_348_n N_A_1864_47#_c_1856_n 0.0104855f $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_449 N_A_27_47#_c_359_n N_A_1864_47#_c_1856_n 0.00169636f $X=9.26 $Y=1.87
+ $X2=0 $Y2=0
cc_450 N_A_27_47#_c_362_n N_A_1864_47#_c_1856_n 0.00161459f $X=9.195 $Y=1.74
+ $X2=0 $Y2=0
cc_451 N_A_27_47#_M1046_g N_A_1864_47#_c_1859_n 0.0128856f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_452 N_A_27_47#_M1046_g N_A_1864_47#_c_1847_n 0.0108297f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_453 N_A_27_47#_M1046_g N_A_1864_47#_c_1849_n 0.00157629f $X=9.885 $Y=0.415
+ $X2=0 $Y2=0
cc_454 N_A_27_47#_c_463_p N_VPWR_M1008_d 7.61525e-19 $X=0.77 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_455 N_A_27_47#_c_356_n N_VPWR_M1008_d 0.00206123f $X=0.885 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_456 N_A_27_47#_c_357_n N_VPWR_M1026_d 0.00710907f $X=9.115 $Y=1.87 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_c_345_n N_VPWR_c_2028_n 0.00869689f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_351_n N_VPWR_c_2028_n 0.00677095f $X=0.655 $Y=1.88 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_463_p N_VPWR_c_2028_n 0.0134205f $X=0.77 $Y=1.795 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_c_354_n N_VPWR_c_2028_n 0.0247016f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_355_n N_VPWR_c_2028_n 2.78216e-19 $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_356_n N_VPWR_c_2028_n 0.00350579f $X=0.885 $Y=1.87 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_345_n N_VPWR_c_2029_n 0.00590576f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_345_n N_VPWR_c_2030_n 0.00239371f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_465 N_A_27_47#_c_355_n N_VPWR_c_2030_n 0.0167602f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_355_n N_VPWR_c_2031_n 0.00472704f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_357_n N_VPWR_c_2032_n 0.00161496f $X=9.115 $Y=1.87 $X2=0
+ $Y2=0
cc_468 N_A_27_47#_c_357_n N_VPWR_c_2033_n 0.0137936f $X=9.115 $Y=1.87 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_c_351_n N_VPWR_c_2039_n 0.00180073f $X=0.655 $Y=1.88 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_354_n N_VPWR_c_2039_n 0.0123893f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_471 N_A_27_47#_c_346_n N_VPWR_c_2040_n 0.00440543f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_c_348_n N_VPWR_c_2042_n 0.00509845f $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_362_n N_VPWR_c_2042_n 0.00254851f $X=9.195 $Y=1.74 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_345_n N_VPWR_c_2027_n 0.00667006f $X=0.965 $Y=1.74 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_346_n N_VPWR_c_2027_n 0.00644068f $X=5.435 $Y=1.99 $X2=0
+ $Y2=0
cc_476 N_A_27_47#_c_348_n N_VPWR_c_2027_n 0.00749179f $X=9.28 $Y=1.99 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_351_n N_VPWR_c_2027_n 0.00415297f $X=0.655 $Y=1.88 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_354_n N_VPWR_c_2027_n 0.00665993f $X=0.26 $Y=1.96 $X2=0
+ $Y2=0
cc_479 N_A_27_47#_c_355_n N_VPWR_c_2027_n 0.202503f $X=5.085 $Y=1.87 $X2=0 $Y2=0
cc_480 N_A_27_47#_c_356_n N_VPWR_c_2027_n 0.0144885f $X=0.885 $Y=1.87 $X2=0
+ $Y2=0
cc_481 N_A_27_47#_c_357_n N_VPWR_c_2027_n 0.175811f $X=9.115 $Y=1.87 $X2=0 $Y2=0
cc_482 N_A_27_47#_c_358_n N_VPWR_c_2027_n 0.0160213f $X=5.375 $Y=1.87 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_c_359_n N_VPWR_c_2027_n 0.0147655f $X=9.26 $Y=1.87 $X2=0 $Y2=0
cc_484 N_A_27_47#_c_361_n N_VPWR_c_2027_n 0.00113432f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_c_362_n N_VPWR_c_2027_n 0.00133703f $X=9.195 $Y=1.74 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_c_355_n A_409_363# 0.00326461f $X=5.085 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_487 N_A_27_47#_c_355_n N_A_483_47#_c_2248_n 0.0182434f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_c_355_n N_A_483_47#_c_2249_n 0.0104101f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_c_355_n N_A_483_47#_c_2242_n 0.00714524f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_490 N_A_27_47#_c_355_n N_A_483_47#_c_2243_n 0.0567945f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_355_n N_A_483_47#_c_2244_n 0.0128797f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_492 N_A_27_47#_c_355_n N_A_483_47#_c_2245_n 0.00118055f $X=5.085 $Y=1.87
+ $X2=0 $Y2=0
cc_493 N_A_27_47#_c_341_n N_A_483_47#_c_2246_n 0.00752556f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_494 N_A_27_47#_c_355_n N_A_483_47#_c_2246_n 0.0136396f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_334_n N_A_483_47#_c_2247_n 0.0047291f $X=4.94 $Y=0.705 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_341_n N_A_483_47#_c_2247_n 0.0617482f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_497 N_A_27_47#_c_355_n N_A_483_47#_c_2247_n 0.0147343f $X=5.085 $Y=1.87 $X2=0
+ $Y2=0
cc_498 N_A_27_47#_c_358_n N_A_483_47#_c_2247_n 0.00171417f $X=5.375 $Y=1.87
+ $X2=0 $Y2=0
cc_499 N_A_27_47#_c_361_n N_A_483_47#_c_2247_n 0.0280654f $X=5.44 $Y=1.74 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_357_n A_1469_329# 0.00136307f $X=9.115 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_501 N_A_27_47#_c_357_n A_1710_329# 0.0068742f $X=9.115 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_502 N_A_27_47#_c_338_n N_VGND_M1033_d 0.00225291f $X=0.655 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_503 N_A_27_47#_M1001_g N_VGND_c_2427_n 0.00585385f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_504 N_A_27_47#_M1001_g N_VGND_c_2428_n 0.00328499f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_505 N_A_27_47#_M1046_g N_VGND_c_2431_n 0.00126551f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_506 N_A_27_47#_c_334_n N_VGND_c_2434_n 0.00556304f $X=4.94 $Y=0.705 $X2=0
+ $Y2=0
cc_507 N_A_27_47#_c_341_n N_VGND_c_2434_n 0.00175476f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_508 N_A_27_47#_c_342_n N_VGND_c_2434_n 3.93869e-19 $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_509 N_A_27_47#_M1046_g N_VGND_c_2436_n 0.00359964f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_510 N_A_27_47#_c_576_p N_VGND_c_2438_n 0.00747191f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_c_338_n N_VGND_c_2438_n 0.00244154f $X=0.655 $Y=0.72 $X2=0
+ $Y2=0
cc_512 N_A_27_47#_M1033_s N_VGND_c_2444_n 0.00419975f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_M1001_g N_VGND_c_2444_n 0.0120602f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_334_n N_VGND_c_2444_n 0.00688389f $X=4.94 $Y=0.705 $X2=0
+ $Y2=0
cc_515 N_A_27_47#_M1046_g N_VGND_c_2444_n 0.00588101f $X=9.885 $Y=0.415 $X2=0
+ $Y2=0
cc_516 N_A_27_47#_c_576_p N_VGND_c_2444_n 0.00626856f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_517 N_A_27_47#_c_338_n N_VGND_c_2444_n 0.00622643f $X=0.655 $Y=0.72 $X2=0
+ $Y2=0
cc_518 N_A_27_47#_c_341_n N_VGND_c_2444_n 0.00170297f $X=5.07 $Y=0.87 $X2=0
+ $Y2=0
cc_519 N_A_27_47#_M1001_g N_VGND_c_2445_n 0.00176556f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_520 N_A_27_47#_c_576_p N_VGND_c_2445_n 0.00897766f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_338_n N_VGND_c_2445_n 0.0228386f $X=0.655 $Y=0.72 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_343_n N_VGND_c_2445_n 6.84395e-19 $X=0.99 $Y=1.235 $X2=0
+ $Y2=0
cc_523 N_SCD_c_591_n N_A_453_315#_c_634_n 0.0477472f $X=1.955 $Y=1.74 $X2=0
+ $Y2=0
cc_524 N_SCD_c_594_n N_A_453_315#_c_636_n 0.011013f $X=1.955 $Y=1.532 $X2=0
+ $Y2=0
cc_525 N_SCD_M1023_g N_SCE_c_737_n 0.0613403f $X=1.98 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_526 N_SCD_M1023_g N_SCE_c_757_n 0.00942128f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_527 N_SCD_M1023_g SCE 0.0111793f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_528 N_SCD_M1023_g SCE 0.0100631f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_529 SCD SCE 0.0500109f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_530 N_SCD_c_594_n SCE 0.0166287f $X=1.955 $Y=1.532 $X2=0 $Y2=0
cc_531 N_SCD_M1023_g N_A_211_363#_c_901_n 0.00398443f $X=1.98 $Y=0.445 $X2=0
+ $Y2=0
cc_532 SCD N_A_211_363#_c_901_n 0.010483f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_533 N_SCD_c_594_n N_A_211_363#_c_901_n 0.00310261f $X=1.955 $Y=1.532 $X2=0
+ $Y2=0
cc_534 N_SCD_M1023_g N_A_211_363#_c_902_n 0.00174175f $X=1.98 $Y=0.445 $X2=0
+ $Y2=0
cc_535 N_SCD_c_591_n N_A_211_363#_c_910_n 0.00304814f $X=1.955 $Y=1.74 $X2=0
+ $Y2=0
cc_536 N_SCD_M1023_g N_A_211_363#_c_910_n 0.00519945f $X=1.98 $Y=0.445 $X2=0
+ $Y2=0
cc_537 SCD N_A_211_363#_c_910_n 0.0522928f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_538 N_SCD_c_594_n N_A_211_363#_c_910_n 0.00238852f $X=1.955 $Y=1.532 $X2=0
+ $Y2=0
cc_539 N_SCD_c_591_n N_VPWR_c_2030_n 0.0156798f $X=1.955 $Y=1.74 $X2=0 $Y2=0
cc_540 SCD N_VPWR_c_2030_n 0.0127353f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_541 N_SCD_c_594_n N_VPWR_c_2030_n 0.00430073f $X=1.955 $Y=1.532 $X2=0 $Y2=0
cc_542 N_SCD_c_591_n N_VPWR_c_2035_n 0.00590576f $X=1.955 $Y=1.74 $X2=0 $Y2=0
cc_543 N_SCD_c_591_n N_VPWR_c_2027_n 0.0055323f $X=1.955 $Y=1.74 $X2=0 $Y2=0
cc_544 N_SCD_c_591_n N_A_483_47#_c_2248_n 0.00161423f $X=1.955 $Y=1.74 $X2=0
+ $Y2=0
cc_545 N_SCD_c_594_n N_A_483_47#_c_2249_n 0.00111228f $X=1.955 $Y=1.532 $X2=0
+ $Y2=0
cc_546 N_SCD_M1023_g N_A_483_47#_c_2242_n 9.19442e-19 $X=1.98 $Y=0.445 $X2=0
+ $Y2=0
cc_547 N_SCD_M1023_g N_VGND_c_2428_n 0.00782772f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_548 SCD N_VGND_c_2428_n 0.0053442f $X=1.525 $Y=1.105 $X2=0 $Y2=0
cc_549 N_SCD_c_594_n N_VGND_c_2428_n 0.00193326f $X=1.955 $Y=1.532 $X2=0 $Y2=0
cc_550 N_SCD_M1023_g N_VGND_c_2439_n 0.00436871f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_551 N_SCD_M1023_g N_VGND_c_2444_n 0.00685866f $X=1.98 $Y=0.445 $X2=0 $Y2=0
cc_552 N_A_453_315#_c_635_n N_SCE_c_738_n 0.00587794f $X=2.895 $Y=1.65 $X2=0
+ $Y2=0
cc_553 N_A_453_315#_c_638_n N_SCE_c_738_n 3.99161e-19 $X=3.725 $Y=1.66 $X2=0
+ $Y2=0
cc_554 N_A_453_315#_c_629_n N_SCE_c_738_n 0.00225992f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_555 N_A_453_315#_c_630_n N_SCE_c_738_n 0.00806346f $X=3.325 $Y=0.71 $X2=0
+ $Y2=0
cc_556 N_A_453_315#_c_635_n N_SCE_c_739_n 0.0214586f $X=2.895 $Y=1.65 $X2=0
+ $Y2=0
cc_557 N_A_453_315#_c_638_n N_SCE_c_739_n 0.0141257f $X=3.725 $Y=1.66 $X2=0
+ $Y2=0
cc_558 N_A_453_315#_c_632_n N_SCE_c_739_n 0.0107851f $X=3.81 $Y=1.575 $X2=0
+ $Y2=0
cc_559 N_A_453_315#_c_640_n N_SCE_c_739_n 0.00343121f $X=3.105 $Y=1.66 $X2=0
+ $Y2=0
cc_560 N_A_453_315#_c_637_n N_SCE_c_747_n 0.0135447f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_561 N_A_453_315#_c_628_n N_SCE_c_740_n 0.0106714f $X=4.045 $Y=0.765 $X2=0
+ $Y2=0
cc_562 N_A_453_315#_c_659_p N_SCE_c_740_n 0.00974544f $X=3.24 $Y=0.47 $X2=0
+ $Y2=0
cc_563 N_A_453_315#_c_629_n N_SCE_c_740_n 0.00847366f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_564 N_A_453_315#_c_638_n N_SCE_c_748_n 0.00717517f $X=3.725 $Y=1.66 $X2=0
+ $Y2=0
cc_565 N_A_453_315#_c_629_n N_SCE_c_741_n 0.00656532f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_566 N_A_453_315#_c_631_n N_SCE_c_741_n 0.0062658f $X=3.81 $Y=1.095 $X2=0
+ $Y2=0
cc_567 N_A_453_315#_c_633_n N_SCE_c_741_n 0.0209712f $X=4.045 $Y=0.93 $X2=0
+ $Y2=0
cc_568 N_A_453_315#_c_637_n N_SCE_c_750_n 0.00327215f $X=3.18 $Y=2.3 $X2=0 $Y2=0
cc_569 N_A_453_315#_c_636_n N_SCE_c_742_n 0.0015675f $X=2.465 $Y=1.65 $X2=0
+ $Y2=0
cc_570 N_A_453_315#_c_636_n SCE 0.00130778f $X=2.465 $Y=1.65 $X2=0 $Y2=0
cc_571 N_A_453_315#_c_636_n N_SCE_c_745_n 0.00966517f $X=2.465 $Y=1.65 $X2=0
+ $Y2=0
cc_572 N_A_453_315#_c_638_n N_D_c_847_n 6.30122e-19 $X=3.725 $Y=1.66 $X2=0 $Y2=0
cc_573 N_A_453_315#_c_628_n N_D_M1035_g 0.0493339f $X=4.045 $Y=0.765 $X2=0 $Y2=0
cc_574 N_A_453_315#_c_631_n N_D_M1035_g 0.00125372f $X=3.81 $Y=1.095 $X2=0 $Y2=0
cc_575 N_A_453_315#_c_632_n N_D_M1035_g 0.00450276f $X=3.81 $Y=1.575 $X2=0 $Y2=0
cc_576 N_A_453_315#_c_638_n N_D_c_850_n 0.0108667f $X=3.725 $Y=1.66 $X2=0 $Y2=0
cc_577 N_A_453_315#_c_632_n N_D_c_850_n 0.0137443f $X=3.81 $Y=1.575 $X2=0 $Y2=0
cc_578 N_A_453_315#_c_638_n N_D_c_851_n 5.53153e-19 $X=3.725 $Y=1.66 $X2=0 $Y2=0
cc_579 N_A_453_315#_c_632_n N_D_c_851_n 0.0021836f $X=3.81 $Y=1.575 $X2=0 $Y2=0
cc_580 N_A_453_315#_c_633_n N_D_c_851_n 0.00265425f $X=4.045 $Y=0.93 $X2=0 $Y2=0
cc_581 N_A_453_315#_c_629_n N_A_211_363#_c_901_n 0.0158576f $X=3.725 $Y=0.71
+ $X2=0 $Y2=0
cc_582 N_A_453_315#_c_630_n N_A_211_363#_c_901_n 0.00794081f $X=3.325 $Y=0.71
+ $X2=0 $Y2=0
cc_583 N_A_453_315#_c_631_n N_A_211_363#_c_901_n 0.0233655f $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_584 N_A_453_315#_c_633_n N_A_211_363#_c_901_n 0.00194022f $X=4.045 $Y=0.93
+ $X2=0 $Y2=0
cc_585 N_A_453_315#_c_634_n N_VPWR_c_2030_n 0.00263268f $X=2.365 $Y=1.74 $X2=0
+ $Y2=0
cc_586 N_A_453_315#_c_637_n N_VPWR_c_2031_n 0.0140911f $X=3.18 $Y=2.3 $X2=0
+ $Y2=0
cc_587 N_A_453_315#_c_638_n N_VPWR_c_2031_n 0.00573442f $X=3.725 $Y=1.66 $X2=0
+ $Y2=0
cc_588 N_A_453_315#_c_634_n N_VPWR_c_2035_n 0.00573288f $X=2.365 $Y=1.74 $X2=0
+ $Y2=0
cc_589 N_A_453_315#_c_637_n N_VPWR_c_2035_n 0.0118139f $X=3.18 $Y=2.3 $X2=0
+ $Y2=0
cc_590 N_A_453_315#_M1011_s N_VPWR_c_2027_n 0.00347325f $X=3.055 $Y=2.065 $X2=0
+ $Y2=0
cc_591 N_A_453_315#_c_634_n N_VPWR_c_2027_n 0.00756413f $X=2.365 $Y=1.74 $X2=0
+ $Y2=0
cc_592 N_A_453_315#_c_635_n N_VPWR_c_2027_n 2.96327e-19 $X=2.895 $Y=1.65 $X2=0
+ $Y2=0
cc_593 N_A_453_315#_c_637_n N_VPWR_c_2027_n 0.00308197f $X=3.18 $Y=2.3 $X2=0
+ $Y2=0
cc_594 N_A_453_315#_c_640_n N_VPWR_c_2027_n 0.00196684f $X=3.105 $Y=1.66 $X2=0
+ $Y2=0
cc_595 N_A_453_315#_c_659_p N_A_483_47#_c_2240_n 0.00220866f $X=3.24 $Y=0.47
+ $X2=0 $Y2=0
cc_596 N_A_453_315#_c_630_n N_A_483_47#_c_2240_n 0.0136508f $X=3.325 $Y=0.71
+ $X2=0 $Y2=0
cc_597 N_A_453_315#_c_634_n N_A_483_47#_c_2248_n 0.0125435f $X=2.365 $Y=1.74
+ $X2=0 $Y2=0
cc_598 N_A_453_315#_c_635_n N_A_483_47#_c_2248_n 0.00245011f $X=2.895 $Y=1.65
+ $X2=0 $Y2=0
cc_599 N_A_453_315#_c_636_n N_A_483_47#_c_2248_n 2.71208e-19 $X=2.465 $Y=1.65
+ $X2=0 $Y2=0
cc_600 N_A_453_315#_c_637_n N_A_483_47#_c_2248_n 0.0233473f $X=3.18 $Y=2.3 $X2=0
+ $Y2=0
cc_601 N_A_453_315#_c_634_n N_A_483_47#_c_2249_n 0.0028028f $X=2.365 $Y=1.74
+ $X2=0 $Y2=0
cc_602 N_A_453_315#_c_635_n N_A_483_47#_c_2249_n 0.017747f $X=2.895 $Y=1.65
+ $X2=0 $Y2=0
cc_603 N_A_453_315#_c_636_n N_A_483_47#_c_2249_n 3.92738e-19 $X=2.465 $Y=1.65
+ $X2=0 $Y2=0
cc_604 N_A_453_315#_c_640_n N_A_483_47#_c_2249_n 0.0225927f $X=3.105 $Y=1.66
+ $X2=0 $Y2=0
cc_605 N_A_453_315#_c_659_p N_A_483_47#_c_2241_n 0.0232736f $X=3.24 $Y=0.47
+ $X2=0 $Y2=0
cc_606 N_A_453_315#_c_635_n N_A_483_47#_c_2242_n 0.00532216f $X=2.895 $Y=1.65
+ $X2=0 $Y2=0
cc_607 N_A_453_315#_c_640_n N_A_483_47#_c_2242_n 6.00227e-19 $X=3.105 $Y=1.66
+ $X2=0 $Y2=0
cc_608 N_A_453_315#_c_638_n N_A_483_47#_c_2243_n 0.00918036f $X=3.725 $Y=1.66
+ $X2=0 $Y2=0
cc_609 N_A_453_315#_c_629_n N_A_483_47#_c_2243_n 0.00373551f $X=3.725 $Y=0.71
+ $X2=0 $Y2=0
cc_610 N_A_453_315#_c_631_n N_A_483_47#_c_2243_n 0.00542999f $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_611 N_A_453_315#_c_632_n N_A_483_47#_c_2243_n 0.017493f $X=3.81 $Y=1.575
+ $X2=0 $Y2=0
cc_612 N_A_453_315#_c_633_n N_A_483_47#_c_2243_n 3.73132e-19 $X=4.045 $Y=0.93
+ $X2=0 $Y2=0
cc_613 N_A_453_315#_c_638_n N_A_483_47#_c_2244_n 0.00169392f $X=3.725 $Y=1.66
+ $X2=0 $Y2=0
cc_614 N_A_453_315#_c_630_n N_A_483_47#_c_2244_n 0.00141688f $X=3.325 $Y=0.71
+ $X2=0 $Y2=0
cc_615 N_A_453_315#_c_631_n N_A_483_47#_c_2244_n 5.39866e-19 $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_616 N_A_453_315#_c_632_n N_A_483_47#_c_2244_n 0.00177774f $X=3.81 $Y=1.575
+ $X2=0 $Y2=0
cc_617 N_A_453_315#_c_640_n N_A_483_47#_c_2244_n 9.72289e-19 $X=3.105 $Y=1.66
+ $X2=0 $Y2=0
cc_618 N_A_453_315#_c_635_n N_A_483_47#_c_2245_n 0.00101345f $X=2.895 $Y=1.65
+ $X2=0 $Y2=0
cc_619 N_A_453_315#_c_638_n N_A_483_47#_c_2245_n 5.57877e-19 $X=3.725 $Y=1.66
+ $X2=0 $Y2=0
cc_620 N_A_453_315#_c_630_n N_A_483_47#_c_2245_n 0.00610396f $X=3.325 $Y=0.71
+ $X2=0 $Y2=0
cc_621 N_A_453_315#_c_631_n N_A_483_47#_c_2245_n 4.87843e-19 $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_622 N_A_453_315#_c_632_n N_A_483_47#_c_2245_n 0.00788805f $X=3.81 $Y=1.575
+ $X2=0 $Y2=0
cc_623 N_A_453_315#_c_640_n N_A_483_47#_c_2245_n 0.0185169f $X=3.105 $Y=1.66
+ $X2=0 $Y2=0
cc_624 N_A_453_315#_c_631_n N_A_483_47#_c_2246_n 4.58758e-19 $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_625 N_A_453_315#_c_631_n N_A_483_47#_c_2247_n 0.0075454f $X=3.81 $Y=1.095
+ $X2=0 $Y2=0
cc_626 N_A_453_315#_c_629_n N_VGND_M1003_d 8.04166e-19 $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_627 N_A_453_315#_c_631_n N_VGND_M1003_d 0.00224031f $X=3.81 $Y=1.095 $X2=0
+ $Y2=0
cc_628 N_A_453_315#_c_628_n N_VGND_c_2429_n 0.00322018f $X=4.045 $Y=0.765 $X2=0
+ $Y2=0
cc_629 N_A_453_315#_c_629_n N_VGND_c_2429_n 0.0051618f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_630 N_A_453_315#_c_631_n N_VGND_c_2429_n 0.0138714f $X=3.81 $Y=1.095 $X2=0
+ $Y2=0
cc_631 N_A_453_315#_c_633_n N_VGND_c_2429_n 7.64617e-19 $X=4.045 $Y=0.93 $X2=0
+ $Y2=0
cc_632 N_A_453_315#_c_628_n N_VGND_c_2434_n 0.00585385f $X=4.045 $Y=0.765 $X2=0
+ $Y2=0
cc_633 N_A_453_315#_c_659_p N_VGND_c_2439_n 0.0102832f $X=3.24 $Y=0.47 $X2=0
+ $Y2=0
cc_634 N_A_453_315#_c_629_n N_VGND_c_2439_n 0.00440669f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_635 N_A_453_315#_M1003_s N_VGND_c_2444_n 0.00248159f $X=3.115 $Y=0.235 $X2=0
+ $Y2=0
cc_636 N_A_453_315#_c_628_n N_VGND_c_2444_n 0.00602844f $X=4.045 $Y=0.765 $X2=0
+ $Y2=0
cc_637 N_A_453_315#_c_659_p N_VGND_c_2444_n 0.00346716f $X=3.24 $Y=0.47 $X2=0
+ $Y2=0
cc_638 N_A_453_315#_c_629_n N_VGND_c_2444_n 0.00360146f $X=3.725 $Y=0.71 $X2=0
+ $Y2=0
cc_639 N_A_453_315#_c_631_n N_VGND_c_2444_n 0.00312535f $X=3.81 $Y=1.095 $X2=0
+ $Y2=0
cc_640 N_SCE_c_748_n N_D_c_847_n 0.0076628f $X=3.86 $Y=1.91 $X2=0 $Y2=0
cc_641 N_SCE_c_749_n N_D_c_848_n 0.0259336f $X=3.96 $Y=1.99 $X2=0 $Y2=0
cc_642 N_SCE_c_739_n N_D_c_850_n 0.00246325f $X=3.49 $Y=1.835 $X2=0 $Y2=0
cc_643 N_SCE_c_748_n N_D_c_850_n 0.00351115f $X=3.86 $Y=1.91 $X2=0 $Y2=0
cc_644 N_SCE_c_749_n N_D_c_850_n 0.00710371f $X=3.96 $Y=1.99 $X2=0 $Y2=0
cc_645 N_SCE_c_739_n N_D_c_851_n 0.00482288f $X=3.49 $Y=1.835 $X2=0 $Y2=0
cc_646 N_SCE_c_738_n N_A_211_363#_c_901_n 0.00520043f $X=3.39 $Y=0.81 $X2=0
+ $Y2=0
cc_647 N_SCE_c_739_n N_A_211_363#_c_901_n 0.00295637f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_648 N_SCE_c_741_n N_A_211_363#_c_901_n 4.50186e-19 $X=3.49 $Y=0.81 $X2=0
+ $Y2=0
cc_649 N_SCE_c_742_n N_A_211_363#_c_901_n 0.0260043f $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_650 N_SCE_c_757_n N_A_211_363#_c_901_n 0.033409f $X=2.095 $Y=0.887 $X2=0
+ $Y2=0
cc_651 N_SCE_c_757_n N_A_211_363#_c_902_n 0.0014863f $X=2.095 $Y=0.887 $X2=0
+ $Y2=0
cc_652 SCE N_A_211_363#_c_902_n 5.29693e-19 $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_653 N_SCE_c_757_n N_A_211_363#_c_910_n 0.00445267f $X=2.095 $Y=0.887 $X2=0
+ $Y2=0
cc_654 SCE N_A_211_363#_c_910_n 0.003009f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_655 SCE N_A_211_363#_c_910_n 5.60605e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_656 N_SCE_c_747_n N_VPWR_c_2031_n 0.012739f $X=3.49 $Y=1.99 $X2=0 $Y2=0
cc_657 N_SCE_c_748_n N_VPWR_c_2031_n 0.00537624f $X=3.86 $Y=1.91 $X2=0 $Y2=0
cc_658 N_SCE_c_749_n N_VPWR_c_2031_n 0.00922413f $X=3.96 $Y=1.99 $X2=0 $Y2=0
cc_659 N_SCE_c_747_n N_VPWR_c_2035_n 0.00427505f $X=3.49 $Y=1.99 $X2=0 $Y2=0
cc_660 N_SCE_c_750_n N_VPWR_c_2035_n 2.07025e-19 $X=3.49 $Y=1.912 $X2=0 $Y2=0
cc_661 N_SCE_c_749_n N_VPWR_c_2040_n 0.00622633f $X=3.96 $Y=1.99 $X2=0 $Y2=0
cc_662 N_SCE_c_747_n N_VPWR_c_2027_n 0.00550264f $X=3.49 $Y=1.99 $X2=0 $Y2=0
cc_663 N_SCE_c_749_n N_VPWR_c_2027_n 0.00581056f $X=3.96 $Y=1.99 $X2=0 $Y2=0
cc_664 N_SCE_c_737_n N_A_483_47#_c_2240_n 0.00247913f $X=2.34 $Y=0.735 $X2=0
+ $Y2=0
cc_665 N_SCE_c_738_n N_A_483_47#_c_2240_n 0.0130093f $X=3.39 $Y=0.81 $X2=0 $Y2=0
cc_666 N_SCE_c_739_n N_A_483_47#_c_2240_n 0.00472997f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_667 N_SCE_c_740_n N_A_483_47#_c_2240_n 4.40509e-19 $X=3.515 $Y=0.735 $X2=0
+ $Y2=0
cc_668 N_SCE_c_742_n N_A_483_47#_c_2240_n 0.0174977f $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_669 SCE N_A_483_47#_c_2240_n 0.00460399f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_670 SCE N_A_483_47#_c_2240_n 0.00210109f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_671 N_SCE_c_745_n N_A_483_47#_c_2240_n 0.00236655f $X=2.585 $Y=0.915 $X2=0
+ $Y2=0
cc_672 N_SCE_c_739_n N_A_483_47#_c_2249_n 0.00475402f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_673 SCE N_A_483_47#_c_2249_n 0.0175986f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_674 N_SCE_c_737_n N_A_483_47#_c_2241_n 0.00868007f $X=2.34 $Y=0.735 $X2=0
+ $Y2=0
cc_675 N_SCE_c_738_n N_A_483_47#_c_2241_n 9.34339e-19 $X=3.39 $Y=0.81 $X2=0
+ $Y2=0
cc_676 N_SCE_c_740_n N_A_483_47#_c_2241_n 0.00110088f $X=3.515 $Y=0.735 $X2=0
+ $Y2=0
cc_677 N_SCE_c_742_n N_A_483_47#_c_2241_n 0.00361707f $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_678 N_SCE_c_745_n N_A_483_47#_c_2241_n 0.00650464f $X=2.585 $Y=0.915 $X2=0
+ $Y2=0
cc_679 N_SCE_c_738_n N_A_483_47#_c_2242_n 0.00119558f $X=3.39 $Y=0.81 $X2=0
+ $Y2=0
cc_680 N_SCE_c_742_n N_A_483_47#_c_2242_n 0.00424618f $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_681 SCE N_A_483_47#_c_2242_n 0.0151057f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_682 N_SCE_c_745_n N_A_483_47#_c_2242_n 9.23968e-19 $X=2.585 $Y=0.915 $X2=0
+ $Y2=0
cc_683 N_SCE_c_739_n N_A_483_47#_c_2243_n 0.00876769f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_684 N_SCE_c_748_n N_A_483_47#_c_2243_n 8.04245e-19 $X=3.86 $Y=1.91 $X2=0
+ $Y2=0
cc_685 N_SCE_c_738_n N_A_483_47#_c_2244_n 9.94869e-19 $X=3.39 $Y=0.81 $X2=0
+ $Y2=0
cc_686 N_SCE_c_739_n N_A_483_47#_c_2244_n 0.00239145f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_687 N_SCE_c_738_n N_A_483_47#_c_2245_n 0.0056856f $X=3.39 $Y=0.81 $X2=0 $Y2=0
cc_688 N_SCE_c_739_n N_A_483_47#_c_2245_n 0.0067276f $X=3.49 $Y=1.835 $X2=0
+ $Y2=0
cc_689 SCE N_VGND_c_2428_n 0.0217684f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_690 N_SCE_c_740_n N_VGND_c_2429_n 0.00315767f $X=3.515 $Y=0.735 $X2=0 $Y2=0
cc_691 N_SCE_c_737_n N_VGND_c_2439_n 0.00585385f $X=2.34 $Y=0.735 $X2=0 $Y2=0
cc_692 N_SCE_c_738_n N_VGND_c_2439_n 0.00335269f $X=3.39 $Y=0.81 $X2=0 $Y2=0
cc_693 N_SCE_c_740_n N_VGND_c_2439_n 0.0042361f $X=3.515 $Y=0.735 $X2=0 $Y2=0
cc_694 N_SCE_c_757_n N_VGND_c_2439_n 5.49067e-19 $X=2.095 $Y=0.887 $X2=0 $Y2=0
cc_695 SCE N_VGND_c_2439_n 0.010028f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_696 N_SCE_c_745_n N_VGND_c_2439_n 9.57457e-19 $X=2.585 $Y=0.915 $X2=0 $Y2=0
cc_697 N_SCE_c_737_n N_VGND_c_2444_n 0.00701375f $X=2.34 $Y=0.735 $X2=0 $Y2=0
cc_698 N_SCE_c_740_n N_VGND_c_2444_n 0.00702835f $X=3.515 $Y=0.735 $X2=0 $Y2=0
cc_699 N_SCE_c_742_n N_VGND_c_2444_n 0.00573209f $X=2.4 $Y=0.93 $X2=0 $Y2=0
cc_700 N_SCE_c_757_n N_VGND_c_2444_n 4.11623e-19 $X=2.095 $Y=0.887 $X2=0 $Y2=0
cc_701 SCE N_VGND_c_2444_n 0.0046728f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_702 N_SCE_c_745_n N_VGND_c_2444_n 0.00280721f $X=2.585 $Y=0.915 $X2=0 $Y2=0
cc_703 SCE A_411_47# 0.00112971f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_704 N_D_c_851_n N_A_211_363#_c_911_n 0.00804097f $X=4.455 $Y=1.49 $X2=0 $Y2=0
cc_705 N_D_c_847_n N_A_211_363#_c_912_n 0.00804097f $X=4.43 $Y=1.89 $X2=0 $Y2=0
cc_706 N_D_c_848_n N_A_211_363#_c_912_n 0.0130205f $X=4.43 $Y=1.99 $X2=0 $Y2=0
cc_707 N_D_M1035_g N_A_211_363#_c_894_n 0.00804097f $X=4.455 $Y=0.445 $X2=0
+ $Y2=0
cc_708 N_D_M1035_g N_A_211_363#_c_901_n 0.00651273f $X=4.455 $Y=0.445 $X2=0
+ $Y2=0
cc_709 N_D_c_848_n N_VPWR_c_2031_n 0.00158845f $X=4.43 $Y=1.99 $X2=0 $Y2=0
cc_710 N_D_c_850_n N_VPWR_c_2031_n 0.00890764f $X=4.24 $Y=1.49 $X2=0 $Y2=0
cc_711 N_D_c_848_n N_VPWR_c_2040_n 0.00538468f $X=4.43 $Y=1.99 $X2=0 $Y2=0
cc_712 N_D_c_850_n N_VPWR_c_2040_n 0.0126704f $X=4.24 $Y=1.49 $X2=0 $Y2=0
cc_713 N_D_c_848_n N_VPWR_c_2027_n 0.00683789f $X=4.43 $Y=1.99 $X2=0 $Y2=0
cc_714 N_D_c_850_n N_VPWR_c_2027_n 0.00524645f $X=4.24 $Y=1.49 $X2=0 $Y2=0
cc_715 N_D_M1035_g N_A_483_47#_c_2243_n 0.00815329f $X=4.455 $Y=0.445 $X2=0
+ $Y2=0
cc_716 N_D_c_850_n N_A_483_47#_c_2243_n 0.0132195f $X=4.24 $Y=1.49 $X2=0 $Y2=0
cc_717 N_D_c_851_n N_A_483_47#_c_2243_n 9.29241e-19 $X=4.455 $Y=1.49 $X2=0 $Y2=0
cc_718 N_D_M1035_g N_A_483_47#_c_2246_n 0.00191251f $X=4.455 $Y=0.445 $X2=0
+ $Y2=0
cc_719 N_D_c_848_n N_A_483_47#_c_2247_n 0.00478382f $X=4.43 $Y=1.99 $X2=0 $Y2=0
cc_720 N_D_M1035_g N_A_483_47#_c_2247_n 0.0256605f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_721 N_D_c_850_n N_A_483_47#_c_2247_n 0.0770577f $X=4.24 $Y=1.49 $X2=0 $Y2=0
cc_722 N_D_c_850_n A_810_413# 0.00495052f $X=4.24 $Y=1.49 $X2=-0.19 $Y2=-0.24
cc_723 N_D_M1035_g N_VGND_c_2434_n 0.00585385f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_724 N_D_M1035_g N_VGND_c_2444_n 0.00662578f $X=4.455 $Y=0.445 $X2=0 $Y2=0
cc_725 N_A_211_363#_M1019_g N_A_1197_21#_M1025_g 0.0207562f $X=5.53 $Y=0.415
+ $X2=0 $Y2=0
cc_726 N_A_211_363#_c_896_n N_A_1197_21#_M1025_g 0.0106463f $X=5.555 $Y=1.245
+ $X2=0 $Y2=0
cc_727 N_A_211_363#_c_904_n N_A_1197_21#_M1025_g 7.74803e-19 $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_728 N_A_211_363#_c_906_n N_A_1197_21#_M1025_g 0.00643317f $X=5.74 $Y=0.85
+ $X2=0 $Y2=0
cc_729 N_A_211_363#_c_908_n N_A_1197_21#_M1025_g 0.020124f $X=5.64 $Y=0.93 $X2=0
+ $Y2=0
cc_730 N_A_211_363#_c_909_n N_A_1197_21#_M1025_g 0.00197683f $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_731 N_A_211_363#_c_897_n N_A_1197_21#_c_1124_n 0.0188661f $X=9.245 $Y=0.705
+ $X2=0 $Y2=0
cc_732 N_A_211_363#_c_898_n N_A_1197_21#_c_1124_n 0.00171392f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_733 N_A_211_363#_c_904_n N_A_1197_21#_c_1134_n 0.00213216f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_734 N_A_211_363#_c_904_n N_A_1197_21#_c_1146_n 0.00443375f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_735 N_A_211_363#_c_904_n N_A_1197_21#_c_1125_n 0.00237294f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_736 N_A_211_363#_c_904_n N_A_1197_21#_c_1126_n 0.0167544f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_737 N_A_211_363#_c_904_n N_A_1197_21#_c_1127_n 0.00983915f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_738 N_A_211_363#_c_904_n N_A_1197_21#_c_1136_n 9.88695e-19 $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_739 N_A_211_363#_c_904_n N_A_1197_21#_c_1148_n 6.83984e-19 $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_740 N_A_211_363#_c_898_n N_A_1197_21#_c_1128_n 0.0114934f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_741 N_A_211_363#_c_899_n N_A_1197_21#_c_1128_n 9.54644e-19 $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_742 N_A_211_363#_c_900_n N_A_1197_21#_c_1128_n 0.00465767f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_743 N_A_211_363#_c_904_n N_A_1197_21#_c_1128_n 0.018108f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_744 N_A_211_363#_c_907_n N_A_1197_21#_c_1128_n 0.00130689f $X=9.26 $Y=1.19
+ $X2=0 $Y2=0
cc_745 N_A_211_363#_c_898_n N_A_1197_21#_c_1129_n 5.16236e-19 $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_746 N_A_211_363#_c_899_n N_A_1197_21#_c_1129_n 0.0188661f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_747 N_A_211_363#_c_900_n N_A_1197_21#_c_1129_n 0.00177719f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_748 N_A_211_363#_c_904_n N_A_1197_21#_c_1129_n 0.00431259f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_749 N_A_211_363#_c_907_n N_A_1197_21#_c_1129_n 6.96061e-19 $X=9.26 $Y=1.19
+ $X2=0 $Y2=0
cc_750 N_A_211_363#_c_904_n N_SET_B_c_1270_n 0.00124936f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_751 N_A_211_363#_c_898_n N_SET_B_c_1274_n 0.0224082f $X=9.37 $Y=0.87 $X2=0
+ $Y2=0
cc_752 N_A_211_363#_c_899_n N_SET_B_c_1274_n 0.00240552f $X=9.37 $Y=0.87 $X2=0
+ $Y2=0
cc_753 N_A_211_363#_c_900_n N_SET_B_c_1274_n 0.00615829f $X=9.762 $Y=1.305 $X2=0
+ $Y2=0
cc_754 N_A_211_363#_c_904_n N_SET_B_c_1274_n 0.181037f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_755 N_A_211_363#_c_907_n N_SET_B_c_1274_n 0.0254944f $X=9.26 $Y=1.19 $X2=0
+ $Y2=0
cc_756 N_A_211_363#_c_904_n N_SET_B_c_1275_n 0.026199f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_757 N_A_211_363#_c_904_n N_SET_B_c_1278_n 0.00418383f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_758 N_A_211_363#_c_904_n N_SET_B_c_1280_n 0.00534011f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_759 N_A_211_363#_c_904_n N_A_1003_47#_c_1400_n 0.00500977f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_760 N_A_211_363#_c_904_n N_A_1003_47#_M1013_g 0.00180419f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_761 N_A_211_363#_c_912_n N_A_1003_47#_c_1409_n 0.00253304f $X=4.965 $Y=1.99
+ $X2=0 $Y2=0
cc_762 N_A_211_363#_M1019_g N_A_1003_47#_c_1414_n 0.00912698f $X=5.53 $Y=0.415
+ $X2=0 $Y2=0
cc_763 N_A_211_363#_c_901_n N_A_1003_47#_c_1414_n 0.00594291f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_764 N_A_211_363#_c_906_n N_A_1003_47#_c_1414_n 0.00259674f $X=5.74 $Y=0.85
+ $X2=0 $Y2=0
cc_765 N_A_211_363#_c_908_n N_A_1003_47#_c_1414_n 7.85233e-19 $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_766 N_A_211_363#_c_909_n N_A_1003_47#_c_1414_n 0.0228193f $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_767 N_A_211_363#_c_911_n N_A_1003_47#_c_1406_n 8.38684e-19 $X=4.965 $Y=1.89
+ $X2=0 $Y2=0
cc_768 N_A_211_363#_c_905_n N_A_1003_47#_c_1406_n 3.03433e-19 $X=5.885 $Y=1.19
+ $X2=0 $Y2=0
cc_769 N_A_211_363#_M1019_g N_A_1003_47#_c_1402_n 0.00114556f $X=5.53 $Y=0.415
+ $X2=0 $Y2=0
cc_770 N_A_211_363#_c_896_n N_A_1003_47#_c_1402_n 8.84907e-19 $X=5.555 $Y=1.245
+ $X2=0 $Y2=0
cc_771 N_A_211_363#_c_904_n N_A_1003_47#_c_1402_n 0.0176753f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_772 N_A_211_363#_c_906_n N_A_1003_47#_c_1402_n 0.0140632f $X=5.74 $Y=0.85
+ $X2=0 $Y2=0
cc_773 N_A_211_363#_c_908_n N_A_1003_47#_c_1402_n 7.77832e-19 $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_774 N_A_211_363#_c_909_n N_A_1003_47#_c_1402_n 0.0249836f $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_775 N_A_211_363#_c_904_n N_A_1003_47#_c_1403_n 0.0403444f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_776 N_A_211_363#_c_896_n N_A_1003_47#_c_1404_n 0.00285126f $X=5.555 $Y=1.245
+ $X2=0 $Y2=0
cc_777 N_A_211_363#_c_904_n N_A_1003_47#_c_1404_n 0.0122211f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_778 N_A_211_363#_c_905_n N_A_1003_47#_c_1404_n 0.00672421f $X=5.885 $Y=1.19
+ $X2=0 $Y2=0
cc_779 N_A_211_363#_c_908_n N_A_1003_47#_c_1404_n 5.70846e-19 $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_780 N_A_211_363#_c_909_n N_A_1003_47#_c_1404_n 0.0053097f $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_781 N_A_211_363#_c_904_n N_A_1525_21#_M1021_g 0.00150419f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_782 N_A_211_363#_c_904_n N_A_1525_21#_c_1512_n 0.0123496f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_783 N_A_211_363#_c_915_n N_A_1525_21#_c_1521_n 0.00190553f $X=9.75 $Y=1.99
+ $X2=0 $Y2=0
cc_784 N_A_211_363#_c_900_n N_A_1525_21#_c_1521_n 0.00861532f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_785 N_A_211_363#_c_916_n N_A_1525_21#_c_1521_n 0.0195275f $X=9.755 $Y=1.74
+ $X2=0 $Y2=0
cc_786 N_A_211_363#_c_904_n N_A_1525_21#_c_1521_n 0.014133f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_787 N_A_211_363#_c_907_n N_A_1525_21#_c_1521_n 0.0273727f $X=9.26 $Y=1.19
+ $X2=0 $Y2=0
cc_788 N_A_211_363#_c_904_n N_A_1525_21#_c_1522_n 0.0276968f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_789 N_A_211_363#_c_904_n N_A_1525_21#_c_1523_n 0.00715543f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_790 N_A_211_363#_c_904_n N_A_1525_21#_c_1513_n 0.00696846f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_791 N_A_211_363#_c_916_n N_A_2058_21#_M1014_g 3.61532e-19 $X=9.755 $Y=1.74
+ $X2=0 $Y2=0
cc_792 N_A_211_363#_c_915_n N_A_2058_21#_c_1674_n 0.0246929f $X=9.75 $Y=1.99
+ $X2=0 $Y2=0
cc_793 N_A_211_363#_c_915_n N_A_1864_47#_c_1856_n 0.0139989f $X=9.75 $Y=1.99
+ $X2=0 $Y2=0
cc_794 N_A_211_363#_c_916_n N_A_1864_47#_c_1856_n 0.00816556f $X=9.755 $Y=1.74
+ $X2=0 $Y2=0
cc_795 N_A_211_363#_c_897_n N_A_1864_47#_c_1859_n 0.00643454f $X=9.245 $Y=0.705
+ $X2=0 $Y2=0
cc_796 N_A_211_363#_c_898_n N_A_1864_47#_c_1859_n 0.0044092f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_797 N_A_211_363#_c_899_n N_A_1864_47#_c_1859_n 0.00178491f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_798 N_A_211_363#_c_900_n N_A_1864_47#_c_1859_n 0.00363475f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_799 N_A_211_363#_c_898_n N_A_1864_47#_c_1847_n 0.0112759f $X=9.37 $Y=0.87
+ $X2=0 $Y2=0
cc_800 N_A_211_363#_c_900_n N_A_1864_47#_c_1847_n 0.00871242f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_801 N_A_211_363#_c_915_n N_A_1864_47#_c_1852_n 0.00960954f $X=9.75 $Y=1.99
+ $X2=0 $Y2=0
cc_802 N_A_211_363#_c_916_n N_A_1864_47#_c_1852_n 0.0367913f $X=9.755 $Y=1.74
+ $X2=0 $Y2=0
cc_803 N_A_211_363#_c_900_n N_A_1864_47#_c_1849_n 0.00613391f $X=9.762 $Y=1.305
+ $X2=0 $Y2=0
cc_804 N_A_211_363#_c_916_n N_A_1864_47#_c_1849_n 0.00832639f $X=9.755 $Y=1.74
+ $X2=0 $Y2=0
cc_805 N_A_211_363#_c_910_n N_VPWR_c_2028_n 0.0204951f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_806 N_A_211_363#_c_910_n N_VPWR_c_2029_n 0.0145541f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_807 N_A_211_363#_c_910_n N_VPWR_c_2030_n 0.0356956f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_808 N_A_211_363#_c_912_n N_VPWR_c_2040_n 0.00694062f $X=4.965 $Y=1.99 $X2=0
+ $Y2=0
cc_809 N_A_211_363#_c_915_n N_VPWR_c_2042_n 0.00440543f $X=9.75 $Y=1.99 $X2=0
+ $Y2=0
cc_810 N_A_211_363#_c_912_n N_VPWR_c_2027_n 0.00741367f $X=4.965 $Y=1.99 $X2=0
+ $Y2=0
cc_811 N_A_211_363#_c_915_n N_VPWR_c_2027_n 0.00650106f $X=9.75 $Y=1.99 $X2=0
+ $Y2=0
cc_812 N_A_211_363#_c_910_n N_VPWR_c_2027_n 0.00372404f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_813 N_A_211_363#_c_901_n N_A_483_47#_c_2240_n 0.0187351f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_814 N_A_211_363#_c_901_n N_A_483_47#_c_2241_n 0.00340984f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_815 N_A_211_363#_c_901_n N_A_483_47#_c_2242_n 0.00571441f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_816 N_A_211_363#_c_901_n N_A_483_47#_c_2243_n 0.100923f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_817 N_A_211_363#_c_901_n N_A_483_47#_c_2244_n 0.0279145f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_818 N_A_211_363#_c_901_n N_A_483_47#_c_2245_n 0.00550979f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_819 N_A_211_363#_c_894_n N_A_483_47#_c_2246_n 0.00100977f $X=5.065 $Y=1.32
+ $X2=0 $Y2=0
cc_820 N_A_211_363#_c_901_n N_A_483_47#_c_2246_n 0.0262326f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_821 N_A_211_363#_c_912_n N_A_483_47#_c_2247_n 0.00719081f $X=4.965 $Y=1.99
+ $X2=0 $Y2=0
cc_822 N_A_211_363#_c_894_n N_A_483_47#_c_2247_n 0.00661068f $X=5.065 $Y=1.32
+ $X2=0 $Y2=0
cc_823 N_A_211_363#_c_901_n N_A_483_47#_c_2247_n 0.0142672f $X=5.595 $Y=0.85
+ $X2=0 $Y2=0
cc_824 N_A_211_363#_c_909_n N_A_483_47#_c_2247_n 0.00193662f $X=5.64 $Y=0.93
+ $X2=0 $Y2=0
cc_825 N_A_211_363#_c_910_n N_VGND_c_2427_n 0.00888183f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_826 N_A_211_363#_c_901_n N_VGND_c_2428_n 0.0050337f $X=5.595 $Y=0.85 $X2=0
+ $Y2=0
cc_827 N_A_211_363#_c_910_n N_VGND_c_2428_n 0.0177642f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_828 N_A_211_363#_c_901_n N_VGND_c_2429_n 0.00134454f $X=5.595 $Y=0.85 $X2=0
+ $Y2=0
cc_829 N_A_211_363#_M1019_g N_VGND_c_2434_n 0.00359964f $X=5.53 $Y=0.415 $X2=0
+ $Y2=0
cc_830 N_A_211_363#_c_897_n N_VGND_c_2436_n 0.00435972f $X=9.245 $Y=0.705 $X2=0
+ $Y2=0
cc_831 N_A_211_363#_c_898_n N_VGND_c_2436_n 0.00363141f $X=9.37 $Y=0.87 $X2=0
+ $Y2=0
cc_832 N_A_211_363#_c_899_n N_VGND_c_2436_n 4.01089e-19 $X=9.37 $Y=0.87 $X2=0
+ $Y2=0
cc_833 N_A_211_363#_M1001_d N_VGND_c_2444_n 0.00285751f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_834 N_A_211_363#_M1019_g N_VGND_c_2444_n 0.00584425f $X=5.53 $Y=0.415 $X2=0
+ $Y2=0
cc_835 N_A_211_363#_c_897_n N_VGND_c_2444_n 0.00634051f $X=9.245 $Y=0.705 $X2=0
+ $Y2=0
cc_836 N_A_211_363#_c_898_n N_VGND_c_2444_n 0.00282859f $X=9.37 $Y=0.87 $X2=0
+ $Y2=0
cc_837 N_A_211_363#_c_901_n N_VGND_c_2444_n 0.199819f $X=5.595 $Y=0.85 $X2=0
+ $Y2=0
cc_838 N_A_211_363#_c_902_n N_VGND_c_2444_n 0.0152682f $X=1.38 $Y=0.85 $X2=0
+ $Y2=0
cc_839 N_A_211_363#_c_906_n N_VGND_c_2444_n 0.0154004f $X=5.74 $Y=0.85 $X2=0
+ $Y2=0
cc_840 N_A_211_363#_c_910_n N_VGND_c_2444_n 0.00339196f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_841 N_A_211_363#_c_909_n A_1121_47# 0.00109936f $X=5.64 $Y=0.93 $X2=-0.19
+ $Y2=-0.24
cc_842 N_A_1197_21#_M1025_g N_SET_B_c_1270_n 0.0119034f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_843 N_A_1197_21#_c_1131_n N_SET_B_c_1270_n 0.0204283f $X=6.085 $Y=1.99 $X2=0
+ $Y2=0
cc_844 N_A_1197_21#_c_1134_n N_SET_B_c_1270_n 0.00844926f $X=6.935 $Y=1.91 $X2=0
+ $Y2=0
cc_845 N_A_1197_21#_c_1136_n N_SET_B_c_1270_n 0.00488436f $X=6.17 $Y=1.74 $X2=0
+ $Y2=0
cc_846 N_A_1197_21#_c_1131_n N_SET_B_c_1282_n 0.0152518f $X=6.085 $Y=1.99 $X2=0
+ $Y2=0
cc_847 N_A_1197_21#_c_1134_n N_SET_B_c_1282_n 0.0108028f $X=6.935 $Y=1.91 $X2=0
+ $Y2=0
cc_848 N_A_1197_21#_c_1181_p N_SET_B_c_1282_n 0.00521779f $X=7.02 $Y=2.21 $X2=0
+ $Y2=0
cc_849 N_A_1197_21#_M1025_g N_SET_B_M1009_g 0.0119041f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_850 N_A_1197_21#_c_1125_n N_SET_B_M1009_g 7.24899e-19 $X=7.5 $Y=1.065 $X2=0
+ $Y2=0
cc_851 N_A_1197_21#_M1013_d N_SET_B_c_1274_n 3.84553e-19 $X=7.355 $Y=0.235 $X2=0
+ $Y2=0
cc_852 N_A_1197_21#_c_1124_n N_SET_B_c_1274_n 0.00525024f $X=8.77 $Y=0.985 $X2=0
+ $Y2=0
cc_853 N_A_1197_21#_c_1125_n N_SET_B_c_1274_n 0.0228791f $X=7.5 $Y=1.065 $X2=0
+ $Y2=0
cc_854 N_A_1197_21#_c_1127_n N_SET_B_c_1274_n 0.0217267f $X=8.445 $Y=0.98 $X2=0
+ $Y2=0
cc_855 N_A_1197_21#_c_1128_n N_SET_B_c_1274_n 0.0142323f $X=8.66 $Y=0.98 $X2=0
+ $Y2=0
cc_856 N_A_1197_21#_c_1125_n N_SET_B_c_1275_n 0.00207888f $X=7.5 $Y=1.065 $X2=0
+ $Y2=0
cc_857 N_A_1197_21#_M1025_g N_SET_B_c_1278_n 0.0148943f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_858 N_A_1197_21#_M1025_g N_SET_B_c_1280_n 0.0010314f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_859 N_A_1197_21#_c_1125_n N_SET_B_c_1280_n 0.00756919f $X=7.5 $Y=1.065 $X2=0
+ $Y2=0
cc_860 N_A_1197_21#_c_1146_n N_A_1003_47#_c_1400_n 0.0149923f $X=7.415 $Y=1.91
+ $X2=0 $Y2=0
cc_861 N_A_1197_21#_c_1126_n N_A_1003_47#_c_1400_n 0.00507662f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_862 N_A_1197_21#_c_1148_n N_A_1003_47#_c_1400_n 9.36723e-19 $X=7.02 $Y=1.87
+ $X2=0 $Y2=0
cc_863 N_A_1197_21#_c_1125_n N_A_1003_47#_M1013_g 0.00991255f $X=7.5 $Y=1.065
+ $X2=0 $Y2=0
cc_864 N_A_1197_21#_c_1126_n N_A_1003_47#_M1013_g 0.00661765f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_865 N_A_1197_21#_c_1131_n N_A_1003_47#_c_1409_n 0.00211032f $X=6.085 $Y=1.99
+ $X2=0 $Y2=0
cc_866 N_A_1197_21#_M1025_g N_A_1003_47#_c_1414_n 0.009343f $X=6.06 $Y=0.445
+ $X2=0 $Y2=0
cc_867 N_A_1197_21#_M1025_g N_A_1003_47#_c_1406_n 0.0103777f $X=6.06 $Y=0.445
+ $X2=0 $Y2=0
cc_868 N_A_1197_21#_c_1131_n N_A_1003_47#_c_1406_n 0.00523372f $X=6.085 $Y=1.99
+ $X2=0 $Y2=0
cc_869 N_A_1197_21#_c_1136_n N_A_1003_47#_c_1406_n 0.0333383f $X=6.17 $Y=1.74
+ $X2=0 $Y2=0
cc_870 N_A_1197_21#_M1025_g N_A_1003_47#_c_1402_n 0.0210093f $X=6.06 $Y=0.445
+ $X2=0 $Y2=0
cc_871 N_A_1197_21#_c_1134_n N_A_1003_47#_c_1403_n 0.0153662f $X=6.935 $Y=1.91
+ $X2=0 $Y2=0
cc_872 N_A_1197_21#_c_1146_n N_A_1003_47#_c_1403_n 0.00200144f $X=7.415 $Y=1.91
+ $X2=0 $Y2=0
cc_873 N_A_1197_21#_c_1126_n N_A_1003_47#_c_1403_n 0.0198741f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_874 N_A_1197_21#_c_1148_n N_A_1003_47#_c_1403_n 0.00666603f $X=7.02 $Y=1.87
+ $X2=0 $Y2=0
cc_875 N_A_1197_21#_M1025_g N_A_1003_47#_c_1404_n 0.0112214f $X=6.06 $Y=0.445
+ $X2=0 $Y2=0
cc_876 N_A_1197_21#_c_1131_n N_A_1003_47#_c_1404_n 0.00155337f $X=6.085 $Y=1.99
+ $X2=0 $Y2=0
cc_877 N_A_1197_21#_c_1136_n N_A_1003_47#_c_1404_n 0.0204654f $X=6.17 $Y=1.74
+ $X2=0 $Y2=0
cc_878 N_A_1197_21#_c_1125_n N_A_1525_21#_M1021_g 0.00976299f $X=7.5 $Y=1.065
+ $X2=0 $Y2=0
cc_879 N_A_1197_21#_c_1126_n N_A_1525_21#_M1021_g 0.00666631f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_880 N_A_1197_21#_c_1127_n N_A_1525_21#_M1021_g 0.00924448f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_881 N_A_1197_21#_c_1128_n N_A_1525_21#_M1021_g 6.32302e-19 $X=8.66 $Y=0.98
+ $X2=0 $Y2=0
cc_882 N_A_1197_21#_c_1129_n N_A_1525_21#_M1021_g 0.00316536f $X=8.77 $Y=1.15
+ $X2=0 $Y2=0
cc_883 N_A_1197_21#_c_1133_n N_A_1525_21#_c_1516_n 0.0134641f $X=8.46 $Y=1.57
+ $X2=0 $Y2=0
cc_884 N_A_1197_21#_c_1146_n N_A_1525_21#_c_1516_n 0.00225739f $X=7.415 $Y=1.91
+ $X2=0 $Y2=0
cc_885 N_A_1197_21#_c_1126_n N_A_1525_21#_c_1516_n 0.00124086f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_886 N_A_1197_21#_c_1126_n N_A_1525_21#_c_1512_n 0.0253829f $X=7.5 $Y=1.785
+ $X2=0 $Y2=0
cc_887 N_A_1197_21#_c_1127_n N_A_1525_21#_c_1512_n 0.0205705f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_888 N_A_1197_21#_c_1129_n N_A_1525_21#_c_1512_n 0.00386043f $X=8.77 $Y=1.15
+ $X2=0 $Y2=0
cc_889 N_A_1197_21#_c_1128_n N_A_1525_21#_c_1522_n 9.59092e-19 $X=8.66 $Y=0.98
+ $X2=0 $Y2=0
cc_890 N_A_1197_21#_c_1129_n N_A_1525_21#_c_1522_n 0.00358318f $X=8.77 $Y=1.15
+ $X2=0 $Y2=0
cc_891 N_A_1197_21#_c_1132_n N_A_1525_21#_c_1523_n 0.00552706f $X=8.46 $Y=1.47
+ $X2=0 $Y2=0
cc_892 N_A_1197_21#_c_1133_n N_A_1525_21#_c_1523_n 0.0118271f $X=8.46 $Y=1.57
+ $X2=0 $Y2=0
cc_893 N_A_1197_21#_c_1127_n N_A_1525_21#_c_1523_n 0.00743994f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_894 N_A_1197_21#_c_1128_n N_A_1525_21#_c_1523_n 0.0266532f $X=8.66 $Y=0.98
+ $X2=0 $Y2=0
cc_895 N_A_1197_21#_c_1129_n N_A_1525_21#_c_1523_n 0.00756441f $X=8.77 $Y=1.15
+ $X2=0 $Y2=0
cc_896 N_A_1197_21#_c_1133_n N_A_1525_21#_c_1513_n 0.00144809f $X=8.46 $Y=1.57
+ $X2=0 $Y2=0
cc_897 N_A_1197_21#_c_1127_n N_A_1525_21#_c_1513_n 0.00706066f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_898 N_A_1197_21#_c_1128_n N_A_1525_21#_c_1513_n 7.22512e-19 $X=8.66 $Y=0.98
+ $X2=0 $Y2=0
cc_899 N_A_1197_21#_c_1129_n N_A_1525_21#_c_1513_n 0.017057f $X=8.77 $Y=1.15
+ $X2=0 $Y2=0
cc_900 N_A_1197_21#_c_1131_n N_VPWR_c_2032_n 0.00403064f $X=6.085 $Y=1.99 $X2=0
+ $Y2=0
cc_901 N_A_1197_21#_c_1134_n N_VPWR_c_2032_n 0.0125643f $X=6.935 $Y=1.91 $X2=0
+ $Y2=0
cc_902 N_A_1197_21#_c_1181_p N_VPWR_c_2032_n 0.00728058f $X=7.02 $Y=2.21 $X2=0
+ $Y2=0
cc_903 N_A_1197_21#_c_1136_n N_VPWR_c_2032_n 0.0129312f $X=6.17 $Y=1.74 $X2=0
+ $Y2=0
cc_904 N_A_1197_21#_c_1133_n N_VPWR_c_2033_n 0.0163727f $X=8.46 $Y=1.57 $X2=0
+ $Y2=0
cc_905 N_A_1197_21#_c_1146_n N_VPWR_c_2033_n 6.52334e-19 $X=7.415 $Y=1.91 $X2=0
+ $Y2=0
cc_906 N_A_1197_21#_c_1131_n N_VPWR_c_2040_n 0.00635673f $X=6.085 $Y=1.99 $X2=0
+ $Y2=0
cc_907 N_A_1197_21#_c_1136_n N_VPWR_c_2040_n 0.0019176f $X=6.17 $Y=1.74 $X2=0
+ $Y2=0
cc_908 N_A_1197_21#_c_1134_n N_VPWR_c_2041_n 0.00550916f $X=6.935 $Y=1.91 $X2=0
+ $Y2=0
cc_909 N_A_1197_21#_c_1181_p N_VPWR_c_2041_n 0.00738128f $X=7.02 $Y=2.21 $X2=0
+ $Y2=0
cc_910 N_A_1197_21#_c_1146_n N_VPWR_c_2041_n 0.00678412f $X=7.415 $Y=1.91 $X2=0
+ $Y2=0
cc_911 N_A_1197_21#_c_1133_n N_VPWR_c_2042_n 0.00702461f $X=8.46 $Y=1.57 $X2=0
+ $Y2=0
cc_912 N_A_1197_21#_M1012_d N_VPWR_c_2027_n 0.00335282f $X=6.755 $Y=2.065 $X2=0
+ $Y2=0
cc_913 N_A_1197_21#_c_1131_n N_VPWR_c_2027_n 0.00769239f $X=6.085 $Y=1.99 $X2=0
+ $Y2=0
cc_914 N_A_1197_21#_c_1133_n N_VPWR_c_2027_n 0.00873182f $X=8.46 $Y=1.57 $X2=0
+ $Y2=0
cc_915 N_A_1197_21#_c_1134_n N_VPWR_c_2027_n 0.00438899f $X=6.935 $Y=1.91 $X2=0
+ $Y2=0
cc_916 N_A_1197_21#_c_1181_p N_VPWR_c_2027_n 0.0029026f $X=7.02 $Y=2.21 $X2=0
+ $Y2=0
cc_917 N_A_1197_21#_c_1146_n N_VPWR_c_2027_n 0.0055933f $X=7.415 $Y=1.91 $X2=0
+ $Y2=0
cc_918 N_A_1197_21#_c_1136_n N_VPWR_c_2027_n 0.00183442f $X=6.17 $Y=1.74 $X2=0
+ $Y2=0
cc_919 N_A_1197_21#_c_1146_n A_1469_329# 0.00432757f $X=7.415 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_920 N_A_1197_21#_c_1126_n A_1469_329# 0.00194122f $X=7.5 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_921 N_A_1197_21#_M1025_g N_VGND_c_2430_n 0.00336814f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_922 N_A_1197_21#_M1025_g N_VGND_c_2434_n 0.0035977f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_923 N_A_1197_21#_c_1124_n N_VGND_c_2436_n 0.00585385f $X=8.77 $Y=0.985 $X2=0
+ $Y2=0
cc_924 N_A_1197_21#_c_1124_n N_VGND_c_2440_n 0.00944167f $X=8.77 $Y=0.985 $X2=0
+ $Y2=0
cc_925 N_A_1197_21#_c_1127_n N_VGND_c_2440_n 0.00400251f $X=8.445 $Y=0.98 $X2=0
+ $Y2=0
cc_926 N_A_1197_21#_c_1128_n N_VGND_c_2440_n 0.00551479f $X=8.66 $Y=0.98 $X2=0
+ $Y2=0
cc_927 N_A_1197_21#_c_1129_n N_VGND_c_2440_n 0.00165636f $X=8.77 $Y=1.15 $X2=0
+ $Y2=0
cc_928 N_A_1197_21#_M1013_d N_VGND_c_2444_n 0.00178362f $X=7.355 $Y=0.235 $X2=0
+ $Y2=0
cc_929 N_A_1197_21#_M1025_g N_VGND_c_2444_n 0.00602697f $X=6.06 $Y=0.445 $X2=0
+ $Y2=0
cc_930 N_A_1197_21#_c_1124_n N_VGND_c_2444_n 0.00777927f $X=8.77 $Y=0.985 $X2=0
+ $Y2=0
cc_931 N_A_1197_21#_M1013_d N_A_1353_47#_c_2647_n 0.00301726f $X=7.355 $Y=0.235
+ $X2=0 $Y2=0
cc_932 N_A_1197_21#_c_1125_n N_A_1353_47#_c_2647_n 0.0179348f $X=7.5 $Y=1.065
+ $X2=0 $Y2=0
cc_933 N_A_1197_21#_c_1127_n N_A_1353_47#_c_2647_n 0.00305646f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_934 N_A_1197_21#_c_1124_n N_A_1353_47#_c_2650_n 0.00535152f $X=8.77 $Y=0.985
+ $X2=0 $Y2=0
cc_935 N_A_1197_21#_c_1125_n N_A_1353_47#_c_2650_n 0.00817558f $X=7.5 $Y=1.065
+ $X2=0 $Y2=0
cc_936 N_A_1197_21#_c_1127_n N_A_1353_47#_c_2650_n 0.01244f $X=8.445 $Y=0.98
+ $X2=0 $Y2=0
cc_937 N_SET_B_c_1270_n N_A_1003_47#_c_1400_n 0.0321902f $X=6.665 $Y=1.89 $X2=0
+ $Y2=0
cc_938 N_SET_B_c_1282_n N_A_1003_47#_c_1400_n 0.0115765f $X=6.665 $Y=1.99 $X2=0
+ $Y2=0
cc_939 N_SET_B_M1009_g N_A_1003_47#_M1013_g 0.0235453f $X=6.69 $Y=0.445 $X2=0
+ $Y2=0
cc_940 N_SET_B_c_1274_n N_A_1003_47#_M1013_g 0.00514187f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_941 N_SET_B_c_1275_n N_A_1003_47#_M1013_g 0.00124772f $X=6.815 $Y=0.85 $X2=0
+ $Y2=0
cc_942 N_SET_B_c_1280_n N_A_1003_47#_M1013_g 0.00217911f $X=6.67 $Y=0.85 $X2=0
+ $Y2=0
cc_943 N_SET_B_c_1270_n N_A_1003_47#_c_1402_n 6.37306e-19 $X=6.665 $Y=1.89 $X2=0
+ $Y2=0
cc_944 N_SET_B_M1009_g N_A_1003_47#_c_1402_n 0.00392982f $X=6.69 $Y=0.445 $X2=0
+ $Y2=0
cc_945 N_SET_B_c_1275_n N_A_1003_47#_c_1402_n 0.0012341f $X=6.815 $Y=0.85 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1278_n N_A_1003_47#_c_1402_n 0.00235335f $X=6.55 $Y=0.98 $X2=0
+ $Y2=0
cc_947 N_SET_B_c_1280_n N_A_1003_47#_c_1402_n 0.0249073f $X=6.67 $Y=0.85 $X2=0
+ $Y2=0
cc_948 N_SET_B_c_1270_n N_A_1003_47#_c_1403_n 0.0155987f $X=6.665 $Y=1.89 $X2=0
+ $Y2=0
cc_949 N_SET_B_c_1274_n N_A_1003_47#_c_1403_n 0.00423591f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_950 N_SET_B_c_1275_n N_A_1003_47#_c_1403_n 4.90254e-19 $X=6.815 $Y=0.85 $X2=0
+ $Y2=0
cc_951 N_SET_B_c_1278_n N_A_1003_47#_c_1403_n 0.0028803f $X=6.55 $Y=0.98 $X2=0
+ $Y2=0
cc_952 N_SET_B_c_1280_n N_A_1003_47#_c_1403_n 0.026111f $X=6.67 $Y=0.85 $X2=0
+ $Y2=0
cc_953 N_SET_B_c_1270_n N_A_1003_47#_c_1404_n 5.39722e-19 $X=6.665 $Y=1.89 $X2=0
+ $Y2=0
cc_954 N_SET_B_c_1274_n N_A_1525_21#_M1021_g 0.00317213f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_955 N_SET_B_c_1274_n N_A_1525_21#_c_1512_n 5.29205e-19 $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_956 N_SET_B_c_1272_n N_A_1525_21#_c_1521_n 0.00716241f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_957 N_SET_B_c_1274_n N_A_1525_21#_c_1521_n 0.0557598f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_958 N_SET_B_c_1276_n N_A_1525_21#_c_1521_n 0.0134169f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1272_n N_A_2058_21#_M1014_g 0.0118142f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_960 N_SET_B_M1000_g N_A_2058_21#_M1014_g 0.0128509f $X=11.005 $Y=0.445 $X2=0
+ $Y2=0
cc_961 N_SET_B_c_1274_n N_A_2058_21#_M1014_g 0.00649356f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_962 N_SET_B_c_1276_n N_A_2058_21#_M1014_g 0.00137705f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1277_n N_A_2058_21#_M1014_g 0.00244823f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_964 N_SET_B_c_1279_n N_A_2058_21#_M1014_g 0.0167241f $X=11.005 $Y=0.98 $X2=0
+ $Y2=0
cc_965 N_SET_B_c_1272_n N_A_2058_21#_c_1674_n 0.0200963f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_966 N_SET_B_c_1284_n N_A_2058_21#_c_1674_n 0.0197678f $X=10.98 $Y=1.99 $X2=0
+ $Y2=0
cc_967 N_SET_B_c_1272_n N_A_2058_21#_c_1679_n 0.00741526f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1284_n N_A_2058_21#_c_1680_n 0.0169103f $X=10.98 $Y=1.99 $X2=0
+ $Y2=0
cc_969 N_SET_B_c_1284_n N_A_2058_21#_c_1698_n 0.00492021f $X=10.98 $Y=1.99 $X2=0
+ $Y2=0
cc_970 N_SET_B_c_1277_n N_A_2058_21#_c_1671_n 0.00677427f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_971 N_SET_B_M1000_g N_A_2058_21#_c_1700_n 7.06195e-19 $X=11.005 $Y=0.445
+ $X2=0 $Y2=0
cc_972 N_SET_B_c_1276_n N_A_2058_21#_c_1700_n 4.03497e-19 $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_973 N_SET_B_c_1277_n N_A_2058_21#_c_1700_n 0.00231197f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_974 N_SET_B_c_1272_n N_A_1864_47#_c_1845_n 0.0234391f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_975 N_SET_B_c_1284_n N_A_1864_47#_c_1845_n 0.0146106f $X=10.98 $Y=1.99 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1279_n N_A_1864_47#_c_1845_n 0.0216199f $X=11.005 $Y=0.98 $X2=0
+ $Y2=0
cc_977 N_SET_B_M1000_g N_A_1864_47#_M1040_g 0.0259143f $X=11.005 $Y=0.445 $X2=0
+ $Y2=0
cc_978 N_SET_B_c_1277_n N_A_1864_47#_M1040_g 0.00128343f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1274_n N_A_1864_47#_c_1859_n 0.00949836f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_980 N_SET_B_c_1274_n N_A_1864_47#_c_1847_n 0.0181691f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_981 N_SET_B_c_1276_n N_A_1864_47#_c_1847_n 0.00218964f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_982 N_SET_B_c_1277_n N_A_1864_47#_c_1847_n 0.010555f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1272_n N_A_1864_47#_c_1848_n 0.0145354f $X=10.98 $Y=1.89 $X2=0
+ $Y2=0
cc_984 N_SET_B_c_1274_n N_A_1864_47#_c_1848_n 0.0103288f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_985 N_SET_B_c_1276_n N_A_1864_47#_c_1848_n 9.69765e-19 $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_986 N_SET_B_c_1277_n N_A_1864_47#_c_1848_n 0.0281583f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_987 N_SET_B_c_1279_n N_A_1864_47#_c_1848_n 0.00455716f $X=11.005 $Y=0.98
+ $X2=0 $Y2=0
cc_988 N_SET_B_c_1279_n N_A_1864_47#_c_1850_n 0.00113254f $X=11.005 $Y=0.98
+ $X2=0 $Y2=0
cc_989 N_SET_B_c_1282_n N_VPWR_c_2032_n 0.0133526f $X=6.665 $Y=1.99 $X2=0 $Y2=0
cc_990 N_SET_B_c_1282_n N_VPWR_c_2041_n 0.00492591f $X=6.665 $Y=1.99 $X2=0 $Y2=0
cc_991 N_SET_B_c_1282_n N_VPWR_c_2027_n 0.0055272f $X=6.665 $Y=1.99 $X2=0 $Y2=0
cc_992 N_SET_B_c_1284_n N_VPWR_c_2027_n 0.00563515f $X=10.98 $Y=1.99 $X2=0 $Y2=0
cc_993 N_SET_B_c_1284_n N_VPWR_c_2051_n 0.0117343f $X=10.98 $Y=1.99 $X2=0 $Y2=0
cc_994 N_SET_B_c_1284_n N_VPWR_c_2052_n 0.0048505f $X=10.98 $Y=1.99 $X2=0 $Y2=0
cc_995 N_SET_B_c_1274_n N_VGND_M1037_s 0.00316071f $X=10.655 $Y=0.85 $X2=0 $Y2=0
cc_996 N_SET_B_M1009_g N_VGND_c_2430_n 0.00519315f $X=6.69 $Y=0.445 $X2=0 $Y2=0
cc_997 N_SET_B_c_1278_n N_VGND_c_2430_n 8.75675e-19 $X=6.55 $Y=0.98 $X2=0 $Y2=0
cc_998 N_SET_B_c_1280_n N_VGND_c_2430_n 0.0109479f $X=6.67 $Y=0.85 $X2=0 $Y2=0
cc_999 N_SET_B_M1000_g N_VGND_c_2431_n 0.00598296f $X=11.005 $Y=0.445 $X2=0
+ $Y2=0
cc_1000 N_SET_B_c_1274_n N_VGND_c_2431_n 0.00808121f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_1001 N_SET_B_c_1276_n N_VGND_c_2431_n 3.46255e-19 $X=10.8 $Y=0.85 $X2=0 $Y2=0
cc_1002 N_SET_B_c_1277_n N_VGND_c_2431_n 0.00367619f $X=10.8 $Y=0.85 $X2=0 $Y2=0
cc_1003 N_SET_B_M1009_g N_VGND_c_2440_n 0.00439071f $X=6.69 $Y=0.445 $X2=0 $Y2=0
cc_1004 N_SET_B_c_1274_n N_VGND_c_2440_n 0.00480627f $X=10.655 $Y=0.85 $X2=0
+ $Y2=0
cc_1005 N_SET_B_c_1280_n N_VGND_c_2440_n 0.00287774f $X=6.67 $Y=0.85 $X2=0 $Y2=0
cc_1006 N_SET_B_M1000_g N_VGND_c_2441_n 0.00384942f $X=11.005 $Y=0.445 $X2=0
+ $Y2=0
cc_1007 N_SET_B_c_1277_n N_VGND_c_2441_n 0.00387176f $X=10.8 $Y=0.85 $X2=0 $Y2=0
cc_1008 N_SET_B_M1009_g N_VGND_c_2444_n 0.00632764f $X=6.69 $Y=0.445 $X2=0 $Y2=0
cc_1009 N_SET_B_M1000_g N_VGND_c_2444_n 0.00623252f $X=11.005 $Y=0.445 $X2=0
+ $Y2=0
cc_1010 N_SET_B_c_1274_n N_VGND_c_2444_n 0.187375f $X=10.655 $Y=0.85 $X2=0 $Y2=0
cc_1011 N_SET_B_c_1275_n N_VGND_c_2444_n 0.0144468f $X=6.815 $Y=0.85 $X2=0 $Y2=0
cc_1012 N_SET_B_c_1276_n N_VGND_c_2444_n 0.0144219f $X=10.8 $Y=0.85 $X2=0 $Y2=0
cc_1013 N_SET_B_c_1277_n N_VGND_c_2444_n 0.00242766f $X=10.8 $Y=0.85 $X2=0 $Y2=0
cc_1014 N_SET_B_c_1280_n N_VGND_c_2444_n 0.00212631f $X=6.67 $Y=0.85 $X2=0 $Y2=0
cc_1015 N_SET_B_c_1274_n N_A_1353_47#_M1009_d 0.0030671f $X=10.655 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_1016 N_SET_B_c_1274_n N_A_1353_47#_M1021_d 0.00218405f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_1017 N_SET_B_c_1274_n N_A_1353_47#_c_2647_n 0.00669858f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_1018 N_SET_B_c_1274_n N_A_1353_47#_c_2650_n 0.00269828f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_1019 N_SET_B_c_1274_n N_A_1353_47#_c_2657_n 0.00779132f $X=10.655 $Y=0.85
+ $X2=0 $Y2=0
cc_1020 N_SET_B_c_1275_n N_A_1353_47#_c_2657_n 6.90415e-19 $X=6.815 $Y=0.85
+ $X2=0 $Y2=0
cc_1021 N_SET_B_c_1274_n A_1769_47# 0.00369541f $X=10.655 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_1022 N_SET_B_M1000_g N_A_2216_47#_c_2675_n 0.00625795f $X=11.005 $Y=0.445
+ $X2=0 $Y2=0
cc_1023 N_SET_B_c_1277_n N_A_2216_47#_c_2675_n 0.00449237f $X=10.8 $Y=0.85 $X2=0
+ $Y2=0
cc_1024 N_A_1003_47#_M1013_g N_A_1525_21#_M1021_g 0.0246977f $X=7.28 $Y=0.555
+ $X2=0 $Y2=0
cc_1025 N_A_1003_47#_c_1400_n N_A_1525_21#_c_1516_n 0.0435094f $X=7.255 $Y=1.57
+ $X2=0 $Y2=0
cc_1026 N_A_1003_47#_c_1400_n N_A_1525_21#_c_1513_n 0.0246977f $X=7.255 $Y=1.57
+ $X2=0 $Y2=0
cc_1027 N_A_1003_47#_c_1400_n N_VPWR_c_2032_n 0.00125978f $X=7.255 $Y=1.57 $X2=0
+ $Y2=0
cc_1028 N_A_1003_47#_c_1409_n N_VPWR_c_2040_n 0.0401746f $X=5.745 $Y=2.335 $X2=0
+ $Y2=0
cc_1029 N_A_1003_47#_c_1400_n N_VPWR_c_2041_n 0.00518775f $X=7.255 $Y=1.57 $X2=0
+ $Y2=0
cc_1030 N_A_1003_47#_M1020_d N_VPWR_c_2027_n 0.00186203f $X=5.055 $Y=2.065 $X2=0
+ $Y2=0
cc_1031 N_A_1003_47#_c_1400_n N_VPWR_c_2027_n 0.00691464f $X=7.255 $Y=1.57 $X2=0
+ $Y2=0
cc_1032 N_A_1003_47#_c_1409_n N_VPWR_c_2027_n 0.0140322f $X=5.745 $Y=2.335 $X2=0
+ $Y2=0
cc_1033 N_A_1003_47#_c_1409_n N_A_483_47#_c_2247_n 0.0108107f $X=5.745 $Y=2.335
+ $X2=0 $Y2=0
cc_1034 N_A_1003_47#_c_1409_n A_1105_413# 0.00898117f $X=5.745 $Y=2.335
+ $X2=-0.19 $Y2=-0.24
cc_1035 N_A_1003_47#_c_1406_n A_1105_413# 0.00585254f $X=5.83 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_1036 N_A_1003_47#_c_1414_n N_VGND_M1025_d 0.00212485f $X=5.995 $Y=0.365 $X2=0
+ $Y2=0
cc_1037 N_A_1003_47#_c_1402_n N_VGND_M1025_d 0.0024324f $X=6.105 $Y=1.195 $X2=0
+ $Y2=0
cc_1038 N_A_1003_47#_c_1414_n N_VGND_c_2430_n 0.0162715f $X=5.995 $Y=0.365 $X2=0
+ $Y2=0
cc_1039 N_A_1003_47#_c_1402_n N_VGND_c_2430_n 0.00440605f $X=6.105 $Y=1.195
+ $X2=0 $Y2=0
cc_1040 N_A_1003_47#_c_1414_n N_VGND_c_2434_n 0.0613692f $X=5.995 $Y=0.365 $X2=0
+ $Y2=0
cc_1041 N_A_1003_47#_M1013_g N_VGND_c_2440_n 0.00357877f $X=7.28 $Y=0.555 $X2=0
+ $Y2=0
cc_1042 N_A_1003_47#_M1027_d N_VGND_c_2444_n 0.00313914f $X=5.015 $Y=0.235 $X2=0
+ $Y2=0
cc_1043 N_A_1003_47#_M1013_g N_VGND_c_2444_n 0.00564328f $X=7.28 $Y=0.555 $X2=0
+ $Y2=0
cc_1044 N_A_1003_47#_c_1414_n N_VGND_c_2444_n 0.0246489f $X=5.995 $Y=0.365 $X2=0
+ $Y2=0
cc_1045 N_A_1003_47#_c_1414_n A_1121_47# 0.00680543f $X=5.995 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1046 N_A_1003_47#_M1013_g N_A_1353_47#_c_2647_n 0.0105513f $X=7.28 $Y=0.555
+ $X2=0 $Y2=0
cc_1047 N_A_1003_47#_c_1400_n N_A_1353_47#_c_2657_n 0.00160442f $X=7.255 $Y=1.57
+ $X2=0 $Y2=0
cc_1048 N_A_1003_47#_M1013_g N_A_1353_47#_c_2657_n 0.00107318f $X=7.28 $Y=0.555
+ $X2=0 $Y2=0
cc_1049 N_A_1525_21#_c_1521_n N_A_2058_21#_M1014_g 0.0042168f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1050 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1674_n 0.0072227f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1051 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1679_n 0.0181818f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1052 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1680_n 0.0114488f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1053 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1707_n 0.0113591f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1054 N_A_1525_21#_c_1517_n N_A_2058_21#_c_1671_n 0.0121855f $X=11.92 $Y=1.57
+ $X2=0 $Y2=0
cc_1055 N_A_1525_21#_M1007_g N_A_2058_21#_c_1671_n 0.00436862f $X=12 $Y=0.555
+ $X2=0 $Y2=0
cc_1056 N_A_1525_21#_c_1510_n N_A_2058_21#_c_1671_n 0.003526f $X=12.345 $Y=0.84
+ $X2=0 $Y2=0
cc_1057 N_A_1525_21#_c_1518_n N_A_2058_21#_c_1671_n 0.0102646f $X=12.345 $Y=1.66
+ $X2=0 $Y2=0
cc_1058 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1671_n 0.0279253f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1059 N_A_1525_21#_c_1524_n N_A_2058_21#_c_1671_n 0.0023592f $X=12.25 $Y=1.53
+ $X2=0 $Y2=0
cc_1060 N_A_1525_21#_c_1514_n N_A_2058_21#_c_1671_n 0.00794288f $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1061 N_A_1525_21#_c_1515_n N_A_2058_21#_c_1671_n 0.0387608f $X=12.215 $Y=1.32
+ $X2=0 $Y2=0
cc_1062 N_A_1525_21#_M1017_s N_A_2058_21#_c_1682_n 0.00508931f $X=12.605
+ $Y=1.505 $X2=0 $Y2=0
cc_1063 N_A_1525_21#_c_1517_n N_A_2058_21#_c_1682_n 0.00875687f $X=11.92 $Y=1.57
+ $X2=0 $Y2=0
cc_1064 N_A_1525_21#_c_1518_n N_A_2058_21#_c_1682_n 0.0165227f $X=12.345 $Y=1.66
+ $X2=0 $Y2=0
cc_1065 N_A_1525_21#_c_1519_n N_A_2058_21#_c_1682_n 0.0367299f $X=12.73 $Y=1.66
+ $X2=0 $Y2=0
cc_1066 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1682_n 0.00675942f $X=12.105
+ $Y=1.53 $X2=0 $Y2=0
cc_1067 N_A_1525_21#_c_1524_n N_A_2058_21#_c_1682_n 0.00263694f $X=12.25 $Y=1.53
+ $X2=0 $Y2=0
cc_1068 N_A_1525_21#_c_1514_n N_A_2058_21#_c_1682_n 0.00278434f $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1069 N_A_1525_21#_c_1519_n N_A_2058_21#_c_1683_n 0.0074661f $X=12.73 $Y=1.66
+ $X2=0 $Y2=0
cc_1070 N_A_1525_21#_c_1521_n N_A_2058_21#_c_1724_n 0.00453864f $X=12.105
+ $Y=1.53 $X2=0 $Y2=0
cc_1071 N_A_1525_21#_c_1514_n N_A_2058_21#_c_1700_n 2.03871e-19 $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1072 N_A_1525_21#_c_1517_n N_A_2058_21#_c_1726_n 0.00494816f $X=11.92 $Y=1.57
+ $X2=0 $Y2=0
cc_1073 N_A_1525_21#_c_1517_n N_A_1864_47#_c_1845_n 0.0590405f $X=11.92 $Y=1.57
+ $X2=0 $Y2=0
cc_1074 N_A_1525_21#_c_1521_n N_A_1864_47#_c_1845_n 0.00993001f $X=12.105
+ $Y=1.53 $X2=0 $Y2=0
cc_1075 N_A_1525_21#_c_1514_n N_A_1864_47#_c_1845_n 0.0311052f $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1076 N_A_1525_21#_M1007_g N_A_1864_47#_M1040_g 0.0160528f $X=12 $Y=0.555
+ $X2=0 $Y2=0
cc_1077 N_A_1525_21#_c_1521_n N_A_1864_47#_c_1852_n 0.0219541f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1078 N_A_1525_21#_c_1521_n N_A_1864_47#_c_1848_n 0.0248947f $X=12.105 $Y=1.53
+ $X2=0 $Y2=0
cc_1079 N_A_1525_21#_c_1521_n N_A_1864_47#_c_1850_n 0.00714757f $X=12.105
+ $Y=1.53 $X2=0 $Y2=0
cc_1080 N_A_1525_21#_M1007_g N_RESET_B_c_1940_n 0.00205214f $X=12 $Y=0.555
+ $X2=-0.19 $Y2=-0.24
cc_1081 N_A_1525_21#_c_1509_n N_RESET_B_c_1940_n 0.00512123f $X=12.615 $Y=0.84
+ $X2=-0.19 $Y2=-0.24
cc_1082 N_A_1525_21#_c_1519_n N_RESET_B_c_1940_n 0.00880997f $X=12.73 $Y=1.66
+ $X2=-0.19 $Y2=-0.24
cc_1083 N_A_1525_21#_c_1524_n N_RESET_B_c_1940_n 0.0025409f $X=12.25 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_1084 N_A_1525_21#_c_1514_n N_RESET_B_c_1940_n 0.0125484f $X=12 $Y=1.362
+ $X2=-0.19 $Y2=-0.24
cc_1085 N_A_1525_21#_c_1515_n N_RESET_B_c_1940_n 0.00419321f $X=12.215 $Y=1.32
+ $X2=-0.19 $Y2=-0.24
cc_1086 N_A_1525_21#_c_1509_n N_RESET_B_M1028_g 0.00647724f $X=12.615 $Y=0.84
+ $X2=0 $Y2=0
cc_1087 N_A_1525_21#_c_1511_n N_RESET_B_M1028_g 0.00441411f $X=12.73 $Y=0.43
+ $X2=0 $Y2=0
cc_1088 N_A_1525_21#_c_1515_n N_RESET_B_M1028_g 0.00206571f $X=12.215 $Y=1.32
+ $X2=0 $Y2=0
cc_1089 N_A_1525_21#_c_1509_n N_RESET_B_c_1942_n 0.0240868f $X=12.615 $Y=0.84
+ $X2=0 $Y2=0
cc_1090 N_A_1525_21#_c_1519_n N_RESET_B_c_1942_n 0.0197121f $X=12.73 $Y=1.66
+ $X2=0 $Y2=0
cc_1091 N_A_1525_21#_c_1514_n N_RESET_B_c_1942_n 0.00118349f $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1092 N_A_1525_21#_c_1515_n N_RESET_B_c_1942_n 0.0186459f $X=12.215 $Y=1.32
+ $X2=0 $Y2=0
cc_1093 N_A_1525_21#_c_1512_n N_VPWR_M1026_d 0.00308755f $X=7.97 $Y=1.32 $X2=0
+ $Y2=0
cc_1094 N_A_1525_21#_c_1523_n N_VPWR_M1026_d 0.00234234f $X=8.8 $Y=1.53 $X2=0
+ $Y2=0
cc_1095 N_A_1525_21#_c_1518_n N_VPWR_M1036_d 0.00323917f $X=12.345 $Y=1.66 $X2=0
+ $Y2=0
cc_1096 N_A_1525_21#_c_1524_n N_VPWR_M1036_d 2.3265e-19 $X=12.25 $Y=1.53 $X2=0
+ $Y2=0
cc_1097 N_A_1525_21#_c_1516_n N_VPWR_c_2033_n 0.0035996f $X=7.725 $Y=1.57 $X2=0
+ $Y2=0
cc_1098 N_A_1525_21#_c_1512_n N_VPWR_c_2033_n 0.011839f $X=7.97 $Y=1.32 $X2=0
+ $Y2=0
cc_1099 N_A_1525_21#_c_1523_n N_VPWR_c_2033_n 7.83548e-19 $X=8.8 $Y=1.53 $X2=0
+ $Y2=0
cc_1100 N_A_1525_21#_c_1513_n N_VPWR_c_2033_n 0.00112189f $X=7.725 $Y=1.362
+ $X2=0 $Y2=0
cc_1101 N_A_1525_21#_c_1516_n N_VPWR_c_2041_n 0.00702461f $X=7.725 $Y=1.57 $X2=0
+ $Y2=0
cc_1102 N_A_1525_21#_c_1517_n N_VPWR_c_2043_n 0.0138544f $X=11.92 $Y=1.57 $X2=0
+ $Y2=0
cc_1103 N_A_1525_21#_c_1516_n N_VPWR_c_2027_n 0.0077967f $X=7.725 $Y=1.57 $X2=0
+ $Y2=0
cc_1104 N_A_1525_21#_c_1517_n N_VPWR_c_2027_n 0.00360784f $X=11.92 $Y=1.57 $X2=0
+ $Y2=0
cc_1105 N_A_1525_21#_c_1517_n N_VPWR_c_2052_n 0.00310943f $X=11.92 $Y=1.57 $X2=0
+ $Y2=0
cc_1106 N_A_1525_21#_c_1523_n A_1710_329# 0.00353943f $X=8.8 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1107 N_A_1525_21#_c_1509_n N_VGND_c_2432_n 0.00307931f $X=12.615 $Y=0.84
+ $X2=0 $Y2=0
cc_1108 N_A_1525_21#_c_1511_n N_VGND_c_2432_n 0.015455f $X=12.73 $Y=0.43 $X2=0
+ $Y2=0
cc_1109 N_A_1525_21#_M1021_g N_VGND_c_2440_n 0.00664108f $X=7.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1110 N_A_1525_21#_M1007_g N_VGND_c_2441_n 0.00357877f $X=12 $Y=0.555 $X2=0
+ $Y2=0
cc_1111 N_A_1525_21#_c_1509_n N_VGND_c_2441_n 0.00387343f $X=12.615 $Y=0.84
+ $X2=0 $Y2=0
cc_1112 N_A_1525_21#_c_1510_n N_VGND_c_2441_n 7.06816e-19 $X=12.345 $Y=0.84
+ $X2=0 $Y2=0
cc_1113 N_A_1525_21#_c_1511_n N_VGND_c_2441_n 0.0130551f $X=12.73 $Y=0.43 $X2=0
+ $Y2=0
cc_1114 N_A_1525_21#_M1028_s N_VGND_c_2444_n 0.00602329f $X=12.605 $Y=0.235
+ $X2=0 $Y2=0
cc_1115 N_A_1525_21#_M1021_g N_VGND_c_2444_n 0.00661646f $X=7.7 $Y=0.555 $X2=0
+ $Y2=0
cc_1116 N_A_1525_21#_M1007_g N_VGND_c_2444_n 0.00669047f $X=12 $Y=0.555 $X2=0
+ $Y2=0
cc_1117 N_A_1525_21#_c_1509_n N_VGND_c_2444_n 0.00696043f $X=12.615 $Y=0.84
+ $X2=0 $Y2=0
cc_1118 N_A_1525_21#_c_1510_n N_VGND_c_2444_n 0.00161396f $X=12.345 $Y=0.84
+ $X2=0 $Y2=0
cc_1119 N_A_1525_21#_c_1511_n N_VGND_c_2444_n 0.0075831f $X=12.73 $Y=0.43 $X2=0
+ $Y2=0
cc_1120 N_A_1525_21#_M1021_g N_A_1353_47#_c_2647_n 0.0106345f $X=7.7 $Y=0.555
+ $X2=0 $Y2=0
cc_1121 N_A_1525_21#_c_1510_n N_A_2216_47#_M1007_d 0.00390488f $X=12.345 $Y=0.84
+ $X2=0 $Y2=0
cc_1122 N_A_1525_21#_M1007_g N_A_2216_47#_c_2678_n 0.0123888f $X=12 $Y=0.555
+ $X2=0 $Y2=0
cc_1123 N_A_1525_21#_c_1510_n N_A_2216_47#_c_2678_n 0.0138009f $X=12.345 $Y=0.84
+ $X2=0 $Y2=0
cc_1124 N_A_1525_21#_c_1511_n N_A_2216_47#_c_2678_n 0.0149851f $X=12.73 $Y=0.43
+ $X2=0 $Y2=0
cc_1125 N_A_1525_21#_c_1514_n N_A_2216_47#_c_2678_n 5.45076e-19 $X=12 $Y=1.362
+ $X2=0 $Y2=0
cc_1126 N_A_2058_21#_c_1707_n N_A_1864_47#_c_1845_n 0.0137054f $X=11.73 $Y=2
+ $X2=0 $Y2=0
cc_1127 N_A_2058_21#_c_1671_n N_A_1864_47#_c_1845_n 0.00730958f $X=11.822
+ $Y=1.915 $X2=0 $Y2=0
cc_1128 N_A_2058_21#_c_1724_n N_A_1864_47#_c_1845_n 4.29792e-19 $X=11.275 $Y=2
+ $X2=0 $Y2=0
cc_1129 N_A_2058_21#_c_1671_n N_A_1864_47#_M1040_g 0.00859654f $X=11.822
+ $Y=1.915 $X2=0 $Y2=0
cc_1130 N_A_2058_21#_c_1700_n N_A_1864_47#_M1040_g 0.00809722f $X=11.75 $Y=0.73
+ $X2=0 $Y2=0
cc_1131 N_A_2058_21#_c_1674_n N_A_1864_47#_c_1856_n 0.00223829f $X=10.39 $Y=1.99
+ $X2=0 $Y2=0
cc_1132 N_A_2058_21#_M1014_g N_A_1864_47#_c_1859_n 0.00176841f $X=10.365
+ $Y=0.445 $X2=0 $Y2=0
cc_1133 N_A_2058_21#_M1014_g N_A_1864_47#_c_1847_n 0.0130772f $X=10.365 $Y=0.445
+ $X2=0 $Y2=0
cc_1134 N_A_2058_21#_M1014_g N_A_1864_47#_c_1852_n 0.0099202f $X=10.365 $Y=0.445
+ $X2=0 $Y2=0
cc_1135 N_A_2058_21#_c_1674_n N_A_1864_47#_c_1852_n 0.00510579f $X=10.39 $Y=1.99
+ $X2=0 $Y2=0
cc_1136 N_A_2058_21#_c_1679_n N_A_1864_47#_c_1852_n 0.0251598f $X=10.485 $Y=1.74
+ $X2=0 $Y2=0
cc_1137 N_A_2058_21#_c_1738_p N_A_1864_47#_c_1852_n 0.0135158f $X=10.7 $Y=2
+ $X2=0 $Y2=0
cc_1138 N_A_2058_21#_M1014_g N_A_1864_47#_c_1848_n 0.0117362f $X=10.365 $Y=0.445
+ $X2=0 $Y2=0
cc_1139 N_A_2058_21#_c_1674_n N_A_1864_47#_c_1848_n 0.00161733f $X=10.39 $Y=1.99
+ $X2=0 $Y2=0
cc_1140 N_A_2058_21#_c_1679_n N_A_1864_47#_c_1848_n 0.018607f $X=10.485 $Y=1.74
+ $X2=0 $Y2=0
cc_1141 N_A_2058_21#_c_1680_n N_A_1864_47#_c_1848_n 0.00697334f $X=11.19 $Y=2
+ $X2=0 $Y2=0
cc_1142 N_A_2058_21#_c_1724_n N_A_1864_47#_c_1848_n 0.00162703f $X=11.275 $Y=2
+ $X2=0 $Y2=0
cc_1143 N_A_2058_21#_c_1707_n N_A_1864_47#_c_1850_n 0.0015192f $X=11.73 $Y=2
+ $X2=0 $Y2=0
cc_1144 N_A_2058_21#_c_1671_n N_A_1864_47#_c_1850_n 0.019966f $X=11.822 $Y=1.915
+ $X2=0 $Y2=0
cc_1145 N_A_2058_21#_c_1724_n N_A_1864_47#_c_1850_n 0.00106299f $X=11.275 $Y=2
+ $X2=0 $Y2=0
cc_1146 N_A_2058_21#_c_1663_n N_RESET_B_c_1940_n 0.0280001f $X=13.5 $Y=1.41
+ $X2=-0.19 $Y2=-0.24
cc_1147 N_A_2058_21#_c_1682_n N_RESET_B_c_1940_n 0.0161897f $X=13.26 $Y=2
+ $X2=-0.19 $Y2=-0.24
cc_1148 N_A_2058_21#_c_1683_n N_RESET_B_c_1940_n 0.010093f $X=13.345 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1149 N_A_2058_21#_c_1672_n N_RESET_B_c_1940_n 6.94961e-19 $X=13.44 $Y=1.16
+ $X2=-0.19 $Y2=-0.24
cc_1150 N_A_2058_21#_c_1663_n N_RESET_B_M1028_g 0.0180605f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1151 N_A_2058_21#_c_1664_n N_RESET_B_M1028_g 0.0162962f $X=13.525 $Y=0.995
+ $X2=0 $Y2=0
cc_1152 N_A_2058_21#_c_1672_n N_RESET_B_M1028_g 0.0022133f $X=13.44 $Y=1.16
+ $X2=0 $Y2=0
cc_1153 N_A_2058_21#_c_1663_n N_RESET_B_c_1942_n 7.57946e-19 $X=13.5 $Y=1.41
+ $X2=0 $Y2=0
cc_1154 N_A_2058_21#_c_1682_n N_RESET_B_c_1942_n 0.00426718f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1155 N_A_2058_21#_c_1672_n N_RESET_B_c_1942_n 0.0196794f $X=13.44 $Y=1.16
+ $X2=0 $Y2=0
cc_1156 N_A_2058_21#_c_1666_n N_A_2845_47#_c_1972_n 0.0107367f $X=14.435
+ $Y=1.025 $X2=0 $Y2=0
cc_1157 N_A_2058_21#_c_1667_n N_A_2845_47#_c_1972_n 0.00396981f $X=14.435
+ $Y=1.535 $X2=0 $Y2=0
cc_1158 N_A_2058_21#_c_1677_n N_A_2845_47#_c_1972_n 0.0137907f $X=14.585 $Y=1.69
+ $X2=0 $Y2=0
cc_1159 N_A_2058_21#_c_1678_n N_A_2845_47#_c_1972_n 0.00569695f $X=14.435
+ $Y=1.612 $X2=0 $Y2=0
cc_1160 N_A_2058_21#_c_1666_n N_A_2845_47#_c_1973_n 0.00187884f $X=14.435
+ $Y=1.025 $X2=0 $Y2=0
cc_1161 N_A_2058_21#_c_1668_n N_A_2845_47#_c_1973_n 0.0139892f $X=14.61 $Y=0.73
+ $X2=0 $Y2=0
cc_1162 N_A_2058_21#_c_1665_n N_A_2845_47#_c_1978_n 0.00177826f $X=14.36 $Y=1.16
+ $X2=0 $Y2=0
cc_1163 N_A_2058_21#_c_1677_n N_A_2845_47#_c_1978_n 0.00258107f $X=14.585
+ $Y=1.69 $X2=0 $Y2=0
cc_1164 N_A_2058_21#_c_1677_n N_A_2845_47#_c_1979_n 0.00727682f $X=14.585
+ $Y=1.69 $X2=0 $Y2=0
cc_1165 N_A_2058_21#_c_1666_n N_A_2845_47#_c_1974_n 0.00418753f $X=14.435
+ $Y=1.025 $X2=0 $Y2=0
cc_1166 N_A_2058_21#_c_1668_n N_A_2845_47#_c_1974_n 0.00426998f $X=14.61 $Y=0.73
+ $X2=0 $Y2=0
cc_1167 N_A_2058_21#_c_1669_n N_A_2845_47#_c_1974_n 0.0108096f $X=14.61 $Y=0.805
+ $X2=0 $Y2=0
cc_1168 N_A_2058_21#_c_1669_n N_A_2845_47#_c_1975_n 0.00524474f $X=14.61
+ $Y=0.805 $X2=0 $Y2=0
cc_1169 N_A_2058_21#_c_1678_n N_A_2845_47#_c_1975_n 0.00463915f $X=14.435
+ $Y=1.612 $X2=0 $Y2=0
cc_1170 N_A_2058_21#_c_1667_n N_A_2845_47#_c_1981_n 0.00757432f $X=14.435
+ $Y=1.535 $X2=0 $Y2=0
cc_1171 N_A_2058_21#_c_1677_n N_A_2845_47#_c_1981_n 0.00121925f $X=14.585
+ $Y=1.69 $X2=0 $Y2=0
cc_1172 N_A_2058_21#_c_1678_n N_A_2845_47#_c_1981_n 0.0107605f $X=14.435
+ $Y=1.612 $X2=0 $Y2=0
cc_1173 N_A_2058_21#_c_1665_n N_A_2845_47#_c_1976_n 0.00648764f $X=14.36 $Y=1.16
+ $X2=0 $Y2=0
cc_1174 N_A_2058_21#_c_1666_n N_A_2845_47#_c_1976_n 0.00125393f $X=14.435
+ $Y=1.025 $X2=0 $Y2=0
cc_1175 N_A_2058_21#_c_1667_n N_A_2845_47#_c_1976_n 0.00125393f $X=14.435
+ $Y=1.535 $X2=0 $Y2=0
cc_1176 N_A_2058_21#_c_1670_n N_A_2845_47#_c_1976_n 0.00774835f $X=14.435
+ $Y=1.16 $X2=0 $Y2=0
cc_1177 N_A_2058_21#_c_1680_n N_VPWR_M1029_d 0.00134994f $X=11.19 $Y=2 $X2=0
+ $Y2=0
cc_1178 N_A_2058_21#_c_1738_p N_VPWR_M1029_d 0.0017095f $X=10.7 $Y=2 $X2=0 $Y2=0
cc_1179 N_A_2058_21#_c_1682_n N_VPWR_M1036_d 0.0046603f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1180 N_A_2058_21#_c_1682_n N_VPWR_M1017_d 0.00809741f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1181 N_A_2058_21#_c_1683_n N_VPWR_M1017_d 0.00503162f $X=13.345 $Y=1.915
+ $X2=0 $Y2=0
cc_1182 N_A_2058_21#_c_1677_n N_VPWR_c_2034_n 0.00820678f $X=14.585 $Y=1.69
+ $X2=0 $Y2=0
cc_1183 N_A_2058_21#_c_1663_n N_VPWR_c_2038_n 0.0103271f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1184 N_A_2058_21#_c_1682_n N_VPWR_c_2038_n 0.00920797f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1185 N_A_2058_21#_c_1674_n N_VPWR_c_2042_n 0.00640896f $X=10.39 $Y=1.99 $X2=0
+ $Y2=0
cc_1186 N_A_2058_21#_c_1738_p N_VPWR_c_2042_n 0.00180198f $X=10.7 $Y=2 $X2=0
+ $Y2=0
cc_1187 N_A_2058_21#_c_1698_n N_VPWR_c_2043_n 0.00353321f $X=11.275 $Y=2.21
+ $X2=0 $Y2=0
cc_1188 N_A_2058_21#_c_1682_n N_VPWR_c_2043_n 0.091697f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1189 N_A_2058_21#_c_1663_n N_VPWR_c_2044_n 0.00622633f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1190 N_A_2058_21#_c_1677_n N_VPWR_c_2044_n 0.00579366f $X=14.585 $Y=1.69
+ $X2=0 $Y2=0
cc_1191 N_A_2058_21#_M1002_d N_VPWR_c_2027_n 0.00350614f $X=11.07 $Y=2.065 $X2=0
+ $Y2=0
cc_1192 N_A_2058_21#_c_1674_n N_VPWR_c_2027_n 0.0109362f $X=10.39 $Y=1.99 $X2=0
+ $Y2=0
cc_1193 N_A_2058_21#_c_1663_n N_VPWR_c_2027_n 0.0117622f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1194 N_A_2058_21#_c_1677_n N_VPWR_c_2027_n 0.0115044f $X=14.585 $Y=1.69 $X2=0
+ $Y2=0
cc_1195 N_A_2058_21#_c_1680_n N_VPWR_c_2027_n 0.0082738f $X=11.19 $Y=2 $X2=0
+ $Y2=0
cc_1196 N_A_2058_21#_c_1738_p N_VPWR_c_2027_n 0.00403319f $X=10.7 $Y=2 $X2=0
+ $Y2=0
cc_1197 N_A_2058_21#_c_1698_n N_VPWR_c_2027_n 0.00608739f $X=11.275 $Y=2.21
+ $X2=0 $Y2=0
cc_1198 N_A_2058_21#_c_1707_n N_VPWR_c_2027_n 0.00955121f $X=11.73 $Y=2 $X2=0
+ $Y2=0
cc_1199 N_A_2058_21#_c_1682_n N_VPWR_c_2027_n 0.00720077f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1200 N_A_2058_21#_c_1726_n N_VPWR_c_2027_n 0.0051168f $X=11.822 $Y=2 $X2=0
+ $Y2=0
cc_1201 N_A_2058_21#_c_1674_n N_VPWR_c_2051_n 0.00535636f $X=10.39 $Y=1.99 $X2=0
+ $Y2=0
cc_1202 N_A_2058_21#_c_1680_n N_VPWR_c_2051_n 0.0107574f $X=11.19 $Y=2 $X2=0
+ $Y2=0
cc_1203 N_A_2058_21#_c_1738_p N_VPWR_c_2051_n 0.0134619f $X=10.7 $Y=2 $X2=0
+ $Y2=0
cc_1204 N_A_2058_21#_c_1698_n N_VPWR_c_2051_n 0.0059431f $X=11.275 $Y=2.21 $X2=0
+ $Y2=0
cc_1205 N_A_2058_21#_c_1680_n N_VPWR_c_2052_n 0.00443454f $X=11.19 $Y=2 $X2=0
+ $Y2=0
cc_1206 N_A_2058_21#_c_1698_n N_VPWR_c_2052_n 0.00725596f $X=11.275 $Y=2.21
+ $X2=0 $Y2=0
cc_1207 N_A_2058_21#_c_1707_n N_VPWR_c_2052_n 0.00535373f $X=11.73 $Y=2 $X2=0
+ $Y2=0
cc_1208 N_A_2058_21#_c_1682_n N_VPWR_c_2052_n 3.92726e-19 $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1209 N_A_2058_21#_c_1726_n N_VPWR_c_2052_n 0.00289943f $X=11.822 $Y=2 $X2=0
+ $Y2=0
cc_1210 N_A_2058_21#_c_1707_n A_2320_329# 0.00234722f $X=11.73 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1211 N_A_2058_21#_c_1671_n A_2320_329# 0.00307681f $X=11.822 $Y=1.915
+ $X2=-0.19 $Y2=-0.24
cc_1212 N_A_2058_21#_c_1726_n A_2320_329# 7.67806e-19 $X=11.822 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_1213 N_A_2058_21#_c_1663_n N_Q_N_c_2380_n 0.0276916f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1214 N_A_2058_21#_c_1665_n N_Q_N_c_2380_n 0.00383439f $X=14.36 $Y=1.16 $X2=0
+ $Y2=0
cc_1215 N_A_2058_21#_c_1667_n N_Q_N_c_2380_n 0.00199673f $X=14.435 $Y=1.535
+ $X2=0 $Y2=0
cc_1216 N_A_2058_21#_c_1677_n N_Q_N_c_2380_n 0.00246924f $X=14.585 $Y=1.69 $X2=0
+ $Y2=0
cc_1217 N_A_2058_21#_c_1682_n N_Q_N_c_2380_n 0.0095008f $X=13.26 $Y=2 $X2=0
+ $Y2=0
cc_1218 N_A_2058_21#_c_1683_n N_Q_N_c_2380_n 0.024475f $X=13.345 $Y=1.915 $X2=0
+ $Y2=0
cc_1219 N_A_2058_21#_c_1664_n Q_N 0.0104384f $X=13.525 $Y=0.995 $X2=0 $Y2=0
cc_1220 N_A_2058_21#_c_1665_n Q_N 0.00368855f $X=14.36 $Y=1.16 $X2=0 $Y2=0
cc_1221 N_A_2058_21#_c_1663_n Q_N 0.00173083f $X=13.5 $Y=1.41 $X2=0 $Y2=0
cc_1222 N_A_2058_21#_c_1664_n Q_N 0.00912135f $X=13.525 $Y=0.995 $X2=0 $Y2=0
cc_1223 N_A_2058_21#_c_1665_n Q_N 0.0308894f $X=14.36 $Y=1.16 $X2=0 $Y2=0
cc_1224 N_A_2058_21#_c_1667_n Q_N 5.09084e-19 $X=14.435 $Y=1.535 $X2=0 $Y2=0
cc_1225 N_A_2058_21#_c_1669_n Q_N 0.00189912f $X=14.61 $Y=0.805 $X2=0 $Y2=0
cc_1226 N_A_2058_21#_c_1683_n Q_N 0.00191463f $X=13.345 $Y=1.915 $X2=0 $Y2=0
cc_1227 N_A_2058_21#_c_1672_n Q_N 0.0157374f $X=13.44 $Y=1.16 $X2=0 $Y2=0
cc_1228 N_A_2058_21#_M1014_g N_VGND_c_2431_n 0.00910937f $X=10.365 $Y=0.445
+ $X2=0 $Y2=0
cc_1229 N_A_2058_21#_c_1663_n N_VGND_c_2432_n 0.00282689f $X=13.5 $Y=1.41 $X2=0
+ $Y2=0
cc_1230 N_A_2058_21#_c_1664_n N_VGND_c_2432_n 0.00322756f $X=13.525 $Y=0.995
+ $X2=0 $Y2=0
cc_1231 N_A_2058_21#_c_1672_n N_VGND_c_2432_n 0.0115066f $X=13.44 $Y=1.16 $X2=0
+ $Y2=0
cc_1232 N_A_2058_21#_c_1668_n N_VGND_c_2433_n 0.00446058f $X=14.61 $Y=0.73 $X2=0
+ $Y2=0
cc_1233 N_A_2058_21#_M1014_g N_VGND_c_2436_n 0.0046653f $X=10.365 $Y=0.445 $X2=0
+ $Y2=0
cc_1234 N_A_2058_21#_c_1664_n N_VGND_c_2442_n 0.00585385f $X=13.525 $Y=0.995
+ $X2=0 $Y2=0
cc_1235 N_A_2058_21#_c_1668_n N_VGND_c_2442_n 0.00585385f $X=14.61 $Y=0.73 $X2=0
+ $Y2=0
cc_1236 N_A_2058_21#_c_1669_n N_VGND_c_2442_n 6.23112e-19 $X=14.61 $Y=0.805
+ $X2=0 $Y2=0
cc_1237 N_A_2058_21#_M1040_d N_VGND_c_2444_n 0.00252169f $X=11.61 $Y=0.235 $X2=0
+ $Y2=0
cc_1238 N_A_2058_21#_M1014_g N_VGND_c_2444_n 0.00461364f $X=10.365 $Y=0.445
+ $X2=0 $Y2=0
cc_1239 N_A_2058_21#_c_1664_n N_VGND_c_2444_n 0.0121987f $X=13.525 $Y=0.995
+ $X2=0 $Y2=0
cc_1240 N_A_2058_21#_c_1668_n N_VGND_c_2444_n 0.0122913f $X=14.61 $Y=0.73 $X2=0
+ $Y2=0
cc_1241 N_A_2058_21#_c_1669_n N_VGND_c_2444_n 3.45313e-19 $X=14.61 $Y=0.805
+ $X2=0 $Y2=0
cc_1242 N_A_2058_21#_M1040_d N_A_2216_47#_c_2678_n 0.00428432f $X=11.61 $Y=0.235
+ $X2=0 $Y2=0
cc_1243 N_A_2058_21#_c_1700_n N_A_2216_47#_c_2678_n 0.0148333f $X=11.75 $Y=0.73
+ $X2=0 $Y2=0
cc_1244 N_A_1864_47#_c_1856_n N_VPWR_c_2042_n 0.0425549f $X=10.06 $Y=2.335 $X2=0
+ $Y2=0
cc_1245 N_A_1864_47#_c_1845_n N_VPWR_c_2043_n 0.00213368f $X=11.51 $Y=1.57 $X2=0
+ $Y2=0
cc_1246 N_A_1864_47#_M1042_d N_VPWR_c_2027_n 0.00228605f $X=9.37 $Y=2.065 $X2=0
+ $Y2=0
cc_1247 N_A_1864_47#_c_1845_n N_VPWR_c_2027_n 0.00687753f $X=11.51 $Y=1.57 $X2=0
+ $Y2=0
cc_1248 N_A_1864_47#_c_1856_n N_VPWR_c_2027_n 0.0306792f $X=10.06 $Y=2.335 $X2=0
+ $Y2=0
cc_1249 N_A_1864_47#_c_1845_n N_VPWR_c_2051_n 0.00132483f $X=11.51 $Y=1.57 $X2=0
+ $Y2=0
cc_1250 N_A_1864_47#_c_1845_n N_VPWR_c_2052_n 0.00510113f $X=11.51 $Y=1.57 $X2=0
+ $Y2=0
cc_1251 N_A_1864_47#_c_1856_n A_1968_413# 0.011644f $X=10.06 $Y=2.335 $X2=-0.19
+ $Y2=-0.24
cc_1252 N_A_1864_47#_c_1852_n A_1968_413# 0.00579594f $X=10.145 $Y=2.25
+ $X2=-0.19 $Y2=-0.24
cc_1253 N_A_1864_47#_c_1859_n N_VGND_c_2431_n 0.0157316f $X=10.06 $Y=0.365 $X2=0
+ $Y2=0
cc_1254 N_A_1864_47#_c_1847_n N_VGND_c_2431_n 0.00418333f $X=10.145 $Y=1.235
+ $X2=0 $Y2=0
cc_1255 N_A_1864_47#_c_1859_n N_VGND_c_2436_n 0.0467275f $X=10.06 $Y=0.365 $X2=0
+ $Y2=0
cc_1256 N_A_1864_47#_M1040_g N_VGND_c_2441_n 0.00357877f $X=11.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1257 N_A_1864_47#_M1010_d N_VGND_c_2444_n 0.00351839f $X=9.32 $Y=0.235 $X2=0
+ $Y2=0
cc_1258 N_A_1864_47#_M1040_g N_VGND_c_2444_n 0.00568762f $X=11.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1259 N_A_1864_47#_c_1859_n N_VGND_c_2444_n 0.0138052f $X=10.06 $Y=0.365 $X2=0
+ $Y2=0
cc_1260 N_A_1864_47#_c_1859_n A_1992_47# 0.00548351f $X=10.06 $Y=0.365 $X2=-0.19
+ $Y2=-0.24
cc_1261 N_A_1864_47#_c_1847_n A_1992_47# 0.00500854f $X=10.145 $Y=1.235
+ $X2=-0.19 $Y2=-0.24
cc_1262 N_A_1864_47#_c_1845_n N_A_2216_47#_c_2678_n 2.09367e-19 $X=11.51 $Y=1.57
+ $X2=0 $Y2=0
cc_1263 N_A_1864_47#_M1040_g N_A_2216_47#_c_2678_n 0.0120232f $X=11.535 $Y=0.555
+ $X2=0 $Y2=0
cc_1264 N_A_1864_47#_c_1850_n N_A_2216_47#_c_2678_n 0.00242255f $X=11.425
+ $Y=1.24 $X2=0 $Y2=0
cc_1265 N_A_1864_47#_c_1845_n N_A_2216_47#_c_2687_n 4.61885e-19 $X=11.51 $Y=1.57
+ $X2=0 $Y2=0
cc_1266 N_A_1864_47#_M1040_g N_A_2216_47#_c_2687_n 0.00111354f $X=11.535
+ $Y=0.555 $X2=0 $Y2=0
cc_1267 N_A_1864_47#_c_1850_n N_A_2216_47#_c_2687_n 0.00244558f $X=11.425
+ $Y=1.24 $X2=0 $Y2=0
cc_1268 N_RESET_B_c_1940_n N_VPWR_c_2037_n 0.00774065f $X=12.965 $Y=1.43 $X2=0
+ $Y2=0
cc_1269 N_RESET_B_M1028_g N_VGND_c_2432_n 0.00721493f $X=12.99 $Y=0.445 $X2=0
+ $Y2=0
cc_1270 N_RESET_B_M1028_g N_VGND_c_2441_n 0.00585385f $X=12.99 $Y=0.445 $X2=0
+ $Y2=0
cc_1271 N_RESET_B_M1028_g N_VGND_c_2444_n 0.012196f $X=12.99 $Y=0.445 $X2=0
+ $Y2=0
cc_1272 N_A_2845_47#_c_1972_n N_VPWR_c_2034_n 0.0177905f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1273 N_A_2845_47#_c_1978_n N_VPWR_c_2034_n 0.0395619f $X=14.392 $Y=1.852
+ $X2=0 $Y2=0
cc_1274 N_A_2845_47#_c_1975_n N_VPWR_c_2034_n 0.0107904f $X=15.005 $Y=1.16 $X2=0
+ $Y2=0
cc_1275 N_A_2845_47#_c_1979_n N_VPWR_c_2044_n 0.0136982f $X=14.35 $Y=1.91 $X2=0
+ $Y2=0
cc_1276 N_A_2845_47#_c_1972_n N_VPWR_c_2045_n 0.00622633f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1277 N_A_2845_47#_c_1972_n N_VPWR_c_2027_n 0.0114577f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1278 N_A_2845_47#_c_1979_n N_VPWR_c_2027_n 0.00938744f $X=14.35 $Y=1.91 $X2=0
+ $Y2=0
cc_1279 N_A_2845_47#_c_1978_n N_Q_N_c_2380_n 0.0560009f $X=14.392 $Y=1.852 $X2=0
+ $Y2=0
cc_1280 N_A_2845_47#_c_1981_n N_Q_N_c_2380_n 0.0242286f $X=14.392 $Y=1.725 $X2=0
+ $Y2=0
cc_1281 N_A_2845_47#_c_1974_n Q_N 0.0527371f $X=14.4 $Y=0.51 $X2=0 $Y2=0
cc_1282 N_A_2845_47#_c_1981_n Q_N 0.0033402f $X=14.392 $Y=1.725 $X2=0 $Y2=0
cc_1283 N_A_2845_47#_c_1976_n Q_N 0.0234515f $X=14.417 $Y=1.16 $X2=0 $Y2=0
cc_1284 N_A_2845_47#_c_1972_n N_Q_c_2413_n 0.00882117f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1285 N_A_2845_47#_c_1972_n N_Q_c_2411_n 0.00751577f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1286 N_A_2845_47#_c_1973_n N_Q_c_2411_n 0.0182741f $X=15.135 $Y=0.995 $X2=0
+ $Y2=0
cc_1287 N_A_2845_47#_c_1975_n N_Q_c_2411_n 0.0220839f $X=15.005 $Y=1.16 $X2=0
+ $Y2=0
cc_1288 N_A_2845_47#_c_1972_n N_VGND_c_2433_n 0.00317666f $X=15.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1289 N_A_2845_47#_c_1973_n N_VGND_c_2433_n 0.00317237f $X=15.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1290 N_A_2845_47#_c_1975_n N_VGND_c_2433_n 0.0108565f $X=15.005 $Y=1.16 $X2=0
+ $Y2=0
cc_1291 N_A_2845_47#_c_1974_n N_VGND_c_2442_n 0.0128467f $X=14.4 $Y=0.51 $X2=0
+ $Y2=0
cc_1292 N_A_2845_47#_c_1973_n N_VGND_c_2443_n 0.00585385f $X=15.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1293 N_A_2845_47#_M1043_s N_VGND_c_2444_n 0.00585424f $X=14.225 $Y=0.235
+ $X2=0 $Y2=0
cc_1294 N_A_2845_47#_c_1973_n N_VGND_c_2444_n 0.0118254f $X=15.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1295 N_A_2845_47#_c_1974_n N_VGND_c_2444_n 0.00781789f $X=14.4 $Y=0.51 $X2=0
+ $Y2=0
cc_1296 N_VPWR_c_2027_n N_A_483_47#_M1044_d 0.00374021f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1297 N_VPWR_c_2030_n N_A_483_47#_c_2248_n 0.0148576f $X=1.72 $Y=1.97 $X2=0
+ $Y2=0
cc_1298 N_VPWR_c_2035_n N_A_483_47#_c_2248_n 0.0160506f $X=3.51 $Y=2.72 $X2=0
+ $Y2=0
cc_1299 N_VPWR_c_2027_n N_A_483_47#_c_2248_n 0.00641613f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1300 N_VPWR_c_2040_n N_A_483_47#_c_2247_n 0.0118139f $X=6.205 $Y=2.72 $X2=0
+ $Y2=0
cc_1301 N_VPWR_c_2027_n N_A_483_47#_c_2247_n 0.00308197f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1302 N_VPWR_c_2027_n A_810_413# 0.00275601f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1303 N_VPWR_c_2027_n A_1105_413# 0.00374905f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1304 N_VPWR_c_2027_n A_1469_329# 0.00291655f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1305 N_VPWR_c_2027_n A_1710_329# 0.00874151f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1306 N_VPWR_c_2027_n A_1968_413# 0.00595f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1307 N_VPWR_c_2027_n A_2320_329# 0.00268452f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1308 N_VPWR_c_2027_n N_Q_N_M1039_d 0.00733619f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1309 N_VPWR_c_2034_n N_Q_N_c_2380_n 0.00161771f $X=14.875 $Y=1.94 $X2=0 $Y2=0
cc_1310 N_VPWR_c_2038_n N_Q_N_c_2380_n 0.0116804f $X=13.43 $Y=2.53 $X2=0 $Y2=0
cc_1311 N_VPWR_c_2044_n N_Q_N_c_2380_n 0.0267723f $X=14.745 $Y=2.72 $X2=0 $Y2=0
cc_1312 N_VPWR_c_2027_n N_Q_N_c_2380_n 0.0145574f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1313 N_VPWR_c_2027_n N_Q_M1016_d 0.00430086f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1314 N_VPWR_c_2034_n Q 0.0437047f $X=14.875 $Y=1.94 $X2=0 $Y2=0
cc_1315 N_VPWR_c_2045_n Q 0.0200025f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1316 N_VPWR_c_2027_n Q 0.0108988f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1317 N_A_483_47#_c_2247_n N_VGND_c_2434_n 0.00877567f $X=4.73 $Y=0.47 $X2=0
+ $Y2=0
cc_1318 N_A_483_47#_c_2241_n N_VGND_c_2439_n 0.0254868f $X=2.87 $Y=0.43 $X2=0
+ $Y2=0
cc_1319 N_A_483_47#_M1024_d N_VGND_c_2444_n 0.00273222f $X=2.415 $Y=0.235 $X2=0
+ $Y2=0
cc_1320 N_A_483_47#_M1035_d N_VGND_c_2444_n 0.00352561f $X=4.53 $Y=0.235 $X2=0
+ $Y2=0
cc_1321 N_A_483_47#_c_2241_n N_VGND_c_2444_n 0.00710198f $X=2.87 $Y=0.43 $X2=0
+ $Y2=0
cc_1322 N_A_483_47#_c_2247_n N_VGND_c_2444_n 0.00300364f $X=4.73 $Y=0.47 $X2=0
+ $Y2=0
cc_1323 Q_N N_VGND_c_2442_n 0.0280021f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1324 N_Q_N_M1005_d N_VGND_c_2444_n 0.00690705f $X=13.6 $Y=0.235 $X2=0 $Y2=0
cc_1325 Q_N N_VGND_c_2444_n 0.0152879f $X=13.945 $Y=0.425 $X2=0 $Y2=0
cc_1326 Q N_VGND_c_2443_n 0.0197547f $X=15.325 $Y=0.425 $X2=0 $Y2=0
cc_1327 N_Q_M1047_d N_VGND_c_2444_n 0.00387172f $X=15.21 $Y=0.235 $X2=0 $Y2=0
cc_1328 Q N_VGND_c_2444_n 0.0108902f $X=15.325 $Y=0.425 $X2=0 $Y2=0
cc_1329 N_VGND_c_2444_n A_411_47# 0.00145468f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1330 N_VGND_c_2444_n A_824_47# 0.00373999f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1331 N_VGND_c_2444_n A_1121_47# 0.0025914f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1332 N_VGND_c_2444_n N_A_1353_47#_M1009_d 0.00292724f $X=15.41 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1333 N_VGND_c_2444_n N_A_1353_47#_M1021_d 0.00201692f $X=15.41 $Y=0 $X2=0
+ $Y2=0
cc_1334 N_VGND_c_2440_n N_A_1353_47#_c_2647_n 0.0247845f $X=8.29 $Y=0 $X2=0
+ $Y2=0
cc_1335 N_VGND_c_2444_n N_A_1353_47#_c_2647_n 0.00350344f $X=15.41 $Y=0 $X2=0
+ $Y2=0
cc_1336 N_VGND_c_2440_n N_A_1353_47#_c_2650_n 0.00242553f $X=8.29 $Y=0 $X2=0
+ $Y2=0
cc_1337 N_VGND_c_2440_n N_A_1353_47#_c_2657_n 0.0600502f $X=8.29 $Y=0 $X2=0
+ $Y2=0
cc_1338 N_VGND_c_2444_n N_A_1353_47#_c_2657_n 0.017744f $X=15.41 $Y=0 $X2=0
+ $Y2=0
cc_1339 N_VGND_c_2444_n A_1769_47# 0.00467499f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1340 N_VGND_c_2444_n A_1992_47# 0.00264886f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1341 N_VGND_c_2444_n N_A_2216_47#_M1000_d 0.00304369f $X=15.41 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_1342 N_VGND_c_2444_n N_A_2216_47#_M1007_d 0.00224765f $X=15.41 $Y=0 $X2=0
+ $Y2=0
cc_1343 N_VGND_c_2431_n N_A_2216_47#_c_2675_n 0.0121987f $X=10.635 $Y=0.36 $X2=0
+ $Y2=0
cc_1344 N_VGND_c_2441_n N_A_2216_47#_c_2675_n 0.0642117f $X=13.1 $Y=0 $X2=0
+ $Y2=0
cc_1345 N_VGND_c_2444_n N_A_2216_47#_c_2675_n 0.0407459f $X=15.41 $Y=0 $X2=0
+ $Y2=0
cc_1346 N_VGND_c_2441_n N_A_2216_47#_c_2678_n 0.0113648f $X=13.1 $Y=0 $X2=0
+ $Y2=0
cc_1347 N_VGND_c_2444_n N_A_2216_47#_c_2678_n 0.00654393f $X=15.41 $Y=0 $X2=0
+ $Y2=0
