# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.125000 0.995000 0.435000 1.615000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 0.995000 1.080000 1.325000 ;
    END
  END B
  PIN X
    ANTENNADIFFAREA  1.061500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.680000 0.515000 1.870000 0.615000 ;
        RECT 1.680000 0.615000 3.570000 0.845000 ;
        RECT 1.680000 1.535000 3.570000 1.760000 ;
        RECT 1.680000 1.760000 1.870000 2.465000 ;
        RECT 2.640000 0.255000 2.830000 0.615000 ;
        RECT 2.640000 1.760000 3.570000 1.765000 ;
        RECT 2.640000 1.765000 2.830000 2.465000 ;
        RECT 3.290000 0.845000 3.570000 1.535000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.095000  0.255000 0.425000 0.615000 ;
      RECT 0.095000  0.615000 1.460000 0.805000 ;
      RECT 0.095000  1.880000 0.425000 2.635000 ;
      RECT 0.655000  1.580000 1.460000 1.750000 ;
      RECT 0.655000  1.750000 0.835000 2.465000 ;
      RECT 1.055000  0.085000 1.385000 0.445000 ;
      RECT 1.090000  1.935000 1.420000 2.635000 ;
      RECT 1.250000  0.805000 1.460000 1.020000 ;
      RECT 1.250000  1.020000 2.935000 1.355000 ;
      RECT 1.250000  1.355000 1.460000 1.580000 ;
      RECT 2.040000  0.085000 2.420000 0.445000 ;
      RECT 2.040000  1.935000 2.420000 2.635000 ;
      RECT 3.000000  0.085000 3.380000 0.445000 ;
      RECT 3.000000  1.935000 3.380000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and2_4
