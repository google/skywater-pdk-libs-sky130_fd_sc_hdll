* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_12 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_27_47# A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_117_297# a_973_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_597_297# A0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# A1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_973_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_119_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_973_297# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_27_47# A0 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_117_297# A1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_597_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_119_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# A1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_1163_47# a_973_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# A0 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR a_973_297# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_27_47# A0 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_117_297# a_973_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_27_47# A0 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_119_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 VPWR S a_973_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 a_27_47# A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VGND a_973_297# a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_1163_47# a_973_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_597_297# A0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VGND S a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 a_1163_47# A0 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_119_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 VPWR S a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X45 VGND a_973_297# a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 a_117_297# A1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 VGND S a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 a_1163_47# A0 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X52 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X53 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 VPWR a_973_297# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 VGND S a_973_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_597_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
