* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
X0 a_80_21# A2 a_1202_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VPWR B1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_1202_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_524_47# B1 a_607_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_80_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_1010_297# A2 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 X a_80_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_80_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_80_21# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR A1 a_1010_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VGND A1 a_524_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_80_21# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VPWR C1 a_80_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_607_47# C1 a_80_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_524_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_818_47# B1 a_524_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND A2 a_524_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND a_80_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_80_21# C1 a_818_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_524_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
