* File: sky130_fd_sc_hdll__and4bb_1.spice
* Created: Wed Sep  2 08:23:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4bb_1.pex.spice"
.subckt sky130_fd_sc_hdll__and4bb_1  VNB VPB A_N B_N C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B_N	B_N
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_A_N_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.1344 PD=0.8 PS=1.48 NRD=12.852 NRS=15.708 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_225_413#_M1007_d N_B_N_M1007_g N_VGND_M1008_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0798 PD=1.36 PS=0.8 NRD=0 NRS=15.708 M=1 R=2.8
+ SA=75000.8 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_425_93# N_A_27_47#_M1000_g N_A_339_93#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1003 A_511_93# N_A_225_413#_M1003_g A_425_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0588 PD=0.79 PS=0.7 NRD=37.14 NRS=24.276 M=1 R=2.8 SA=75000.6
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1001 A_615_93# N_C_M1001_g A_511_93# VNB NSHORT L=0.15 W=0.42 AD=0.0945
+ AS=0.0777 PD=0.87 PS=0.79 NRD=48.564 NRS=37.14 M=1 R=2.8 SA=75001.2 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_D_M1009_g A_615_93# VNB NSHORT L=0.15 W=0.42
+ AD=0.0889065 AS=0.0945 PD=0.804673 PS=0.87 NRD=44.76 NRS=48.564 M=1 R=2.8
+ SA=75001.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1013 N_X_M1013_d N_A_339_93#_M1013_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.137593 PD=1.82 PS=1.24533 NRD=0 NRS=2.76 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_A_N_M1011_g N_A_27_47#_M1011_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.063 AS=0.1386 PD=0.72 PS=1.5 NRD=2.3443 NRS=30.4759 M=1 R=2.33333
+ SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1004 N_A_225_413#_M1004_d N_B_N_M1004_g N_VPWR_M1011_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.063 PD=1.38 PS=0.72 NRD=2.3443 NRS=7.0329 M=1 R=2.33333
+ SA=90000.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1012 N_A_339_93#_M1012_d N_A_27_47#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.063 AS=0.1134 PD=0.72 PS=1.38 NRD=7.0329 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_225_413#_M1005_g N_A_339_93#_M1012_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0714 AS=0.063 PD=0.76 PS=0.72 NRD=14.0658 NRS=2.3443 M=1
+ R=2.33333 SA=90000.7 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1002 N_A_339_93#_M1002_d N_C_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0777 AS=0.0714 PD=0.79 PS=0.76 NRD=18.7544 NRS=14.0658 M=1 R=2.33333
+ SA=90001.2 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_D_M1006_g N_A_339_93#_M1002_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0874606 AS=0.0777 PD=0.795634 PS=0.79 NRD=28.1316 NRS=23.443 M=1
+ R=2.33333 SA=90001.7 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1010 N_X_M1010_d N_A_339_93#_M1010_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.208239 PD=2.54 PS=1.89437 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hdll__and4bb_1.pxi.spice"
*
.ends
*
*
