* NGSPICE file created from sky130_fd_sc_hdll__a31o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
M1000 a_27_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.47e+12p pd=1.294e+07u as=1.76e+12p ps=1.552e+07u
M1001 a_213_47# A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.08e+11p ps=1.94e+06u
M1002 a_27_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 X a_297_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=0p ps=0u
M1004 VGND a_297_47# X VNB nshort w=650000u l=150000u
+  ad=1.404e+12p pd=1.082e+07u as=4.16e+11p ps=3.88e+06u
M1005 a_297_47# A1 a_213_47# VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1006 VPWR a_297_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A3 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_297_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_27_297# B1 a_297_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1010 VGND a_297_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR A2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND B1 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_297_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_495_47# A2 a_401_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u
M1015 a_27_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_119_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_401_47# A1 a_297_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_297_47# B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A3 a_495_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_297_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_297_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR A1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_297_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

