* File: sky130_fd_sc_hdll__a21o_1.pxi.spice
* Created: Wed Sep  2 08:17:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21O_1%A_81_21# N_A_81_21#_M1001_d N_A_81_21#_M1005_s
+ N_A_81_21#_c_43_n N_A_81_21#_M1000_g N_A_81_21#_c_46_n N_A_81_21#_M1003_g
+ N_A_81_21#_c_44_n N_A_81_21#_c_52_p N_A_81_21#_c_84_p N_A_81_21#_c_48_n
+ N_A_81_21#_c_49_n N_A_81_21#_c_57_p N_A_81_21#_c_45_n
+ PM_SKY130_FD_SC_HDLL__A21O_1%A_81_21#
x_PM_SKY130_FD_SC_HDLL__A21O_1%B1 N_B1_c_99_n N_B1_M1005_g N_B1_c_100_n
+ N_B1_M1001_g B1 N_B1_c_101_n B1 PM_SKY130_FD_SC_HDLL__A21O_1%B1
x_PM_SKY130_FD_SC_HDLL__A21O_1%A1 N_A1_c_128_n N_A1_M1002_g N_A1_c_129_n
+ N_A1_M1007_g A1 A1 A1 A1 PM_SKY130_FD_SC_HDLL__A21O_1%A1
x_PM_SKY130_FD_SC_HDLL__A21O_1%A2 N_A2_c_166_n N_A2_M1004_g N_A2_c_167_n
+ N_A2_M1006_g A2 A2 PM_SKY130_FD_SC_HDLL__A21O_1%A2
x_PM_SKY130_FD_SC_HDLL__A21O_1%X N_X_M1000_s N_X_M1003_s X X X X X X
+ PM_SKY130_FD_SC_HDLL__A21O_1%X
x_PM_SKY130_FD_SC_HDLL__A21O_1%VPWR N_VPWR_M1003_d N_VPWR_M1002_d N_VPWR_c_200_n
+ N_VPWR_c_201_n VPWR N_VPWR_c_202_n N_VPWR_c_203_n N_VPWR_c_204_n
+ N_VPWR_c_199_n N_VPWR_c_206_n N_VPWR_c_207_n PM_SKY130_FD_SC_HDLL__A21O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A21O_1%A_317_297# N_A_317_297#_M1005_d
+ N_A_317_297#_M1006_d N_A_317_297#_c_244_n N_A_317_297#_c_241_n
+ N_A_317_297#_c_243_n N_A_317_297#_c_242_n
+ PM_SKY130_FD_SC_HDLL__A21O_1%A_317_297#
x_PM_SKY130_FD_SC_HDLL__A21O_1%VGND N_VGND_M1000_d N_VGND_M1004_d N_VGND_c_260_n
+ N_VGND_c_261_n N_VGND_c_262_n VGND N_VGND_c_263_n N_VGND_c_264_n
+ N_VGND_c_265_n N_VGND_c_266_n PM_SKY130_FD_SC_HDLL__A21O_1%VGND
cc_1 VNB N_A_81_21#_c_43_n 0.0231009f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_2 VNB N_A_81_21#_c_44_n 0.0039428f $X=-0.19 $Y=-0.24 $X2=0.745 $Y2=1.16
cc_3 VNB N_A_81_21#_c_45_n 0.0380336f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_4 VNB N_B1_c_99_n 0.0218982f $X=-0.19 $Y=-0.24 $X2=1.595 $Y2=0.235
cc_5 VNB N_B1_c_100_n 0.0208706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_B1_c_101_n 0.00675582f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.985
cc_7 VNB N_A1_c_128_n 0.022529f $X=-0.19 $Y=-0.24 $X2=1.595 $Y2=0.235
cc_8 VNB N_A1_c_129_n 0.0165174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A1 0.00158898f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_10 VNB A1 0.0042505f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.56
cc_11 VNB N_A2_c_166_n 0.0222885f $X=-0.19 $Y=-0.24 $X2=1.595 $Y2=0.235
cc_12 VNB N_A2_c_167_n 0.040215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB X 0.0456623f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=0.995
cc_14 VNB N_VPWR_c_199_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_260_n 0.0290013f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.985
cc_16 VNB N_VGND_c_261_n 0.0341424f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.505
cc_17 VNB N_VGND_c_262_n 0.00557808f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.16
cc_18 VNB N_VGND_c_263_n 0.0134401f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.55
cc_19 VNB N_VGND_c_264_n 0.191361f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.615
cc_20 VNB N_VGND_c_265_n 0.0203949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_266_n 0.0204472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A_81_21#_c_46_n 0.0213798f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_23 VPB N_A_81_21#_c_44_n 0.00273801f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.16
cc_24 VPB N_A_81_21#_c_48_n 0.0126267f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=1.725
cc_25 VPB N_A_81_21#_c_49_n 0.00794157f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.81
cc_26 VPB N_A_81_21#_c_45_n 0.0166338f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.202
cc_27 VPB N_B1_c_99_n 0.0310193f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=0.235
cc_28 VPB N_B1_c_101_n 0.00274273f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_29 VPB N_A1_c_128_n 0.0246804f $X=-0.19 $Y=1.305 $X2=1.595 $Y2=0.235
cc_30 VPB A1 0.00179665f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_31 VPB N_A2_c_167_n 0.0350041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB X 0.0465488f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.995
cc_33 VPB N_VPWR_c_200_n 0.0088519f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=0.56
cc_34 VPB N_VPWR_c_201_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.715 $Y2=0.835
cc_35 VPB N_VPWR_c_202_n 0.0154228f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.16
cc_36 VPB N_VPWR_c_203_n 0.0289996f $X=-0.19 $Y=1.305 $X2=1.26 $Y2=1.81
cc_37 VPB N_VPWR_c_204_n 0.0252876f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=1.615
cc_38 VPB N_VPWR_c_199_n 0.0628982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_206_n 0.0059962f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.202
cc_40 VPB N_VPWR_c_207_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_317_297#_c_241_n 0.0117588f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.985
cc_42 VPB N_A_317_297#_c_242_n 0.0269742f $X=-0.19 $Y=1.305 $X2=0.715 $Y2=1.16
cc_43 N_A_81_21#_c_44_n N_B1_c_99_n 0.00587993f $X=0.745 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_44 N_A_81_21#_c_52_p N_B1_c_99_n 0.00312161f $X=1.515 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_45 N_A_81_21#_c_48_n N_B1_c_99_n 0.00119195f $X=1.23 $Y=1.725 $X2=-0.19
+ $Y2=-0.24
cc_46 N_A_81_21#_c_45_n N_B1_c_99_n 0.00824467f $X=0.505 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_47 N_A_81_21#_c_44_n N_B1_c_100_n 0.00394282f $X=0.745 $Y=1.16 $X2=0 $Y2=0
cc_48 N_A_81_21#_c_52_p N_B1_c_100_n 0.0121994f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_49 N_A_81_21#_c_57_p N_B1_c_100_n 0.0129081f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_50 N_A_81_21#_c_44_n N_B1_c_101_n 0.0257617f $X=0.745 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_81_21#_c_52_p N_B1_c_101_n 0.0373758f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_52 N_A_81_21#_c_48_n N_B1_c_101_n 0.0219963f $X=1.23 $Y=1.725 $X2=0 $Y2=0
cc_53 N_A_81_21#_c_45_n N_B1_c_101_n 0.00130368f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_54 N_A_81_21#_c_52_p N_A1_c_129_n 0.00155471f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_55 N_A_81_21#_c_57_p N_A1_c_129_n 0.00464411f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_56 N_A_81_21#_c_52_p A1 0.01611f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_57 N_A_81_21#_c_57_p A1 0.0194705f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_58 N_A_81_21#_c_52_p A1 0.00283874f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_59 N_A_81_21#_c_43_n X 0.0183412f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A_81_21#_c_46_n X 0.0118809f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_81_21#_c_44_n X 0.0459364f $X=0.745 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_81_21#_c_48_n X 0.016194f $X=1.23 $Y=1.725 $X2=0 $Y2=0
cc_63 N_A_81_21#_c_44_n N_VPWR_M1003_d 6.29821e-19 $X=0.745 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_81_21#_c_48_n N_VPWR_M1003_d 0.00389372f $X=1.23 $Y=1.725 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_81_21#_c_46_n N_VPWR_c_200_n 0.0182157f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_81_21#_c_48_n N_VPWR_c_200_n 0.0245714f $X=1.23 $Y=1.725 $X2=0 $Y2=0
cc_67 N_A_81_21#_c_49_n N_VPWR_c_200_n 0.0438938f $X=1.26 $Y=1.81 $X2=0 $Y2=0
cc_68 N_A_81_21#_c_46_n N_VPWR_c_202_n 0.00427505f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_81_21#_c_49_n N_VPWR_c_203_n 0.017241f $X=1.26 $Y=1.81 $X2=0 $Y2=0
cc_70 N_A_81_21#_M1005_s N_VPWR_c_199_n 0.0036094f $X=1.135 $Y=1.485 $X2=0 $Y2=0
cc_71 N_A_81_21#_c_46_n N_VPWR_c_199_n 0.00836369f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_81_21#_c_49_n N_VPWR_c_199_n 0.0102724f $X=1.26 $Y=1.81 $X2=0 $Y2=0
cc_73 N_A_81_21#_c_52_p N_A_317_297#_c_243_n 0.0041884f $X=1.515 $Y=0.735 $X2=0
+ $Y2=0
cc_74 N_A_81_21#_c_44_n N_VGND_M1000_d 8.64196e-19 $X=0.745 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_81_21#_c_52_p N_VGND_M1000_d 0.0165754f $X=1.515 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_81_21#_c_84_p N_VGND_M1000_d 0.00486568f $X=0.885 $Y=0.735 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_81_21#_c_52_p N_VGND_c_261_n 0.00263609f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_78 N_A_81_21#_c_57_p N_VGND_c_261_n 0.0174683f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_79 N_A_81_21#_M1001_d N_VGND_c_264_n 0.00671976f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_80 N_A_81_21#_c_43_n N_VGND_c_264_n 0.0128603f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_81_21#_c_52_p N_VGND_c_264_n 0.00685568f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_82 N_A_81_21#_c_84_p N_VGND_c_264_n 0.00470238f $X=0.885 $Y=0.735 $X2=0 $Y2=0
cc_83 N_A_81_21#_c_57_p N_VGND_c_264_n 0.0110045f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_84 N_A_81_21#_c_43_n N_VGND_c_265_n 0.00574689f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_81_21#_c_84_p N_VGND_c_265_n 0.0017532f $X=0.885 $Y=0.735 $X2=0 $Y2=0
cc_86 N_A_81_21#_c_43_n N_VGND_c_266_n 0.010052f $X=0.48 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_81_21#_c_52_p N_VGND_c_266_n 0.0327754f $X=1.515 $Y=0.735 $X2=0 $Y2=0
cc_88 N_A_81_21#_c_84_p N_VGND_c_266_n 0.0175141f $X=0.885 $Y=0.735 $X2=0 $Y2=0
cc_89 N_A_81_21#_c_57_p N_VGND_c_266_n 0.0148149f $X=1.665 $Y=0.635 $X2=0 $Y2=0
cc_90 N_A_81_21#_c_45_n N_VGND_c_266_n 7.85384e-19 $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_91 N_B1_c_99_n N_A1_c_128_n 0.0436964f $X=1.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_92 N_B1_c_101_n N_A1_c_128_n 0.00103342f $X=1.445 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_93 N_B1_c_100_n N_A1_c_129_n 0.0234635f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B1_c_100_n A1 0.00114693f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B1_c_99_n A1 0.00102824f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B1_c_101_n A1 0.0274393f $X=1.445 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B1_c_99_n N_VPWR_c_200_n 0.00376087f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B1_c_99_n N_VPWR_c_201_n 0.00131852f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B1_c_99_n N_VPWR_c_203_n 0.00702461f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B1_c_99_n N_VPWR_c_199_n 0.0141576f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B1_c_100_n N_VGND_c_261_n 0.00391752f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_102 N_B1_c_100_n N_VGND_c_264_n 0.00710481f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_103 N_B1_c_100_n N_VGND_c_266_n 0.00962689f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A1_c_129_n N_A2_c_166_n 0.0281841f $X=2.005 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_105 A1 N_A2_c_166_n 0.00789404f $X=2.015 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_106 N_A1_c_128_n N_A2_c_167_n 0.0513214f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_107 A1 N_A2_c_167_n 0.00230712f $X=2.015 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A1_c_128_n A2 3.11313e-19 $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_109 A1 A2 0.00129754f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_110 A1 A2 0.0222472f $X=2.015 $Y=1.105 $X2=0 $Y2=0
cc_111 N_A1_c_128_n N_VPWR_c_201_n 0.0150175f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A1_c_128_n N_VPWR_c_203_n 0.00447018f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A1_c_128_n N_VPWR_c_199_n 0.00777771f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A1_c_128_n N_A_317_297#_c_244_n 0.00563789f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A1_c_128_n N_A_317_297#_c_241_n 0.0182788f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_116 A1 N_A_317_297#_c_241_n 0.0240264f $X=2.015 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A1_c_128_n N_A_317_297#_c_243_n 3.47712e-19 $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_118 A1 N_A_317_297#_c_243_n 0.00366311f $X=2.015 $Y=1.105 $X2=0 $Y2=0
cc_119 A1 N_VGND_c_260_n 0.0195781f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_120 N_A1_c_129_n N_VGND_c_261_n 0.00457622f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_121 A1 N_VGND_c_261_n 0.00774909f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_122 N_A1_c_129_n N_VGND_c_264_n 0.00763114f $X=2.005 $Y=0.995 $X2=0 $Y2=0
cc_123 A1 N_VGND_c_264_n 0.00774184f $X=2.015 $Y=0.425 $X2=0 $Y2=0
cc_124 A1 A_416_47# 0.00681055f $X=2.015 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_125 N_A2_c_167_n N_VPWR_c_201_n 0.0123594f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_167_n N_VPWR_c_204_n 0.00642146f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A2_c_167_n N_VPWR_c_199_n 0.0119091f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_167_n N_A_317_297#_c_241_n 0.0247047f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_129 A2 N_A_317_297#_c_241_n 0.016027f $X=2.545 $Y=1.19 $X2=0 $Y2=0
cc_130 N_A2_c_166_n N_VGND_c_260_n 0.0136567f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A2_c_167_n N_VGND_c_260_n 0.00414539f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_132 A2 N_VGND_c_260_n 0.00663626f $X=2.545 $Y=1.19 $X2=0 $Y2=0
cc_133 N_A2_c_166_n N_VGND_c_261_n 0.00585385f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_166_n N_VGND_c_264_n 0.0119735f $X=2.435 $Y=0.995 $X2=0 $Y2=0
cc_135 X N_VPWR_c_200_n 0.0424564f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_136 X N_VPWR_c_202_n 0.017115f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_137 N_X_M1003_s N_VPWR_c_199_n 0.00430346f $X=0.145 $Y=1.485 $X2=0 $Y2=0
cc_138 X N_VPWR_c_199_n 0.00988906f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_139 N_X_M1000_s N_VGND_c_264_n 0.00387432f $X=0.145 $Y=0.235 $X2=0 $Y2=0
cc_140 X N_VGND_c_264_n 0.00988906f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_141 X N_VGND_c_265_n 0.0169196f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_142 N_VPWR_c_199_n N_A_317_297#_M1005_d 0.00512507f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_143 N_VPWR_c_199_n N_A_317_297#_M1006_d 0.004171f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_144 N_VPWR_c_201_n N_A_317_297#_c_244_n 0.0387104f $X=2.22 $Y=2.02 $X2=0
+ $Y2=0
cc_145 N_VPWR_c_203_n N_A_317_297#_c_244_n 0.0135675f $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_146 N_VPWR_c_199_n N_A_317_297#_c_244_n 0.00873917f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_147 N_VPWR_M1002_d N_A_317_297#_c_241_n 0.00690516f $X=2.07 $Y=1.485 $X2=0
+ $Y2=0
cc_148 N_VPWR_c_201_n N_A_317_297#_c_241_n 0.0205755f $X=2.22 $Y=2.02 $X2=0
+ $Y2=0
cc_149 N_VPWR_c_204_n N_A_317_297#_c_242_n 0.0170688f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_150 N_VPWR_c_199_n N_A_317_297#_c_242_n 0.00988367f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_151 N_VGND_c_264_n A_416_47# 0.0073888f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
