* File: sky130_fd_sc_hdll__buf_2.pex.spice
* Created: Thu Aug 27 19:00:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_2%A 2 3 5 8 10 17
r35 16 17 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r36 13 16 39.3438 $w=3.3e-07 $l=2.25e-07 $layer=POLY_cond $X=0.27 $Y=1.16
+ $X2=0.495 $Y2=1.16
r37 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r38 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r39 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r40 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.73
+ $X2=0.495 $Y2=2.125
r41 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.63 $X2=0.495
+ $Y2=1.73
r42 1 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r43 1 2 101.131 $w=2e-07 $l=3.05e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_2%A_27_47# 1 2 7 9 10 12 13 14 15 17 18 20 21
+ 24 28 30 31 32 33 37 39 41
r81 44 45 3.14621 $w=3.83e-07 $l=2.5e-08 $layer=POLY_cond $X=0.995 $Y=1.202
+ $X2=1.02 $Y2=1.202
r82 40 44 6.92167 $w=3.83e-07 $l=5.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.995 $Y2=1.202
r83 39 42 8.48463 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=0.875 $Y2=1.325
r84 39 41 7.28133 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=0.875 $Y=1.16
+ $X2=0.875 $Y2=0.995
r85 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r86 37 42 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.81 $Y=1.535
+ $X2=0.81 $Y2=1.325
r87 34 41 10.1844 $w=2.13e-07 $l=1.9e-07 $layer=LI1_cond $X=0.832 $Y=0.805
+ $X2=0.832 $Y2=0.995
r88 32 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.725 $Y=1.62
+ $X2=0.81 $Y2=1.535
r89 32 33 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.725 $Y=1.62
+ $X2=0.345 $Y2=1.62
r90 30 34 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=0.725 $Y=0.72
+ $X2=0.832 $Y2=0.805
r91 30 31 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.725 $Y=0.72
+ $X2=0.345 $Y2=0.72
r92 26 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=1.705
+ $X2=0.345 $Y2=1.62
r93 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=1.705
+ $X2=0.26 $Y2=1.96
r94 22 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r95 22 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.445
r96 18 21 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.62 $Y=0.995
+ $X2=1.595 $Y2=1.202
r97 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.62 $Y=0.995
+ $X2=1.62 $Y2=0.56
r98 15 21 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.595 $Y=1.41
+ $X2=1.595 $Y2=1.202
r99 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.595 $Y=1.41
+ $X2=1.595 $Y2=1.985
r100 14 45 13.6412 $w=3.83e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.12 $Y=1.16
+ $X2=1.02 $Y2=1.202
r101 13 21 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.595 $Y2=1.202
r102 13 14 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=1.495 $Y=1.16
+ $X2=1.12 $Y2=1.16
r103 10 45 20.4303 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.202
r104 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r105 7 44 24.8035 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=1.202
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=0.56
r107 2 28 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.805 $X2=0.26 $Y2=1.96
r108 1 24 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_2%VPWR 1 2 9 11 13 17 19 21 27 33 37
r29 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r33 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 28 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=0.765 $Y2=2.72
r35 28 30 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.93 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 27 36 4.02327 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=2.082 $Y2=2.72
r37 27 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 21 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.765 $Y2=2.72
r39 19 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r40 17 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=0.6
+ $Y2=2.72
r41 17 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 13 16 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=1.995 $Y=1.66
+ $X2=1.995 $Y2=2.34
r43 11 36 3.18895 $w=2.6e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.995 $Y=2.635
+ $X2=2.082 $Y2=2.72
r44 11 16 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=1.995 $Y=2.635
+ $X2=1.995 $Y2=2.34
r45 7 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=2.72
r46 7 9 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.765 $Y=2.635
+ $X2=0.765 $Y2=1.96
r47 2 16 400 $w=1.7e-07 $l=9.7857e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.485 $X2=1.95 $Y2=2.34
r48 2 13 400 $w=1.7e-07 $l=3.41467e-07 $layer=licon1_PDIFF $count=1 $X=1.685
+ $Y=1.485 $X2=1.95 $Y2=1.66
r49 1 9 300 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.805 $X2=0.765 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_2%X 1 2 7 8 9 10 11 12
r22 11 12 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.482 $Y=1.87
+ $X2=1.482 $Y2=2.21
r23 11 31 1.4914 $w=4.23e-07 $l=5.5e-08 $layer=LI1_cond $X=1.482 $Y=1.87
+ $X2=1.482 $Y2=1.815
r24 10 31 7.72815 $w=4.23e-07 $l=2.85e-07 $layer=LI1_cond $X=1.482 $Y=1.53
+ $X2=1.482 $Y2=1.815
r25 9 10 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.482 $Y=1.19
+ $X2=1.482 $Y2=1.53
r26 8 9 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=1.482 $Y=0.85
+ $X2=1.482 $Y2=1.19
r27 8 23 8.67722 $w=4.23e-07 $l=3.2e-07 $layer=LI1_cond $X=1.482 $Y=0.85
+ $X2=1.482 $Y2=0.53
r28 7 23 0.542326 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=1.482 $Y=0.51
+ $X2=1.482 $Y2=0.53
r29 2 31 300 $w=1.7e-07 $l=4.35603e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.485 $X2=1.355 $Y2=1.815
r30 1 23 182 $w=1.7e-07 $l=4.13642e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.355 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_2%VGND 1 2 9 11 13 15 17 19 24 26 30
r32 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r34 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.61 $Y=0 $X2=0.775
+ $Y2=0
r35 23 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r36 23 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r37 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r38 20 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=0.775
+ $Y2=0
r39 20 22 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.94 $Y=0 $X2=1.61
+ $Y2=0
r40 19 29 4.02327 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=2.082
+ $Y2=0
r41 19 22 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.865 $Y=0 $X2=1.61
+ $Y2=0
r42 17 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 15 24 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.61
+ $Y2=0
r44 11 29 3.18895 $w=2.6e-07 $l=1.22327e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=2.082 $Y2=0
r45 11 13 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.995 $Y=0.085
+ $X2=1.995 $Y2=0.4
r46 7 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.085
+ $X2=0.775 $Y2=0
r47 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.775 $Y=0.085
+ $X2=0.775 $Y2=0.38
r48 2 13 91 $w=1.7e-07 $l=3.27261e-07 $layer=licon1_NDIFF $count=2 $X=1.695
+ $Y=0.235 $X2=1.95 $Y2=0.4
r49 1 9 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.775 $Y2=0.38
.ends

