* File: sky130_fd_sc_hdll__or4bb_2.spice
* Created: Wed Sep  2 08:50:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4bb_2.pex.spice"
.subckt sky130_fd_sc_hdll__or4bb_2  VNB VPB C_N D_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_C_N_M1001_g N_A_27_410#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1302 PD=0.715 PS=1.46 NRD=5.712 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_216_93#_M1003_d N_D_N_M1003_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.06195 PD=1.46 PS=0.715 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_A_336_413#_M1002_d N_A_216_93#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.07035 AS=0.1386 PD=0.755 PS=1.5 NRD=0 NRS=18.564 M=1 R=2.8
+ SA=75000.3 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1015 N_VGND_M1015_d N_A_27_410#_M1015_g N_A_336_413#_M1002_d VNB NSHORT L=0.15
+ W=0.42 AD=0.06405 AS=0.07035 PD=0.725 PS=0.755 NRD=0 NRS=17.136 M=1 R=2.8
+ SA=75000.7 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1012 N_A_336_413#_M1012_d N_B_M1012_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07035 AS=0.06405 PD=0.755 PS=0.725 NRD=2.856 NRS=8.568 M=1 R=2.8
+ SA=75001.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_A_336_413#_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.07035 PD=0.816449 PS=0.755 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1007_d N_A_336_413#_M1013_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.143516 AS=0.104 PD=1.26355 PS=0.97 NRD=11.988 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1014_d N_A_336_413#_M1014_g N_X_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.104 PD=1.87 PS=0.97 NRD=3.684 NRS=8.304 M=1 R=4.33333 SA=75002
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_C_N_M1010_g N_A_27_410#_M1010_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.126812 AS=0.1134 PD=1.34 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1011 N_A_216_93#_M1011_d N_D_N_M1011_g N_VPWR_M1010_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1218 AS=0.126812 PD=1.42 PS=1.34 NRD=2.3443 NRS=115.816 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1008 A_426_413# N_A_216_93#_M1008_g N_A_336_413#_M1008_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1257 AS=0.1134 PD=1.35 PS=1.38 NRD=114.575 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1006 A_532_297# N_A_27_410#_M1006_g A_426_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.1257 PD=0.65 PS=1.35 NRD=28.1316 NRS=114.575 M=1 R=2.33333
+ SA=90000.2 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1009 A_614_297# N_B_M1009_g A_532_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.06405
+ AS=0.0483 PD=0.725 PS=0.65 NRD=45.7237 NRS=28.1316 M=1 R=2.33333 SA=90000.6
+ SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_614_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.06405 PD=0.804507 PS=0.725 NRD=76.83 NRS=45.7237 M=1
+ R=2.33333 SA=90001.1 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1000_d N_A_336_413#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.218803 AS=0.145 PD=1.91549 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90000.8 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_336_413#_M1005_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.145 PD=2.59 PS=1.29 NRD=5.91 NRS=0.9653 M=1 R=5.55556 SA=90001.3
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX17_noxref noxref_16 D_N D_N PROBETYPE=1
pX18_noxref noxref_17 A A PROBETYPE=1
pX19_noxref noxref_18 B B PROBETYPE=1
c_95 VPB 0 1.99056e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or4bb_2.pxi.spice"
*
.ends
*
*
