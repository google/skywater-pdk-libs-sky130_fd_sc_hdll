# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand4bb_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  10.58000 BY  2.720000 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 0.995000 0.330000 1.615000 ;
    END
  END A_N
  PIN B_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.585000 0.995000 1.025000 1.615000 ;
    END
  END B_N
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.045000 1.075000 7.985000 1.275000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.395000 1.075000 10.340000 1.275000 ;
    END
  END D
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.736000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.355000 0.655000 4.015000 0.905000 ;
        RECT 2.355000 1.445000 9.865000 1.665000 ;
        RECT 2.355000 1.665000 2.655000 2.465000 ;
        RECT 3.295000 1.665000 3.675000 2.465000 ;
        RECT 3.665000 0.905000 4.015000 1.445000 ;
        RECT 4.235000 1.665000 4.615000 2.465000 ;
        RECT 5.175000 1.665000 5.555000 2.465000 ;
        RECT 6.665000 1.665000 7.045000 2.465000 ;
        RECT 7.605000 1.665000 7.985000 2.465000 ;
        RECT 8.545000 1.665000 8.925000 2.465000 ;
        RECT 9.485000 1.665000 9.865000 2.465000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.085000  0.255000  0.345000 0.635000 ;
      RECT  0.085000  0.635000  1.505000 0.805000 ;
      RECT  0.085000  1.785000  1.505000 1.980000 ;
      RECT  0.085000  1.980000  0.370000 2.440000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.540000  2.195000  0.815000 2.635000 ;
      RECT  0.985000  2.150000  1.845000 2.465000 ;
      RECT  1.115000  0.255000  1.845000 0.465000 ;
      RECT  1.195000  0.805000  1.505000 1.785000 ;
      RECT  1.675000  0.465000  1.845000 1.075000 ;
      RECT  1.675000  1.075000  2.025000 1.305000 ;
      RECT  1.675000  1.305000  1.845000 2.150000 ;
      RECT  2.015000  0.255000  6.025000 0.485000 ;
      RECT  2.015000  0.485000  2.185000 0.905000 ;
      RECT  2.015000  1.495000  2.185000 2.635000 ;
      RECT  2.355000  1.075000  3.200000 1.245000 ;
      RECT  2.825000  1.835000  3.125000 2.635000 ;
      RECT  3.895000  1.835000  4.065000 2.635000 ;
      RECT  4.185000  1.075000  5.555000 1.275000 ;
      RECT  4.235000  0.655000  8.010000 0.905000 ;
      RECT  4.835000  1.835000  5.005000 2.635000 ;
      RECT  5.825000  1.835000  6.465000 2.635000 ;
      RECT  6.265000  0.255000  8.375000 0.485000 ;
      RECT  7.265000  1.835000  7.435000 2.635000 ;
      RECT  8.205000  0.485000  8.375000 0.655000 ;
      RECT  8.205000  0.655000 10.285000 0.825000 ;
      RECT  8.205000  1.835000  8.375000 2.635000 ;
      RECT  8.595000  0.085000  8.925000 0.485000 ;
      RECT  9.145000  1.835000  9.315000 2.635000 ;
      RECT  9.535000  0.085000  9.865000 0.485000 ;
      RECT 10.085000  1.445000 10.360000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.795000  1.105000  1.965000 1.275000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.330000  1.105000  4.500000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
    LAYER met1 ;
      RECT 1.735000 1.075000 2.025000 1.120000 ;
      RECT 1.735000 1.120000 4.575000 1.260000 ;
      RECT 1.735000 1.260000 2.025000 1.305000 ;
      RECT 4.235000 1.075000 4.575000 1.120000 ;
      RECT 4.235000 1.260000 4.575000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4bb_4
