* File: sky130_fd_sc_hdll__and2_4.pex.spice
* Created: Thu Aug 27 18:56:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2_4%A 1 3 4 6 7 11
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.16 $X2=0.35 $Y2=1.16
r24 7 11 13.755 $w=3.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.28 $Y=1.53 $X2=0.28
+ $Y2=1.16
r25 4 10 38.7502 $w=3.47e-07 $l=2.1609e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.407 $Y2=1.16
r26 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.56
r27 1 10 45.8462 $w=3.47e-07 $l=2.92831e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.407 $Y2=1.16
r28 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_4%B 1 3 4 6 7 11 13
c33 4 0 1.95678e-19 $X=0.98 $Y=1.41
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.16 $X2=0.945 $Y2=1.16
r35 7 11 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.74 $Y=1.16
+ $X2=0.945 $Y2=1.16
r36 7 13 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.74 $Y=1.16 $X2=0.69
+ $Y2=1.16
r37 4 10 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.97 $Y2=1.16
r38 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41 $X2=0.98
+ $Y2=1.985
r39 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.885 $Y=0.995
+ $X2=0.97 $Y2=1.16
r40 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.885 $Y=0.995
+ $X2=0.885 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_4%A_27_47# 1 2 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 35 39 41 42 44 46 52 57 66
c110 66 0 1.13405e-19 $X=2.975 $Y=1.202
c111 44 0 1.95678e-19 $X=1.355 $Y=1.02
r112 66 67 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.975 $Y=1.202
+ $X2=3 $Y2=1.202
r113 63 64 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.47 $Y=1.202
+ $X2=2.495 $Y2=1.202
r114 62 63 59.1132 $w=3.71e-07 $l=4.55e-07 $layer=POLY_cond $X=2.015 $Y=1.202
+ $X2=2.47 $Y2=1.202
r115 61 62 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r116 58 59 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.535 $Y2=1.202
r117 53 66 26.6334 $w=3.71e-07 $l=2.05e-07 $layer=POLY_cond $X=2.77 $Y=1.202
+ $X2=2.975 $Y2=1.202
r118 53 64 35.7278 $w=3.71e-07 $l=2.75e-07 $layer=POLY_cond $X=2.77 $Y=1.202
+ $X2=2.495 $Y2=1.202
r119 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.77
+ $Y=1.16 $X2=2.77 $Y2=1.16
r120 50 61 50.6685 $w=3.71e-07 $l=3.9e-07 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=1.99 $Y2=1.202
r121 50 59 8.44474 $w=3.71e-07 $l=6.5e-08 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=1.535 $Y2=1.202
r122 49 52 40.2495 $w=3.33e-07 $l=1.17e-06 $layer=LI1_cond $X=1.6 $Y=1.187
+ $X2=2.77 $Y2=1.187
r123 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r124 47 57 0.271299 $w=3.35e-07 $l=1.05e-07 $layer=LI1_cond $X=1.46 $Y=1.187
+ $X2=1.355 $Y2=1.187
r125 47 49 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=1.46 $Y=1.187
+ $X2=1.6 $Y2=1.187
r126 45 57 7.47207 $w=2.1e-07 $l=1.68e-07 $layer=LI1_cond $X=1.355 $Y=1.355
+ $X2=1.355 $Y2=1.187
r127 45 46 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=1.355 $Y=1.355
+ $X2=1.355 $Y2=1.58
r128 44 57 7.47207 $w=2.1e-07 $l=1.67e-07 $layer=LI1_cond $X=1.355 $Y=1.02
+ $X2=1.355 $Y2=1.187
r129 43 44 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.355 $Y2=1.02
r130 41 46 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.25 $Y=1.665
+ $X2=1.355 $Y2=1.58
r131 41 42 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.25 $Y=1.665
+ $X2=0.835 $Y2=1.665
r132 37 42 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.745 $Y=1.75
+ $X2=0.835 $Y2=1.665
r133 37 39 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.745 $Y=1.75
+ $X2=0.745 $Y2=1.96
r134 36 56 4.74669 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=0.71
+ $X2=0.26 $Y2=0.71
r135 35 43 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=1.25 $Y=0.71
+ $X2=1.355 $Y2=0.805
r136 35 36 48.1579 $w=1.88e-07 $l=8.25e-07 $layer=LI1_cond $X=1.25 $Y=0.71
+ $X2=0.425 $Y2=0.71
r137 31 56 2.73294 $w=3.3e-07 $l=9.5e-08 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.71
r138 31 33 8.20679 $w=3.28e-07 $l=2.35e-07 $layer=LI1_cond $X=0.26 $Y=0.615
+ $X2=0.26 $Y2=0.38
r139 28 67 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3 $Y=0.995 $X2=3
+ $Y2=1.202
r140 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3 $Y=0.995 $X2=3
+ $Y2=0.56
r141 25 66 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.202
r142 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.985
r143 22 64 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=1.202
r144 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=1.985
r145 19 63 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=1.202
r146 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.47 $Y=0.995
+ $X2=2.47 $Y2=0.56
r147 16 62 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.202
r148 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.015 $Y=1.41
+ $X2=2.015 $Y2=1.985
r149 13 61 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=1.202
r150 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=0.56
r151 10 59 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.202
r152 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.985
r153 7 58 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r154 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r155 2 39 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.96
r156 1 56 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
r157 1 33 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_4%VPWR 1 2 3 4 13 15 17 21 23 27 31 34 35 36
+ 43 44 50 53
r56 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r57 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r59 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r60 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 41 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 38 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.42 $Y=2.72 $X2=2.23
+ $Y2=2.72
r64 38 40 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.99 $Y2=2.72
r65 36 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 36 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 34 40 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3 $Y=2.72 $X2=2.99
+ $Y2=2.72
r68 34 35 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3 $Y=2.72 $X2=3.19
+ $Y2=2.72
r69 33 43 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.38 $Y=2.72 $X2=3.45
+ $Y2=2.72
r70 33 35 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.38 $Y=2.72 $X2=3.19
+ $Y2=2.72
r71 29 35 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.19 $Y=2.635
+ $X2=3.19 $Y2=2.72
r72 29 31 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=3.19 $Y=2.635
+ $X2=3.19 $Y2=2.02
r73 25 53 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=2.635
+ $X2=2.23 $Y2=2.72
r74 25 27 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=2.23 $Y=2.635
+ $X2=2.23 $Y2=2.02
r75 24 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.42 $Y=2.72
+ $X2=1.255 $Y2=2.72
r76 23 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.04 $Y=2.72 $X2=2.23
+ $Y2=2.72
r77 23 24 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.04 $Y=2.72
+ $X2=1.42 $Y2=2.72
r78 19 50 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=2.72
r79 19 21 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=1.255 $Y=2.635
+ $X2=1.255 $Y2=2.02
r80 18 47 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r81 17 50 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=1.255 $Y2=2.72
r82 17 18 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=0.425 $Y2=2.72
r83 13 47 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r84 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2
r85 4 31 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.215 $Y2=2.02
r86 3 27 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.105
+ $Y=1.485 $X2=2.255 $Y2=2.02
r87 2 21 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.255 $Y2=2.02
r88 1 15 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_4%X 1 2 3 4 15 17 19 20 23 27 29 31 36 38 40
+ 42 45 47
c61 29 0 1.13405e-19 $X=3.29 $Y=0.73
r62 45 47 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=3.43 $Y=0.845
+ $X2=3.43 $Y2=0.85
r63 42 45 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=3.43 $Y=0.73
+ $X2=3.43 $Y2=0.845
r64 42 47 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=3.43 $Y=0.89 $X2=3.43
+ $Y2=0.85
r65 41 42 26.5473 $w=2.78e-07 $l=6.45e-07 $layer=LI1_cond $X=3.43 $Y=1.535
+ $X2=3.43 $Y2=0.89
r66 34 36 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.775 $Y=0.68
+ $X2=1.87 $Y2=0.68
r67 32 40 4.43576 $w=2.27e-07 $l=9.5e-08 $layer=LI1_cond $X=2.83 $Y=1.65
+ $X2=2.735 $Y2=1.65
r68 31 41 6.90206 $w=2.3e-07 $l=1.88944e-07 $layer=LI1_cond $X=3.29 $Y=1.65
+ $X2=3.43 $Y2=1.535
r69 31 32 23.0489 $w=2.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.29 $Y=1.65
+ $X2=2.83 $Y2=1.65
r70 30 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.83 $Y=0.73
+ $X2=2.735 $Y2=0.73
r71 29 42 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=3.29 $Y=0.73 $X2=3.43
+ $Y2=0.73
r72 29 30 23.0489 $w=2.28e-07 $l=4.6e-07 $layer=LI1_cond $X=3.29 $Y=0.73
+ $X2=2.83 $Y2=0.73
r73 25 40 1.99853 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.735 $Y=1.765
+ $X2=2.735 $Y2=1.65
r74 25 27 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.735 $Y=1.765
+ $X2=2.735 $Y2=1.96
r75 21 38 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=2.735 $Y=0.615
+ $X2=2.735 $Y2=0.73
r76 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=2.735 $Y=0.615
+ $X2=2.735 $Y2=0.42
r77 19 40 4.43576 $w=2.27e-07 $l=9.64883e-08 $layer=LI1_cond $X=2.64 $Y=1.647
+ $X2=2.735 $Y2=1.65
r78 19 20 39.4392 $w=2.23e-07 $l=7.7e-07 $layer=LI1_cond $X=2.64 $Y=1.647
+ $X2=1.87 $Y2=1.647
r79 17 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=2.64 $Y=0.73
+ $X2=2.735 $Y2=0.73
r80 17 36 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=2.64 $Y=0.73
+ $X2=1.87 $Y2=0.73
r81 13 20 6.87974 $w=2.25e-07 $l=1.5331e-07 $layer=LI1_cond $X=1.775 $Y=1.76
+ $X2=1.87 $Y2=1.647
r82 13 15 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=1.775 $Y=1.76
+ $X2=1.775 $Y2=1.96
r83 4 40 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.485 $X2=2.735 $Y2=1.62
r84 4 27 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=2.585
+ $Y=1.485 $X2=2.735 $Y2=1.96
r85 3 15 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=1.485 $X2=1.775 $Y2=1.96
r86 2 38 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.235 $X2=2.735 $Y2=0.76
r87 2 23 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=2.545
+ $Y=0.235 $X2=2.735 $Y2=0.42
r88 1 34 182 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.775 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_4%VGND 1 2 3 12 14 16 17 23 25 35 36 39 43
r61 43 46 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.23 $Y=0 $X2=2.23
+ $Y2=0.36
r62 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r64 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r66 33 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r67 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r68 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r69 30 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.23
+ $Y2=0
r70 30 32 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.42 $Y=0 $X2=2.99
+ $Y2=0
r71 28 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r72 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r73 25 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r74 25 27 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.69
+ $Y2=0
r75 23 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.38 $Y=0 $X2=3.45
+ $Y2=0
r77 17 32 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=3 $Y=0 $X2=2.99 $Y2=0
r78 16 21 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.19
+ $Y2=0.36
r79 16 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3.38
+ $Y2=0
r80 16 17 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.19 $Y=0 $X2=3 $Y2=0
r81 15 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r82 14 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=2.23
+ $Y2=0
r83 14 15 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.04 $Y=0 $X2=1.385
+ $Y2=0
r84 10 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r85 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.36
r86 3 21 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.235 $X2=3.215 $Y2=0.36
r87 2 46 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.255 $Y2=0.36
r88 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=0.96
+ $Y=0.235 $X2=1.22 $Y2=0.36
.ends

