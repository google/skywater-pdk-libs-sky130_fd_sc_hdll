* File: sky130_fd_sc_hdll__o221a_1.pxi.spice
* Created: Thu Aug 27 19:20:17 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221A_1%C1 N_C1_c_65_n N_C1_M1011_g N_C1_c_62_n
+ N_C1_M1010_g C1 N_C1_c_64_n PM_SKY130_FD_SC_HDLL__O221A_1%C1
x_PM_SKY130_FD_SC_HDLL__O221A_1%B1 N_B1_c_91_n N_B1_M1003_g N_B1_c_92_n
+ N_B1_M1008_g B1 B1 PM_SKY130_FD_SC_HDLL__O221A_1%B1
x_PM_SKY130_FD_SC_HDLL__O221A_1%B2 N_B2_c_127_n N_B2_M1005_g N_B2_c_128_n
+ N_B2_M1000_g B2 B2 B2 PM_SKY130_FD_SC_HDLL__O221A_1%B2
x_PM_SKY130_FD_SC_HDLL__O221A_1%A2 N_A2_c_161_n N_A2_M1004_g N_A2_c_162_n
+ N_A2_M1007_g N_A2_c_163_n A2 A2 N_A2_c_165_n PM_SKY130_FD_SC_HDLL__O221A_1%A2
x_PM_SKY130_FD_SC_HDLL__O221A_1%A1 N_A1_c_199_n N_A1_M1001_g N_A1_c_200_n
+ N_A1_M1002_g A1 A1 PM_SKY130_FD_SC_HDLL__O221A_1%A1
x_PM_SKY130_FD_SC_HDLL__O221A_1%A_27_297# N_A_27_297#_M1010_s
+ N_A_27_297#_M1011_s N_A_27_297#_M1005_d N_A_27_297#_c_231_n
+ N_A_27_297#_M1006_g N_A_27_297#_c_232_n N_A_27_297#_M1009_g
+ N_A_27_297#_c_238_n N_A_27_297#_c_233_n N_A_27_297#_c_234_n
+ N_A_27_297#_c_261_n N_A_27_297#_c_249_n N_A_27_297#_c_250_n
+ N_A_27_297#_c_278_n N_A_27_297#_c_289_n N_A_27_297#_c_240_n
+ N_A_27_297#_c_241_n N_A_27_297#_c_235_n N_A_27_297#_c_243_n
+ N_A_27_297#_c_236_n N_A_27_297#_c_274_n N_A_27_297#_c_267_n
+ PM_SKY130_FD_SC_HDLL__O221A_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O221A_1%VPWR N_VPWR_M1011_d N_VPWR_M1001_d
+ N_VPWR_c_348_n N_VPWR_c_349_n VPWR N_VPWR_c_350_n N_VPWR_c_351_n
+ N_VPWR_c_352_n N_VPWR_c_347_n N_VPWR_c_354_n N_VPWR_c_355_n
+ PM_SKY130_FD_SC_HDLL__O221A_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O221A_1%X N_X_M1006_d N_X_M1009_d N_X_c_407_n X X
+ PM_SKY130_FD_SC_HDLL__O221A_1%X
x_PM_SKY130_FD_SC_HDLL__O221A_1%A_124_47# N_A_124_47#_M1010_d
+ N_A_124_47#_M1000_d N_A_124_47#_c_425_n
+ PM_SKY130_FD_SC_HDLL__O221A_1%A_124_47#
x_PM_SKY130_FD_SC_HDLL__O221A_1%A_230_47# N_A_230_47#_M1008_d
+ N_A_230_47#_M1007_d N_A_230_47#_c_443_n N_A_230_47#_c_453_n
+ N_A_230_47#_c_456_n PM_SKY130_FD_SC_HDLL__O221A_1%A_230_47#
x_PM_SKY130_FD_SC_HDLL__O221A_1%VGND N_VGND_M1007_s N_VGND_M1002_d
+ N_VGND_c_474_n N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ N_VGND_c_479_n VGND N_VGND_c_480_n N_VGND_c_481_n
+ PM_SKY130_FD_SC_HDLL__O221A_1%VGND
cc_1 VNB N_C1_c_62_n 0.0224786f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_2 VNB C1 0.0164091f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C1_c_64_n 0.0397886f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_4 VNB N_B1_c_91_n 0.0221664f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_5 VNB N_B1_c_92_n 0.0170614f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_6 VNB B1 0.00268992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B2_c_127_n 0.0246007f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_8 VNB N_B2_c_128_n 0.0222253f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_9 VNB B2 0.00467014f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_A2_c_161_n 0.0233486f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_11 VNB N_A2_c_162_n 0.0224885f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_12 VNB N_A2_c_163_n 0.00385613f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_13 VNB A2 0.00106613f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_14 VNB N_A2_c_165_n 0.00656239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_199_n 0.0251948f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_16 VNB N_A1_c_200_n 0.016947f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_17 VNB A1 0.00207995f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_A_27_297#_c_231_n 0.0196341f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_19 VNB N_A_27_297#_c_232_n 0.024368f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.202
cc_20 VNB N_A_27_297#_c_233_n 0.0154614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_297#_c_234_n 0.00289488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_297#_c_235_n 6.45819e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_297#_c_236_n 0.00771092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_347_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_407_n 0.028684f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_26 VNB X 0.0262028f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_27 VNB N_A_124_47#_c_425_n 0.00242915f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_28 VNB N_A_230_47#_c_443_n 0.0103861f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_29 VNB N_VGND_c_474_n 0.00860609f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_30 VNB N_VGND_c_475_n 0.00462888f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.202
cc_31 VNB N_VGND_c_476_n 0.0533489f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_477_n 0.00650718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_478_n 0.0177863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_479_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_480_n 0.0242908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_481_n 0.22706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_C1_c_65_n 0.0202619f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_38 VPB N_C1_c_64_n 0.0173392f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_39 VPB N_B1_c_91_n 0.0248124f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_40 VPB B1 9.0173e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B2_c_127_n 0.0288626f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_42 VPB B2 0.00141303f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_43 VPB N_A2_c_161_n 0.0279851f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_44 VPB A2 0.00434359f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_45 VPB N_A1_c_199_n 0.0254415f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_46 VPB N_A_27_297#_c_232_n 0.0301245f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.202
cc_47 VPB N_A_27_297#_c_238_n 0.0290449f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_27_297#_c_234_n 0.00181441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_27_297#_c_240_n 0.00848573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_297#_c_241_n 0.00260609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_235_n 0.00118507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_243_n 0.0142826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_348_n 0.00254116f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.202
cc_54 VPB N_VPWR_c_349_n 0.00281864f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.202
cc_55 VPB N_VPWR_c_350_n 0.0163015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_351_n 0.0526033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_352_n 0.0236039f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_347_n 0.0468928f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_354_n 0.00438518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_355_n 0.00580052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.0576226f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_62 N_C1_c_65_n N_B1_c_91_n 0.0275594f $X=0.52 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_63 N_C1_c_62_n N_B1_c_91_n 0.0158089f $X=0.545 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_64 N_C1_c_64_n N_B1_c_91_n 0.00283116f $X=0.52 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_65 N_C1_c_62_n N_B1_c_92_n 0.0211798f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_66 N_C1_c_62_n B1 3.13122e-19 $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_67 N_C1_c_62_n N_A_27_297#_c_233_n 0.0066915f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_68 N_C1_c_65_n N_A_27_297#_c_234_n 0.00225468f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_69 N_C1_c_62_n N_A_27_297#_c_234_n 0.0085797f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_70 C1 N_A_27_297#_c_234_n 0.0207096f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_C1_c_64_n N_A_27_297#_c_234_n 0.0132323f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_72 N_C1_c_65_n N_A_27_297#_c_249_n 5.56577e-19 $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C1_c_65_n N_A_27_297#_c_250_n 6.08578e-19 $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C1_c_65_n N_A_27_297#_c_243_n 0.0198337f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_75 C1 N_A_27_297#_c_243_n 0.0255124f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_76 N_C1_c_64_n N_A_27_297#_c_243_n 0.00770852f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_77 N_C1_c_62_n N_A_27_297#_c_236_n 0.0103596f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_78 C1 N_A_27_297#_c_236_n 0.0180213f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_79 N_C1_c_64_n N_A_27_297#_c_236_n 0.00172493f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_80 N_C1_c_65_n N_VPWR_c_348_n 0.0127807f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_81 N_C1_c_65_n N_VPWR_c_350_n 0.00505556f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_82 N_C1_c_65_n N_VPWR_c_347_n 0.00949224f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_83 N_C1_c_62_n N_A_124_47#_c_425_n 0.00159062f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_84 N_C1_c_62_n N_VGND_c_476_n 0.00413245f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_85 N_C1_c_62_n N_VGND_c_481_n 0.0070422f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_86 N_B1_c_91_n N_B2_c_127_n 0.0919199f $X=1.05 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_87 B1 N_B2_c_127_n 0.00196695f $X=1.09 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_88 N_B1_c_92_n N_B2_c_128_n 0.0245684f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_89 N_B1_c_91_n B2 0.00120316f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_90 B1 B2 0.027089f $X=1.09 $Y=1.19 $X2=0 $Y2=0
cc_91 N_B1_c_92_n N_A_27_297#_c_233_n 5.34835e-19 $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_92 N_B1_c_91_n N_A_27_297#_c_234_n 0.00351822f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B1_c_92_n N_A_27_297#_c_234_n 0.00316216f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_94 B1 N_A_27_297#_c_234_n 0.0254059f $X=1.09 $Y=1.19 $X2=0 $Y2=0
cc_95 N_B1_c_91_n N_A_27_297#_c_261_n 0.0154974f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_96 B1 N_A_27_297#_c_261_n 0.020653f $X=1.09 $Y=1.19 $X2=0 $Y2=0
cc_97 N_B1_c_91_n N_A_27_297#_c_249_n 0.00477003f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B1_c_91_n N_A_27_297#_c_250_n 0.00881639f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B1_c_91_n N_A_27_297#_c_243_n 5.04145e-19 $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B1_c_92_n N_A_27_297#_c_236_n 0.00155254f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_101 N_B1_c_91_n N_A_27_297#_c_267_n 0.00135561f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B1_c_91_n N_VPWR_c_348_n 0.00656953f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B1_c_91_n N_VPWR_c_351_n 0.00589065f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B1_c_91_n N_VPWR_c_347_n 0.00916603f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B1_c_91_n N_A_124_47#_c_425_n 0.002429f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B1_c_92_n N_A_124_47#_c_425_n 0.00844544f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_107 B1 N_A_124_47#_c_425_n 0.00245026f $X=1.09 $Y=1.19 $X2=0 $Y2=0
cc_108 N_B1_c_92_n N_A_230_47#_c_443_n 0.0062585f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_109 B1 N_A_230_47#_c_443_n 0.0127702f $X=1.09 $Y=1.19 $X2=0 $Y2=0
cc_110 N_B1_c_92_n N_VGND_c_476_n 0.00368123f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_111 N_B1_c_92_n N_VGND_c_481_n 0.00561117f $X=1.075 $Y=0.985 $X2=0 $Y2=0
cc_112 N_B2_c_127_n N_A2_c_161_n 0.00332761f $X=1.46 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_113 B2 N_A2_c_161_n 5.81844e-19 $X=1.45 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_114 N_B2_c_127_n A2 0.00188387f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_115 B2 A2 0.0343559f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B2_c_127_n N_A2_c_165_n 8.98273e-19 $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_117 B2 N_A2_c_165_n 0.0222031f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_118 B2 N_A_27_297#_M1005_d 0.00493019f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_119 B2 N_A_27_297#_c_234_n 0.00356744f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B2_c_127_n N_A_27_297#_c_261_n 0.00176803f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_121 B2 N_A_27_297#_c_261_n 0.0175308f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B2_c_127_n N_A_27_297#_c_249_n 0.00336143f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_123 B2 N_A_27_297#_c_243_n 0.0011718f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B2_c_127_n N_A_27_297#_c_274_n 0.00964897f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_125 B2 N_A_27_297#_c_274_n 0.0275369f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_126 N_B2_c_127_n N_A_27_297#_c_267_n 0.0110383f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B2_c_127_n N_VPWR_c_351_n 0.00492735f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B2_c_127_n N_VPWR_c_347_n 0.0078319f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B2_c_128_n N_A_124_47#_c_425_n 0.00805977f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B2_c_127_n N_A_230_47#_c_443_n 0.00155179f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B2_c_128_n N_A_230_47#_c_443_n 0.0104553f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_132 B2 N_A_230_47#_c_443_n 0.0274086f $X=1.45 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B2_c_128_n N_VGND_c_474_n 0.00309694f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_134 N_B2_c_128_n N_VGND_c_476_n 0.00368123f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B2_c_128_n N_VGND_c_481_n 0.00666343f $X=1.52 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_c_161_n N_A1_c_199_n 0.0912336f $X=2.485 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_137 N_A2_c_163_n N_A1_c_199_n 0.00325949f $X=2.45 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_138 N_A2_c_162_n N_A1_c_200_n 0.0104671f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A2_c_163_n N_A1_c_200_n 2.10122e-19 $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_140 N_A2_c_161_n A1 3.2427e-19 $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_163_n A1 0.0132665f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_142 A2 A1 0.00100098f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_143 A2 N_A_27_297#_M1005_d 0.0120391f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A2_c_161_n N_A_27_297#_c_278_n 0.0131521f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_161_n N_A_27_297#_c_241_n 0.00210828f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_163_n N_A_27_297#_c_241_n 0.00303383f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_147 A2 N_A_27_297#_c_241_n 0.0101491f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A2_c_161_n N_A_27_297#_c_267_n 0.00105956f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_163_n N_A_27_297#_c_267_n 0.00566529f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_150 A2 N_A_27_297#_c_267_n 0.0296998f $X=1.98 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A2_c_161_n N_VPWR_c_349_n 0.00266957f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A2_c_161_n N_VPWR_c_351_n 0.00517074f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_161_n N_VPWR_c_347_n 0.00806399f $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_161_n N_A_230_47#_c_443_n 7.117e-19 $X=2.485 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A2_c_162_n N_A_230_47#_c_443_n 0.0118967f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_163_n N_A_230_47#_c_443_n 0.0184096f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_165_n N_A_230_47#_c_443_n 0.0281754f $X=2.147 $Y=1.255 $X2=0 $Y2=0
cc_158 N_A2_c_162_n N_VGND_c_474_n 0.00492082f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_162_n N_VGND_c_478_n 0.00426565f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_162_n N_VGND_c_481_n 0.00706326f $X=2.51 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_200_n N_A_27_297#_c_231_n 0.0251965f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A1_c_199_n N_A_27_297#_c_232_n 0.0512444f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_163 A1 N_A_27_297#_c_232_n 0.00128773f $X=2.85 $Y=1.105 $X2=0 $Y2=0
cc_164 N_A1_c_199_n N_A_27_297#_c_278_n 0.00126993f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A1_c_199_n N_A_27_297#_c_289_n 0.00443178f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A1_c_199_n N_A_27_297#_c_240_n 0.0189729f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_167 A1 N_A_27_297#_c_240_n 0.023452f $X=2.85 $Y=1.105 $X2=0 $Y2=0
cc_168 N_A1_c_199_n N_A_27_297#_c_235_n 0.00174f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_169 A1 N_A_27_297#_c_235_n 0.0125888f $X=2.85 $Y=1.105 $X2=0 $Y2=0
cc_170 N_A1_c_199_n N_VPWR_c_349_n 0.02004f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_199_n N_VPWR_c_351_n 0.00427505f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A1_c_199_n N_VPWR_c_347_n 0.00727648f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_200_n N_X_c_407_n 6.69442e-19 $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_199_n N_A_230_47#_c_453_n 0.00291749f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A1_c_200_n N_A_230_47#_c_453_n 0.00347266f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_176 A1 N_A_230_47#_c_453_n 0.0048882f $X=2.85 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A1_c_200_n N_A_230_47#_c_456_n 0.00412835f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A1_c_200_n N_VGND_c_475_n 0.00291373f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_179 A1 N_VGND_c_475_n 0.00149698f $X=2.85 $Y=1.105 $X2=0 $Y2=0
cc_180 N_A1_c_200_n N_VGND_c_478_n 0.00541964f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_200_n N_VGND_c_481_n 0.00967482f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_261_n N_VPWR_M1011_d 0.00849478f $X=1.03 $Y=1.607 $X2=-0.19
+ $Y2=-0.24
cc_183 N_A_27_297#_c_243_n N_VPWR_M1011_d 0.0015192f $X=0.755 $Y=1.587 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A_27_297#_c_240_n N_VPWR_M1001_d 0.00250873f $X=3.375 $Y=1.54 $X2=0
+ $Y2=0
cc_185 N_A_27_297#_c_238_n N_VPWR_c_348_n 0.0260202f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_243_n N_VPWR_c_348_n 0.0112132f $X=0.755 $Y=1.587 $X2=0
+ $Y2=0
cc_187 N_A_27_297#_c_267_n N_VPWR_c_348_n 0.0107633f $X=2.355 $Y=2.17 $X2=0
+ $Y2=0
cc_188 N_A_27_297#_c_232_n N_VPWR_c_349_n 0.00689479f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_c_278_n N_VPWR_c_349_n 0.0141783f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_c_289_n N_VPWR_c_349_n 0.00593609f $X=2.66 $Y=1.875 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_c_240_n N_VPWR_c_349_n 0.0244146f $X=3.375 $Y=1.54 $X2=0
+ $Y2=0
cc_192 N_A_27_297#_c_238_n N_VPWR_c_350_n 0.0196165f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_193 N_A_27_297#_c_250_n N_VPWR_c_351_n 0.00294834f $X=1.235 $Y=1.96 $X2=0
+ $Y2=0
cc_194 N_A_27_297#_c_278_n N_VPWR_c_351_n 0.00551866f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_195 N_A_27_297#_c_274_n N_VPWR_c_351_n 0.00368324f $X=1.5 $Y=2.17 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_267_n N_VPWR_c_351_n 0.0564672f $X=2.355 $Y=2.17 $X2=0
+ $Y2=0
cc_197 N_A_27_297#_c_232_n N_VPWR_c_352_n 0.00628074f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_M1011_s N_VPWR_c_347_n 0.00463664f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_M1005_d N_VPWR_c_347_n 0.0070165f $X=1.55 $Y=1.485 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_232_n N_VPWR_c_347_n 0.0119903f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_238_n N_VPWR_c_347_n 0.0107063f $X=0.28 $Y=1.96 $X2=0 $Y2=0
cc_202 N_A_27_297#_c_250_n N_VPWR_c_347_n 0.00536598f $X=1.235 $Y=1.96 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_278_n N_VPWR_c_347_n 0.0100174f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_274_n N_VPWR_c_347_n 0.00661985f $X=1.5 $Y=2.17 $X2=0 $Y2=0
cc_205 N_A_27_297#_c_267_n N_VPWR_c_347_n 0.0324864f $X=2.355 $Y=2.17 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_261_n A_228_297# 0.00242967f $X=1.03 $Y=1.607 $X2=-0.19
+ $Y2=-0.24
cc_207 N_A_27_297#_c_249_n A_228_297# 0.00177676f $X=1.132 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_208 N_A_27_297#_c_250_n A_228_297# 7.2151e-19 $X=1.235 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_209 N_A_27_297#_c_274_n A_228_297# 0.00434223f $X=1.5 $Y=2.17 $X2=-0.19
+ $Y2=-0.24
cc_210 N_A_27_297#_c_278_n A_515_297# 0.00359193f $X=2.575 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_27_297#_c_289_n A_515_297# 0.0025022f $X=2.66 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_27_297#_c_231_n N_X_c_407_n 0.00780351f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_27_297#_c_232_n N_X_c_407_n 0.00256506f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_27_297#_c_235_n N_X_c_407_n 0.00577617f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_231_n X 0.00393278f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_27_297#_c_232_n X 0.0253785f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_27_297#_c_240_n X 0.0111565f $X=3.375 $Y=1.54 $X2=0 $Y2=0
cc_218 N_A_27_297#_c_235_n X 0.0350488f $X=3.46 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_27_297#_c_234_n N_A_124_47#_M1010_d 9.62153e-19 $X=0.67 $Y=1.455
+ $X2=-0.19 $Y2=-0.24
cc_220 N_A_27_297#_c_236_n N_A_124_47#_M1010_d 0.00317792f $X=0.67 $Y=0.735
+ $X2=-0.19 $Y2=-0.24
cc_221 N_A_27_297#_c_233_n N_A_124_47#_c_425_n 0.0122361f $X=0.335 $Y=0.39 $X2=0
+ $Y2=0
cc_222 N_A_27_297#_c_236_n N_A_124_47#_c_425_n 0.00381329f $X=0.67 $Y=0.735
+ $X2=0 $Y2=0
cc_223 N_A_27_297#_c_236_n N_A_230_47#_c_443_n 0.00986579f $X=0.67 $Y=0.735
+ $X2=0 $Y2=0
cc_224 N_A_27_297#_c_231_n N_A_230_47#_c_453_n 4.97148e-19 $X=3.4 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_27_297#_c_240_n N_A_230_47#_c_453_n 0.00211033f $X=3.375 $Y=1.54
+ $X2=0 $Y2=0
cc_226 N_A_27_297#_c_241_n N_A_230_47#_c_453_n 0.00400266f $X=2.745 $Y=1.54
+ $X2=0 $Y2=0
cc_227 N_A_27_297#_c_231_n N_VGND_c_475_n 0.00291373f $X=3.4 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_27_297#_c_233_n N_VGND_c_476_n 0.0202909f $X=0.335 $Y=0.39 $X2=0
+ $Y2=0
cc_229 N_A_27_297#_c_236_n N_VGND_c_476_n 0.00289823f $X=0.67 $Y=0.735 $X2=0
+ $Y2=0
cc_230 N_A_27_297#_c_231_n N_VGND_c_480_n 0.00541763f $X=3.4 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_27_297#_M1010_s N_VGND_c_481_n 0.00209319f $X=0.21 $Y=0.235 $X2=0
+ $Y2=0
cc_232 N_A_27_297#_c_231_n N_VGND_c_481_n 0.0106607f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_27_297#_c_233_n N_VGND_c_481_n 0.0122524f $X=0.335 $Y=0.39 $X2=0
+ $Y2=0
cc_234 N_A_27_297#_c_236_n N_VGND_c_481_n 0.00519685f $X=0.67 $Y=0.735 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_347_n A_228_297# 0.00281856f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_236 N_VPWR_c_347_n A_515_297# 0.00464656f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_237 N_VPWR_c_347_n N_X_M1009_d 0.00233913f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_c_352_n X 0.0376376f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_239 N_VPWR_c_347_n X 0.0213505f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_240 N_X_c_407_n N_A_230_47#_c_453_n 0.00575354f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_241 N_X_c_407_n N_VGND_c_480_n 0.0366863f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_242 N_X_M1006_d N_VGND_c_481_n 0.00267115f $X=3.475 $Y=0.235 $X2=0 $Y2=0
cc_243 N_X_c_407_n N_VGND_c_481_n 0.0220874f $X=3.66 $Y=0.39 $X2=0 $Y2=0
cc_244 N_A_124_47#_c_425_n N_A_230_47#_M1008_d 0.00378684f $X=1.73 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_245 N_A_124_47#_M1000_d N_A_230_47#_c_443_n 0.00680324f $X=1.595 $Y=0.235
+ $X2=0 $Y2=0
cc_246 N_A_124_47#_c_425_n N_A_230_47#_c_443_n 0.0470756f $X=1.73 $Y=0.39 $X2=0
+ $Y2=0
cc_247 N_A_124_47#_c_425_n N_VGND_c_474_n 0.0143014f $X=1.73 $Y=0.39 $X2=0 $Y2=0
cc_248 N_A_124_47#_c_425_n N_VGND_c_476_n 0.0527563f $X=1.73 $Y=0.39 $X2=0 $Y2=0
cc_249 N_A_124_47#_M1010_d N_VGND_c_481_n 0.0033767f $X=0.62 $Y=0.235 $X2=0
+ $Y2=0
cc_250 N_A_124_47#_M1000_d N_VGND_c_481_n 0.0021262f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_124_47#_c_425_n N_VGND_c_481_n 0.0419716f $X=1.73 $Y=0.39 $X2=0 $Y2=0
cc_252 N_A_230_47#_c_443_n N_VGND_M1007_s 0.0063498f $X=2.605 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_230_47#_c_443_n N_VGND_c_474_n 0.0224613f $X=2.605 $Y=0.73 $X2=0
+ $Y2=0
cc_254 N_A_230_47#_c_443_n N_VGND_c_476_n 0.0032114f $X=2.605 $Y=0.73 $X2=0
+ $Y2=0
cc_255 N_A_230_47#_c_443_n N_VGND_c_478_n 0.00266837f $X=2.605 $Y=0.73 $X2=0
+ $Y2=0
cc_256 N_A_230_47#_c_456_n N_VGND_c_478_n 0.0177776f $X=2.77 $Y=0.39 $X2=0 $Y2=0
cc_257 N_A_230_47#_M1008_d N_VGND_c_481_n 0.00240642f $X=1.15 $Y=0.235 $X2=0
+ $Y2=0
cc_258 N_A_230_47#_M1007_d N_VGND_c_481_n 0.0026238f $X=2.585 $Y=0.235 $X2=0
+ $Y2=0
cc_259 N_A_230_47#_c_443_n N_VGND_c_481_n 0.012346f $X=2.605 $Y=0.73 $X2=0 $Y2=0
cc_260 N_A_230_47#_c_456_n N_VGND_c_481_n 0.0122607f $X=2.77 $Y=0.39 $X2=0 $Y2=0
