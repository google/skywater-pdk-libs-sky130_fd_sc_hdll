* File: sky130_fd_sc_hdll__inputiso0n_1.pxi.spice
* Created: Thu Aug 27 19:08:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A N_A_c_48_n N_A_c_49_n N_A_M1002_g
+ N_A_M1005_g A A N_A_c_46_n N_A_c_47_n PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%SLEEP_B N_SLEEP_B_M1003_g N_SLEEP_B_c_80_n
+ N_SLEEP_B_c_81_n N_SLEEP_B_M1004_g SLEEP_B N_SLEEP_B_c_78_n SLEEP_B
+ PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%SLEEP_B
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A_27_75# N_A_27_75#_M1005_s
+ N_A_27_75#_M1002_d N_A_27_75#_c_117_n N_A_27_75#_M1001_g N_A_27_75#_c_118_n
+ N_A_27_75#_M1000_g N_A_27_75#_c_119_n N_A_27_75#_c_120_n N_A_27_75#_c_121_n
+ N_A_27_75#_c_124_n N_A_27_75#_c_125_n N_A_27_75#_c_126_n N_A_27_75#_c_122_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%A_27_75#
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VPWR N_VPWR_M1002_s N_VPWR_M1004_d
+ N_VPWR_c_187_n N_VPWR_c_188_n N_VPWR_c_189_n N_VPWR_c_190_n N_VPWR_c_191_n
+ VPWR N_VPWR_c_192_n N_VPWR_c_186_n PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VPWR
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%X N_X_M1001_d N_X_M1000_d N_X_c_216_n X X X
+ X X X N_X_c_218_n X PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%X
x_PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VGND N_VGND_M1003_d N_VGND_c_240_n
+ N_VGND_c_241_n N_VGND_c_242_n VGND N_VGND_c_243_n N_VGND_c_244_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO0N_1%VGND
cc_1 VNB N_A_M1005_g 0.0275859f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_2 VNB N_A_c_46_n 0.0314472f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.16
cc_3 VNB N_A_c_47_n 0.01147f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.16
cc_4 VNB N_SLEEP_B_M1003_g 0.0219754f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.78
cc_5 VNB N_SLEEP_B_c_78_n 0.021383f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB SLEEP_B 0.00466194f $X=-0.19 $Y=-0.24 $X2=0.232 $Y2=1.53
cc_7 VNB N_A_27_75#_c_117_n 0.0233006f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_8 VNB N_A_27_75#_c_118_n 0.0263222f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_9 VNB N_A_27_75#_c_119_n 0.0167511f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.16
cc_10 VNB N_A_27_75#_c_120_n 0.0092701f $X=-0.19 $Y=-0.24 $X2=0.452 $Y2=0.995
cc_11 VNB N_A_27_75#_c_121_n 0.0108744f $X=-0.19 $Y=-0.24 $X2=0.452 $Y2=1.325
cc_12 VNB N_A_27_75#_c_122_n 9.57069e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_186_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.425 $Y2=1.2
cc_14 VNB N_X_c_216_n 0.0037621f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_15 VNB X 0.0405607f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_16 VNB N_X_c_218_n 0.0160773f $X=-0.19 $Y=-0.24 $X2=0.232 $Y2=1.2
cc_17 VNB N_VGND_c_240_n 0.00686176f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_18 VNB N_VGND_c_241_n 0.0342604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_242_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_20 VNB N_VGND_c_243_n 0.0235029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_244_n 0.15801f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_22 VPB N_A_c_48_n 0.021869f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.68
cc_23 VPB N_A_c_49_n 0.0289159f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.78
cc_24 VPB A 0.0221615f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_25 VPB N_A_c_46_n 0.00561185f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_26 VPB N_A_c_47_n 0.00128319f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_27 VPB N_SLEEP_B_c_80_n 0.0211694f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_28 VPB N_SLEEP_B_c_81_n 0.0232003f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.585
cc_29 VPB N_SLEEP_B_c_78_n 0.00288282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB SLEEP_B 0.00187008f $X=-0.19 $Y=1.305 $X2=0.232 $Y2=1.53
cc_31 VPB N_A_27_75#_c_118_n 0.0331469f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_A_27_75#_c_124_n 0.0041724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_75#_c_125_n 0.00335032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_75#_c_126_n 0.00569323f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_75#_c_122_n 0.00170982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_187_n 0.0115481f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.585
cc_37 VPB N_VPWR_c_188_n 0.0305804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_189_n 0.00727093f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_190_n 0.0224301f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_40 VPB N_VPWR_c_191_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0.452 $Y2=0.995
cc_41 VPB N_VPWR_c_192_n 0.0220863f $X=-0.19 $Y=1.305 $X2=0.232 $Y2=1.2
cc_42 VPB N_VPWR_c_186_n 0.0599671f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.2
cc_43 VPB X 0.0275926f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_44 VPB X 0.0260164f $X=-0.19 $Y=1.305 $X2=0.425 $Y2=1.16
cc_45 N_A_M1005_g N_SLEEP_B_M1003_g 0.0182346f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_46 N_A_c_48_n N_SLEEP_B_c_80_n 0.0182346f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_47 N_A_c_49_n N_SLEEP_B_c_81_n 0.0295651f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_48 N_A_c_46_n N_SLEEP_B_c_78_n 0.0182346f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A_c_47_n N_SLEEP_B_c_78_n 2.91318e-19 $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A_c_46_n SLEEP_B 0.00171024f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_51 N_A_c_47_n SLEEP_B 0.0148844f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_M1005_g N_A_27_75#_c_119_n 8.59843e-19 $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_A_27_75#_c_120_n 0.015115f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_54 N_A_c_46_n N_A_27_75#_c_120_n 2.87475e-19 $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_c_47_n N_A_27_75#_c_120_n 0.00950835f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_c_46_n N_A_27_75#_c_121_n 0.00437359f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_57 N_A_c_47_n N_A_27_75#_c_121_n 0.0274862f $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_c_49_n N_A_27_75#_c_124_n 0.00361973f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_59 N_A_c_48_n N_A_27_75#_c_126_n 0.00322503f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_60 A N_A_27_75#_c_126_n 0.00710367f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_61 N_A_c_49_n N_VPWR_c_188_n 0.0052997f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_62 A N_VPWR_c_188_n 0.014564f $X=0.145 $Y=1.445 $X2=0 $Y2=0
cc_63 N_A_c_46_n N_VPWR_c_188_n 8.04075e-19 $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_c_47_n N_VPWR_c_188_n 5.44174e-19 $X=0.425 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_c_49_n N_VPWR_c_190_n 0.00628791f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_66 N_A_c_49_n N_VPWR_c_186_n 0.00622823f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_67 N_A_M1005_g N_VGND_c_241_n 0.0044865f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_VGND_c_244_n 0.00541051f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_69 N_SLEEP_B_M1003_g N_A_27_75#_c_117_n 0.0150079f $X=0.96 $Y=0.585 $X2=0
+ $Y2=0
cc_70 N_SLEEP_B_c_80_n N_A_27_75#_c_118_n 0.0139718f $X=0.985 $Y=1.68 $X2=0
+ $Y2=0
cc_71 N_SLEEP_B_c_81_n N_A_27_75#_c_118_n 0.00784135f $X=0.985 $Y=1.78 $X2=0
+ $Y2=0
cc_72 N_SLEEP_B_c_78_n N_A_27_75#_c_118_n 0.0123365f $X=1.02 $Y=1.16 $X2=0 $Y2=0
cc_73 SLEEP_B N_A_27_75#_c_118_n 0.00190545f $X=1.1 $Y=1.19 $X2=0 $Y2=0
cc_74 N_SLEEP_B_M1003_g N_A_27_75#_c_120_n 0.0135049f $X=0.96 $Y=0.585 $X2=0
+ $Y2=0
cc_75 N_SLEEP_B_c_78_n N_A_27_75#_c_120_n 0.00318062f $X=1.02 $Y=1.16 $X2=0
+ $Y2=0
cc_76 SLEEP_B N_A_27_75#_c_120_n 0.0312046f $X=1.1 $Y=1.19 $X2=0 $Y2=0
cc_77 N_SLEEP_B_c_81_n N_A_27_75#_c_124_n 0.011278f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_78 N_SLEEP_B_c_80_n N_A_27_75#_c_125_n 0.00579938f $X=0.985 $Y=1.68 $X2=0
+ $Y2=0
cc_79 N_SLEEP_B_c_81_n N_A_27_75#_c_125_n 0.00869312f $X=0.985 $Y=1.78 $X2=0
+ $Y2=0
cc_80 N_SLEEP_B_c_78_n N_A_27_75#_c_125_n 0.00148643f $X=1.02 $Y=1.16 $X2=0
+ $Y2=0
cc_81 SLEEP_B N_A_27_75#_c_125_n 0.0190066f $X=1.1 $Y=1.19 $X2=0 $Y2=0
cc_82 N_SLEEP_B_c_80_n N_A_27_75#_c_126_n 0.00207597f $X=0.985 $Y=1.68 $X2=0
+ $Y2=0
cc_83 N_SLEEP_B_c_81_n N_A_27_75#_c_126_n 8.61603e-19 $X=0.985 $Y=1.78 $X2=0
+ $Y2=0
cc_84 SLEEP_B N_A_27_75#_c_126_n 0.0043027f $X=1.1 $Y=1.19 $X2=0 $Y2=0
cc_85 N_SLEEP_B_M1003_g N_A_27_75#_c_122_n 4.56649e-19 $X=0.96 $Y=0.585 $X2=0
+ $Y2=0
cc_86 N_SLEEP_B_c_80_n N_A_27_75#_c_122_n 0.00137971f $X=0.985 $Y=1.68 $X2=0
+ $Y2=0
cc_87 N_SLEEP_B_c_78_n N_A_27_75#_c_122_n 7.29826e-19 $X=1.02 $Y=1.16 $X2=0
+ $Y2=0
cc_88 SLEEP_B N_A_27_75#_c_122_n 0.0144024f $X=1.1 $Y=1.19 $X2=0 $Y2=0
cc_89 N_SLEEP_B_c_81_n N_VPWR_c_189_n 0.00670958f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_90 N_SLEEP_B_c_81_n N_VPWR_c_190_n 0.00601158f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_91 N_SLEEP_B_c_81_n N_VPWR_c_186_n 0.00622823f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_92 N_SLEEP_B_M1003_g N_VGND_c_240_n 0.0074433f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_93 N_SLEEP_B_M1003_g N_VGND_c_241_n 0.0044865f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_94 N_SLEEP_B_M1003_g N_VGND_c_244_n 0.00541051f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_95 N_A_27_75#_c_125_n N_VPWR_M1004_d 0.0079285f $X=1.525 $Y=1.66 $X2=0 $Y2=0
cc_96 N_A_27_75#_c_124_n N_VPWR_c_188_n 0.00129362f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_97 N_A_27_75#_c_118_n N_VPWR_c_189_n 0.0138671f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_27_75#_c_124_n N_VPWR_c_189_n 0.0218238f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_99 N_A_27_75#_c_125_n N_VPWR_c_189_n 0.0219076f $X=1.525 $Y=1.66 $X2=0 $Y2=0
cc_100 N_A_27_75#_c_124_n N_VPWR_c_190_n 0.0101858f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_101 N_A_27_75#_c_118_n N_VPWR_c_192_n 0.00622633f $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_102 N_A_27_75#_c_118_n N_VPWR_c_186_n 0.011586f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_27_75#_c_124_n N_VPWR_c_186_n 0.0103957f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_104 N_A_27_75#_c_120_n N_X_M1001_d 0.00242723f $X=1.525 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_105 N_A_27_75#_c_117_n N_X_c_216_n 0.0037431f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_27_75#_c_118_n N_X_c_216_n 0.0016869f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_27_75#_c_120_n N_X_c_216_n 0.00329134f $X=1.525 $Y=0.81 $X2=0 $Y2=0
cc_108 N_A_27_75#_c_117_n X 0.00633727f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_27_75#_c_118_n X 0.0153137f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_27_75#_c_120_n X 0.0119205f $X=1.525 $Y=0.81 $X2=0 $Y2=0
cc_111 N_A_27_75#_c_122_n X 0.0346586f $X=1.61 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_27_75#_c_118_n X 0.0131756f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_27_75#_c_120_n A_123_75# 0.00297727f $X=1.525 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_114 N_A_27_75#_c_120_n N_VGND_M1003_d 0.00484777f $X=1.525 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_27_75#_c_117_n N_VGND_c_240_n 0.0044954f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_27_75#_c_120_n N_VGND_c_240_n 0.0190303f $X=1.525 $Y=0.81 $X2=0 $Y2=0
cc_117 N_A_27_75#_c_119_n N_VGND_c_241_n 0.0141462f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_118 N_A_27_75#_c_120_n N_VGND_c_241_n 0.00912453f $X=1.525 $Y=0.81 $X2=0
+ $Y2=0
cc_119 N_A_27_75#_c_117_n N_VGND_c_243_n 0.00420701f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_120 N_A_27_75#_c_120_n N_VGND_c_243_n 0.00212778f $X=1.525 $Y=0.81 $X2=0
+ $Y2=0
cc_121 N_A_27_75#_c_117_n N_VGND_c_244_n 0.00816627f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_27_75#_c_119_n N_VGND_c_244_n 0.0118806f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_123 N_A_27_75#_c_120_n N_VGND_c_244_n 0.02414f $X=1.525 $Y=0.81 $X2=0 $Y2=0
cc_124 N_VPWR_c_186_n N_X_M1000_d 0.00581497f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_125 N_VPWR_c_189_n X 0.0336344f $X=1.34 $Y=2 $X2=0 $Y2=0
cc_126 N_VPWR_c_192_n X 0.0322136f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_127 N_VPWR_c_186_n X 0.0175942f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_128 N_X_c_216_n N_VGND_c_243_n 0.021889f $X=1.955 $Y=0.4 $X2=0 $Y2=0
cc_129 N_X_c_218_n N_VGND_c_243_n 0.0179238f $X=2.08 $Y=0.545 $X2=0 $Y2=0
cc_130 N_X_M1001_d N_VGND_c_244_n 0.00209344f $X=1.625 $Y=0.235 $X2=0 $Y2=0
cc_131 N_X_c_216_n N_VGND_c_244_n 0.0133552f $X=1.955 $Y=0.4 $X2=0 $Y2=0
cc_132 N_X_c_218_n N_VGND_c_244_n 0.00962794f $X=2.08 $Y=0.545 $X2=0 $Y2=0
