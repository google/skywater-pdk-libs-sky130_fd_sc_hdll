* File: sky130_fd_sc_hdll__and2_2.pxi.spice
* Created: Wed Sep  2 08:21:23 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2_2%A N_A_c_60_n N_A_c_61_n N_A_M1002_g N_A_M1007_g
+ N_A_c_57_n N_A_c_58_n A A N_A_c_59_n A PM_SKY130_FD_SC_HDLL__AND2_2%A
x_PM_SKY130_FD_SC_HDLL__AND2_2%B N_B_M1004_g N_B_c_96_n N_B_c_97_n N_B_M1006_g B
+ N_B_c_95_n PM_SKY130_FD_SC_HDLL__AND2_2%B
x_PM_SKY130_FD_SC_HDLL__AND2_2%A_27_75# N_A_27_75#_M1007_s N_A_27_75#_M1002_d
+ N_A_27_75#_c_134_n N_A_27_75#_M1001_g N_A_27_75#_c_143_n N_A_27_75#_M1000_g
+ N_A_27_75#_c_135_n N_A_27_75#_c_145_n N_A_27_75#_M1005_g N_A_27_75#_c_136_n
+ N_A_27_75#_M1003_g N_A_27_75#_c_137_n N_A_27_75#_c_138_n N_A_27_75#_c_139_n
+ N_A_27_75#_c_140_n N_A_27_75#_c_147_n N_A_27_75#_c_148_n N_A_27_75#_c_149_n
+ N_A_27_75#_c_141_n N_A_27_75#_c_151_n N_A_27_75#_c_142_n
+ PM_SKY130_FD_SC_HDLL__AND2_2%A_27_75#
x_PM_SKY130_FD_SC_HDLL__AND2_2%VPWR N_VPWR_M1002_s N_VPWR_M1006_d N_VPWR_M1005_s
+ N_VPWR_c_233_n N_VPWR_c_234_n N_VPWR_c_235_n N_VPWR_c_236_n N_VPWR_c_237_n
+ N_VPWR_c_238_n N_VPWR_c_239_n VPWR N_VPWR_c_240_n N_VPWR_c_232_n
+ PM_SKY130_FD_SC_HDLL__AND2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2_2%X N_X_M1001_d N_X_M1000_d N_X_c_272_n X X X X X X
+ N_X_c_289_n X PM_SKY130_FD_SC_HDLL__AND2_2%X
x_PM_SKY130_FD_SC_HDLL__AND2_2%VGND N_VGND_M1004_d N_VGND_M1003_s N_VGND_c_303_n
+ N_VGND_c_304_n N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n VGND
+ N_VGND_c_308_n N_VGND_c_309_n PM_SKY130_FD_SC_HDLL__AND2_2%VGND
cc_1 VNB N_A_M1007_g 0.0275861f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_2 VNB N_A_c_57_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_3 VNB N_A_c_58_n 0.0314655f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_4 VNB N_A_c_59_n 0.0114036f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=1.325
cc_5 VNB N_B_M1004_g 0.0219663f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.78
cc_6 VNB B 0.00287878f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.2
cc_7 VNB N_B_c_95_n 0.0261505f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_8 VNB N_A_27_75#_c_134_n 0.0206551f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_9 VNB N_A_27_75#_c_135_n 0.0217584f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_10 VNB N_A_27_75#_c_136_n 0.0232526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_75#_c_137_n 0.0237142f $X=-0.19 $Y=-0.24 $X2=0.44 $Y2=1.325
cc_12 VNB N_A_27_75#_c_138_n 0.016877f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.51
cc_13 VNB N_A_27_75#_c_139_n 0.00756005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_75#_c_140_n 0.0108802f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=1.2
cc_15 VNB N_A_27_75#_c_141_n 0.00398033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_75#_c_142_n 0.00972688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_232_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB X 9.00734e-19 $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.2
cc_19 VNB N_VGND_c_303_n 0.00686176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_304_n 0.0108057f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.2
cc_21 VNB N_VGND_c_305_n 0.0352669f $X=-0.19 $Y=-0.24 $X2=0.45 $Y2=1.16
cc_22 VNB N_VGND_c_306_n 0.0342225f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.465
cc_23 VNB N_VGND_c_307_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_308_n 0.0235355f $X=-0.19 $Y=-0.24 $X2=0.222 $Y2=1.2
cc_25 VNB N_VGND_c_309_n 0.174029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_A_c_60_n 0.0213057f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.68
cc_27 VPB N_A_c_61_n 0.0264279f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.78
cc_28 VPB N_A_c_57_n 0.00118048f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_29 VPB N_A_c_58_n 0.0065078f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_30 VPB N_A_c_59_n 7.65169e-19 $X=-0.19 $Y=1.305 $X2=0.222 $Y2=1.325
cc_31 VPB A 0.0250781f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.51
cc_32 VPB N_B_c_96_n 0.0211451f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_33 VPB N_B_c_97_n 0.0232012f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.585
cc_34 VPB B 2.38851e-19 $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.2
cc_35 VPB N_B_c_95_n 0.0058252f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_36 VPB N_A_27_75#_c_143_n 0.0188367f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.2
cc_37 VPB N_A_27_75#_c_135_n 0.0125467f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_38 VPB N_A_27_75#_c_145_n 0.0216209f $X=-0.19 $Y=1.305 $X2=0.13 $Y2=1.105
cc_39 VPB N_A_27_75#_c_137_n 0.00976233f $X=-0.19 $Y=1.305 $X2=0.44 $Y2=1.325
cc_40 VPB N_A_27_75#_c_147_n 0.00426034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_75#_c_148_n 0.00331537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_75#_c_149_n 0.00422225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_75#_c_141_n 0.00302901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_75#_c_151_n 0.00176402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_75#_c_142_n 0.00652517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_233_n 0.0112292f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.2
cc_47 VPB N_VPWR_c_234_n 0.0307832f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.16
cc_48 VPB N_VPWR_c_235_n 0.00741355f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.465
cc_49 VPB N_VPWR_c_236_n 0.0107802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_237_n 0.0447066f $X=-0.19 $Y=1.305 $X2=0.44 $Y2=0.995
cc_51 VPB N_VPWR_c_238_n 0.0224301f $X=-0.19 $Y=1.305 $X2=0.222 $Y2=1.55
cc_52 VPB N_VPWR_c_239_n 0.00533035f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_240_n 0.0221069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_232_n 0.0576203f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB X 0.00127749f $X=-0.19 $Y=1.305 $X2=0.45 $Y2=1.2
cc_56 N_A_M1007_g N_B_M1004_g 0.0185917f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_57 N_A_c_60_n N_B_c_96_n 0.0185917f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_58 N_A_c_61_n N_B_c_97_n 0.0299216f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_59 N_A_c_57_n B 0.0210606f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_60 N_A_c_58_n B 2.63054e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_c_57_n N_B_c_95_n 9.57478e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_c_58_n N_B_c_95_n 0.0185917f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_M1007_g N_A_27_75#_c_138_n 8.50375e-19 $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_64 N_A_M1007_g N_A_27_75#_c_139_n 0.0143648f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_65 N_A_c_57_n N_A_27_75#_c_139_n 0.0198329f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_58_n N_A_27_75#_c_139_n 5.77599e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_67 N_A_c_57_n N_A_27_75#_c_140_n 0.00768785f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_c_58_n N_A_27_75#_c_140_n 0.00471094f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_59_n N_A_27_75#_c_140_n 0.0213112f $X=0.222 $Y=1.325 $X2=0 $Y2=0
cc_70 N_A_c_61_n N_A_27_75#_c_147_n 0.00331967f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_71 A N_A_27_75#_c_147_n 0.00115835f $X=0.23 $Y=1.51 $X2=0 $Y2=0
cc_72 N_A_c_60_n N_A_27_75#_c_149_n 0.00192164f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_73 N_A_c_57_n N_A_27_75#_c_149_n 0.00665152f $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_74 A N_A_27_75#_c_149_n 0.00998682f $X=0.23 $Y=1.51 $X2=0 $Y2=0
cc_75 N_A_c_61_n N_VPWR_c_234_n 0.00524062f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_76 N_A_c_57_n N_VPWR_c_234_n 8.11503e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_c_58_n N_VPWR_c_234_n 9.06381e-19 $X=0.45 $Y=1.16 $X2=0 $Y2=0
cc_78 A N_VPWR_c_234_n 0.0190809f $X=0.23 $Y=1.51 $X2=0 $Y2=0
cc_79 N_A_c_61_n N_VPWR_c_238_n 0.00628791f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_80 N_A_c_61_n N_VPWR_c_232_n 0.00622823f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_81 N_A_M1007_g N_VGND_c_306_n 0.0044865f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_82 N_A_M1007_g N_VGND_c_309_n 0.00541051f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_83 N_B_M1004_g N_A_27_75#_c_134_n 0.014501f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_84 N_B_c_96_n N_A_27_75#_c_143_n 0.010202f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_85 N_B_c_97_n N_A_27_75#_c_143_n 0.00782704f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_86 N_B_M1004_g N_A_27_75#_c_139_n 0.0135049f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_87 B N_A_27_75#_c_139_n 0.0276376f $X=0.965 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B_c_95_n N_A_27_75#_c_139_n 0.0058992f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_97_n N_A_27_75#_c_147_n 0.0108082f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_90 N_B_c_96_n N_A_27_75#_c_148_n 0.00606455f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_91 N_B_c_97_n N_A_27_75#_c_148_n 0.0091817f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_92 B N_A_27_75#_c_148_n 0.0184909f $X=0.965 $Y=1.105 $X2=0 $Y2=0
cc_93 N_B_c_95_n N_A_27_75#_c_148_n 0.00382224f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_94 N_B_c_96_n N_A_27_75#_c_149_n 0.00199388f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_95 N_B_c_97_n N_A_27_75#_c_149_n 9.22061e-19 $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_96 B N_A_27_75#_c_149_n 0.0017303f $X=0.965 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B_M1004_g N_A_27_75#_c_141_n 0.00151853f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_98 B N_A_27_75#_c_141_n 0.0200245f $X=0.965 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B_c_95_n N_A_27_75#_c_141_n 0.00271118f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B_c_96_n N_A_27_75#_c_151_n 0.00312673f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_101 N_B_c_96_n N_A_27_75#_c_142_n 0.00231465f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_102 B N_A_27_75#_c_142_n 2.82256e-19 $X=0.965 $Y=1.105 $X2=0 $Y2=0
cc_103 N_B_c_95_n N_A_27_75#_c_142_n 0.0213755f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B_c_97_n N_VPWR_c_235_n 0.00685081f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_105 N_B_c_97_n N_VPWR_c_238_n 0.00610687f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_106 N_B_c_97_n N_VPWR_c_232_n 0.00622823f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_107 N_B_M1004_g N_VGND_c_303_n 0.0074433f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_108 N_B_M1004_g N_VGND_c_306_n 0.0044865f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_109 N_B_M1004_g N_VGND_c_309_n 0.00541051f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_110 N_A_27_75#_c_148_n N_VPWR_M1006_d 0.00742181f $X=1.435 $Y=1.66 $X2=0
+ $Y2=0
cc_111 N_A_27_75#_c_147_n N_VPWR_c_234_n 0.00129362f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_112 N_A_27_75#_c_143_n N_VPWR_c_235_n 0.0132785f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_27_75#_c_145_n N_VPWR_c_235_n 8.4585e-19 $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_27_75#_c_147_n N_VPWR_c_235_n 0.021875f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_115 N_A_27_75#_c_148_n N_VPWR_c_235_n 0.022882f $X=1.435 $Y=1.66 $X2=0 $Y2=0
cc_116 N_A_27_75#_c_145_n N_VPWR_c_237_n 0.0254686f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_27_75#_c_147_n N_VPWR_c_238_n 0.0102131f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_118 N_A_27_75#_c_143_n N_VPWR_c_240_n 0.00622633f $X=1.575 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_27_75#_c_145_n N_VPWR_c_240_n 0.00506625f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_27_75#_c_143_n N_VPWR_c_232_n 0.0107643f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_27_75#_c_145_n N_VPWR_c_232_n 0.00925586f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_122 N_A_27_75#_c_147_n N_VPWR_c_232_n 0.0104052f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_123 N_A_27_75#_c_134_n N_X_c_272_n 0.00393211f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_27_75#_c_135_n N_X_c_272_n 0.00532927f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_27_75#_c_141_n N_X_c_272_n 0.00539009f $X=1.52 $Y=1.325 $X2=0 $Y2=0
cc_126 N_A_27_75#_c_134_n X 0.00551225f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_27_75#_c_143_n X 0.0061861f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_27_75#_c_135_n X 0.0138062f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_75#_c_145_n X 0.0159358f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_75#_c_136_n X 0.0157252f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_27_75#_c_137_n X 0.0227954f $X=2.165 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_27_75#_c_148_n X 0.00827169f $X=1.435 $Y=1.66 $X2=0 $Y2=0
cc_133 N_A_27_75#_c_141_n X 0.0378745f $X=1.52 $Y=1.325 $X2=0 $Y2=0
cc_134 N_A_27_75#_c_151_n X 0.0111494f $X=1.52 $Y=1.575 $X2=0 $Y2=0
cc_135 N_A_27_75#_c_142_n X 6.59779e-19 $X=1.64 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_27_75#_c_143_n X 0.00567252f $X=1.575 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_27_75#_c_135_n X 0.00483998f $X=2.065 $Y=1.16 $X2=0 $Y2=0
cc_138 N_A_27_75#_c_145_n X 0.0112391f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_27_75#_c_141_n X 5.8182e-19 $X=1.52 $Y=1.325 $X2=0 $Y2=0
cc_140 N_A_27_75#_c_136_n N_X_c_289_n 0.0103106f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_27_75#_c_139_n A_123_75# 0.00297727f $X=1.435 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_27_75#_c_139_n N_VGND_M1004_d 0.00484777f $X=1.435 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_27_75#_c_134_n N_VGND_c_303_n 0.0044954f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_27_75#_c_139_n N_VGND_c_303_n 0.0190303f $X=1.435 $Y=0.81 $X2=0 $Y2=0
cc_145 N_A_27_75#_c_136_n N_VGND_c_305_n 0.00620633f $X=2.19 $Y=0.995 $X2=0
+ $Y2=0
cc_146 N_A_27_75#_c_138_n N_VGND_c_306_n 0.0141462f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_147 N_A_27_75#_c_139_n N_VGND_c_306_n 0.00920408f $X=1.435 $Y=0.81 $X2=0
+ $Y2=0
cc_148 N_A_27_75#_c_134_n N_VGND_c_308_n 0.00420655f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_27_75#_c_136_n N_VGND_c_308_n 0.00448754f $X=2.19 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_27_75#_c_141_n N_VGND_c_308_n 0.00212733f $X=1.52 $Y=1.325 $X2=0
+ $Y2=0
cc_151 N_A_27_75#_c_134_n N_VGND_c_309_n 0.00750763f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_27_75#_c_136_n N_VGND_c_309_n 0.0089406f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_27_75#_c_138_n N_VGND_c_309_n 0.0118806f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_154 N_A_27_75#_c_139_n N_VGND_c_309_n 0.0204503f $X=1.435 $Y=0.81 $X2=0 $Y2=0
cc_155 N_A_27_75#_c_141_n N_VGND_c_309_n 0.00390104f $X=1.52 $Y=1.325 $X2=0
+ $Y2=0
cc_156 N_VPWR_c_232_n N_X_M1000_d 0.0061046f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_237_n X 0.0751153f $X=2.46 $Y=1.66 $X2=0 $Y2=0
cc_158 N_VPWR_c_235_n X 0.0337061f $X=1.34 $Y=2 $X2=0 $Y2=0
cc_159 N_VPWR_c_240_n X 0.0297082f $X=2.375 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_232_n X 0.0169361f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_237_n N_VGND_c_305_n 0.0101475f $X=2.46 $Y=1.66 $X2=0 $Y2=0
cc_162 X N_VGND_c_305_n 0.0257094f $X=1.965 $Y=0.425 $X2=0 $Y2=0
cc_163 N_X_c_289_n N_VGND_c_305_n 0.023475f $X=2.07 $Y=0.545 $X2=0 $Y2=0
cc_164 N_X_c_272_n N_VGND_c_308_n 0.0204947f $X=1.935 $Y=0.4 $X2=0 $Y2=0
cc_165 N_X_c_289_n N_VGND_c_308_n 0.0168081f $X=2.07 $Y=0.545 $X2=0 $Y2=0
cc_166 N_X_M1001_d N_VGND_c_309_n 0.00394877f $X=1.625 $Y=0.235 $X2=0 $Y2=0
cc_167 N_X_c_272_n N_VGND_c_309_n 0.0126015f $X=1.935 $Y=0.4 $X2=0 $Y2=0
cc_168 N_X_c_289_n N_VGND_c_309_n 0.00998659f $X=2.07 $Y=0.545 $X2=0 $Y2=0
