* File: sky130_fd_sc_hdll__nor3_1.pex.spice
* Created: Thu Aug 27 19:16:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%C 1 3 4 6 7 12
r30 12 13 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r31 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r33 4 13 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 12 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%B 1 3 4 6 11 14 15
c37 14 0 7.51322e-20 $X=0.695 $Y=1.53
r38 14 15 13.7484 $w=2.83e-07 $l=3.4e-07 $layer=LI1_cond $X=0.737 $Y=1.53
+ $X2=0.737 $Y2=1.87
r39 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r40 8 14 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.737 $Y=1.325
+ $X2=0.737 $Y2=1.53
r41 7 11 7.08927 $w=3.28e-07 $l=2.03e-07 $layer=LI1_cond $X=0.737 $Y=1.16
+ $X2=0.94 $Y2=1.16
r42 7 8 1.61437 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=0.737 $Y=1.16
+ $X2=0.737 $Y2=1.325
r43 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.965 $Y2=1.16
r44 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r45 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r46 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%A 1 3 4 6 7 8 9 14
c31 14 0 7.51322e-20 $X=1.435 $Y=1.202
r32 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.83
+ $Y=1.16 $X2=1.83 $Y2=1.16
r33 14 16 53.4803 $w=3.56e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.83 $Y2=1.202
r34 13 14 3.38483 $w=3.56e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r35 8 9 8.74552 $w=4.63e-07 $l=3.4e-07 $layer=LI1_cond $X=1.972 $Y=1.19
+ $X2=1.972 $Y2=1.53
r36 8 17 0.771663 $w=4.63e-07 $l=3e-08 $layer=LI1_cond $X=1.972 $Y=1.19
+ $X2=1.972 $Y2=1.16
r37 7 17 7.97386 $w=4.63e-07 $l=3.1e-07 $layer=LI1_cond $X=1.972 $Y=0.85
+ $X2=1.972 $Y2=1.16
r38 4 14 18.7059 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r40 1 13 23.0368 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%Y 1 2 3 10 12 14 15 17 24 27 29 33
r56 27 33 2.40809 $w=3.33e-07 $l=7e-08 $layer=LI1_cond $X=0.257 $Y=2.28
+ $X2=0.257 $Y2=2.21
r57 24 27 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=2.365
+ $X2=0.257 $Y2=2.28
r58 24 33 0.27521 $w=3.33e-07 $l=8e-09 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=2.21
r59 24 29 18.6455 $w=3.33e-07 $l=5.42e-07 $layer=LI1_cond $X=0.257 $Y=2.202
+ $X2=0.257 $Y2=1.66
r60 22 23 10.5364 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.265 $Y=0.55
+ $X2=1.265 $Y2=0.74
r61 17 19 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=0.217 $Y=0.55
+ $X2=0.217 $Y2=0.74
r62 14 23 5.37557 $w=2.2e-07 $l=1.12916e-07 $layer=LI1_cond $X=1.33 $Y=0.825
+ $X2=1.265 $Y2=0.74
r63 14 15 94.9251 $w=1.68e-07 $l=1.455e-06 $layer=LI1_cond $X=1.33 $Y=0.825
+ $X2=1.33 $Y2=2.28
r64 13 24 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=0.425 $Y=2.365
+ $X2=0.257 $Y2=2.365
r65 12 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.245 $Y=2.365
+ $X2=1.33 $Y2=2.28
r66 12 13 53.4973 $w=1.68e-07 $l=8.2e-07 $layer=LI1_cond $X=1.245 $Y=2.365
+ $X2=0.425 $Y2=2.365
r67 11 19 3.11056 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.217 $Y2=0.74
r68 10 23 2.2496 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.115 $Y=0.74
+ $X2=1.265 $Y2=0.74
r69 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.74
+ $X2=0.345 $Y2=0.74
r70 3 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r71 3 29 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r72 2 22 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.55
r73 1 17 182 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%VPWR 1 4 6 8 10 17
r24 17 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r25 16 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r26 16 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r27 10 16 7.05937 $w=1.7e-07 $l=3.57e-07 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=1.942 $Y2=2.72
r28 10 12 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r29 8 19 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 8 12 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r31 4 16 2.9068 $w=5.9e-07 $l=1.11781e-07 $layer=LI1_cond $X=1.88 $Y=2.635
+ $X2=1.942 $Y2=2.72
r32 4 6 12.873 $w=5.88e-07 $l=6.35e-07 $layer=LI1_cond $X=1.88 $Y=2.635 $X2=1.88
+ $Y2=2
r33 1 6 150 $w=1.7e-07 $l=7.17635e-07 $layer=licon1_PDIFF $count=4 $X=1.525
+ $Y=1.485 $X2=2.01 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_1%VGND 1 2 9 11 13 18 24 30 33
r32 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 30 32 1.43529 $w=5.1e-07 $l=6e-08 $layer=LI1_cond $X=2.01 $Y=0.2 $X2=2.07
+ $Y2=0.2
r34 28 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r35 27 30 9.56863 $w=5.1e-07 $l=4e-07 $layer=LI1_cond $X=1.61 $Y=0.2 $X2=2.01
+ $Y2=0.2
r36 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r37 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r38 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r39 22 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r40 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r41 19 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r42 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r43 18 27 9.53121 $w=5.1e-07 $l=2.66458e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.61 $Y2=0.2
r44 18 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.15
+ $Y2=0
r45 13 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r46 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r47 11 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r48 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r49 7 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r50 7 9 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.39
r51 2 30 91 $w=1.7e-07 $l=5.97495e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=2.01 $Y2=0.39
r52 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

