* File: sky130_fd_sc_hdll__a2bb2oi_4.pxi.spice
* Created: Thu Aug 27 18:55:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B1 N_B1_c_151_n N_B1_M1011_g N_B1_c_160_n
+ N_B1_M1000_g N_B1_c_152_n N_B1_M1012_g N_B1_c_161_n N_B1_M1002_g N_B1_c_162_n
+ N_B1_M1018_g N_B1_c_153_n N_B1_M1033_g N_B1_c_154_n N_B1_M1032_g N_B1_c_155_n
+ N_B1_M1038_g N_B1_c_156_n N_B1_c_165_n N_B1_c_166_n N_B1_c_157_n N_B1_c_158_n
+ B1 N_B1_c_159_n B1 PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B2 N_B2_c_278_n N_B2_M1014_g N_B2_c_284_n
+ N_B2_M1005_g N_B2_c_279_n N_B2_M1030_g N_B2_c_285_n N_B2_M1010_g N_B2_c_280_n
+ N_B2_M1031_g N_B2_c_286_n N_B2_M1020_g N_B2_c_287_n N_B2_M1026_g N_B2_c_281_n
+ N_B2_M1034_g B2 N_B2_c_282_n N_B2_c_283_n B2
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_4%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_831_21# N_A_831_21#_M1001_s
+ N_A_831_21#_M1019_s N_A_831_21#_M1015_d N_A_831_21#_M1037_d
+ N_A_831_21#_M1007_d N_A_831_21#_M1022_d N_A_831_21#_c_345_n
+ N_A_831_21#_M1006_g N_A_831_21#_c_363_n N_A_831_21#_M1004_g
+ N_A_831_21#_c_346_n N_A_831_21#_M1008_g N_A_831_21#_c_364_n
+ N_A_831_21#_M1009_g N_A_831_21#_c_347_n N_A_831_21#_M1017_g
+ N_A_831_21#_c_365_n N_A_831_21#_M1023_g N_A_831_21#_c_366_n
+ N_A_831_21#_M1029_g N_A_831_21#_c_348_n N_A_831_21#_M1035_g
+ N_A_831_21#_c_349_n N_A_831_21#_c_350_n N_A_831_21#_c_351_n
+ N_A_831_21#_c_352_n N_A_831_21#_c_380_p N_A_831_21#_c_353_n
+ N_A_831_21#_c_384_p N_A_831_21#_c_354_n N_A_831_21#_c_391_p
+ N_A_831_21#_c_367_n N_A_831_21#_c_355_n N_A_831_21#_c_408_p
+ N_A_831_21#_c_368_n N_A_831_21#_c_356_n N_A_831_21#_c_357_n
+ N_A_831_21#_c_358_n N_A_831_21#_c_359_n N_A_831_21#_c_360_n
+ N_A_831_21#_c_370_n N_A_831_21#_c_361_n N_A_831_21#_c_371_n
+ N_A_831_21#_c_362_n PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_831_21#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A1_N N_A1_N_c_559_n N_A1_N_M1001_g
+ N_A1_N_c_565_n N_A1_N_M1013_g N_A1_N_c_560_n N_A1_N_M1003_g N_A1_N_c_566_n
+ N_A1_N_M1021_g N_A1_N_c_561_n N_A1_N_M1019_g N_A1_N_c_567_n N_A1_N_M1027_g
+ N_A1_N_c_568_n N_A1_N_M1028_g N_A1_N_c_562_n N_A1_N_M1024_g A1_N
+ N_A1_N_c_563_n N_A1_N_c_564_n A1_N PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A2_N N_A2_N_c_640_n N_A2_N_M1015_g
+ N_A2_N_c_645_n N_A2_N_M1007_g N_A2_N_c_641_n N_A2_N_M1025_g N_A2_N_c_646_n
+ N_A2_N_M1016_g N_A2_N_c_642_n N_A2_N_M1037_g N_A2_N_c_647_n N_A2_N_M1022_g
+ N_A2_N_c_648_n N_A2_N_M1036_g N_A2_N_c_643_n N_A2_N_M1039_g A2_N
+ N_A2_N_c_668_n N_A2_N_c_644_n A2_N PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_27_297# N_A_27_297#_M1000_d
+ N_A_27_297#_M1002_d N_A_27_297#_M1005_s N_A_27_297#_M1020_s
+ N_A_27_297#_M1032_d N_A_27_297#_M1009_d N_A_27_297#_M1029_d
+ N_A_27_297#_c_716_n N_A_27_297#_c_717_n N_A_27_297#_c_718_n
+ N_A_27_297#_c_719_n N_A_27_297#_c_738_n N_A_27_297#_c_742_n
+ N_A_27_297#_c_743_n N_A_27_297#_c_746_n N_A_27_297#_c_753_n
+ N_A_27_297#_c_782_p N_A_27_297#_c_810_p N_A_27_297#_c_755_n
+ N_A_27_297#_c_720_n N_A_27_297#_c_721_n N_A_27_297#_c_770_p
+ N_A_27_297#_c_747_n N_A_27_297#_c_748_n N_A_27_297#_c_785_p
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VPWR N_VPWR_M1000_s N_VPWR_M1018_s
+ N_VPWR_M1010_d N_VPWR_M1026_d N_VPWR_M1013_d N_VPWR_M1027_d N_VPWR_c_818_n
+ N_VPWR_c_819_n N_VPWR_c_820_n N_VPWR_c_821_n N_VPWR_c_822_n N_VPWR_c_823_n
+ N_VPWR_c_824_n N_VPWR_c_825_n N_VPWR_c_826_n N_VPWR_c_827_n N_VPWR_c_828_n
+ N_VPWR_c_829_n N_VPWR_c_830_n VPWR N_VPWR_c_831_n N_VPWR_c_817_n
+ N_VPWR_c_833_n N_VPWR_c_834_n N_VPWR_c_835_n N_VPWR_c_836_n VPWR
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%Y N_Y_M1014_s N_Y_M1031_s N_Y_M1006_s
+ N_Y_M1017_s N_Y_M1004_s N_Y_M1023_s N_Y_c_963_n N_Y_c_964_n N_Y_c_965_n
+ N_Y_c_980_n N_Y_c_1025_n N_Y_c_970_n N_Y_c_971_n Y N_Y_c_966_n N_Y_c_1011_n
+ N_Y_c_967_n N_Y_c_968_n Y Y N_Y_c_1021_n PM_SKY130_FD_SC_HDLL__A2BB2OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_1259_297# N_A_1259_297#_M1013_s
+ N_A_1259_297#_M1021_s N_A_1259_297#_M1028_s N_A_1259_297#_M1016_s
+ N_A_1259_297#_M1036_s N_A_1259_297#_c_1060_n N_A_1259_297#_c_1061_n
+ N_A_1259_297#_c_1062_n N_A_1259_297#_c_1116_n N_A_1259_297#_c_1063_n
+ N_A_1259_297#_c_1064_n N_A_1259_297#_c_1120_n N_A_1259_297#_c_1074_n
+ N_A_1259_297#_c_1077_n N_A_1259_297#_c_1081_n N_A_1259_297#_c_1065_n
+ N_A_1259_297#_c_1082_n PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_1259_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VGND N_VGND_M1011_d N_VGND_M1012_d
+ N_VGND_M1038_d N_VGND_M1008_d N_VGND_M1035_d N_VGND_M1003_d N_VGND_M1024_d
+ N_VGND_M1025_s N_VGND_M1039_s N_VGND_c_1128_n N_VGND_c_1129_n N_VGND_c_1130_n
+ N_VGND_c_1131_n N_VGND_c_1132_n N_VGND_c_1133_n N_VGND_c_1134_n
+ N_VGND_c_1135_n N_VGND_c_1136_n N_VGND_c_1137_n N_VGND_c_1138_n
+ N_VGND_c_1139_n N_VGND_c_1140_n N_VGND_c_1141_n N_VGND_c_1142_n
+ N_VGND_c_1143_n N_VGND_c_1144_n N_VGND_c_1145_n N_VGND_c_1146_n
+ N_VGND_c_1147_n N_VGND_c_1148_n N_VGND_c_1149_n VGND N_VGND_c_1150_n
+ N_VGND_c_1151_n N_VGND_c_1152_n N_VGND_c_1153_n N_VGND_c_1154_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_109_47# N_A_109_47#_M1011_s
+ N_A_109_47#_M1033_s N_A_109_47#_M1030_d N_A_109_47#_M1034_d
+ N_A_109_47#_c_1296_n N_A_109_47#_c_1293_n N_A_109_47#_c_1294_n
+ N_A_109_47#_c_1307_n N_A_109_47#_c_1295_n N_A_109_47#_c_1312_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_4%A_109_47#
cc_1 VNB N_B1_c_151_n 0.0221045f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B1_c_152_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_B1_c_153_n 0.0169194f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_B1_c_154_n 0.021894f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_5 VNB N_B1_c_155_n 0.0166524f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_6 VNB N_B1_c_156_n 3.4661e-19 $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.445
cc_7 VNB N_B1_c_157_n 0.0210139f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.18
cc_8 VNB N_B1_c_158_n 0.00348417f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.16
cc_9 VNB N_B1_c_159_n 0.0614014f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_10 VNB N_B2_c_278_n 0.0166285f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_B2_c_279_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_12 VNB N_B2_c_280_n 0.017207f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_13 VNB N_B2_c_281_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_14 VNB N_B2_c_282_n 0.0014172f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_15 VNB N_B2_c_283_n 0.0738529f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_16 VNB N_A_831_21#_c_345_n 0.0155668f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_17 VNB N_A_831_21#_c_346_n 0.0167431f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.285
cc_18 VNB N_A_831_21#_c_347_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.16
cc_19 VNB N_A_831_21#_c_348_n 0.0206044f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.202
cc_20 VNB N_A_831_21#_c_349_n 0.0209354f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=1.202
cc_21 VNB N_A_831_21#_c_350_n 0.00467747f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_22 VNB N_A_831_21#_c_351_n 0.00345181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_831_21#_c_352_n 3.42463e-19 $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.18
cc_24 VNB N_A_831_21#_c_353_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_831_21#_c_354_n 0.00447396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_831_21#_c_355_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_831_21#_c_356_n 0.0116369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_831_21#_c_357_n 0.0220401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_831_21#_c_358_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_831_21#_c_359_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_831_21#_c_360_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_831_21#_c_361_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_831_21#_c_362_n 0.0776706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A1_N_c_559_n 0.0197939f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_35 VNB N_A1_N_c_560_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_36 VNB N_A1_N_c_561_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_37 VNB N_A1_N_c_562_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_38 VNB N_A1_N_c_563_n 0.00310534f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_39 VNB N_A1_N_c_564_n 0.0795074f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_40 VNB N_A2_N_c_640_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_41 VNB N_A2_N_c_641_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_42 VNB N_A2_N_c_642_n 0.017199f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_43 VNB N_A2_N_c_643_n 0.0200893f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_44 VNB N_A2_N_c_644_n 0.0777999f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_45 VNB N_VPWR_c_817_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_963_n 0.00686188f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_47 VNB N_Y_c_964_n 0.01006f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.285
cc_48 VNB N_Y_c_965_n 0.00410882f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=1.53
cc_49 VNB N_Y_c_966_n 0.00533617f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.16
cc_50 VNB N_Y_c_967_n 8.91652e-19 $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_51 VNB N_Y_c_968_n 0.00227901f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.202
cc_52 VNB N_VGND_c_1128_n 0.0110498f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=1.53
cc_53 VNB N_VGND_c_1129_n 0.00674759f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.16
cc_54 VNB N_VGND_c_1130_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.16
cc_55 VNB N_VGND_c_1131_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_56 VNB N_VGND_c_1132_n 0.00467422f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.202
cc_57 VNB N_VGND_c_1133_n 0.00468725f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_58 VNB N_VGND_c_1134_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_59 VNB N_VGND_c_1135_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_60 VNB N_VGND_c_1136_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.335 $Y2=1.18
cc_61 VNB N_VGND_c_1137_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_1138_n 0.0609029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1139_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1140_n 0.0195522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_1141_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1142_n 0.019187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1143_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1144_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1145_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1146_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1147_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1148_n 0.0193072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1149_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1150_n 0.0114597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1151_n 0.48942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1152_n 0.00323927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1153_n 0.0203792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1154_n 0.0208752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_109_47#_c_1293_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_80 VNB N_A_109_47#_c_1294_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_81 VNB N_A_109_47#_c_1295_n 0.00248542f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_82 VPB N_B1_c_160_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_83 VPB N_B1_c_161_n 0.0159725f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_84 VPB N_B1_c_162_n 0.0164061f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_85 VPB N_B1_c_154_n 0.0247298f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_86 VPB N_B1_c_156_n 0.00253726f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.445
cc_87 VPB N_B1_c_165_n 0.0104448f $X=-0.19 $Y=1.305 $X2=3.595 $Y2=1.53
cc_88 VPB N_B1_c_166_n 3.61527e-19 $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.53
cc_89 VPB N_B1_c_158_n 0.00267987f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.16
cc_90 VPB N_B1_c_159_n 0.0357538f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.202
cc_91 VPB N_B2_c_284_n 0.0159745f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_92 VPB N_B2_c_285_n 0.0158724f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_93 VPB N_B2_c_286_n 0.0158907f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_94 VPB N_B2_c_287_n 0.0159964f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_95 VPB N_B2_c_283_n 0.0449676f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_96 VPB N_A_831_21#_c_363_n 0.0155159f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.995
cc_97 VPB N_A_831_21#_c_364_n 0.015551f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.53
cc_98 VPB N_A_831_21#_c_365_n 0.0155647f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.53
cc_99 VPB N_A_831_21#_c_366_n 0.0203762f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_831_21#_c_367_n 0.00196649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_831_21#_c_368_n 0.0147349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_831_21#_c_357_n 0.00837143f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_831_21#_c_370_n 0.00180098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_831_21#_c_371_n 0.00152372f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_831_21#_c_362_n 0.0488332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A1_N_c_565_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_107 VPB N_A1_N_c_566_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_108 VPB N_A1_N_c_567_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_109 VPB N_A1_N_c_568_n 0.0161064f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_110 VPB N_A1_N_c_564_n 0.0483911f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_111 VPB N_A2_N_c_645_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_112 VPB N_A2_N_c_646_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_113 VPB N_A2_N_c_647_n 0.0159557f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_114 VPB N_A2_N_c_648_n 0.0191521f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_115 VPB N_A2_N_c_644_n 0.0464475f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_116 VPB N_A_27_297#_c_716_n 0.0332602f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.56
cc_117 VPB N_A_27_297#_c_717_n 0.0018222f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.53
cc_118 VPB N_A_27_297#_c_718_n 0.0107748f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.18
cc_119 VPB N_A_27_297#_c_719_n 0.00169605f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.16
cc_120 VPB N_A_27_297#_c_720_n 0.00183227f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.18
cc_121 VPB N_A_27_297#_c_721_n 0.0107114f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.18
cc_122 VPB N_VPWR_c_818_n 0.00495424f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.56
cc_123 VPB N_VPWR_c_819_n 0.018841f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.285
cc_124 VPB N_VPWR_c_820_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.18
cc_125 VPB N_VPWR_c_821_n 0.0180033f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.16
cc_126 VPB N_VPWR_c_822_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_823_n 0.0180033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_824_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.16
cc_129 VPB N_VPWR_c_825_n 0.00495424f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.202
cc_130 VPB N_VPWR_c_826_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.202
cc_131 VPB N_VPWR_c_827_n 0.0745755f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_132 VPB N_VPWR_c_828_n 0.00401341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_829_n 0.0196545f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.18
cc_134 VPB N_VPWR_c_830_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.335 $Y2=1.18
cc_135 VPB N_VPWR_c_831_n 0.0650397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_817_n 0.0600649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_833_n 0.0233763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_834_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_835_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_836_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_Y_c_965_n 0.00175631f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.53
cc_142 VPB N_Y_c_970_n 0.00180551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_Y_c_971_n 0.00226581f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_144 VPB Y 0.00206711f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_1259_297#_c_1060_n 0.00778987f $X=-0.19 $Y=1.305 $X2=1.46
+ $Y2=0.56
cc_146 VPB N_A_1259_297#_c_1061_n 0.00188366f $X=-0.19 $Y=1.305 $X2=3.81
+ $Y2=0.995
cc_147 VPB N_A_1259_297#_c_1062_n 0.00594968f $X=-0.19 $Y=1.305 $X2=3.81
+ $Y2=0.56
cc_148 VPB N_A_1259_297#_c_1063_n 0.00210846f $X=-0.19 $Y=1.305 $X2=1.705
+ $Y2=1.53
cc_149 VPB N_A_1259_297#_c_1064_n 0.00419265f $X=-0.19 $Y=1.305 $X2=3.785
+ $Y2=1.16
cc_150 VPB N_A_1259_297#_c_1065_n 0.00147495f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.202
cc_151 N_B1_c_153_n N_B2_c_278_n 0.0163834f $X=1.46 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_152 N_B1_c_162_n N_B2_c_284_n 0.0354803f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B1_c_156_n N_B2_c_284_n 7.66774e-19 $X=1.62 $Y=1.445 $X2=0 $Y2=0
cc_154 N_B1_c_165_n N_B2_c_284_n 0.0134805f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_155 N_B1_c_165_n N_B2_c_285_n 0.0119837f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_156 N_B1_c_165_n N_B2_c_286_n 0.0119406f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_157 N_B1_c_154_n N_B2_c_287_n 0.0372348f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B1_c_165_n N_B2_c_287_n 0.0113577f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B1_c_158_n N_B2_c_287_n 0.00101445f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_155_n N_B2_c_281_n 0.022365f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B1_c_154_n N_B2_c_282_n 6.98835e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B1_c_165_n N_B2_c_282_n 0.109756f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_163 N_B1_c_157_n N_B2_c_282_n 0.0176509f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_164 N_B1_c_158_n N_B2_c_282_n 0.0176873f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_154_n N_B2_c_283_n 0.0263635f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B1_c_156_n N_B2_c_283_n 0.00286998f $X=1.62 $Y=1.445 $X2=0 $Y2=0
cc_167 N_B1_c_165_n N_B2_c_283_n 0.0233215f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_168 N_B1_c_157_n N_B2_c_283_n 0.00212345f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_169 N_B1_c_158_n N_B2_c_283_n 0.0039261f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_170 N_B1_c_159_n N_B2_c_283_n 0.0163834f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_171 N_B1_c_155_n N_A_831_21#_c_345_n 0.0257803f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_154_n N_A_831_21#_c_363_n 0.0220261f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B1_c_158_n N_A_831_21#_c_363_n 6.99641e-19 $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_154_n N_A_831_21#_c_362_n 0.0253366f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_158_n N_A_831_21#_c_362_n 0.00111783f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_176 N_B1_c_165_n N_A_27_297#_M1005_s 0.00191634f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_177 N_B1_c_165_n N_A_27_297#_M1020_s 0.00191634f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_178 N_B1_c_158_n N_A_27_297#_M1032_d 0.00158474f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_179 N_B1_c_160_n N_A_27_297#_c_716_n 0.0113204f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_161_n N_A_27_297#_c_716_n 6.54437e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B1_c_160_n N_A_27_297#_c_717_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B1_c_161_n N_A_27_297#_c_717_n 0.0155617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B1_c_157_n N_A_27_297#_c_717_n 0.0458726f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_184 N_B1_c_159_n N_A_27_297#_c_717_n 0.00807006f $X=1.435 $Y=1.202 $X2=0
+ $Y2=0
cc_185 N_B1_c_160_n N_A_27_297#_c_718_n 0.00118933f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B1_c_157_n N_A_27_297#_c_718_n 0.0276437f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_187 N_B1_c_159_n N_A_27_297#_c_718_n 3.16729e-19 $X=1.435 $Y=1.202 $X2=0
+ $Y2=0
cc_188 N_B1_c_162_n N_A_27_297#_c_719_n 2.91946e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B1_c_166_n N_A_27_297#_c_719_n 0.00226125f $X=1.705 $Y=1.53 $X2=0 $Y2=0
cc_190 N_B1_c_157_n N_A_27_297#_c_719_n 0.0196329f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_191 N_B1_c_159_n N_A_27_297#_c_719_n 0.0060737f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_192 N_B1_c_162_n N_A_27_297#_c_738_n 0.0140073f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B1_c_165_n N_A_27_297#_c_738_n 0.0152761f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_194 N_B1_c_166_n N_A_27_297#_c_738_n 0.00941049f $X=1.705 $Y=1.53 $X2=0 $Y2=0
cc_195 N_B1_c_157_n N_A_27_297#_c_738_n 0.00560053f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_196 N_B1_c_165_n N_A_27_297#_c_742_n 0.0354946f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_197 N_B1_c_154_n N_A_27_297#_c_743_n 0.0122041f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_165_n N_A_27_297#_c_743_n 0.0208798f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_199 N_B1_c_158_n N_A_27_297#_c_743_n 0.0160249f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B1_c_158_n N_A_27_297#_c_746_n 0.00356241f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_201 N_B1_c_165_n N_A_27_297#_c_747_n 0.0137032f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_202 N_B1_c_165_n N_A_27_297#_c_748_n 0.0137032f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_203 N_B1_c_165_n N_VPWR_M1018_s 5.67527e-19 $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_204 N_B1_c_166_n N_VPWR_M1018_s 0.00176937f $X=1.705 $Y=1.53 $X2=0 $Y2=0
cc_205 N_B1_c_165_n N_VPWR_M1010_d 0.00192086f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_206 N_B1_c_165_n N_VPWR_M1026_d 0.00175772f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_207 N_B1_c_158_n N_VPWR_M1026_d 7.87733e-19 $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B1_c_160_n N_VPWR_c_818_n 0.00553644f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_161_n N_VPWR_c_818_n 0.00295479f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B1_c_161_n N_VPWR_c_819_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B1_c_162_n N_VPWR_c_819_n 0.0053025f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B1_c_162_n N_VPWR_c_820_n 0.00300743f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B1_c_154_n N_VPWR_c_824_n 0.00300743f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B1_c_154_n N_VPWR_c_827_n 0.0053025f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B1_c_160_n N_VPWR_c_817_n 0.0127552f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_161_n N_VPWR_c_817_n 0.0124092f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B1_c_162_n N_VPWR_c_817_n 0.00693014f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B1_c_154_n N_VPWR_c_817_n 0.00695535f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B1_c_160_n N_VPWR_c_833_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_220 N_B1_c_154_n N_Y_c_964_n 0.00437722f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_221 N_B1_c_155_n N_Y_c_964_n 0.0126966f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_165_n N_Y_c_964_n 0.00577176f $X=3.595 $Y=1.53 $X2=0 $Y2=0
cc_223 N_B1_c_158_n N_Y_c_964_n 0.0294729f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_224 N_B1_c_154_n N_Y_c_965_n 0.00260377f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B1_c_155_n N_Y_c_965_n 0.00172919f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B1_c_158_n N_Y_c_965_n 0.0277636f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B1_c_155_n N_Y_c_980_n 8.53746e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_228 N_B1_c_154_n N_Y_c_971_n 3.08554e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B1_c_158_n N_Y_c_971_n 0.0114244f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B1_c_155_n N_Y_c_967_n 3.78735e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B1_c_151_n N_VGND_c_1129_n 0.00460404f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B1_c_157_n N_VGND_c_1129_n 0.0138247f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_233 N_B1_c_151_n N_VGND_c_1130_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B1_c_152_n N_VGND_c_1130_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B1_c_152_n N_VGND_c_1131_n 0.00385467f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B1_c_153_n N_VGND_c_1131_n 0.00365101f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B1_c_155_n N_VGND_c_1132_n 0.00268723f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B1_c_153_n N_VGND_c_1138_n 0.00395087f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B1_c_155_n N_VGND_c_1138_n 0.00437852f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B1_c_151_n N_VGND_c_1151_n 0.0105827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B1_c_152_n N_VGND_c_1151_n 0.00620835f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B1_c_153_n N_VGND_c_1151_n 0.0058395f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B1_c_155_n N_VGND_c_1151_n 0.00605933f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B1_c_151_n N_A_109_47#_c_1296_n 0.00539651f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_B1_c_152_n N_A_109_47#_c_1296_n 0.00693563f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_B1_c_153_n N_A_109_47#_c_1296_n 5.34196e-19 $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_B1_c_152_n N_A_109_47#_c_1293_n 0.00929182f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_248 N_B1_c_153_n N_A_109_47#_c_1293_n 0.00650032f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_B1_c_157_n N_A_109_47#_c_1293_n 0.0400808f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_250 N_B1_c_159_n N_A_109_47#_c_1293_n 0.00468948f $X=1.435 $Y=1.202 $X2=0
+ $Y2=0
cc_251 N_B1_c_151_n N_A_109_47#_c_1294_n 0.00302596f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_B1_c_152_n N_A_109_47#_c_1294_n 0.00116636f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_B1_c_157_n N_A_109_47#_c_1294_n 0.0307014f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_254 N_B1_c_159_n N_A_109_47#_c_1294_n 0.00358305f $X=1.435 $Y=1.202 $X2=0
+ $Y2=0
cc_255 N_B1_c_153_n N_A_109_47#_c_1307_n 0.00374999f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_B1_c_152_n N_A_109_47#_c_1295_n 5.13362e-19 $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_B1_c_153_n N_A_109_47#_c_1295_n 0.0074807f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_258 N_B1_c_165_n N_A_109_47#_c_1295_n 0.00186641f $X=3.595 $Y=1.53 $X2=0
+ $Y2=0
cc_259 N_B1_c_157_n N_A_109_47#_c_1295_n 0.0217292f $X=1.535 $Y=1.18 $X2=0 $Y2=0
cc_260 N_B2_c_284_n N_A_27_297#_c_738_n 0.01205f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B2_c_285_n N_A_27_297#_c_742_n 0.0120931f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B2_c_286_n N_A_27_297#_c_742_n 0.0120931f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B2_c_287_n N_A_27_297#_c_743_n 0.01205f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B2_c_284_n N_VPWR_c_820_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B2_c_284_n N_VPWR_c_821_n 0.0053025f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B2_c_285_n N_VPWR_c_821_n 0.0053025f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B2_c_285_n N_VPWR_c_822_n 0.00300743f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B2_c_286_n N_VPWR_c_822_n 0.00300743f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B2_c_286_n N_VPWR_c_823_n 0.0053025f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B2_c_287_n N_VPWR_c_823_n 0.0053025f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B2_c_287_n N_VPWR_c_824_n 0.00300743f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B2_c_284_n N_VPWR_c_817_n 0.00693014f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B2_c_285_n N_VPWR_c_817_n 0.00690493f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B2_c_286_n N_VPWR_c_817_n 0.00690493f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B2_c_287_n N_VPWR_c_817_n 0.00693014f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B2_c_278_n N_Y_c_963_n 0.00375858f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B2_c_279_n N_Y_c_963_n 0.0114491f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B2_c_280_n N_Y_c_963_n 0.0114769f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B2_c_282_n N_Y_c_963_n 0.110141f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B2_c_283_n N_Y_c_963_n 0.0117061f $X=3.315 $Y=1.202 $X2=0 $Y2=0
cc_281 N_B2_c_281_n N_Y_c_964_n 0.00793017f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B2_c_281_n N_Y_c_967_n 0.00321762f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B2_c_278_n N_VGND_c_1138_n 0.00357877f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B2_c_279_n N_VGND_c_1138_n 0.00357877f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B2_c_280_n N_VGND_c_1138_n 0.00357877f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B2_c_281_n N_VGND_c_1138_n 0.00357877f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_278_n N_VGND_c_1151_n 0.00538422f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_279_n N_VGND_c_1151_n 0.00548399f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B2_c_280_n N_VGND_c_1151_n 0.00560377f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B2_c_281_n N_VGND_c_1151_n 0.00562222f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B2_c_278_n N_A_109_47#_c_1312_n 0.0121897f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_279_n N_A_109_47#_c_1312_n 0.00931157f $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_B2_c_280_n N_A_109_47#_c_1312_n 0.00964761f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_B2_c_281_n N_A_109_47#_c_1312_n 0.0100245f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B2_c_282_n N_A_109_47#_c_1312_n 0.00123352f $X=3.21 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_831_21#_c_350_n N_A1_N_c_559_n 0.00595356f $X=6.24 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_297 N_A_831_21#_c_351_n N_A1_N_c_559_n 0.0101683f $X=6.675 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_298 N_A_831_21#_c_380_p N_A1_N_c_559_n 0.0110728f $X=6.89 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_831_21#_c_358_n N_A1_N_c_559_n 0.00161382f $X=6.865 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_300 N_A_831_21#_c_380_p N_A1_N_c_560_n 0.00686626f $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_301 N_A_831_21#_c_353_n N_A1_N_c_560_n 0.00901745f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_302 N_A_831_21#_c_384_p N_A1_N_c_560_n 5.24597e-19 $X=7.83 $Y=0.39 $X2=0
+ $Y2=0
cc_303 N_A_831_21#_c_358_n N_A1_N_c_560_n 0.00116636f $X=6.865 $Y=0.815 $X2=0
+ $Y2=0
cc_304 N_A_831_21#_c_380_p N_A1_N_c_561_n 5.45498e-19 $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_305 N_A_831_21#_c_353_n N_A1_N_c_561_n 0.00901745f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_306 N_A_831_21#_c_384_p N_A1_N_c_561_n 0.00651696f $X=7.83 $Y=0.39 $X2=0
+ $Y2=0
cc_307 N_A_831_21#_c_359_n N_A1_N_c_561_n 0.00119564f $X=7.805 $Y=0.815 $X2=0
+ $Y2=0
cc_308 N_A_831_21#_c_354_n N_A1_N_c_562_n 0.0117701f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_309 N_A_831_21#_c_391_p N_A1_N_c_562_n 5.32212e-19 $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_310 N_A_831_21#_c_349_n N_A1_N_c_563_n 0.0131912f $X=6.155 $Y=1.16 $X2=0
+ $Y2=0
cc_311 N_A_831_21#_c_351_n N_A1_N_c_563_n 0.00896514f $X=6.675 $Y=0.82 $X2=0
+ $Y2=0
cc_312 N_A_831_21#_c_353_n N_A1_N_c_563_n 0.0397461f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_313 N_A_831_21#_c_354_n N_A1_N_c_563_n 0.00520815f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_314 N_A_831_21#_c_358_n N_A1_N_c_563_n 0.0306016f $X=6.865 $Y=0.815 $X2=0
+ $Y2=0
cc_315 N_A_831_21#_c_359_n N_A1_N_c_563_n 0.0307352f $X=7.805 $Y=0.815 $X2=0
+ $Y2=0
cc_316 N_A_831_21#_c_349_n N_A1_N_c_564_n 0.00125151f $X=6.155 $Y=1.16 $X2=0
+ $Y2=0
cc_317 N_A_831_21#_c_353_n N_A1_N_c_564_n 0.00345541f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_318 N_A_831_21#_c_358_n N_A1_N_c_564_n 0.00358305f $X=6.865 $Y=0.815 $X2=0
+ $Y2=0
cc_319 N_A_831_21#_c_359_n N_A1_N_c_564_n 0.00486271f $X=7.805 $Y=0.815 $X2=0
+ $Y2=0
cc_320 N_A_831_21#_c_354_n N_A2_N_c_640_n 0.00879863f $X=8.555 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_321 N_A_831_21#_c_391_p N_A2_N_c_640_n 0.00644736f $X=8.77 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_322 N_A_831_21#_c_360_n N_A2_N_c_640_n 0.00116636f $X=8.745 $Y=0.815
+ $X2=-0.19 $Y2=-0.24
cc_323 N_A_831_21#_c_370_n N_A2_N_c_645_n 2.98195e-19 $X=8.77 $Y=1.62 $X2=0
+ $Y2=0
cc_324 N_A_831_21#_c_391_p N_A2_N_c_641_n 0.00686626f $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_325 N_A_831_21#_c_355_n N_A2_N_c_641_n 0.00901745f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_326 N_A_831_21#_c_408_p N_A2_N_c_641_n 5.24597e-19 $X=9.71 $Y=0.39 $X2=0
+ $Y2=0
cc_327 N_A_831_21#_c_360_n N_A2_N_c_641_n 0.00116636f $X=8.745 $Y=0.815 $X2=0
+ $Y2=0
cc_328 N_A_831_21#_c_367_n N_A2_N_c_646_n 0.0128924f $X=9.585 $Y=1.54 $X2=0
+ $Y2=0
cc_329 N_A_831_21#_c_391_p N_A2_N_c_642_n 5.45498e-19 $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_330 N_A_831_21#_c_355_n N_A2_N_c_642_n 0.00901745f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_331 N_A_831_21#_c_408_p N_A2_N_c_642_n 0.00651696f $X=9.71 $Y=0.39 $X2=0
+ $Y2=0
cc_332 N_A_831_21#_c_361_n N_A2_N_c_642_n 0.00119564f $X=9.685 $Y=0.815 $X2=0
+ $Y2=0
cc_333 N_A_831_21#_c_367_n N_A2_N_c_647_n 0.0129531f $X=9.585 $Y=1.54 $X2=0
+ $Y2=0
cc_334 N_A_831_21#_c_368_n N_A2_N_c_648_n 0.0153339f $X=10.135 $Y=1.54 $X2=0
+ $Y2=0
cc_335 N_A_831_21#_c_357_n N_A2_N_c_648_n 0.00179194f $X=10.297 $Y=1.455 $X2=0
+ $Y2=0
cc_336 N_A_831_21#_c_356_n N_A2_N_c_643_n 0.0130523f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_337 N_A_831_21#_c_357_n N_A2_N_c_643_n 0.0193229f $X=10.297 $Y=1.455 $X2=0
+ $Y2=0
cc_338 N_A_831_21#_c_354_n N_A2_N_c_668_n 0.00789367f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_339 N_A_831_21#_c_367_n N_A2_N_c_668_n 0.0464102f $X=9.585 $Y=1.54 $X2=0
+ $Y2=0
cc_340 N_A_831_21#_c_355_n N_A2_N_c_668_n 0.0397461f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_341 N_A_831_21#_c_368_n N_A2_N_c_668_n 0.00856241f $X=10.135 $Y=1.54 $X2=0
+ $Y2=0
cc_342 N_A_831_21#_c_356_n N_A2_N_c_668_n 0.00621501f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_343 N_A_831_21#_c_357_n N_A2_N_c_668_n 0.0165945f $X=10.297 $Y=1.455 $X2=0
+ $Y2=0
cc_344 N_A_831_21#_c_360_n N_A2_N_c_668_n 0.0306016f $X=8.745 $Y=0.815 $X2=0
+ $Y2=0
cc_345 N_A_831_21#_c_370_n N_A2_N_c_668_n 0.0195033f $X=8.77 $Y=1.62 $X2=0 $Y2=0
cc_346 N_A_831_21#_c_361_n N_A2_N_c_668_n 0.0307352f $X=9.685 $Y=0.815 $X2=0
+ $Y2=0
cc_347 N_A_831_21#_c_371_n N_A2_N_c_668_n 0.0195033f $X=9.71 $Y=1.62 $X2=0 $Y2=0
cc_348 N_A_831_21#_c_367_n N_A2_N_c_644_n 0.00869222f $X=9.585 $Y=1.54 $X2=0
+ $Y2=0
cc_349 N_A_831_21#_c_355_n N_A2_N_c_644_n 0.00345541f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_350 N_A_831_21#_c_368_n N_A2_N_c_644_n 9.36362e-19 $X=10.135 $Y=1.54 $X2=0
+ $Y2=0
cc_351 N_A_831_21#_c_360_n N_A2_N_c_644_n 0.00358305f $X=8.745 $Y=0.815 $X2=0
+ $Y2=0
cc_352 N_A_831_21#_c_370_n N_A2_N_c_644_n 0.00659607f $X=8.77 $Y=1.62 $X2=0
+ $Y2=0
cc_353 N_A_831_21#_c_361_n N_A2_N_c_644_n 0.00486271f $X=9.685 $Y=0.815 $X2=0
+ $Y2=0
cc_354 N_A_831_21#_c_371_n N_A2_N_c_644_n 0.00639012f $X=9.71 $Y=1.62 $X2=0
+ $Y2=0
cc_355 N_A_831_21#_c_363_n N_A_27_297#_c_753_n 0.0143578f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_356 N_A_831_21#_c_364_n N_A_27_297#_c_753_n 0.0143578f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_357 N_A_831_21#_c_365_n N_A_27_297#_c_755_n 0.0131651f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_358 N_A_831_21#_c_366_n N_A_27_297#_c_755_n 0.00955151f $X=5.665 $Y=1.41
+ $X2=0 $Y2=0
cc_359 N_A_831_21#_c_366_n N_A_27_297#_c_720_n 0.00169565f $X=5.665 $Y=1.41
+ $X2=0 $Y2=0
cc_360 N_A_831_21#_c_365_n N_A_27_297#_c_721_n 6.83928e-19 $X=5.195 $Y=1.41
+ $X2=0 $Y2=0
cc_361 N_A_831_21#_c_366_n N_A_27_297#_c_721_n 0.0148745f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_362 N_A_831_21#_c_349_n N_A_27_297#_c_721_n 0.0268831f $X=6.155 $Y=1.16 $X2=0
+ $Y2=0
cc_363 N_A_831_21#_c_362_n N_A_27_297#_c_721_n 3.25111e-19 $X=5.665 $Y=1.202
+ $X2=0 $Y2=0
cc_364 N_A_831_21#_c_363_n N_VPWR_c_827_n 0.00429453f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_365 N_A_831_21#_c_364_n N_VPWR_c_827_n 0.00429453f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_366 N_A_831_21#_c_365_n N_VPWR_c_827_n 0.00429453f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_367 N_A_831_21#_c_366_n N_VPWR_c_827_n 0.00429355f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_368 N_A_831_21#_M1007_d N_VPWR_c_817_n 0.00232895f $X=8.625 $Y=1.485 $X2=0
+ $Y2=0
cc_369 N_A_831_21#_M1022_d N_VPWR_c_817_n 0.00232895f $X=9.565 $Y=1.485 $X2=0
+ $Y2=0
cc_370 N_A_831_21#_c_363_n N_VPWR_c_817_n 0.00609021f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_371 N_A_831_21#_c_364_n N_VPWR_c_817_n 0.00606499f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_372 N_A_831_21#_c_365_n N_VPWR_c_817_n 0.00606499f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_373 N_A_831_21#_c_366_n N_VPWR_c_817_n 0.00734727f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_374 N_A_831_21#_c_345_n N_Y_c_965_n 0.00200554f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A_831_21#_c_363_n N_Y_c_965_n 6.35261e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_831_21#_c_346_n N_Y_c_965_n 0.00176907f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A_831_21#_c_349_n N_Y_c_965_n 0.0130288f $X=6.155 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_831_21#_c_362_n N_Y_c_965_n 0.0208386f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_379 N_A_831_21#_c_345_n N_Y_c_980_n 0.00635652f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_831_21#_c_346_n N_Y_c_980_n 0.0066581f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_831_21#_c_347_n N_Y_c_980_n 5.38967e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A_831_21#_c_364_n N_Y_c_970_n 0.017098f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A_831_21#_c_365_n N_Y_c_970_n 0.0132091f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_384 N_A_831_21#_c_362_n N_Y_c_970_n 0.00820504f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_385 N_A_831_21#_c_363_n N_Y_c_971_n 0.0135627f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A_831_21#_c_349_n N_Y_c_971_n 0.0501494f $X=6.155 $Y=1.16 $X2=0 $Y2=0
cc_387 N_A_831_21#_c_362_n N_Y_c_971_n 0.00825408f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_388 N_A_831_21#_c_346_n N_Y_c_966_n 0.00901745f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_389 N_A_831_21#_c_347_n N_Y_c_966_n 0.0101784f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_390 N_A_831_21#_c_348_n N_Y_c_966_n 3.33825e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_391 N_A_831_21#_c_349_n N_Y_c_966_n 0.0695917f $X=6.155 $Y=1.16 $X2=0 $Y2=0
cc_392 N_A_831_21#_c_352_n N_Y_c_966_n 0.00355122f $X=6.325 $Y=0.82 $X2=0 $Y2=0
cc_393 N_A_831_21#_c_362_n N_Y_c_966_n 0.00831339f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_394 N_A_831_21#_c_346_n N_Y_c_1011_n 5.19459e-19 $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_395 N_A_831_21#_c_347_n N_Y_c_1011_n 0.00633209f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_396 N_A_831_21#_c_345_n N_Y_c_968_n 0.00785496f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_397 N_A_831_21#_c_346_n N_Y_c_968_n 0.00116579f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_398 N_A_831_21#_c_349_n N_Y_c_968_n 0.00948654f $X=6.155 $Y=1.16 $X2=0 $Y2=0
cc_399 N_A_831_21#_c_362_n N_Y_c_968_n 0.00436011f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_400 N_A_831_21#_c_365_n Y 0.00195641f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_401 N_A_831_21#_c_366_n Y 0.00201624f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_402 N_A_831_21#_c_349_n Y 0.0216824f $X=6.155 $Y=1.16 $X2=0 $Y2=0
cc_403 N_A_831_21#_c_362_n Y 0.006151f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_404 N_A_831_21#_c_364_n N_Y_c_1021_n 5.74067e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_405 N_A_831_21#_c_365_n N_Y_c_1021_n 0.00820799f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_406 N_A_831_21#_c_367_n N_A_1259_297#_M1016_s 0.00187091f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_407 N_A_831_21#_c_368_n N_A_1259_297#_M1036_s 0.00394616f $X=10.135 $Y=1.54
+ $X2=0 $Y2=0
cc_408 N_A_831_21#_c_366_n N_A_1259_297#_c_1062_n 3.82164e-19 $X=5.665 $Y=1.41
+ $X2=0 $Y2=0
cc_409 N_A_831_21#_c_349_n N_A_1259_297#_c_1062_n 0.00552702f $X=6.155 $Y=1.16
+ $X2=0 $Y2=0
cc_410 N_A_831_21#_c_351_n N_A_1259_297#_c_1062_n 0.0081926f $X=6.675 $Y=0.82
+ $X2=0 $Y2=0
cc_411 N_A_831_21#_c_354_n N_A_1259_297#_c_1063_n 0.00282032f $X=8.555 $Y=0.815
+ $X2=0 $Y2=0
cc_412 N_A_831_21#_c_354_n N_A_1259_297#_c_1064_n 0.00936521f $X=8.555 $Y=0.815
+ $X2=0 $Y2=0
cc_413 N_A_831_21#_c_370_n N_A_1259_297#_c_1064_n 0.00226124f $X=8.77 $Y=1.62
+ $X2=0 $Y2=0
cc_414 N_A_831_21#_M1007_d N_A_1259_297#_c_1074_n 0.00352392f $X=8.625 $Y=1.485
+ $X2=0 $Y2=0
cc_415 N_A_831_21#_c_367_n N_A_1259_297#_c_1074_n 0.00385532f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_416 N_A_831_21#_c_370_n N_A_1259_297#_c_1074_n 0.013395f $X=8.77 $Y=1.62
+ $X2=0 $Y2=0
cc_417 N_A_831_21#_M1022_d N_A_1259_297#_c_1077_n 0.00352392f $X=9.565 $Y=1.485
+ $X2=0 $Y2=0
cc_418 N_A_831_21#_c_367_n N_A_1259_297#_c_1077_n 0.00385532f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_419 N_A_831_21#_c_368_n N_A_1259_297#_c_1077_n 0.00385532f $X=10.135 $Y=1.54
+ $X2=0 $Y2=0
cc_420 N_A_831_21#_c_371_n N_A_1259_297#_c_1077_n 0.013395f $X=9.71 $Y=1.62
+ $X2=0 $Y2=0
cc_421 N_A_831_21#_c_368_n N_A_1259_297#_c_1081_n 0.0191286f $X=10.135 $Y=1.54
+ $X2=0 $Y2=0
cc_422 N_A_831_21#_c_367_n N_A_1259_297#_c_1082_n 0.0143018f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_423 N_A_831_21#_c_351_n N_VGND_M1035_d 0.00223655f $X=6.675 $Y=0.82 $X2=0
+ $Y2=0
cc_424 N_A_831_21#_c_352_n N_VGND_M1035_d 0.00567948f $X=6.325 $Y=0.82 $X2=0
+ $Y2=0
cc_425 N_A_831_21#_c_353_n N_VGND_M1003_d 0.00251047f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_426 N_A_831_21#_c_354_n N_VGND_M1024_d 0.00162089f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_427 N_A_831_21#_c_355_n N_VGND_M1025_s 0.00251047f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_428 N_A_831_21#_c_356_n N_VGND_M1039_s 0.00324618f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_429 N_A_831_21#_c_345_n N_VGND_c_1132_n 0.00268723f $X=4.23 $Y=0.995 $X2=0
+ $Y2=0
cc_430 N_A_831_21#_c_346_n N_VGND_c_1133_n 0.00410249f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_431 N_A_831_21#_c_347_n N_VGND_c_1133_n 0.00276126f $X=5.17 $Y=0.995 $X2=0
+ $Y2=0
cc_432 N_A_831_21#_c_380_p N_VGND_c_1134_n 0.0183628f $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_433 N_A_831_21#_c_353_n N_VGND_c_1134_n 0.0127273f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_434 N_A_831_21#_c_354_n N_VGND_c_1135_n 0.0122559f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_435 N_A_831_21#_c_391_p N_VGND_c_1136_n 0.0183628f $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_436 N_A_831_21#_c_355_n N_VGND_c_1136_n 0.0127273f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_437 N_A_831_21#_c_356_n N_VGND_c_1137_n 0.0130714f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_438 N_A_831_21#_c_345_n N_VGND_c_1140_n 0.00424029f $X=4.23 $Y=0.995 $X2=0
+ $Y2=0
cc_439 N_A_831_21#_c_346_n N_VGND_c_1140_n 0.00424138f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_440 N_A_831_21#_c_351_n N_VGND_c_1142_n 0.00193763f $X=6.675 $Y=0.82 $X2=0
+ $Y2=0
cc_441 N_A_831_21#_c_380_p N_VGND_c_1142_n 0.0223596f $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_442 N_A_831_21#_c_353_n N_VGND_c_1142_n 0.00266636f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_443 N_A_831_21#_c_353_n N_VGND_c_1144_n 0.00198695f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_444 N_A_831_21#_c_384_p N_VGND_c_1144_n 0.0231806f $X=7.83 $Y=0.39 $X2=0
+ $Y2=0
cc_445 N_A_831_21#_c_354_n N_VGND_c_1144_n 0.00254521f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_446 N_A_831_21#_c_354_n N_VGND_c_1146_n 0.00198695f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_447 N_A_831_21#_c_391_p N_VGND_c_1146_n 0.0223596f $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_448 N_A_831_21#_c_355_n N_VGND_c_1146_n 0.00266636f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_449 N_A_831_21#_c_355_n N_VGND_c_1148_n 0.00198695f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_450 N_A_831_21#_c_408_p N_VGND_c_1148_n 0.0231806f $X=9.71 $Y=0.39 $X2=0
+ $Y2=0
cc_451 N_A_831_21#_c_356_n N_VGND_c_1148_n 0.00248202f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_452 N_A_831_21#_c_356_n N_VGND_c_1150_n 0.00321285f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_453 N_A_831_21#_M1001_s N_VGND_c_1151_n 0.0025535f $X=6.705 $Y=0.235 $X2=0
+ $Y2=0
cc_454 N_A_831_21#_M1019_s N_VGND_c_1151_n 0.00304143f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_455 N_A_831_21#_M1015_d N_VGND_c_1151_n 0.0025535f $X=8.585 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_831_21#_M1037_d N_VGND_c_1151_n 0.00304426f $X=9.525 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_831_21#_c_345_n N_VGND_c_1151_n 0.00586948f $X=4.23 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_A_831_21#_c_346_n N_VGND_c_1151_n 0.00609398f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_A_831_21#_c_347_n N_VGND_c_1151_n 0.00608656f $X=5.17 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_A_831_21#_c_348_n N_VGND_c_1151_n 0.012103f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_461 N_A_831_21#_c_351_n N_VGND_c_1151_n 0.0044874f $X=6.675 $Y=0.82 $X2=0
+ $Y2=0
cc_462 N_A_831_21#_c_352_n N_VGND_c_1151_n 7.23891e-19 $X=6.325 $Y=0.82 $X2=0
+ $Y2=0
cc_463 N_A_831_21#_c_380_p N_VGND_c_1151_n 0.0141302f $X=6.89 $Y=0.39 $X2=0
+ $Y2=0
cc_464 N_A_831_21#_c_353_n N_VGND_c_1151_n 0.00972452f $X=7.615 $Y=0.815 $X2=0
+ $Y2=0
cc_465 N_A_831_21#_c_384_p N_VGND_c_1151_n 0.0143352f $X=7.83 $Y=0.39 $X2=0
+ $Y2=0
cc_466 N_A_831_21#_c_354_n N_VGND_c_1151_n 0.0094839f $X=8.555 $Y=0.815 $X2=0
+ $Y2=0
cc_467 N_A_831_21#_c_391_p N_VGND_c_1151_n 0.0141302f $X=8.77 $Y=0.39 $X2=0
+ $Y2=0
cc_468 N_A_831_21#_c_355_n N_VGND_c_1151_n 0.00972452f $X=9.495 $Y=0.815 $X2=0
+ $Y2=0
cc_469 N_A_831_21#_c_408_p N_VGND_c_1151_n 0.0143352f $X=9.71 $Y=0.39 $X2=0
+ $Y2=0
cc_470 N_A_831_21#_c_356_n N_VGND_c_1151_n 0.0111318f $X=10.135 $Y=0.82 $X2=0
+ $Y2=0
cc_471 N_A_831_21#_c_347_n N_VGND_c_1153_n 0.00424138f $X=5.17 $Y=0.995 $X2=0
+ $Y2=0
cc_472 N_A_831_21#_c_348_n N_VGND_c_1153_n 0.00585385f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_473 N_A_831_21#_c_348_n N_VGND_c_1154_n 0.00481673f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_474 N_A_831_21#_c_349_n N_VGND_c_1154_n 0.0123169f $X=6.155 $Y=1.16 $X2=0
+ $Y2=0
cc_475 N_A_831_21#_c_351_n N_VGND_c_1154_n 0.0128272f $X=6.675 $Y=0.82 $X2=0
+ $Y2=0
cc_476 N_A_831_21#_c_352_n N_VGND_c_1154_n 0.0136696f $X=6.325 $Y=0.82 $X2=0
+ $Y2=0
cc_477 N_A1_N_c_562_n N_A2_N_c_640_n 0.0248009f $X=8.09 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_478 N_A1_N_c_568_n N_A2_N_c_645_n 0.00971598f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_479 N_A1_N_c_563_n N_A2_N_c_668_n 0.00892696f $X=7.515 $Y=1.16 $X2=0 $Y2=0
cc_480 N_A1_N_c_564_n N_A2_N_c_668_n 9.13244e-19 $X=8.065 $Y=1.202 $X2=0 $Y2=0
cc_481 N_A1_N_c_563_n N_A2_N_c_644_n 7.60823e-19 $X=7.515 $Y=1.16 $X2=0 $Y2=0
cc_482 N_A1_N_c_564_n N_A2_N_c_644_n 0.0248009f $X=8.065 $Y=1.202 $X2=0 $Y2=0
cc_483 N_A1_N_c_565_n N_A_27_297#_c_721_n 0.00140438f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_484 N_A1_N_c_565_n N_VPWR_c_825_n 0.00553644f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_485 N_A1_N_c_566_n N_VPWR_c_825_n 0.00295479f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_486 N_A1_N_c_567_n N_VPWR_c_826_n 0.00300743f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_487 N_A1_N_c_568_n N_VPWR_c_826_n 0.00300743f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_488 N_A1_N_c_565_n N_VPWR_c_827_n 0.00673617f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_489 N_A1_N_c_566_n N_VPWR_c_829_n 0.00702461f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_490 N_A1_N_c_567_n N_VPWR_c_829_n 0.00702461f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_491 N_A1_N_c_568_n N_VPWR_c_831_n 0.00702461f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_492 N_A1_N_c_565_n N_VPWR_c_817_n 0.0131262f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A1_N_c_566_n N_VPWR_c_817_n 0.0124092f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_494 N_A1_N_c_567_n N_VPWR_c_817_n 0.0124092f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_495 N_A1_N_c_568_n N_VPWR_c_817_n 0.0124344f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_496 N_A1_N_c_565_n N_A_1259_297#_c_1060_n 0.0113322f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_497 N_A1_N_c_566_n N_A_1259_297#_c_1060_n 6.55571e-19 $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_A1_N_c_565_n N_A_1259_297#_c_1061_n 0.0138566f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_499 N_A1_N_c_566_n N_A_1259_297#_c_1061_n 0.015701f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_500 N_A1_N_c_563_n N_A_1259_297#_c_1061_n 0.0440627f $X=7.515 $Y=1.16 $X2=0
+ $Y2=0
cc_501 N_A1_N_c_564_n N_A_1259_297#_c_1061_n 0.00824911f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_502 N_A1_N_c_565_n N_A_1259_297#_c_1062_n 0.00119373f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_503 N_A1_N_c_563_n N_A_1259_297#_c_1062_n 0.00307248f $X=7.515 $Y=1.16 $X2=0
+ $Y2=0
cc_504 N_A1_N_c_564_n N_A_1259_297#_c_1062_n 3.18853e-19 $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_505 N_A1_N_c_567_n N_A_1259_297#_c_1063_n 0.015701f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_506 N_A1_N_c_568_n N_A_1259_297#_c_1063_n 0.0166579f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_507 N_A1_N_c_563_n N_A_1259_297#_c_1063_n 0.0398335f $X=7.515 $Y=1.16 $X2=0
+ $Y2=0
cc_508 N_A1_N_c_564_n N_A_1259_297#_c_1063_n 0.00839792f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_509 N_A1_N_c_563_n N_A_1259_297#_c_1065_n 0.0187469f $X=7.515 $Y=1.16 $X2=0
+ $Y2=0
cc_510 N_A1_N_c_564_n N_A_1259_297#_c_1065_n 0.00632266f $X=8.065 $Y=1.202 $X2=0
+ $Y2=0
cc_511 N_A1_N_c_560_n N_VGND_c_1134_n 0.00379224f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_512 N_A1_N_c_561_n N_VGND_c_1134_n 0.00276126f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_513 N_A1_N_c_562_n N_VGND_c_1135_n 0.00268723f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A1_N_c_559_n N_VGND_c_1142_n 0.00424416f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A1_N_c_560_n N_VGND_c_1142_n 0.00423334f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_516 N_A1_N_c_561_n N_VGND_c_1144_n 0.00423334f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_517 N_A1_N_c_562_n N_VGND_c_1144_n 0.00437852f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_518 N_A1_N_c_559_n N_VGND_c_1151_n 0.00718664f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_519 N_A1_N_c_560_n N_VGND_c_1151_n 0.006093f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_520 N_A1_N_c_561_n N_VGND_c_1151_n 0.00608558f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_521 N_A1_N_c_562_n N_VGND_c_1151_n 0.00615622f $X=8.09 $Y=0.995 $X2=0 $Y2=0
cc_522 N_A1_N_c_559_n N_VGND_c_1154_n 0.00481673f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_523 N_A2_N_c_645_n N_VPWR_c_831_n 0.00429453f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_524 N_A2_N_c_646_n N_VPWR_c_831_n 0.00429453f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_525 N_A2_N_c_647_n N_VPWR_c_831_n 0.00429453f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_526 N_A2_N_c_648_n N_VPWR_c_831_n 0.00429453f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_527 N_A2_N_c_645_n N_VPWR_c_817_n 0.00609021f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_528 N_A2_N_c_646_n N_VPWR_c_817_n 0.00606499f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_529 N_A2_N_c_647_n N_VPWR_c_817_n 0.00606499f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_530 N_A2_N_c_648_n N_VPWR_c_817_n 0.00708296f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_531 N_A2_N_c_645_n N_A_1259_297#_c_1064_n 2.98195e-19 $X=8.535 $Y=1.41 $X2=0
+ $Y2=0
cc_532 N_A2_N_c_645_n N_A_1259_297#_c_1074_n 0.0143578f $X=8.535 $Y=1.41 $X2=0
+ $Y2=0
cc_533 N_A2_N_c_646_n N_A_1259_297#_c_1074_n 0.01161f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_534 N_A2_N_c_647_n N_A_1259_297#_c_1077_n 0.01161f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_535 N_A2_N_c_648_n N_A_1259_297#_c_1077_n 0.01161f $X=9.945 $Y=1.41 $X2=0
+ $Y2=0
cc_536 N_A2_N_c_640_n N_VGND_c_1135_n 0.00268723f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_537 N_A2_N_c_641_n N_VGND_c_1136_n 0.00379224f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_538 N_A2_N_c_642_n N_VGND_c_1136_n 0.00276126f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_539 N_A2_N_c_643_n N_VGND_c_1137_n 0.00438629f $X=9.97 $Y=0.995 $X2=0 $Y2=0
cc_540 N_A2_N_c_640_n N_VGND_c_1146_n 0.00423334f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_541 N_A2_N_c_641_n N_VGND_c_1146_n 0.00423334f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_542 N_A2_N_c_642_n N_VGND_c_1148_n 0.00423334f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_543 N_A2_N_c_643_n N_VGND_c_1148_n 0.00439206f $X=9.97 $Y=0.995 $X2=0 $Y2=0
cc_544 N_A2_N_c_640_n N_VGND_c_1151_n 0.00587047f $X=8.51 $Y=0.995 $X2=0 $Y2=0
cc_545 N_A2_N_c_641_n N_VGND_c_1151_n 0.006093f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A2_N_c_642_n N_VGND_c_1151_n 0.00608558f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_547 N_A2_N_c_643_n N_VGND_c_1151_n 0.00721763f $X=9.97 $Y=0.995 $X2=0 $Y2=0
cc_548 N_A_27_297#_c_717_n N_VPWR_M1000_s 0.00182839f $X=1.075 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_549 N_A_27_297#_c_738_n N_VPWR_M1018_s 0.00374973f $X=2.015 $Y=1.88 $X2=0
+ $Y2=0
cc_550 N_A_27_297#_c_742_n N_VPWR_M1010_d 0.00351985f $X=2.955 $Y=1.88 $X2=0
+ $Y2=0
cc_551 N_A_27_297#_c_743_n N_VPWR_M1026_d 0.00371333f $X=3.895 $Y=1.88 $X2=0
+ $Y2=0
cc_552 N_A_27_297#_c_716_n N_VPWR_c_818_n 0.0413039f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_553 N_A_27_297#_c_717_n N_VPWR_c_818_n 0.0139937f $X=1.075 $Y=1.54 $X2=0
+ $Y2=0
cc_554 N_A_27_297#_c_738_n N_VPWR_c_819_n 0.00260836f $X=2.015 $Y=1.88 $X2=0
+ $Y2=0
cc_555 N_A_27_297#_c_770_p N_VPWR_c_819_n 0.0145763f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_556 N_A_27_297#_c_738_n N_VPWR_c_820_n 0.0138782f $X=2.015 $Y=1.88 $X2=0
+ $Y2=0
cc_557 N_A_27_297#_c_738_n N_VPWR_c_821_n 0.00253649f $X=2.015 $Y=1.88 $X2=0
+ $Y2=0
cc_558 N_A_27_297#_c_742_n N_VPWR_c_821_n 0.00253649f $X=2.955 $Y=1.88 $X2=0
+ $Y2=0
cc_559 N_A_27_297#_c_747_n N_VPWR_c_821_n 0.0149176f $X=2.14 $Y=1.96 $X2=0 $Y2=0
cc_560 N_A_27_297#_c_742_n N_VPWR_c_822_n 0.0138782f $X=2.955 $Y=1.88 $X2=0
+ $Y2=0
cc_561 N_A_27_297#_c_742_n N_VPWR_c_823_n 0.00253649f $X=2.955 $Y=1.88 $X2=0
+ $Y2=0
cc_562 N_A_27_297#_c_743_n N_VPWR_c_823_n 0.00253649f $X=3.895 $Y=1.88 $X2=0
+ $Y2=0
cc_563 N_A_27_297#_c_748_n N_VPWR_c_823_n 0.0149176f $X=3.08 $Y=1.96 $X2=0 $Y2=0
cc_564 N_A_27_297#_c_743_n N_VPWR_c_824_n 0.0137994f $X=3.895 $Y=1.88 $X2=0
+ $Y2=0
cc_565 N_A_27_297#_c_743_n N_VPWR_c_827_n 0.00253649f $X=3.895 $Y=1.88 $X2=0
+ $Y2=0
cc_566 N_A_27_297#_c_753_n N_VPWR_c_827_n 0.0386815f $X=4.835 $Y=2.38 $X2=0
+ $Y2=0
cc_567 N_A_27_297#_c_782_p N_VPWR_c_827_n 0.0149886f $X=4.145 $Y=2.38 $X2=0
+ $Y2=0
cc_568 N_A_27_297#_c_755_n N_VPWR_c_827_n 0.0340228f $X=5.685 $Y=2.38 $X2=0
+ $Y2=0
cc_569 N_A_27_297#_c_720_n N_VPWR_c_827_n 0.0246084f $X=5.875 $Y=2.295 $X2=0
+ $Y2=0
cc_570 N_A_27_297#_c_785_p N_VPWR_c_827_n 0.0146338f $X=4.955 $Y=2.38 $X2=0
+ $Y2=0
cc_571 N_A_27_297#_M1000_d N_VPWR_c_817_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_572 N_A_27_297#_M1002_d N_VPWR_c_817_n 0.00315605f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_573 N_A_27_297#_M1005_s N_VPWR_c_817_n 0.00250248f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_574 N_A_27_297#_M1020_s N_VPWR_c_817_n 0.00250248f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_575 N_A_27_297#_M1032_d N_VPWR_c_817_n 0.00241559f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_576 N_A_27_297#_M1009_d N_VPWR_c_817_n 0.00231265f $X=4.815 $Y=1.485 $X2=0
+ $Y2=0
cc_577 N_A_27_297#_M1029_d N_VPWR_c_817_n 0.00217517f $X=5.755 $Y=1.485 $X2=0
+ $Y2=0
cc_578 N_A_27_297#_c_716_n N_VPWR_c_817_n 0.0128576f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_579 N_A_27_297#_c_738_n N_VPWR_c_817_n 0.0105426f $X=2.015 $Y=1.88 $X2=0
+ $Y2=0
cc_580 N_A_27_297#_c_742_n N_VPWR_c_817_n 0.0102844f $X=2.955 $Y=1.88 $X2=0
+ $Y2=0
cc_581 N_A_27_297#_c_743_n N_VPWR_c_817_n 0.0102828f $X=3.895 $Y=1.88 $X2=0
+ $Y2=0
cc_582 N_A_27_297#_c_753_n N_VPWR_c_817_n 0.0239144f $X=4.835 $Y=2.38 $X2=0
+ $Y2=0
cc_583 N_A_27_297#_c_782_p N_VPWR_c_817_n 0.00962418f $X=4.145 $Y=2.38 $X2=0
+ $Y2=0
cc_584 N_A_27_297#_c_755_n N_VPWR_c_817_n 0.0213236f $X=5.685 $Y=2.38 $X2=0
+ $Y2=0
cc_585 N_A_27_297#_c_720_n N_VPWR_c_817_n 0.0142419f $X=5.875 $Y=2.295 $X2=0
+ $Y2=0
cc_586 N_A_27_297#_c_770_p N_VPWR_c_817_n 0.0091658f $X=1.2 $Y=1.96 $X2=0 $Y2=0
cc_587 N_A_27_297#_c_747_n N_VPWR_c_817_n 0.00954719f $X=2.14 $Y=1.96 $X2=0
+ $Y2=0
cc_588 N_A_27_297#_c_748_n N_VPWR_c_817_n 0.00954719f $X=3.08 $Y=1.96 $X2=0
+ $Y2=0
cc_589 N_A_27_297#_c_785_p N_VPWR_c_817_n 0.00923924f $X=4.955 $Y=2.38 $X2=0
+ $Y2=0
cc_590 N_A_27_297#_c_716_n N_VPWR_c_833_n 0.0217765f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_591 N_A_27_297#_c_753_n N_Y_M1004_s 0.00352392f $X=4.835 $Y=2.38 $X2=0 $Y2=0
cc_592 N_A_27_297#_c_755_n N_Y_M1023_s 0.00345323f $X=5.685 $Y=2.38 $X2=0 $Y2=0
cc_593 N_A_27_297#_c_753_n N_Y_c_1025_n 0.0131184f $X=4.835 $Y=2.38 $X2=0 $Y2=0
cc_594 N_A_27_297#_M1009_d N_Y_c_970_n 0.00192601f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_595 N_A_27_297#_c_810_p N_Y_c_970_n 0.0138549f $X=4.96 $Y=1.96 $X2=0 $Y2=0
cc_596 N_A_27_297#_c_721_n Y 0.0133966f $X=5.9 $Y=1.65 $X2=0 $Y2=0
cc_597 N_A_27_297#_c_755_n N_Y_c_1021_n 0.0159034f $X=5.685 $Y=2.38 $X2=0 $Y2=0
cc_598 N_A_27_297#_c_721_n N_Y_c_1021_n 0.0393635f $X=5.9 $Y=1.65 $X2=0 $Y2=0
cc_599 N_A_27_297#_c_720_n N_A_1259_297#_c_1060_n 0.0139f $X=5.875 $Y=2.295
+ $X2=0 $Y2=0
cc_600 N_A_27_297#_c_721_n N_A_1259_297#_c_1060_n 0.05207f $X=5.9 $Y=1.65 $X2=0
+ $Y2=0
cc_601 N_A_27_297#_c_721_n N_A_1259_297#_c_1062_n 0.0140417f $X=5.9 $Y=1.65
+ $X2=0 $Y2=0
cc_602 N_VPWR_c_817_n N_Y_M1004_s 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_603 N_VPWR_c_817_n N_Y_M1023_s 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_604 N_VPWR_c_817_n N_A_1259_297#_M1013_s 0.00217517f $X=10.35 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_605 N_VPWR_c_817_n N_A_1259_297#_M1021_s 0.00404839f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_606 N_VPWR_c_817_n N_A_1259_297#_M1028_s 0.00297222f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_607 N_VPWR_c_817_n N_A_1259_297#_M1016_s 0.00231264f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_608 N_VPWR_c_817_n N_A_1259_297#_M1036_s 0.00285989f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_609 N_VPWR_c_825_n N_A_1259_297#_c_1060_n 0.0412102f $X=6.89 $Y=1.96 $X2=0
+ $Y2=0
cc_610 N_VPWR_c_827_n N_A_1259_297#_c_1060_n 0.0210596f $X=6.805 $Y=2.72 $X2=0
+ $Y2=0
cc_611 N_VPWR_c_817_n N_A_1259_297#_c_1060_n 0.0124725f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_612 N_VPWR_M1013_d N_A_1259_297#_c_1061_n 0.00182839f $X=6.745 $Y=1.485 $X2=0
+ $Y2=0
cc_613 N_VPWR_c_825_n N_A_1259_297#_c_1061_n 0.0139937f $X=6.89 $Y=1.96 $X2=0
+ $Y2=0
cc_614 N_VPWR_c_829_n N_A_1259_297#_c_1116_n 0.0145763f $X=7.705 $Y=2.72 $X2=0
+ $Y2=0
cc_615 N_VPWR_c_817_n N_A_1259_297#_c_1116_n 0.0091658f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_616 N_VPWR_M1027_d N_A_1259_297#_c_1063_n 0.00187091f $X=7.685 $Y=1.485 $X2=0
+ $Y2=0
cc_617 N_VPWR_c_826_n N_A_1259_297#_c_1063_n 0.0143191f $X=7.83 $Y=1.96 $X2=0
+ $Y2=0
cc_618 N_VPWR_c_831_n N_A_1259_297#_c_1120_n 0.015002f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_619 N_VPWR_c_817_n N_A_1259_297#_c_1120_n 0.00962794f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_620 N_VPWR_c_831_n N_A_1259_297#_c_1074_n 0.0386815f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_621 N_VPWR_c_817_n N_A_1259_297#_c_1074_n 0.0239144f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_622 N_VPWR_c_831_n N_A_1259_297#_c_1077_n 0.0553066f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_623 N_VPWR_c_817_n N_A_1259_297#_c_1077_n 0.0337249f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_624 N_VPWR_c_831_n N_A_1259_297#_c_1082_n 0.0149886f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_625 N_VPWR_c_817_n N_A_1259_297#_c_1082_n 0.00962421f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_626 N_Y_c_964_n N_VGND_M1038_d 0.00162089f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_627 N_Y_c_966_n N_VGND_M1008_d 0.00251047f $X=5.215 $Y=0.815 $X2=0 $Y2=0
cc_628 N_Y_c_964_n N_VGND_c_1132_n 0.0122559f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_629 N_Y_c_980_n N_VGND_c_1133_n 0.0171386f $X=4.49 $Y=0.39 $X2=0 $Y2=0
cc_630 N_Y_c_966_n N_VGND_c_1133_n 0.0127273f $X=5.215 $Y=0.815 $X2=0 $Y2=0
cc_631 N_Y_c_964_n N_VGND_c_1138_n 0.00255089f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_632 N_Y_c_980_n N_VGND_c_1140_n 0.019813f $X=4.49 $Y=0.39 $X2=0 $Y2=0
cc_633 N_Y_c_966_n N_VGND_c_1140_n 0.00266636f $X=5.215 $Y=0.815 $X2=0 $Y2=0
cc_634 N_Y_c_968_n N_VGND_c_1140_n 0.00185026f $X=4.4 $Y=0.815 $X2=0 $Y2=0
cc_635 N_Y_M1014_s N_VGND_c_1151_n 0.00256987f $X=1.955 $Y=0.235 $X2=0 $Y2=0
cc_636 N_Y_M1031_s N_VGND_c_1151_n 0.00297142f $X=2.895 $Y=0.235 $X2=0 $Y2=0
cc_637 N_Y_M1006_s N_VGND_c_1151_n 0.00256339f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_638 N_Y_M1017_s N_VGND_c_1151_n 0.00366014f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_639 N_Y_c_964_n N_VGND_c_1151_n 0.00765082f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_640 N_Y_c_980_n N_VGND_c_1151_n 0.0139822f $X=4.49 $Y=0.39 $X2=0 $Y2=0
cc_641 N_Y_c_966_n N_VGND_c_1151_n 0.00972452f $X=5.215 $Y=0.815 $X2=0 $Y2=0
cc_642 N_Y_c_1011_n N_VGND_c_1151_n 0.0141809f $X=5.43 $Y=0.39 $X2=0 $Y2=0
cc_643 N_Y_c_968_n N_VGND_c_1151_n 0.00300741f $X=4.4 $Y=0.815 $X2=0 $Y2=0
cc_644 N_Y_c_966_n N_VGND_c_1153_n 0.00198695f $X=5.215 $Y=0.815 $X2=0 $Y2=0
cc_645 N_Y_c_1011_n N_VGND_c_1153_n 0.0205249f $X=5.43 $Y=0.39 $X2=0 $Y2=0
cc_646 N_Y_c_963_n N_A_109_47#_M1030_d 0.00214342f $X=3.165 $Y=0.775 $X2=0 $Y2=0
cc_647 N_Y_c_964_n N_A_109_47#_M1034_d 0.00253211f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_648 N_Y_c_963_n N_A_109_47#_c_1295_n 0.00841895f $X=3.165 $Y=0.775 $X2=0
+ $Y2=0
cc_649 N_Y_M1014_s N_A_109_47#_c_1312_n 0.00400389f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_650 N_Y_M1031_s N_A_109_47#_c_1312_n 0.00507817f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_651 N_Y_c_963_n N_A_109_47#_c_1312_n 0.0727148f $X=3.165 $Y=0.775 $X2=0 $Y2=0
cc_652 N_Y_c_964_n N_A_109_47#_c_1312_n 0.0161283f $X=4.145 $Y=0.815 $X2=0 $Y2=0
cc_653 N_VGND_c_1151_n N_A_109_47#_M1011_s 0.0025535f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_654 N_VGND_c_1151_n N_A_109_47#_M1033_s 0.00215206f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_655 N_VGND_c_1151_n N_A_109_47#_M1030_d 0.00255381f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_656 N_VGND_c_1151_n N_A_109_47#_M1034_d 0.00264825f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_657 N_VGND_c_1130_n N_A_109_47#_c_1296_n 0.0223596f $X=1.115 $Y=0 $X2=0 $Y2=0
cc_658 N_VGND_c_1131_n N_A_109_47#_c_1296_n 0.0183628f $X=1.2 $Y=0.39 $X2=0
+ $Y2=0
cc_659 N_VGND_c_1151_n N_A_109_47#_c_1296_n 0.0141302f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_660 N_VGND_M1012_d N_A_109_47#_c_1293_n 0.00348805f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_661 N_VGND_c_1130_n N_A_109_47#_c_1293_n 0.00266636f $X=1.115 $Y=0 $X2=0
+ $Y2=0
cc_662 N_VGND_c_1131_n N_A_109_47#_c_1293_n 0.0131987f $X=1.2 $Y=0.39 $X2=0
+ $Y2=0
cc_663 N_VGND_c_1138_n N_A_109_47#_c_1293_n 0.00199443f $X=3.935 $Y=0 $X2=0
+ $Y2=0
cc_664 N_VGND_c_1151_n N_A_109_47#_c_1293_n 0.0100158f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_665 N_VGND_c_1129_n N_A_109_47#_c_1294_n 0.00750114f $X=0.26 $Y=0.39 $X2=0
+ $Y2=0
cc_666 N_VGND_c_1131_n N_A_109_47#_c_1307_n 0.0172916f $X=1.2 $Y=0.39 $X2=0
+ $Y2=0
cc_667 N_VGND_c_1138_n N_A_109_47#_c_1307_n 0.0186086f $X=3.935 $Y=0 $X2=0 $Y2=0
cc_668 N_VGND_c_1151_n N_A_109_47#_c_1307_n 0.0111017f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_669 N_VGND_c_1131_n N_A_109_47#_c_1295_n 0.00582645f $X=1.2 $Y=0.39 $X2=0
+ $Y2=0
cc_670 N_VGND_c_1138_n N_A_109_47#_c_1312_n 0.110952f $X=3.935 $Y=0 $X2=0 $Y2=0
cc_671 N_VGND_c_1151_n N_A_109_47#_c_1312_n 0.0703895f $X=10.35 $Y=0 $X2=0 $Y2=0
