* NGSPICE file created from sky130_fd_sc_hdll__or2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or2_2 A B VGND VNB VPB VPWR X
M1000 VPWR A a_129_297# VPB phighvt w=420000u l=180000u
+  ad=5.957e+11p pd=5.29e+06u as=9.66e+10p ps=1.3e+06u
M1001 X a_39_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=0p ps=0u
M1002 a_129_297# B a_39_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 VGND A a_39_297# VNB nshort w=420000u l=150000u
+  ad=5.337e+11p pd=5.39e+06u as=1.134e+11p ps=1.38e+06u
M1004 VGND a_39_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1005 X a_39_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_39_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_39_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

