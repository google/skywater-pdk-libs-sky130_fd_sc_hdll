* File: sky130_fd_sc_hdll__muxb4to1_4.pex.spice
* Created: Wed Sep  2 08:35:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[0] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r83 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.905 $Y2=1.16
r84 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=1.62 $Y=1.16
+ $X2=1.88 $Y2=1.16
r85 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.62
+ $Y=1.16 $X2=1.62 $Y2=1.16
r86 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=1.46 $Y=1.16
+ $X2=1.62 $Y2=1.16
r87 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.16
+ $X2=1.46 $Y2=1.16
r88 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.965 $Y2=1.16
r89 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r90 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=0.52 $Y=1.16 $X2=0.94
+ $Y2=1.16
r91 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r92 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=1.19
+ $X2=1.62 $Y2=1.19
r93 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.28 $Y=1.19
+ $X2=0.94 $Y2=1.19
r94 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.28
+ $Y=1.16 $X2=1.28 $Y2=1.16
r95 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=0.965 $Y2=1.16
r96 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=1.055 $Y=1.16
+ $X2=1.28 $Y2=1.16
r97 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.435 $Y2=1.16
r98 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.28 $Y2=1.16
r99 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.69 $Y=1.19
+ $X2=0.94 $Y2=1.19
r100 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.905 $Y=1.295
+ $X2=1.905 $Y2=1.16
r101 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.905 $Y=1.295
+ $X2=1.905 $Y2=1.985
r102 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.16
r103 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r104 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=1.16
r105 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.46 $Y=1.025
+ $X2=1.46 $Y2=0.56
r106 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.16
r107 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=1.435 $Y=1.295
+ $X2=1.435 $Y2=1.985
r108 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r109 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.985
r110 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.16
r111 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r112 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.16
r113 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r114 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.16
r115 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_559_265# 1 2 7 9 10 11 12 14 15 17 19
+ 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c117 20 0 1.10627e-19 $X=4.215 $Y=1.4
r118 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.585 $Y=1.77
+ $X2=5.585 $Y2=1.605
r119 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=1.395
+ $X2=5.505 $Y2=1.23
r120 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.505 $Y=1.395
+ $X2=5.505 $Y2=1.605
r121 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.505 $Y=1.065
+ $X2=5.505 $Y2=1.23
r122 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.505 $Y=1.065
+ $X2=5.505 $Y2=0.825
r123 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=0.7
+ $X2=5.545 $Y2=0.825
r124 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=0.7
+ $X2=5.545 $Y2=0.445
r125 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=4.875 $Y=1.23
+ $X2=4.625 $Y2=1.23
r126 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.875
+ $Y=1.23 $X2=4.875 $Y2=1.23
r127 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=4.535 $Y=1.285
+ $X2=4.625 $Y2=1.23
r128 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=4.535 $Y=1.23
+ $X2=4.875 $Y2=1.23
r129 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.535
+ $Y=1.23 $X2=4.535 $Y2=1.23
r130 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=1.23
+ $X2=5.505 $Y2=1.23
r131 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=5.42 $Y=1.23
+ $X2=4.875 $Y2=1.23
r132 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.535 $Y2=1.285
r133 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=4.305 $Y=1.475
+ $X2=4.305 $Y2=1.965
r134 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.925 $Y=1.4
+ $X2=3.835 $Y2=1.4
r135 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.215 $Y=1.4
+ $X2=4.305 $Y2=1.475
r136 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.215 $Y=1.4
+ $X2=3.925 $Y2=1.4
r137 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=1.475
+ $X2=3.835 $Y2=1.4
r138 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.835 $Y=1.475
+ $X2=3.835 $Y2=1.965
r139 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.455 $Y=1.4
+ $X2=3.365 $Y2=1.4
r140 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.745 $Y=1.4
+ $X2=3.835 $Y2=1.4
r141 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.745 $Y=1.4
+ $X2=3.455 $Y2=1.4
r142 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.475
+ $X2=3.365 $Y2=1.4
r143 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.365 $Y=1.475
+ $X2=3.365 $Y2=1.965
r144 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.275 $Y=1.4
+ $X2=3.365 $Y2=1.4
r145 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.275 $Y=1.4
+ $X2=2.985 $Y2=1.4
r146 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.895 $Y=1.475
+ $X2=2.985 $Y2=1.4
r147 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.895 $Y=1.475
+ $X2=2.895 $Y2=1.965
r148 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.625 $X2=5.585 $Y2=1.77
r149 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.45
+ $Y=0.235 $X2=5.585 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[0] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c115 11 0 1.3204e-19 $X=3.66 $Y=0.255
r116 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.2
+ $Y=1.16 $X2=6.2 $Y2=1.16
r117 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=5.82 $Y=1.55
+ $X2=6.027 $Y2=1.16
r118 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.82 $Y=1.55
+ $X2=5.82 $Y2=2.035
r119 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.795 $Y=0.735
+ $X2=5.795 $Y2=0.445
r120 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.45 $Y=0.81 $X2=5.35
+ $Y2=0.81
r121 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=6.027 $Y2=1.16
r122 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=5.795 $Y2=0.735
r123 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=5.72 $Y=0.81
+ $X2=5.45 $Y2=0.81
r124 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=5.375 $Y=0.735
+ $X2=5.35 $Y2=0.81
r125 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.375 $Y=0.735
+ $X2=5.375 $Y2=0.445
r126 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=5.35 $Y=1.55
+ $X2=5.35 $Y2=2.035
r127 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.35 $Y=1.45 $X2=5.35
+ $Y2=1.55
r128 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.35 $Y=0.885
+ $X2=5.35 $Y2=0.81
r129 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=5.35 $Y=0.885
+ $X2=5.35 $Y2=1.45
r130 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.25 $Y=0.81 $X2=5.35
+ $Y2=0.81
r131 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.25 $Y=0.81
+ $X2=4.915 $Y2=0.81
r132 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.84 $Y=0.735
+ $X2=4.915 $Y2=0.81
r133 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=4.84 $Y=0.255
+ $X2=4.84 $Y2=0.735
r134 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.155 $Y=0.18
+ $X2=4.08 $Y2=0.18
r135 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.765 $Y=0.18
+ $X2=4.84 $Y2=0.255
r136 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.765 $Y=0.18
+ $X2=4.155 $Y2=0.18
r137 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.08 $Y=0.255
+ $X2=4.08 $Y2=0.18
r138 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.08 $Y=0.255
+ $X2=4.08 $Y2=0.59
r139 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.735 $Y=0.18
+ $X2=3.66 $Y2=0.18
r140 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.005 $Y=0.18
+ $X2=4.08 $Y2=0.18
r141 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.005 $Y=0.18
+ $X2=3.735 $Y2=0.18
r142 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.18
r143 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.66 $Y=0.255
+ $X2=3.66 $Y2=0.59
r144 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.315 $Y=0.18
+ $X2=3.24 $Y2=0.18
r145 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.66 $Y2=0.18
r146 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.585 $Y=0.18
+ $X2=3.315 $Y2=0.18
r147 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.24 $Y=0.255
+ $X2=3.24 $Y2=0.18
r148 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.24 $Y=0.255
+ $X2=3.24 $Y2=0.59
r149 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.165 $Y=0.18
+ $X2=3.24 $Y2=0.18
r150 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.165 $Y=0.18
+ $X2=2.895 $Y2=0.18
r151 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.82 $Y=0.255
+ $X2=2.895 $Y2=0.18
r152 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.82 $Y=0.255
+ $X2=2.82 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[1] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c118 30 0 1.3204e-19 $X=9.22 $Y=0.255
r119 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=6.67 $Y=1.16
+ $X2=7.02 $Y2=1.16
r120 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.06 $Y=0.255
+ $X2=10.06 $Y2=0.59
r121 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.715 $Y=0.18
+ $X2=9.64 $Y2=0.18
r122 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=10.06 $Y2=0.255
r123 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=9.715 $Y2=0.18
r124 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.18
r125 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.59
r126 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.295 $Y=0.18
+ $X2=9.22 $Y2=0.18
r127 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.64 $Y2=0.18
r128 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.295 $Y2=0.18
r129 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.18
r130 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.59
r131 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.875 $Y=0.18
+ $X2=8.8 $Y2=0.18
r132 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=9.22 $Y2=0.18
r133 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=8.875 $Y2=0.18
r134 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.8 $Y=0.255
+ $X2=8.8 $Y2=0.18
r135 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.8 $Y=0.255
+ $X2=8.8 $Y2=0.59
r136 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.725 $Y=0.18
+ $X2=8.8 $Y2=0.18
r137 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=8.725 $Y=0.18
+ $X2=8.115 $Y2=0.18
r138 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.04 $Y=0.255
+ $X2=8.115 $Y2=0.18
r139 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=8.04 $Y=0.255
+ $X2=8.04 $Y2=0.735
r140 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.63 $Y=0.81 $X2=7.53
+ $Y2=0.81
r141 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.965 $Y=0.81
+ $X2=8.04 $Y2=0.735
r142 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.965 $Y=0.81
+ $X2=7.63 $Y2=0.81
r143 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.53 $Y=1.55
+ $X2=7.53 $Y2=2.035
r144 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.53 $Y=1.45 $X2=7.53
+ $Y2=1.55
r145 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=7.53 $Y=0.885
+ $X2=7.53 $Y2=0.81
r146 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=7.53 $Y=0.885
+ $X2=7.53 $Y2=1.45
r147 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.505 $Y=0.735
+ $X2=7.53 $Y2=0.81
r148 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.505 $Y=0.735
+ $X2=7.505 $Y2=0.445
r149 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.16 $Y=0.81 $X2=7.06
+ $Y2=0.81
r150 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=7.43 $Y=0.81 $X2=7.53
+ $Y2=0.81
r151 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=7.43 $Y=0.81
+ $X2=7.16 $Y2=0.81
r152 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=7.085 $Y=0.735
+ $X2=7.06 $Y2=0.81
r153 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.085 $Y=0.735
+ $X2=7.085 $Y2=0.445
r154 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=7.06 $Y=1.55
+ $X2=7.06 $Y2=2.035
r155 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=7.06 $Y=1.16
+ $X2=7.06 $Y2=1.55
r156 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.02
+ $Y=1.16 $X2=7.02 $Y2=1.16
r157 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=7.06 $Y=1.16
+ $X2=7.06 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1430_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c116 20 0 1.74242e-19 $X=9.895 $Y=1.4
r117 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=8.345 $Y=1.285
+ $X2=8.255 $Y2=1.23
r118 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.345
+ $Y=1.23 $X2=8.345 $Y2=1.23
r119 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=8.005 $Y=1.23
+ $X2=8.255 $Y2=1.23
r120 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=8.005 $Y=1.23
+ $X2=8.345 $Y2=1.23
r121 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.005
+ $Y=1.23 $X2=8.005 $Y2=1.23
r122 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=1.23
+ $X2=7.375 $Y2=1.23
r123 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=7.46 $Y=1.23
+ $X2=8.005 $Y2=1.23
r124 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=1.395
+ $X2=7.375 $Y2=1.23
r125 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=7.375 $Y=1.395
+ $X2=7.375 $Y2=1.605
r126 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.375 $Y=1.065
+ $X2=7.375 $Y2=1.23
r127 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=7.375 $Y=1.065
+ $X2=7.375 $Y2=0.825
r128 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=7.335 $Y=0.7
+ $X2=7.335 $Y2=0.825
r129 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=0.7
+ $X2=7.335 $Y2=0.445
r130 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.295 $Y=1.77
+ $X2=7.295 $Y2=1.605
r131 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.985 $Y=1.475
+ $X2=9.985 $Y2=1.965
r132 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.605 $Y=1.4
+ $X2=9.515 $Y2=1.4
r133 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=9.895 $Y=1.4
+ $X2=9.985 $Y2=1.475
r134 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.895 $Y=1.4
+ $X2=9.605 $Y2=1.4
r135 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.515 $Y=1.475
+ $X2=9.515 $Y2=1.4
r136 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.515 $Y=1.475
+ $X2=9.515 $Y2=1.965
r137 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.135 $Y=1.4
+ $X2=9.045 $Y2=1.4
r138 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.425 $Y=1.4
+ $X2=9.515 $Y2=1.4
r139 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.425 $Y=1.4
+ $X2=9.135 $Y2=1.4
r140 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.045 $Y=1.475
+ $X2=9.045 $Y2=1.4
r141 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.045 $Y=1.475
+ $X2=9.045 $Y2=1.965
r142 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=8.955 $Y=1.4
+ $X2=9.045 $Y2=1.4
r143 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.955 $Y=1.4
+ $X2=8.665 $Y2=1.4
r144 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.665 $Y2=1.4
r145 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.345 $Y2=1.285
r146 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=8.575 $Y=1.475
+ $X2=8.575 $Y2=1.965
r147 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.15
+ $Y=1.625 $X2=7.295 $Y2=1.77
r148 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.16
+ $Y=0.235 $X2=7.295 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[1] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r86 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=1.16
+ $X2=12.385 $Y2=1.16
r87 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=12.28 $Y=1.16
+ $X2=12.36 $Y2=1.16
r88 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.28
+ $Y=1.16 $X2=12.28 $Y2=1.16
r89 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=11.94 $Y=1.16
+ $X2=12.28 $Y2=1.16
r90 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=1.16
+ $X2=11.94 $Y2=1.16
r91 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.42 $Y=1.16
+ $X2=11.445 $Y2=1.16
r92 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=11.26 $Y=1.16
+ $X2=11.42 $Y2=1.16
r93 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.26
+ $Y=1.16 $X2=11.26 $Y2=1.16
r94 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=11 $Y=1.16 $X2=11.26
+ $Y2=1.16
r95 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=10.975 $Y=1.16
+ $X2=11 $Y2=1.16
r96 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=11.6 $Y=1.19
+ $X2=11.26 $Y2=1.19
r97 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.6
+ $Y=1.16 $X2=11.6 $Y2=1.16
r98 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.535 $Y=1.16
+ $X2=11.445 $Y2=1.16
r99 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=11.535 $Y=1.16
+ $X2=11.6 $Y2=1.16
r100 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=11.825 $Y=1.16
+ $X2=11.915 $Y2=1.16
r101 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=11.825 $Y=1.16
+ $X2=11.6 $Y2=1.16
r102 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=12.19 $Y=1.19
+ $X2=12.28 $Y2=1.19
r103 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.19 $Y=1.19
+ $X2=11.6 $Y2=1.19
r104 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.16
r105 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.985
r106 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=1.16
r107 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=0.56
r108 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=1.16
r109 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=0.56
r110 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.16
r111 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.985
r112 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.445 $Y=1.295
+ $X2=11.445 $Y2=1.16
r113 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.445 $Y=1.295
+ $X2=11.445 $Y2=1.985
r114 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.42 $Y=1.025
+ $X2=11.42 $Y2=1.16
r115 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.42 $Y=1.025
+ $X2=11.42 $Y2=0.56
r116 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11 $Y=1.025 $X2=11
+ $Y2=1.16
r117 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11 $Y=1.025 $X2=11
+ $Y2=0.56
r118 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.975 $Y=1.295
+ $X2=10.975 $Y2=1.16
r119 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=10.975 $Y=1.295
+ $X2=10.975 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[2] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
r88 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.76 $Y=1.16
+ $X2=14.785 $Y2=1.16
r89 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=14.5 $Y=1.16
+ $X2=14.76 $Y2=1.16
r90 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.5
+ $Y=1.16 $X2=14.5 $Y2=1.16
r91 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=14.34 $Y=1.16
+ $X2=14.5 $Y2=1.16
r92 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=14.315 $Y=1.16
+ $X2=14.34 $Y2=1.16
r93 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=1.16
+ $X2=13.845 $Y2=1.16
r94 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13.82
+ $Y=1.16 $X2=13.82 $Y2=1.16
r95 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=13.4 $Y=1.16
+ $X2=13.82 $Y2=1.16
r96 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=1.16
+ $X2=13.4 $Y2=1.16
r97 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=1.19
+ $X2=14.5 $Y2=1.19
r98 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=14.16 $Y=1.19
+ $X2=13.82 $Y2=1.19
r99 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.16
+ $Y=1.16 $X2=14.16 $Y2=1.16
r100 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=13.935 $Y=1.16
+ $X2=13.845 $Y2=1.16
r101 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=13.935 $Y=1.16
+ $X2=14.16 $Y2=1.16
r102 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=14.225 $Y=1.16
+ $X2=14.315 $Y2=1.16
r103 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=14.225 $Y=1.16
+ $X2=14.16 $Y2=1.16
r104 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.57 $Y=1.19
+ $X2=13.82 $Y2=1.19
r105 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.785 $Y=1.295
+ $X2=14.785 $Y2=1.16
r106 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.785 $Y=1.295
+ $X2=14.785 $Y2=1.985
r107 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.76 $Y=1.025
+ $X2=14.76 $Y2=1.16
r108 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.76 $Y=1.025
+ $X2=14.76 $Y2=0.56
r109 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.34 $Y=1.025
+ $X2=14.34 $Y2=1.16
r110 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=14.34 $Y=1.025
+ $X2=14.34 $Y2=0.56
r111 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.315 $Y=1.295
+ $X2=14.315 $Y2=1.16
r112 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=14.315 $Y=1.295
+ $X2=14.315 $Y2=1.985
r113 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.16
r114 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.985
r115 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=1.16
r116 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=0.56
r117 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=1.16
r118 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=0.56
r119 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.16
r120 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_3135_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c119 20 0 1.10627e-19 $X=17.095 $Y=1.4
c120 11 0 1.74242e-19 $X=15.865 $Y=1.4
r121 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=1.77
+ $X2=18.465 $Y2=1.605
r122 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=1.395
+ $X2=18.385 $Y2=1.23
r123 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=18.385 $Y=1.395
+ $X2=18.385 $Y2=1.605
r124 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.385 $Y=1.065
+ $X2=18.385 $Y2=1.23
r125 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=18.385 $Y=1.065
+ $X2=18.385 $Y2=0.825
r126 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=18.425 $Y=0.7
+ $X2=18.425 $Y2=0.825
r127 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=18.425 $Y=0.7
+ $X2=18.425 $Y2=0.445
r128 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=17.755 $Y=1.23
+ $X2=17.505 $Y2=1.23
r129 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.755
+ $Y=1.23 $X2=17.755 $Y2=1.23
r130 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=17.415
+ $Y=1.285 $X2=17.505 $Y2=1.23
r131 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=17.415 $Y=1.23
+ $X2=17.755 $Y2=1.23
r132 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.415
+ $Y=1.23 $X2=17.415 $Y2=1.23
r133 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.3 $Y=1.23
+ $X2=18.385 $Y2=1.23
r134 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=18.3 $Y=1.23
+ $X2=17.755 $Y2=1.23
r135 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=17.185
+ $Y=1.475 $X2=17.415 $Y2=1.285
r136 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=17.185 $Y=1.475
+ $X2=17.185 $Y2=1.965
r137 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.805 $Y=1.4
+ $X2=16.715 $Y2=1.4
r138 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.095 $Y=1.4
+ $X2=17.185 $Y2=1.475
r139 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.095 $Y=1.4
+ $X2=16.805 $Y2=1.4
r140 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.715 $Y=1.475
+ $X2=16.715 $Y2=1.4
r141 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.715 $Y=1.475
+ $X2=16.715 $Y2=1.965
r142 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.335 $Y=1.4
+ $X2=16.245 $Y2=1.4
r143 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.625 $Y=1.4
+ $X2=16.715 $Y2=1.4
r144 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.625 $Y=1.4
+ $X2=16.335 $Y2=1.4
r145 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=16.245 $Y=1.475
+ $X2=16.245 $Y2=1.4
r146 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=16.245 $Y=1.475
+ $X2=16.245 $Y2=1.965
r147 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=16.155 $Y=1.4
+ $X2=16.245 $Y2=1.4
r148 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=16.155 $Y=1.4
+ $X2=15.865 $Y2=1.4
r149 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=15.775 $Y=1.475
+ $X2=15.865 $Y2=1.4
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.775 $Y=1.475
+ $X2=15.775 $Y2=1.965
r151 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.32
+ $Y=1.625 $X2=18.465 $Y2=1.77
r152 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.33
+ $Y=0.235 $X2=18.465 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[2] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c115 11 0 1.3204e-19 $X=16.54 $Y=0.255
r116 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.08
+ $Y=1.16 $X2=19.08 $Y2=1.16
r117 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=18.7 $Y=1.55
+ $X2=18.907 $Y2=1.16
r118 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.7 $Y=1.55
+ $X2=18.7 $Y2=2.035
r119 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.675 $Y=0.735
+ $X2=18.675 $Y2=0.445
r120 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.33 $Y=0.81
+ $X2=18.23 $Y2=0.81
r121 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.907 $Y2=1.16
r122 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.675 $Y2=0.735
r123 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=18.6 $Y=0.81
+ $X2=18.33 $Y2=0.81
r124 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=18.255 $Y=0.735
+ $X2=18.23 $Y2=0.81
r125 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=18.255 $Y=0.735
+ $X2=18.255 $Y2=0.445
r126 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=18.23 $Y=1.55
+ $X2=18.23 $Y2=2.035
r127 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=18.23 $Y=1.45 $X2=18.23
+ $Y2=1.55
r128 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=18.23 $Y=0.885
+ $X2=18.23 $Y2=0.81
r129 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=18.23 $Y=0.885
+ $X2=18.23 $Y2=1.45
r130 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=18.13 $Y=0.81
+ $X2=18.23 $Y2=0.81
r131 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=18.13 $Y=0.81
+ $X2=17.795 $Y2=0.81
r132 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.72 $Y=0.735
+ $X2=17.795 $Y2=0.81
r133 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=17.72 $Y=0.255
+ $X2=17.72 $Y2=0.735
r134 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.035 $Y=0.18
+ $X2=16.96 $Y2=0.18
r135 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.645 $Y=0.18
+ $X2=17.72 $Y2=0.255
r136 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=17.645 $Y=0.18
+ $X2=17.035 $Y2=0.18
r137 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.96 $Y=0.255
+ $X2=16.96 $Y2=0.18
r138 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.96 $Y=0.255
+ $X2=16.96 $Y2=0.59
r139 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.615 $Y=0.18
+ $X2=16.54 $Y2=0.18
r140 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.885 $Y=0.18
+ $X2=16.96 $Y2=0.18
r141 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.885 $Y=0.18
+ $X2=16.615 $Y2=0.18
r142 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.54 $Y=0.255
+ $X2=16.54 $Y2=0.18
r143 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.54 $Y=0.255
+ $X2=16.54 $Y2=0.59
r144 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.195 $Y=0.18
+ $X2=16.12 $Y2=0.18
r145 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.465 $Y=0.18
+ $X2=16.54 $Y2=0.18
r146 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.465 $Y=0.18
+ $X2=16.195 $Y2=0.18
r147 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.12 $Y=0.255
+ $X2=16.12 $Y2=0.18
r148 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.12 $Y=0.255
+ $X2=16.12 $Y2=0.59
r149 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=16.045 $Y=0.18
+ $X2=16.12 $Y2=0.18
r150 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=16.045 $Y=0.18
+ $X2=15.775 $Y2=0.18
r151 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.7 $Y=0.255
+ $X2=15.775 $Y2=0.18
r152 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.7 $Y=0.255
+ $X2=15.7 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%S[3] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c118 30 0 1.3204e-19 $X=22.1 $Y=0.255
r119 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=19.55 $Y=1.16
+ $X2=19.9 $Y2=1.16
r120 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.94 $Y=0.255
+ $X2=22.94 $Y2=0.59
r121 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.595 $Y=0.18
+ $X2=22.52 $Y2=0.18
r122 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=22.865 $Y=0.18
+ $X2=22.94 $Y2=0.255
r123 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.865 $Y=0.18
+ $X2=22.595 $Y2=0.18
r124 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.52 $Y=0.255
+ $X2=22.52 $Y2=0.18
r125 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.52 $Y=0.255
+ $X2=22.52 $Y2=0.59
r126 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.175 $Y=0.18
+ $X2=22.1 $Y2=0.18
r127 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.445 $Y=0.18
+ $X2=22.52 $Y2=0.18
r128 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.445 $Y=0.18
+ $X2=22.175 $Y2=0.18
r129 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.1 $Y=0.255
+ $X2=22.1 $Y2=0.18
r130 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.1 $Y=0.255
+ $X2=22.1 $Y2=0.59
r131 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.755 $Y=0.18
+ $X2=21.68 $Y2=0.18
r132 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.025 $Y=0.18
+ $X2=22.1 $Y2=0.18
r133 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.025 $Y=0.18
+ $X2=21.755 $Y2=0.18
r134 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.68 $Y=0.255
+ $X2=21.68 $Y2=0.18
r135 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.68 $Y=0.255
+ $X2=21.68 $Y2=0.59
r136 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.605 $Y=0.18
+ $X2=21.68 $Y2=0.18
r137 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=21.605 $Y=0.18
+ $X2=20.995 $Y2=0.18
r138 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.92 $Y=0.255
+ $X2=20.995 $Y2=0.18
r139 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=20.92 $Y=0.255
+ $X2=20.92 $Y2=0.735
r140 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.51 $Y=0.81
+ $X2=20.41 $Y2=0.81
r141 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.845 $Y=0.81
+ $X2=20.92 $Y2=0.735
r142 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=20.845 $Y=0.81
+ $X2=20.51 $Y2=0.81
r143 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=20.41 $Y=1.55
+ $X2=20.41 $Y2=2.035
r144 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=20.41 $Y=1.45 $X2=20.41
+ $Y2=1.55
r145 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=20.41 $Y=0.885
+ $X2=20.41 $Y2=0.81
r146 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=20.41 $Y=0.885
+ $X2=20.41 $Y2=1.45
r147 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=20.385 $Y=0.735
+ $X2=20.41 $Y2=0.81
r148 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=20.385 $Y=0.735
+ $X2=20.385 $Y2=0.445
r149 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.04 $Y=0.81
+ $X2=19.94 $Y2=0.81
r150 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=20.31 $Y=0.81
+ $X2=20.41 $Y2=0.81
r151 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=20.31 $Y=0.81
+ $X2=20.04 $Y2=0.81
r152 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=19.965 $Y=0.735
+ $X2=19.94 $Y2=0.81
r153 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=19.965 $Y=0.735
+ $X2=19.965 $Y2=0.445
r154 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=19.94 $Y=1.55
+ $X2=19.94 $Y2=2.035
r155 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=19.94 $Y=1.16
+ $X2=19.94 $Y2=1.55
r156 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.9
+ $Y=1.16 $X2=19.9 $Y2=1.16
r157 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=19.94 $Y=1.16
+ $X2=19.94 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4006_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
r114 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=21.225
+ $Y=1.285 $X2=21.135 $Y2=1.23
r115 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.225
+ $Y=1.23 $X2=21.225 $Y2=1.23
r116 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=20.885 $Y=1.23
+ $X2=21.135 $Y2=1.23
r117 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=20.885 $Y=1.23
+ $X2=21.225 $Y2=1.23
r118 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.885
+ $Y=1.23 $X2=20.885 $Y2=1.23
r119 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.34 $Y=1.23
+ $X2=20.255 $Y2=1.23
r120 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=20.34 $Y=1.23
+ $X2=20.885 $Y2=1.23
r121 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=1.395
+ $X2=20.255 $Y2=1.23
r122 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=20.255 $Y=1.395
+ $X2=20.255 $Y2=1.605
r123 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.255 $Y=1.065
+ $X2=20.255 $Y2=1.23
r124 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=20.255 $Y=1.065
+ $X2=20.255 $Y2=0.825
r125 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=20.215 $Y=0.7
+ $X2=20.215 $Y2=0.825
r126 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=20.215 $Y=0.7
+ $X2=20.215 $Y2=0.445
r127 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.175 $Y=1.77
+ $X2=20.175 $Y2=1.605
r128 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.865 $Y=1.475
+ $X2=22.865 $Y2=1.965
r129 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.485 $Y=1.4
+ $X2=22.395 $Y2=1.4
r130 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=22.775 $Y=1.4
+ $X2=22.865 $Y2=1.475
r131 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.775 $Y=1.4
+ $X2=22.485 $Y2=1.4
r132 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=22.395 $Y=1.475
+ $X2=22.395 $Y2=1.4
r133 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.395 $Y=1.475
+ $X2=22.395 $Y2=1.965
r134 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.015 $Y=1.4
+ $X2=21.925 $Y2=1.4
r135 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.305 $Y=1.4
+ $X2=22.395 $Y2=1.4
r136 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.305 $Y=1.4
+ $X2=22.015 $Y2=1.4
r137 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=21.925 $Y=1.475
+ $X2=21.925 $Y2=1.4
r138 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.925 $Y=1.475
+ $X2=21.925 $Y2=1.965
r139 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.835 $Y=1.4
+ $X2=21.925 $Y2=1.4
r140 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.835 $Y=1.4
+ $X2=21.545 $Y2=1.4
r141 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.545 $Y2=1.4
r142 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.225 $Y2=1.285
r143 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.455 $Y=1.475
+ $X2=21.455 $Y2=1.965
r144 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.03
+ $Y=1.625 $X2=20.175 $Y2=1.77
r145 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.04
+ $Y=0.235 $X2=20.175 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%D[3] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
r81 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=1.16
+ $X2=25.265 $Y2=1.16
r82 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=25.16 $Y=1.16
+ $X2=25.24 $Y2=1.16
r83 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=25.16
+ $Y=1.16 $X2=25.16 $Y2=1.16
r84 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=24.82 $Y=1.16
+ $X2=25.16 $Y2=1.16
r85 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=1.16
+ $X2=24.82 $Y2=1.16
r86 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.3 $Y=1.16
+ $X2=24.325 $Y2=1.16
r87 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=24.14 $Y=1.16
+ $X2=24.3 $Y2=1.16
r88 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.14
+ $Y=1.16 $X2=24.14 $Y2=1.16
r89 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=23.88 $Y=1.16
+ $X2=24.14 $Y2=1.16
r90 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=23.855 $Y=1.16
+ $X2=23.88 $Y2=1.16
r91 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=24.48 $Y=1.19
+ $X2=24.14 $Y2=1.19
r92 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=24.48
+ $Y=1.16 $X2=24.48 $Y2=1.16
r93 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.415 $Y=1.16
+ $X2=24.325 $Y2=1.16
r94 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=24.415 $Y=1.16
+ $X2=24.48 $Y2=1.16
r95 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=24.705 $Y=1.16
+ $X2=24.795 $Y2=1.16
r96 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=24.705 $Y=1.16
+ $X2=24.48 $Y2=1.16
r97 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=25.07 $Y=1.19
+ $X2=25.16 $Y2=1.19
r98 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=25.07 $Y=1.19
+ $X2=24.48 $Y2=1.19
r99 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.16
r100 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.985
r101 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=1.16
r102 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=0.56
r103 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=1.16
r104 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=0.56
r105 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.16
r106 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.985
r107 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.325 $Y=1.295
+ $X2=24.325 $Y2=1.16
r108 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.325 $Y=1.295
+ $X2=24.325 $Y2=1.985
r109 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.3 $Y=1.025
+ $X2=24.3 $Y2=1.16
r110 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.3 $Y=1.025
+ $X2=24.3 $Y2=0.56
r111 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=23.88 $Y=1.025
+ $X2=23.88 $Y2=1.16
r112 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=23.88 $Y=1.025
+ $X2=23.88 $Y2=0.56
r113 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.855 $Y=1.295
+ $X2=23.855 $Y2=1.16
r114 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=23.855 $Y=1.295
+ $X2=23.855 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 61 63 69 71 75 79 83 85 89 93 97 101 105 109 113 119 121 125
+ 129 133 135 139 143 147 151 153 155 160 161 162 163 165 166 168 169 171 172
+ 173 174 176 177 179 180 181 182 183 184 189 214 218 223 248 252 261 264 267
+ 270 273 276 279 282 285 288
r346 288 289 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=2.72
+ $X2=24.61 $Y2=2.72
r347 285 286 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=2.72
+ $X2=19.55 $Y2=2.72
r348 282 283 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r349 280 283 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=14.95 $Y2=2.72
r350 279 280 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r351 270 271 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r352 267 268 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r353 264 265 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r354 262 265 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r355 261 262 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r356 256 289 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.07 $Y=2.72
+ $X2=24.61 $Y2=2.72
r357 255 256 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=2.72
+ $X2=25.07 $Y2=2.72
r358 253 288 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.695 $Y=2.72
+ $X2=24.56 $Y2=2.72
r359 253 255 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=24.695 $Y=2.72
+ $X2=25.07 $Y2=2.72
r360 252 291 4.17176 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=25.365 $Y=2.72
+ $X2=25.562 $Y2=2.72
r361 252 255 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.365 $Y=2.72
+ $X2=25.07 $Y2=2.72
r362 251 289 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=2.72
+ $X2=24.61 $Y2=2.72
r363 250 251 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=2.72
+ $X2=24.15 $Y2=2.72
r364 248 288 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.425 $Y=2.72
+ $X2=24.56 $Y2=2.72
r365 248 250 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=24.425 $Y=2.72
+ $X2=24.15 $Y2=2.72
r366 247 251 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=2.72
+ $X2=24.15 $Y2=2.72
r367 246 247 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=2.72
+ $X2=23.23 $Y2=2.72
r368 244 247 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=2.72
+ $X2=23.23 $Y2=2.72
r369 243 246 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=2.72
+ $X2=23.23 $Y2=2.72
r370 243 244 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=2.72
+ $X2=20.93 $Y2=2.72
r371 241 244 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=20.93 $Y2=2.72
r372 241 286 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=19.55 $Y2=2.72
r373 240 241 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=2.72
+ $X2=20.47 $Y2=2.72
r374 238 285 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.84 $Y=2.72
+ $X2=19.69 $Y2=2.72
r375 238 240 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=19.84 $Y=2.72
+ $X2=20.47 $Y2=2.72
r376 237 286 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=18.63 $Y=2.72
+ $X2=19.55 $Y2=2.72
r377 236 237 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=2.72
+ $X2=18.63 $Y2=2.72
r378 234 237 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.71 $Y=2.72
+ $X2=18.63 $Y2=2.72
r379 233 234 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=17.71 $Y=2.72
+ $X2=17.71 $Y2=2.72
r380 231 234 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=17.71 $Y2=2.72
r381 231 283 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=14.95 $Y2=2.72
r382 230 233 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=15.41 $Y=2.72
+ $X2=17.71 $Y2=2.72
r383 230 231 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r384 228 282 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.155 $Y=2.72
+ $X2=15.02 $Y2=2.72
r385 228 230 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=15.155 $Y=2.72
+ $X2=15.41 $Y2=2.72
r386 227 280 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r387 226 227 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r388 224 276 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.275 $Y=2.72
+ $X2=13.14 $Y2=2.72
r389 224 226 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.275 $Y=2.72
+ $X2=13.57 $Y2=2.72
r390 223 279 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.945 $Y=2.72
+ $X2=14.08 $Y2=2.72
r391 223 226 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.945 $Y=2.72
+ $X2=13.57 $Y2=2.72
r392 222 271 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=2.72
+ $X2=11.73 $Y2=2.72
r393 221 222 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r394 219 270 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=11.68 $Y2=2.72
r395 219 221 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=2.72
+ $X2=12.19 $Y2=2.72
r396 218 273 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.485 $Y=2.72
+ $X2=12.62 $Y2=2.72
r397 218 221 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.485 $Y=2.72
+ $X2=12.19 $Y2=2.72
r398 217 271 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r399 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r400 214 270 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.545 $Y=2.72
+ $X2=11.68 $Y2=2.72
r401 214 216 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.545 $Y=2.72
+ $X2=11.27 $Y2=2.72
r402 213 217 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r403 212 213 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r404 210 213 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r405 209 212 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=10.35 $Y2=2.72
r406 209 210 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r407 207 210 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r408 207 268 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r409 206 207 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r410 204 267 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=6.81 $Y2=2.72
r411 204 206 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.96 $Y=2.72
+ $X2=7.59 $Y2=2.72
r412 203 268 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r413 202 203 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r414 200 203 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r415 199 200 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r416 197 200 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r417 197 265 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r418 196 199 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r419 196 197 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r420 194 264 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r421 194 196 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.53 $Y2=2.72
r422 193 262 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r423 192 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r424 190 258 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r425 190 192 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r426 189 261 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r427 189 192 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r428 184 256 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=2.72
+ $X2=25.07 $Y2=2.72
r429 184 291 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=2.72
+ $X2=25.53 $Y2=2.72
r430 183 227 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r431 183 276 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r432 182 183 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r433 182 222 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r434 182 273 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r435 181 193 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r436 181 258 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r437 179 246 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=23.485 $Y=2.72
+ $X2=23.23 $Y2=2.72
r438 179 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=23.485 $Y=2.72
+ $X2=23.62 $Y2=2.72
r439 178 250 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=23.755 $Y=2.72
+ $X2=24.15 $Y2=2.72
r440 178 180 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=23.755 $Y=2.72
+ $X2=23.62 $Y2=2.72
r441 176 240 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=20.535 $Y=2.72
+ $X2=20.47 $Y2=2.72
r442 176 177 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=20.535 $Y=2.72
+ $X2=20.672 $Y2=2.72
r443 175 243 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=20.81 $Y=2.72
+ $X2=20.93 $Y2=2.72
r444 175 177 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=20.81 $Y=2.72
+ $X2=20.672 $Y2=2.72
r445 173 236 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=18.8 $Y=2.72
+ $X2=18.63 $Y2=2.72
r446 173 174 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.8 $Y=2.72
+ $X2=18.95 $Y2=2.72
r447 171 233 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=17.83 $Y=2.72
+ $X2=17.71 $Y2=2.72
r448 171 172 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=17.83 $Y=2.72
+ $X2=17.967 $Y2=2.72
r449 170 236 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=18.105 $Y=2.72
+ $X2=18.63 $Y2=2.72
r450 170 172 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=18.105 $Y=2.72
+ $X2=17.967 $Y2=2.72
r451 168 212 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.605 $Y=2.72
+ $X2=10.35 $Y2=2.72
r452 168 169 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.605 $Y=2.72
+ $X2=10.74 $Y2=2.72
r453 167 216 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=11.27 $Y2=2.72
r454 167 169 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.875 $Y=2.72
+ $X2=10.74 $Y2=2.72
r455 165 206 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.655 $Y=2.72
+ $X2=7.59 $Y2=2.72
r456 165 166 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=7.655 $Y=2.72
+ $X2=7.792 $Y2=2.72
r457 164 209 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.93 $Y=2.72
+ $X2=8.05 $Y2=2.72
r458 164 166 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=7.93 $Y=2.72
+ $X2=7.792 $Y2=2.72
r459 162 202 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=5.75 $Y2=2.72
r460 162 163 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.92 $Y=2.72
+ $X2=6.07 $Y2=2.72
r461 160 199 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=4.83 $Y2=2.72
r462 160 161 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=4.95 $Y=2.72
+ $X2=5.087 $Y2=2.72
r463 159 202 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.75 $Y2=2.72
r464 159 161 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.087 $Y2=2.72
r465 155 158 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=25.5 $Y=1.66
+ $X2=25.5 $Y2=2.34
r466 153 291 3.11294 $w=2.7e-07 $l=1.11781e-07 $layer=LI1_cond $X=25.5 $Y=2.635
+ $X2=25.562 $Y2=2.72
r467 153 158 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.5 $Y=2.635
+ $X2=25.5 $Y2=2.34
r468 149 288 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=2.635
+ $X2=24.56 $Y2=2.72
r469 149 151 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=24.56 $Y=2.635
+ $X2=24.56 $Y2=2
r470 145 180 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=23.62 $Y=2.635
+ $X2=23.62 $Y2=2.72
r471 145 147 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=23.62 $Y=2.635
+ $X2=23.62 $Y2=2
r472 141 177 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=20.672 $Y=2.635
+ $X2=20.672 $Y2=2.72
r473 141 143 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=20.672 $Y=2.635
+ $X2=20.672 $Y2=1.77
r474 137 285 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.69 $Y=2.635
+ $X2=19.69 $Y2=2.72
r475 137 139 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=19.69 $Y=2.635
+ $X2=19.69 $Y2=1.77
r476 136 174 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.1 $Y=2.72
+ $X2=18.95 $Y2=2.72
r477 135 285 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.54 $Y=2.72
+ $X2=19.69 $Y2=2.72
r478 135 136 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=19.54 $Y=2.72
+ $X2=19.1 $Y2=2.72
r479 131 174 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.95 $Y=2.635
+ $X2=18.95 $Y2=2.72
r480 131 133 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=18.95 $Y=2.635
+ $X2=18.95 $Y2=1.77
r481 127 172 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=17.967 $Y=2.635
+ $X2=17.967 $Y2=2.72
r482 127 129 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=17.967 $Y=2.635
+ $X2=17.967 $Y2=1.77
r483 123 282 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.02 $Y=2.635
+ $X2=15.02 $Y2=2.72
r484 123 125 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=15.02 $Y=2.635
+ $X2=15.02 $Y2=2
r485 122 279 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.215 $Y=2.72
+ $X2=14.08 $Y2=2.72
r486 121 282 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=15.02 $Y2=2.72
r487 121 122 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=14.215 $Y2=2.72
r488 117 279 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=2.635
+ $X2=14.08 $Y2=2.72
r489 117 119 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.08 $Y=2.635
+ $X2=14.08 $Y2=2
r490 113 116 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.14 $Y=1.66
+ $X2=13.14 $Y2=2.34
r491 111 276 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.14 $Y=2.635
+ $X2=13.14 $Y2=2.72
r492 111 116 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.14 $Y=2.635
+ $X2=13.14 $Y2=2.34
r493 110 273 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.755 $Y=2.72
+ $X2=12.62 $Y2=2.72
r494 109 276 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.005 $Y=2.72
+ $X2=13.14 $Y2=2.72
r495 109 110 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=13.005 $Y=2.72
+ $X2=12.755 $Y2=2.72
r496 105 108 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=12.62 $Y=1.66
+ $X2=12.62 $Y2=2.34
r497 103 273 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.62 $Y=2.635
+ $X2=12.62 $Y2=2.72
r498 103 108 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.62 $Y=2.635
+ $X2=12.62 $Y2=2.34
r499 99 270 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=2.635
+ $X2=11.68 $Y2=2.72
r500 99 101 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.68 $Y=2.635
+ $X2=11.68 $Y2=2
r501 95 169 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.74 $Y=2.635
+ $X2=10.74 $Y2=2.72
r502 95 97 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.74 $Y=2.635
+ $X2=10.74 $Y2=2
r503 91 166 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=7.792 $Y=2.635
+ $X2=7.792 $Y2=2.72
r504 91 93 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=7.792 $Y=2.635
+ $X2=7.792 $Y2=1.77
r505 87 267 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.81 $Y=2.635
+ $X2=6.81 $Y2=2.72
r506 87 89 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=6.81 $Y=2.635
+ $X2=6.81 $Y2=1.77
r507 86 163 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.22 $Y=2.72
+ $X2=6.07 $Y2=2.72
r508 85 267 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.66 $Y=2.72
+ $X2=6.81 $Y2=2.72
r509 85 86 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=6.66 $Y=2.72
+ $X2=6.22 $Y2=2.72
r510 81 163 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=2.635
+ $X2=6.07 $Y2=2.72
r511 81 83 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=6.07 $Y=2.635
+ $X2=6.07 $Y2=1.77
r512 77 161 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=2.72
r513 77 79 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=5.087 $Y=2.635
+ $X2=5.087 $Y2=1.77
r514 73 264 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r515 73 75 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r516 72 261 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r517 71 264 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r518 71 72 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r519 67 261 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r520 67 69 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r521 63 66 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r522 61 258 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.197 $Y2=2.72
r523 61 66 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r524 20 158 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=2.34
r525 20 155 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=1.66
r526 19 151 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=24.415
+ $Y=1.485 $X2=24.56 $Y2=2
r527 18 147 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=23.495
+ $Y=1.485 $X2=23.62 $Y2=2
r528 17 143 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.5
+ $Y=1.625 $X2=20.645 $Y2=1.77
r529 16 139 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=19.58
+ $Y=1.625 $X2=19.705 $Y2=1.77
r530 15 133 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=18.79
+ $Y=1.625 $X2=18.935 $Y2=1.77
r531 14 129 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=17.87
+ $Y=1.625 $X2=17.995 $Y2=1.77
r532 13 125 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=14.875
+ $Y=1.485 $X2=15.02 $Y2=2
r533 12 119 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=13.935
+ $Y=1.485 $X2=14.08 $Y2=2
r534 11 116 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=2.34
r535 11 113 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=1.66
r536 10 108 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=2.34
r537 10 105 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=1.66
r538 9 101 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.535
+ $Y=1.485 $X2=11.68 $Y2=2
r539 8 97 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=10.615
+ $Y=1.485 $X2=10.74 $Y2=2
r540 7 93 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.62
+ $Y=1.625 $X2=7.765 $Y2=1.77
r541 6 89 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=6.7
+ $Y=1.625 $X2=6.825 $Y2=1.77
r542 5 83 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.625 $X2=6.055 $Y2=1.77
r543 4 79 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=1.625 $X2=5.115 $Y2=1.77
r544 3 75 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r545 2 69 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r546 1 66 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r547 1 63 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_117_297# 1 2 3 4 5 16 18 20 24 26 31
+ 32 33 36 38 42 47 48
c89 36 0 1.3204e-19 $X=3.6 $Y=1.7
r90 40 42 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=4.555 $Y=2.295
+ $X2=4.555 $Y2=1.73
r91 39 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=2.38
+ $X2=3.6 $Y2=2.38
r92 38 40 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=4.405 $Y=2.38
+ $X2=4.555 $Y2=2.295
r93 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.405 $Y=2.38
+ $X2=3.735 $Y2=2.38
r94 34 48 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.295 $X2=3.6
+ $Y2=2.38
r95 34 36 25.3964 $w=2.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.6 $Y=2.295
+ $X2=3.6 $Y2=1.7
r96 32 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=2.38
+ $X2=3.6 $Y2=2.38
r97 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.465 $Y=2.38
+ $X2=2.795 $Y2=2.38
r98 29 33 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.645 $Y=2.295
+ $X2=2.795 $Y2=2.38
r99 29 31 22.8568 $w=2.98e-07 $l=5.95e-07 $layer=LI1_cond $X=2.645 $Y=2.295
+ $X2=2.645 $Y2=1.7
r100 28 31 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=2.645 $Y=1.665
+ $X2=2.645 $Y2=1.7
r101 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r102 26 28 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=2.645 $Y2=1.665
r103 26 27 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.495 $Y=1.58
+ $X2=1.835 $Y2=1.58
r104 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r105 22 24 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.34
r106 21 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r107 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r108 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r109 16 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r110 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.34
r111 5 42 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=4.395
+ $Y=1.555 $X2=4.54 $Y2=1.73
r112 4 36 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.555 $X2=3.6 $Y2=1.7
r113 3 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.555 $X2=2.66 $Y2=1.7
r114 2 47 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r115 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r116 1 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r117 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 50 51 55 59 61 64 66 67 71 75 77 80 82 86 88 90 92 94 98 102 104 106 108
+ 110 113 114 115 116 117 118 119 123 127 129 132 133 134 135 136 147 152 157
+ 162 165 168 173 178 181
c416 115 0 3.48484e-19 $X=15.865 $Y=1.87
c417 106 0 1.20815e-19 $X=21.79 $Y=1.215
c418 104 0 1.20815e-19 $X=16.85 $Y=1.215
c419 90 0 1.20815e-19 $X=8.91 $Y=1.215
c420 88 0 1.20815e-19 $X=3.97 $Y=1.215
r421 136 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.69 $Y=1.87
+ $X2=21.69 $Y2=1.87
r422 135 168 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.95 $Y=1.87
+ $X2=16.95 $Y2=1.87
r423 134 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.81 $Y=1.87
+ $X2=8.81 $Y2=1.87
r424 133 181 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=3.925 $Y=1.87
+ $X2=3.275 $Y2=1.87
r425 133 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=1.87
+ $X2=4.07 $Y2=1.87
r426 132 181 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.13 $Y=1.87
+ $X2=3.275 $Y2=1.87
r427 132 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.13 $Y=1.87
+ $X2=3.13 $Y2=1.87
r428 129 178 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.63 $Y=1.87
+ $X2=22.63 $Y2=1.87
r429 127 136 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=22.485 $Y=1.87
+ $X2=21.835 $Y2=1.87
r430 127 129 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.485 $Y=1.87
+ $X2=22.63 $Y2=1.87
r431 125 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.01 $Y=1.87
+ $X2=16.01 $Y2=1.87
r432 123 135 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=16.155 $Y=1.87
+ $X2=16.805 $Y2=1.87
r433 123 125 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.155 $Y=1.87
+ $X2=16.01 $Y2=1.87
r434 121 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.75 $Y=1.87
+ $X2=9.75 $Y2=1.87
r435 119 134 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=9.605 $Y=1.87
+ $X2=8.955 $Y2=1.87
r436 119 121 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.605 $Y=1.87
+ $X2=9.75 $Y2=1.87
r437 118 135 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=17.095 $Y=1.87
+ $X2=16.89 $Y2=1.87
r438 117 136 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.545 $Y=1.87
+ $X2=21.69 $Y2=1.87
r439 117 118 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=21.545 $Y=1.87
+ $X2=17.095 $Y2=1.87
r440 116 121 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.895 $Y=1.87
+ $X2=9.75 $Y2=1.87
r441 115 125 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.865 $Y=1.87
+ $X2=16.01 $Y2=1.87
r442 115 116 7.3886 $w=1.4e-07 $l=5.97e-06 $layer=MET1_cond $X=15.865 $Y=1.87
+ $X2=9.895 $Y2=1.87
r443 114 133 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=4.215 $Y=1.87
+ $X2=4.01 $Y2=1.87
r444 113 134 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.665 $Y=1.87
+ $X2=8.81 $Y2=1.87
r445 113 114 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=8.665 $Y=1.87
+ $X2=4.215 $Y2=1.87
r446 110 112 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=22.73 $Y=0.68
+ $X2=22.73 $Y2=0.885
r447 107 178 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=22.63 $Y=1.365
+ $X2=22.63 $Y2=1.7
r448 107 108 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=22.63 $Y=1.365
+ $X2=22.63 $Y2=1.215
r449 105 173 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=21.69 $Y=1.365
+ $X2=21.69 $Y2=1.7
r450 105 106 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.69 $Y=1.365
+ $X2=21.79 $Y2=1.215
r451 103 168 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=16.95 $Y=1.365
+ $X2=16.95 $Y2=1.7
r452 103 104 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.95 $Y=1.365
+ $X2=16.85 $Y2=1.215
r453 101 165 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=16.01 $Y=1.365
+ $X2=16.01 $Y2=1.7
r454 101 102 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=16.01 $Y=1.365
+ $X2=16.01 $Y2=1.215
r455 98 100 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.91 $Y=0.68
+ $X2=15.91 $Y2=0.885
r456 94 96 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.85 $Y=0.68
+ $X2=9.85 $Y2=0.885
r457 91 162 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.75 $Y=1.365
+ $X2=9.75 $Y2=1.7
r458 91 92 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=9.75 $Y=1.365
+ $X2=9.75 $Y2=1.215
r459 89 157 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.81 $Y=1.365
+ $X2=8.81 $Y2=1.7
r460 89 90 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=8.81 $Y=1.365
+ $X2=8.91 $Y2=1.215
r461 87 152 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.07 $Y=1.365
+ $X2=4.07 $Y2=1.7
r462 87 88 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=4.07 $Y=1.365
+ $X2=3.97 $Y2=1.215
r463 85 147 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.13 $Y=1.365
+ $X2=3.13 $Y2=1.7
r464 85 86 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.13 $Y=1.365
+ $X2=3.13 $Y2=1.215
r465 82 84 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.03 $Y=0.68
+ $X2=3.03 $Y2=0.885
r466 80 108 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=22.68 $Y=1.065
+ $X2=22.63 $Y2=1.215
r467 80 112 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=22.68 $Y=1.065
+ $X2=22.68 $Y2=0.885
r468 78 106 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=22.055 $Y=1.215
+ $X2=21.79 $Y2=1.215
r469 77 108 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=22.465 $Y=1.215
+ $X2=22.63 $Y2=1.215
r470 77 78 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=22.465 $Y=1.215
+ $X2=22.055 $Y2=1.215
r471 73 106 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=21.89 $Y=1.065
+ $X2=21.79 $Y2=1.215
r472 73 75 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=21.89 $Y=1.065
+ $X2=21.89 $Y2=0.68
r473 69 104 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=16.75 $Y=1.065
+ $X2=16.85 $Y2=1.215
r474 69 71 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=16.75 $Y=1.065
+ $X2=16.75 $Y2=0.68
r475 68 102 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=16.175 $Y=1.215
+ $X2=16.01 $Y2=1.215
r476 67 104 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=16.585 $Y=1.215
+ $X2=16.85 $Y2=1.215
r477 67 68 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=16.585 $Y=1.215
+ $X2=16.175 $Y2=1.215
r478 66 102 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=15.96 $Y=1.065
+ $X2=16.01 $Y2=1.215
r479 66 100 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=15.96 $Y=1.065
+ $X2=15.96 $Y2=0.885
r480 64 92 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=9.8 $Y=1.065
+ $X2=9.75 $Y2=1.215
r481 64 96 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.8 $Y=1.065
+ $X2=9.8 $Y2=0.885
r482 62 90 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=9.175 $Y=1.215
+ $X2=8.91 $Y2=1.215
r483 61 92 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.585 $Y=1.215
+ $X2=9.75 $Y2=1.215
r484 61 62 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=9.585 $Y=1.215
+ $X2=9.175 $Y2=1.215
r485 57 90 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.01 $Y=1.065
+ $X2=8.91 $Y2=1.215
r486 57 59 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.01 $Y=1.065
+ $X2=9.01 $Y2=0.68
r487 53 88 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.97 $Y2=1.215
r488 53 55 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=3.87 $Y=1.065
+ $X2=3.87 $Y2=0.68
r489 52 86 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.215
+ $X2=3.13 $Y2=1.215
r490 51 88 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=3.705 $Y=1.215
+ $X2=3.97 $Y2=1.215
r491 51 52 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.705 $Y=1.215
+ $X2=3.295 $Y2=1.215
r492 50 86 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.08 $Y=1.065
+ $X2=3.13 $Y2=1.215
r493 50 84 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.08 $Y=1.065
+ $X2=3.08 $Y2=0.885
r494 16 178 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.485
+ $Y=1.555 $X2=22.63 $Y2=1.7
r495 15 173 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=21.545
+ $Y=1.555 $X2=21.69 $Y2=1.7
r496 14 168 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.805
+ $Y=1.555 $X2=16.95 $Y2=1.7
r497 13 165 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=15.865
+ $Y=1.555 $X2=16.01 $Y2=1.7
r498 12 162 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.605
+ $Y=1.555 $X2=9.75 $Y2=1.7
r499 11 157 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.665
+ $Y=1.555 $X2=8.81 $Y2=1.7
r500 10 152 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.555 $X2=4.07 $Y2=1.7
r501 9 147 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.985
+ $Y=1.555 $X2=3.13 $Y2=1.7
r502 8 110 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=22.595
+ $Y=0.33 $X2=22.73 $Y2=0.68
r503 7 75 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=21.755
+ $Y=0.33 $X2=21.89 $Y2=0.68
r504 6 71 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=16.615
+ $Y=0.33 $X2=16.75 $Y2=0.68
r505 5 98 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=15.775
+ $Y=0.33 $X2=15.91 $Y2=0.68
r506 4 94 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=0.33 $X2=9.85 $Y2=0.68
r507 3 59 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=0.33 $X2=9.01 $Y2=0.68
r508 2 55 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=3.735
+ $Y=0.33 $X2=3.87 $Y2=0.68
r509 1 82 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.33 $X2=3.03 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1643_311# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 40 42 44 46
c105 24 0 1.3204e-19 $X=9.28 $Y=1.7
r106 40 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.15 $Y=1.665
+ $X2=12.15 $Y2=1.58
r107 40 42 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.15 $Y=1.665
+ $X2=12.15 $Y2=2.34
r108 39 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=1.58
+ $X2=11.21 $Y2=1.58
r109 38 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.985 $Y=1.58
+ $X2=12.15 $Y2=1.58
r110 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=1.58
+ $X2=11.375 $Y2=1.58
r111 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=1.665
+ $X2=11.21 $Y2=1.58
r112 34 36 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.21 $Y=1.665
+ $X2=11.21 $Y2=2.34
r113 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=1.58
+ $X2=11.21 $Y2=1.58
r114 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=11.045 $Y=1.58
+ $X2=10.385 $Y2=1.58
r115 29 31 22.8568 $w=2.98e-07 $l=5.95e-07 $layer=LI1_cond $X=10.235 $Y=2.295
+ $X2=10.235 $Y2=1.7
r116 28 33 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.235 $Y=1.665
+ $X2=10.385 $Y2=1.58
r117 28 31 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=10.235 $Y=1.665
+ $X2=10.235 $Y2=1.7
r118 27 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.415 $Y=2.38
+ $X2=9.28 $Y2=2.38
r119 26 29 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.085 $Y=2.38
+ $X2=10.235 $Y2=2.295
r120 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.085 $Y=2.38
+ $X2=9.415 $Y2=2.38
r121 22 44 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=2.295
+ $X2=9.28 $Y2=2.38
r122 22 24 25.3964 $w=2.68e-07 $l=5.95e-07 $layer=LI1_cond $X=9.28 $Y=2.295
+ $X2=9.28 $Y2=1.7
r123 20 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.145 $Y=2.38
+ $X2=9.28 $Y2=2.38
r124 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.145 $Y=2.38
+ $X2=8.475 $Y2=2.38
r125 16 21 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.325 $Y=2.295
+ $X2=8.475 $Y2=2.38
r126 16 18 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=8.325 $Y=2.295
+ $X2=8.325 $Y2=1.73
r127 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=1.66
r128 5 42 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=2.34
r129 4 46 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.485 $X2=11.21 $Y2=1.66
r130 4 36 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.065
+ $Y=1.485 $X2=11.21 $Y2=2.34
r131 3 31 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.075
+ $Y=1.555 $X2=10.22 $Y2=1.7
r132 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.135
+ $Y=1.555 $X2=9.28 $Y2=1.7
r133 1 18 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=8.215
+ $Y=1.555 $X2=8.34 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2693_297# 1 2 3 4 5 16 18 20 24 26 31
+ 32 33 36 38 42 47 48
c102 36 0 1.3204e-19 $X=16.48 $Y=1.7
r103 40 42 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=17.435 $Y=2.295
+ $X2=17.435 $Y2=1.73
r104 39 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.615 $Y=2.38
+ $X2=16.48 $Y2=2.38
r105 38 40 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=17.285 $Y=2.38
+ $X2=17.435 $Y2=2.295
r106 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.285 $Y=2.38
+ $X2=16.615 $Y2=2.38
r107 34 48 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.48 $Y=2.295
+ $X2=16.48 $Y2=2.38
r108 34 36 25.3964 $w=2.68e-07 $l=5.95e-07 $layer=LI1_cond $X=16.48 $Y=2.295
+ $X2=16.48 $Y2=1.7
r109 32 48 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.345 $Y=2.38
+ $X2=16.48 $Y2=2.38
r110 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.345 $Y=2.38
+ $X2=15.675 $Y2=2.38
r111 29 33 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=15.525 $Y=2.295
+ $X2=15.675 $Y2=2.38
r112 29 31 22.8568 $w=2.98e-07 $l=5.95e-07 $layer=LI1_cond $X=15.525 $Y=2.295
+ $X2=15.525 $Y2=1.7
r113 28 31 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=15.525 $Y=1.665
+ $X2=15.525 $Y2=1.7
r114 27 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=1.58
+ $X2=14.55 $Y2=1.58
r115 26 28 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=15.375 $Y=1.58
+ $X2=15.525 $Y2=1.665
r116 26 27 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=15.375 $Y=1.58
+ $X2=14.715 $Y2=1.58
r117 22 47 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.55 $Y=1.665
+ $X2=14.55 $Y2=1.58
r118 22 24 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.55 $Y=1.665
+ $X2=14.55 $Y2=2.34
r119 21 45 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.775 $Y=1.58
+ $X2=13.61 $Y2=1.58
r120 20 47 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=1.58
+ $X2=14.55 $Y2=1.58
r121 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=1.58
+ $X2=13.775 $Y2=1.58
r122 16 45 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.61 $Y=1.665
+ $X2=13.61 $Y2=1.58
r123 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.61 $Y=1.665
+ $X2=13.61 $Y2=2.34
r124 5 42 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=17.275
+ $Y=1.555 $X2=17.42 $Y2=1.73
r125 4 36 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.335
+ $Y=1.555 $X2=16.48 $Y2=1.7
r126 3 31 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=15.415
+ $Y=1.555 $X2=15.54 $Y2=1.7
r127 2 47 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=1.485 $X2=14.55 $Y2=1.66
r128 2 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.405
+ $Y=1.485 $X2=14.55 $Y2=2.34
r129 1 45 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=1.66
r130 1 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4219_311# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 40 42 44 46
c92 24 0 1.3204e-19 $X=22.16 $Y=1.7
r93 40 48 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.03 $Y=1.665
+ $X2=25.03 $Y2=1.58
r94 40 42 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=25.03 $Y=1.665
+ $X2=25.03 $Y2=2.34
r95 39 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=1.58
+ $X2=24.09 $Y2=1.58
r96 38 48 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.865 $Y=1.58
+ $X2=25.03 $Y2=1.58
r97 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=1.58
+ $X2=24.255 $Y2=1.58
r98 34 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=24.09 $Y=1.665
+ $X2=24.09 $Y2=1.58
r99 34 36 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=24.09 $Y=1.665
+ $X2=24.09 $Y2=2.34
r100 32 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=1.58
+ $X2=24.09 $Y2=1.58
r101 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=23.925 $Y=1.58
+ $X2=23.265 $Y2=1.58
r102 29 31 22.8568 $w=2.98e-07 $l=5.95e-07 $layer=LI1_cond $X=23.115 $Y=2.295
+ $X2=23.115 $Y2=1.7
r103 28 33 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=23.115 $Y=1.665
+ $X2=23.265 $Y2=1.58
r104 28 31 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=23.115 $Y=1.665
+ $X2=23.115 $Y2=1.7
r105 27 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=22.295 $Y=2.38
+ $X2=22.16 $Y2=2.38
r106 26 29 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=22.965 $Y=2.38
+ $X2=23.115 $Y2=2.295
r107 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.965 $Y=2.38
+ $X2=22.295 $Y2=2.38
r108 22 44 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.16 $Y=2.295
+ $X2=22.16 $Y2=2.38
r109 22 24 25.3964 $w=2.68e-07 $l=5.95e-07 $layer=LI1_cond $X=22.16 $Y=2.295
+ $X2=22.16 $Y2=1.7
r110 20 44 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=22.025 $Y=2.38
+ $X2=22.16 $Y2=2.38
r111 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.025 $Y=2.38
+ $X2=21.355 $Y2=2.38
r112 16 21 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=21.205 $Y=2.295
+ $X2=21.355 $Y2=2.38
r113 16 18 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=21.205 $Y=2.295
+ $X2=21.205 $Y2=1.73
r114 5 48 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=1.66
r115 5 42 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=2.34
r116 4 46 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=1.485 $X2=24.09 $Y2=1.66
r117 4 36 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=23.945
+ $Y=1.485 $X2=24.09 $Y2=2.34
r118 3 31 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.955
+ $Y=1.555 $X2=23.1 $Y2=1.7
r119 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.015
+ $Y=1.555 $X2=22.16 $Y2=1.7
r120 1 18 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=21.095
+ $Y=1.555 $X2=21.22 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 61 63 67 69 73 77 81 85 89 93 97 101 103 107 111 113 117 121
+ 125 129 133 137 141 143 145 148 149 151 152 154 155 157 158 160 161 163 164
+ 166 167 169 170 172 173 175 176 177 178 179 180 185 212 216 221 248 252 261
+ 264 267 270 273 276 279 282
r340 282 283 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=0
+ $X2=24.61 $Y2=0
r341 279 280 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r342 277 280 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=14.95 $Y2=0
r343 276 277 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r344 267 268 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r345 264 265 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r346 262 265 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r347 261 262 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r348 256 283 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.07 $Y=0
+ $X2=24.61 $Y2=0
r349 255 256 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=0
+ $X2=25.07 $Y2=0
r350 253 282 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.695 $Y=0
+ $X2=24.56 $Y2=0
r351 253 255 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=24.695 $Y=0
+ $X2=25.07 $Y2=0
r352 252 285 3.97515 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=25.365 $Y=0
+ $X2=25.562 $Y2=0
r353 252 255 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=25.365 $Y=0
+ $X2=25.07 $Y2=0
r354 251 283 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=0
+ $X2=24.61 $Y2=0
r355 250 251 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=0
+ $X2=24.15 $Y2=0
r356 248 282 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=24.425 $Y=0
+ $X2=24.56 $Y2=0
r357 248 250 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=24.425 $Y=0
+ $X2=24.15 $Y2=0
r358 247 251 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=0
+ $X2=24.15 $Y2=0
r359 246 247 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=0
+ $X2=23.23 $Y2=0
r360 244 247 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r361 243 246 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r362 243 244 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=0
+ $X2=20.93 $Y2=0
r363 241 244 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=20.93 $Y2=0
r364 240 241 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=0
+ $X2=20.47 $Y2=0
r365 238 241 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=0
+ $X2=20.47 $Y2=0
r366 237 238 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=0
+ $X2=19.55 $Y2=0
r367 235 238 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=18.63 $Y=0
+ $X2=19.55 $Y2=0
r368 234 235 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=0
+ $X2=18.63 $Y2=0
r369 232 235 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=17.71 $Y=0
+ $X2=18.63 $Y2=0
r370 231 232 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=17.71 $Y=0
+ $X2=17.71 $Y2=0
r371 229 232 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=17.71 $Y2=0
r372 229 280 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=14.95 $Y2=0
r373 228 231 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=15.41 $Y=0
+ $X2=17.71 $Y2=0
r374 228 229 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r375 226 279 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.135 $Y=0
+ $X2=15.01 $Y2=0
r376 226 228 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.135 $Y=0
+ $X2=15.41 $Y2=0
r377 225 277 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r378 224 225 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r379 222 273 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.275 $Y=0
+ $X2=13.15 $Y2=0
r380 222 224 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.275 $Y=0
+ $X2=13.57 $Y2=0
r381 221 276 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.945 $Y=0
+ $X2=14.08 $Y2=0
r382 221 224 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=13.945 $Y=0
+ $X2=13.57 $Y2=0
r383 220 268 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.19 $Y=0
+ $X2=11.73 $Y2=0
r384 219 220 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r385 217 267 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.815 $Y=0
+ $X2=11.68 $Y2=0
r386 217 219 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.815 $Y=0
+ $X2=12.19 $Y2=0
r387 216 270 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.485 $Y=0
+ $X2=12.61 $Y2=0
r388 216 219 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.485 $Y=0
+ $X2=12.19 $Y2=0
r389 215 268 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=11.73 $Y2=0
r390 214 215 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r391 212 267 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.68 $Y2=0
r392 212 214 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.545 $Y=0
+ $X2=11.27 $Y2=0
r393 211 215 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r394 210 211 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r395 208 211 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=10.35 $Y2=0
r396 207 210 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.05 $Y=0
+ $X2=10.35 $Y2=0
r397 207 208 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r398 205 208 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r399 204 205 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r400 202 205 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r401 201 202 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r402 199 202 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r403 198 199 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r404 196 199 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r405 195 196 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r406 193 196 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=4.83 $Y2=0
r407 193 265 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=2.07 $Y2=0
r408 192 195 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0
+ $X2=4.83 $Y2=0
r409 192 193 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r410 190 264 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.13 $Y2=0
r411 190 192 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.255 $Y=0
+ $X2=2.53 $Y2=0
r412 189 262 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r413 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r414 186 258 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r415 186 188 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.69 $Y2=0
r416 185 261 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=1.2 $Y2=0
r417 185 188 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=0.69 $Y2=0
r418 180 256 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=0
+ $X2=25.07 $Y2=0
r419 180 285 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=0
+ $X2=25.53 $Y2=0
r420 179 225 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r421 179 273 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r422 178 179 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r423 178 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r424 178 270 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r425 177 189 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r426 177 258 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r427 175 246 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=23.505 $Y=0
+ $X2=23.23 $Y2=0
r428 175 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.505 $Y=0
+ $X2=23.63 $Y2=0
r429 174 250 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=23.755 $Y=0
+ $X2=24.15 $Y2=0
r430 174 176 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=23.755 $Y=0
+ $X2=23.63 $Y2=0
r431 172 240 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=20.51 $Y=0
+ $X2=20.47 $Y2=0
r432 172 173 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.51 $Y=0
+ $X2=20.655 $Y2=0
r433 171 243 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=20.8 $Y=0
+ $X2=20.93 $Y2=0
r434 171 173 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=20.8 $Y=0
+ $X2=20.655 $Y2=0
r435 169 237 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=19.59 $Y=0
+ $X2=19.55 $Y2=0
r436 169 170 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.59 $Y=0
+ $X2=19.735 $Y2=0
r437 168 240 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=19.88 $Y=0
+ $X2=20.47 $Y2=0
r438 168 170 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.88 $Y=0
+ $X2=19.735 $Y2=0
r439 166 234 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=18.76 $Y=0
+ $X2=18.63 $Y2=0
r440 166 167 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.76 $Y=0
+ $X2=18.905 $Y2=0
r441 165 237 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=19.05 $Y=0
+ $X2=19.55 $Y2=0
r442 165 167 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=19.05 $Y=0
+ $X2=18.905 $Y2=0
r443 163 231 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=17.84 $Y=0
+ $X2=17.71 $Y2=0
r444 163 164 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=17.84 $Y=0
+ $X2=17.985 $Y2=0
r445 162 234 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=18.13 $Y=0
+ $X2=18.63 $Y2=0
r446 162 164 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=18.13 $Y=0
+ $X2=17.985 $Y2=0
r447 160 210 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.35 $Y2=0
r448 160 161 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.625 $Y=0
+ $X2=10.75 $Y2=0
r449 159 214 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.875 $Y=0
+ $X2=11.27 $Y2=0
r450 159 161 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.875 $Y=0
+ $X2=10.75 $Y2=0
r451 157 204 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=7.63 $Y=0 $X2=7.59
+ $Y2=0
r452 157 158 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.63 $Y=0
+ $X2=7.775 $Y2=0
r453 156 207 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=8.05 $Y2=0
r454 156 158 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7.92 $Y=0
+ $X2=7.775 $Y2=0
r455 154 201 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=6.71 $Y=0 $X2=6.67
+ $Y2=0
r456 154 155 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.71 $Y=0
+ $X2=6.855 $Y2=0
r457 153 204 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=7 $Y=0 $X2=7.59
+ $Y2=0
r458 153 155 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=7 $Y=0 $X2=6.855
+ $Y2=0
r459 151 198 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.88 $Y=0
+ $X2=5.75 $Y2=0
r460 151 152 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.88 $Y=0
+ $X2=6.025 $Y2=0
r461 150 201 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=6.17 $Y=0 $X2=6.67
+ $Y2=0
r462 150 152 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=6.17 $Y=0
+ $X2=6.025 $Y2=0
r463 148 195 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=4.83 $Y2=0
r464 148 149 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=4.96 $Y=0
+ $X2=5.105 $Y2=0
r465 147 198 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.75
+ $Y2=0
r466 147 149 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=5.25 $Y=0
+ $X2=5.105 $Y2=0
r467 143 285 3.16801 $w=2.5e-07 $l=1.15521e-07 $layer=LI1_cond $X=25.49 $Y=0.085
+ $X2=25.562 $Y2=0
r468 143 145 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=25.49 $Y=0.085
+ $X2=25.49 $Y2=0.38
r469 139 282 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=24.56 $Y=0.085
+ $X2=24.56 $Y2=0
r470 139 141 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=24.56 $Y=0.085
+ $X2=24.56 $Y2=0.38
r471 135 176 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=23.63 $Y=0.085
+ $X2=23.63 $Y2=0
r472 135 137 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=23.63 $Y=0.085
+ $X2=23.63 $Y2=0.38
r473 131 173 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=20.655 $Y=0.085
+ $X2=20.655 $Y2=0
r474 131 133 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=20.655 $Y=0.085
+ $X2=20.655 $Y2=0.445
r475 127 170 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=19.735 $Y=0.085
+ $X2=19.735 $Y2=0
r476 127 129 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=19.735 $Y=0.085
+ $X2=19.735 $Y2=0.445
r477 123 167 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=18.905 $Y=0.085
+ $X2=18.905 $Y2=0
r478 123 125 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=18.905 $Y=0.085
+ $X2=18.905 $Y2=0.445
r479 119 164 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=17.985 $Y=0.085
+ $X2=17.985 $Y2=0
r480 119 121 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=17.985 $Y=0.085
+ $X2=17.985 $Y2=0.445
r481 115 279 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=15.01 $Y=0.085
+ $X2=15.01 $Y2=0
r482 115 117 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=15.01 $Y=0.085
+ $X2=15.01 $Y2=0.38
r483 114 276 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.215 $Y=0
+ $X2=14.08 $Y2=0
r484 113 279 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=15.01 $Y2=0
r485 113 114 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.215 $Y2=0
r486 109 276 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.08 $Y=0.085
+ $X2=14.08 $Y2=0
r487 109 111 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.08 $Y=0.085
+ $X2=14.08 $Y2=0.38
r488 105 273 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.15 $Y=0.085
+ $X2=13.15 $Y2=0
r489 105 107 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=13.15 $Y=0.085
+ $X2=13.15 $Y2=0.38
r490 104 270 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.735 $Y=0
+ $X2=12.61 $Y2=0
r491 103 273 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.025 $Y=0
+ $X2=13.15 $Y2=0
r492 103 104 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.025 $Y=0
+ $X2=12.735 $Y2=0
r493 99 270 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.61 $Y=0.085
+ $X2=12.61 $Y2=0
r494 99 101 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=12.61 $Y=0.085
+ $X2=12.61 $Y2=0.38
r495 95 267 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0
r496 95 97 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.68 $Y=0.085
+ $X2=11.68 $Y2=0.38
r497 91 161 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0
r498 91 93 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.75 $Y=0.085
+ $X2=10.75 $Y2=0.38
r499 87 158 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.775 $Y2=0
r500 87 89 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=7.775 $Y=0.085
+ $X2=7.775 $Y2=0.445
r501 83 155 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.855 $Y=0.085
+ $X2=6.855 $Y2=0
r502 83 85 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.855 $Y=0.085
+ $X2=6.855 $Y2=0.445
r503 79 152 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.025 $Y=0.085
+ $X2=6.025 $Y2=0
r504 79 81 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=6.025 $Y=0.085
+ $X2=6.025 $Y2=0.445
r505 75 149 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0
r506 75 77 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=5.105 $Y=0.085
+ $X2=5.105 $Y2=0.445
r507 71 264 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0
r508 71 73 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.13 $Y=0.085
+ $X2=2.13 $Y2=0.38
r509 70 261 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.2
+ $Y2=0
r510 69 264 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.13 $Y2=0
r511 69 70 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.335 $Y2=0
r512 65 261 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r513 65 67 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.38
r514 61 258 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r515 61 63 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r516 20 145 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=0.235 $X2=25.45 $Y2=0.38
r517 19 141 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=24.375
+ $Y=0.235 $X2=24.56 $Y2=0.38
r518 18 137 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=23.545
+ $Y=0.235 $X2=23.67 $Y2=0.38
r519 17 133 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=20.46
+ $Y=0.235 $X2=20.595 $Y2=0.445
r520 16 129 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=19.63
+ $Y=0.235 $X2=19.755 $Y2=0.445
r521 15 125 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=18.75
+ $Y=0.235 $X2=18.885 $Y2=0.445
r522 14 121 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=17.92
+ $Y=0.235 $X2=18.045 $Y2=0.445
r523 13 117 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=14.835
+ $Y=0.235 $X2=14.97 $Y2=0.38
r524 12 111 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=13.895
+ $Y=0.235 $X2=14.08 $Y2=0.38
r525 11 107 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=0.235 $X2=13.19 $Y2=0.38
r526 10 101 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=0.235 $X2=12.57 $Y2=0.38
r527 9 97 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.495
+ $Y=0.235 $X2=11.68 $Y2=0.38
r528 8 93 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.235 $X2=10.79 $Y2=0.38
r529 7 89 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=7.58
+ $Y=0.235 $X2=7.715 $Y2=0.445
r530 6 85 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=0.235 $X2=6.875 $Y2=0.445
r531 5 81 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.005 $Y2=0.445
r532 4 77 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.165 $Y2=0.445
r533 3 73 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.09 $Y2=0.38
r534 2 67 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r535 1 63 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_119_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=4.29 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=4.33 $Y=0.425
+ $X2=4.33 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.535 $Y=0.34
+ $X2=3.45 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.205 $Y=0.34
+ $X2=4.33 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.205 $Y=0.34
+ $X2=3.535 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=0.425
+ $X2=3.45 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=3.45 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.365 $Y=0.34
+ $X2=2.695 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.56 $Y=0.715
+ $X2=2.56 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.695 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.56 $Y=0.425
+ $X2=2.56 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0.8
+ $X2=1.67 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=2.56 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=1.835 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=0.715
+ $X2=1.67 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.8
+ $X2=1.67 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=0.8
+ $X2=0.895 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.895 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.73 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=4.155
+ $Y=0.33 $X2=4.29 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.315
+ $Y=0.33 $X2=3.45 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.33 $X2=2.61 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_1693_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.15 $Y=0.715
+ $X2=12.15 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.375 $Y=0.8
+ $X2=11.21 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=11.985 $Y=0.8
+ $X2=12.15 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.985 $Y=0.8
+ $X2=11.375 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.21 $Y=0.715
+ $X2=11.21 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.21 $Y=0.715
+ $X2=11.21 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.045 $Y=0.8
+ $X2=11.21 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=11.045 $Y=0.8
+ $X2=10.455 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.32 $Y=0.715
+ $X2=10.455 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=10.32 $Y=0.715
+ $X2=10.32 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.32 $Y=0.425
+ $X2=10.32 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=0.34
+ $X2=9.43 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=10.32 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=9.515 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=9.43 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=8.675 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=8.55 $Y=0.425
+ $X2=8.675 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.55 $Y=0.425
+ $X2=8.55 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.015
+ $Y=0.235 $X2=12.15 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=11.075
+ $Y=0.235 $X2=11.21 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=0.33 $X2=10.27 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.33 $X2=9.43 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.33 $X2=8.59 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_2695_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=17.17 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=17.21 $Y=0.425
+ $X2=17.21 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.415 $Y=0.34
+ $X2=16.33 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=17.085 $Y=0.34
+ $X2=17.21 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.085 $Y=0.34
+ $X2=16.415 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.33 $Y=0.425
+ $X2=16.33 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.33 $Y=0.425
+ $X2=16.33 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.245 $Y=0.34
+ $X2=16.33 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.245 $Y=0.34
+ $X2=15.575 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=15.44 $Y=0.715
+ $X2=15.44 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.44 $Y=0.425
+ $X2=15.575 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.44 $Y=0.425
+ $X2=15.44 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.715 $Y=0.8
+ $X2=14.55 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=15.305 $Y=0.8
+ $X2=15.44 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=15.305 $Y=0.8
+ $X2=14.715 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.55 $Y=0.715
+ $X2=14.55 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.55 $Y=0.715
+ $X2=14.55 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.385 $Y=0.8
+ $X2=14.55 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.385 $Y=0.8
+ $X2=13.775 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.61 $Y=0.715
+ $X2=13.775 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.61 $Y=0.715
+ $X2=13.61 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=17.035
+ $Y=0.33 $X2=17.17 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.195
+ $Y=0.33 $X2=16.33 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.365
+ $Y=0.33 $X2=15.49 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=14.415
+ $Y=0.235 $X2=14.55 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=13.475
+ $Y=0.235 $X2=13.61 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_4%A_4269_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=25.03 $Y=0.715
+ $X2=25.03 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=24.255 $Y=0.8
+ $X2=24.09 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=24.865 $Y=0.8
+ $X2=25.03 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=24.865 $Y=0.8
+ $X2=24.255 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=24.09 $Y=0.715
+ $X2=24.09 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=24.09 $Y=0.715
+ $X2=24.09 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.925 $Y=0.8
+ $X2=24.09 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=23.925 $Y=0.8
+ $X2=23.335 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.2 $Y=0.715
+ $X2=23.335 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=23.2 $Y=0.715
+ $X2=23.2 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=23.2 $Y=0.425
+ $X2=23.2 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.395 $Y=0.34
+ $X2=22.31 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=23.065 $Y=0.34
+ $X2=23.2 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=23.065 $Y=0.34
+ $X2=22.395 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.31 $Y=0.425
+ $X2=22.31 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=22.31 $Y=0.425
+ $X2=22.31 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=22.225 $Y=0.34
+ $X2=22.31 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.225 $Y=0.34
+ $X2=21.555 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=21.43 $Y=0.425
+ $X2=21.555 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=21.43 $Y=0.425
+ $X2=21.43 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=24.895
+ $Y=0.235 $X2=25.03 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=23.955
+ $Y=0.235 $X2=24.09 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=23.015
+ $Y=0.33 $X2=23.15 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.175
+ $Y=0.33 $X2=22.31 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.345
+ $Y=0.33 $X2=21.47 $Y2=0.59
.ends

