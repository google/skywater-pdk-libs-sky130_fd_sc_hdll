* File: sky130_fd_sc_hdll__and3b_1.pxi.spice
* Created: Thu Aug 27 18:58:17 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND3B_1%A_N N_A_N_c_65_n N_A_N_c_66_n N_A_N_M1002_g
+ N_A_N_M1006_g A_N A_N A_N N_A_N_c_63_n N_A_N_c_64_n
+ PM_SKY130_FD_SC_HDLL__AND3B_1%A_N
x_PM_SKY130_FD_SC_HDLL__AND3B_1%A_117_413# N_A_117_413#_M1006_d
+ N_A_117_413#_M1002_d N_A_117_413#_c_87_n N_A_117_413#_M1005_g
+ N_A_117_413#_M1000_g N_A_117_413#_c_89_n N_A_117_413#_c_90_n
+ N_A_117_413#_c_91_n PM_SKY130_FD_SC_HDLL__AND3B_1%A_117_413#
x_PM_SKY130_FD_SC_HDLL__AND3B_1%B N_B_c_128_n N_B_c_131_n N_B_M1003_g
+ N_B_M1007_g B B PM_SKY130_FD_SC_HDLL__AND3B_1%B
x_PM_SKY130_FD_SC_HDLL__AND3B_1%C N_C_M1009_g N_C_c_168_n N_C_M1004_g C C
+ PM_SKY130_FD_SC_HDLL__AND3B_1%C
x_PM_SKY130_FD_SC_HDLL__AND3B_1%A_225_311# N_A_225_311#_M1000_s
+ N_A_225_311#_M1005_s N_A_225_311#_M1003_d N_A_225_311#_c_199_n
+ N_A_225_311#_M1008_g N_A_225_311#_c_200_n N_A_225_311#_M1001_g
+ N_A_225_311#_c_205_n N_A_225_311#_c_201_n N_A_225_311#_c_206_n
+ N_A_225_311#_c_207_n N_A_225_311#_c_202_n N_A_225_311#_c_209_n
+ N_A_225_311#_c_210_n N_A_225_311#_c_203_n N_A_225_311#_c_231_n
+ N_A_225_311#_c_212_n PM_SKY130_FD_SC_HDLL__AND3B_1%A_225_311#
x_PM_SKY130_FD_SC_HDLL__AND3B_1%VPWR N_VPWR_M1002_s N_VPWR_M1005_d
+ N_VPWR_M1004_d N_VPWR_c_281_n N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n
+ N_VPWR_c_299_n N_VPWR_c_285_n N_VPWR_c_286_n VPWR N_VPWR_c_287_n
+ N_VPWR_c_280_n N_VPWR_c_289_n PM_SKY130_FD_SC_HDLL__AND3B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND3B_1%X N_X_M1001_d N_X_M1008_d N_X_c_338_n
+ N_X_c_335_n N_X_c_336_n X X N_X_c_340_n PM_SKY130_FD_SC_HDLL__AND3B_1%X
x_PM_SKY130_FD_SC_HDLL__AND3B_1%VGND N_VGND_M1006_s N_VGND_M1009_d
+ N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n VGND N_VGND_c_354_n
+ N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n
+ PM_SKY130_FD_SC_HDLL__AND3B_1%VGND
cc_1 VNB A_N 0.00882809f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_2 VNB N_A_N_c_63_n 0.0472185f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_3 VNB N_A_N_c_64_n 0.0214835f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=0.995
cc_4 VNB N_A_117_413#_c_87_n 0.0323927f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.675
cc_5 VNB N_A_117_413#_M1000_g 0.0341647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_117_413#_c_89_n 0.0183572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_413#_c_90_n 0.00142667f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_8 VNB N_A_117_413#_c_91_n 0.018353f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_B_c_128_n 0.00693081f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_10 VNB N_B_M1007_g 0.0361971f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.675
cc_11 VNB N_C_M1009_g 0.0278755f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_12 VNB N_C_c_168_n 0.0220248f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_13 VNB C 0.0114747f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.675
cc_14 VNB N_A_225_311#_c_199_n 0.0266281f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_15 VNB N_A_225_311#_c_200_n 0.0217084f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_225_311#_c_201_n 0.00619913f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_17 VNB N_A_225_311#_c_202_n 0.00537442f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_311#_c_203_n 0.00167047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_280_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_335_n 0.0251985f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_21 VNB N_X_c_336_n 0.00489291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.0134195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_351_n 0.0099134f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.675
cc_24 VNB N_VGND_c_352_n 0.0388813f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_25 VNB N_VGND_c_353_n 0.0026508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_354_n 0.0657208f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_27 VNB N_VGND_c_355_n 0.016967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_356_n 0.238978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_357_n 0.00436989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_A_N_c_65_n 0.0138445f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_31 VPB N_A_N_c_66_n 0.0325653f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_32 VPB A_N 0.0279341f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_N_c_63_n 0.0487935f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_34 VPB N_A_117_413#_c_87_n 0.0354257f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.675
cc_35 VPB N_A_117_413#_c_90_n 0.0175788f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_36 VPB N_B_c_128_n 0.00974811f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_37 VPB N_B_c_131_n 0.0506702f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_38 VPB N_B_M1003_g 0.0131193f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_39 VPB B 0.0115079f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_40 VPB N_C_c_168_n 0.0273391f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_41 VPB N_A_225_311#_c_199_n 0.031519f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_42 VPB N_A_225_311#_c_205_n 0.00373964f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=0.995
cc_43 VPB N_A_225_311#_c_206_n 0.00386438f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_225_311#_c_207_n 0.00403783f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.87
cc_45 VPB N_A_225_311#_c_202_n 0.00115659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_225_311#_c_209_n 0.0131678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_225_311#_c_210_n 0.00562457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_225_311#_c_203_n 0.0011804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_225_311#_c_212_n 0.003401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_281_n 0.0098875f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_51 VPB N_VPWR_c_282_n 0.0192177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_283_n 0.0578347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_284_n 0.00498307f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_54 VPB N_VPWR_c_285_n 0.0276399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_286_n 0.00411068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_287_n 0.0209898f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_280_n 0.0623217f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_289_n 0.00146645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_X_c_338_n 0.00497936f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_X_c_335_n 0.0183724f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_61 VPB N_X_c_340_n 0.0216726f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 N_A_N_c_63_n N_A_117_413#_c_87_n 0.00414924f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_63 A_N N_A_117_413#_c_89_n 0.0118403f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_N_c_64_n N_A_117_413#_c_89_n 0.0220735f $X=0.352 $Y=0.995 $X2=0 $Y2=0
cc_65 N_A_N_c_66_n N_A_117_413#_c_90_n 0.00586027f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_66 A_N N_A_117_413#_c_90_n 0.0439765f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_67 N_A_N_c_63_n N_A_117_413#_c_90_n 0.0194016f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_N_c_64_n N_A_225_311#_c_201_n 0.00458211f $X=0.352 $Y=0.995 $X2=0
+ $Y2=0
cc_69 N_A_N_c_66_n N_VPWR_c_282_n 0.00656462f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_70 A_N N_VPWR_c_282_n 0.0230454f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_N_c_63_n N_VPWR_c_282_n 0.00102514f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_N_c_66_n N_VPWR_c_283_n 0.0109746f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_73 N_A_N_c_66_n N_VPWR_c_280_n 0.0148061f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_74 A_N N_VPWR_c_280_n 0.00417076f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_75 A_N N_VGND_c_352_n 0.0231087f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_N_c_63_n N_VGND_c_352_n 0.0069709f $X=0.26 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_N_c_64_n N_VGND_c_352_n 0.0082712f $X=0.352 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_N_c_64_n N_VGND_c_354_n 0.00439675f $X=0.352 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_N_c_64_n N_VGND_c_356_n 0.00512902f $X=0.352 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_117_413#_c_87_n N_B_c_128_n 0.0125342f $X=1.485 $Y=1.48 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_117_413#_c_87_n N_B_c_131_n 8.20148e-19 $X=1.485 $Y=1.48 $X2=0 $Y2=0
cc_82 N_A_117_413#_c_87_n N_B_M1003_g 0.012504f $X=1.485 $Y=1.48 $X2=0 $Y2=0
cc_83 N_A_117_413#_M1000_g N_B_M1007_g 0.0388046f $X=1.51 $Y=0.475 $X2=0 $Y2=0
cc_84 N_A_117_413#_c_90_n N_A_225_311#_c_205_n 0.0193726f $X=0.73 $Y=2.26 $X2=0
+ $Y2=0
cc_85 N_A_117_413#_c_87_n N_A_225_311#_c_201_n 0.00402884f $X=1.485 $Y=1.48
+ $X2=0 $Y2=0
cc_86 N_A_117_413#_M1000_g N_A_225_311#_c_201_n 0.0135153f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_87 N_A_117_413#_c_89_n N_A_225_311#_c_201_n 0.00494617f $X=0.73 $Y=1.245
+ $X2=0 $Y2=0
cc_88 N_A_117_413#_c_91_n N_A_225_311#_c_201_n 0.0139713f $X=1.35 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_117_413#_c_87_n N_A_225_311#_c_206_n 0.0175425f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_90 N_A_117_413#_c_91_n N_A_225_311#_c_206_n 0.0124955f $X=1.35 $Y=1.16 $X2=0
+ $Y2=0
cc_91 N_A_117_413#_c_87_n N_A_225_311#_c_207_n 0.00303382f $X=1.485 $Y=1.48
+ $X2=0 $Y2=0
cc_92 N_A_117_413#_c_90_n N_A_225_311#_c_207_n 0.0103923f $X=0.73 $Y=2.26 $X2=0
+ $Y2=0
cc_93 N_A_117_413#_c_91_n N_A_225_311#_c_207_n 0.0198862f $X=1.35 $Y=1.16 $X2=0
+ $Y2=0
cc_94 N_A_117_413#_M1000_g N_A_225_311#_c_202_n 0.0173781f $X=1.51 $Y=0.475
+ $X2=0 $Y2=0
cc_95 N_A_117_413#_c_91_n N_A_225_311#_c_202_n 0.0204125f $X=1.35 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_117_413#_c_90_n N_VPWR_c_282_n 0.0167876f $X=0.73 $Y=2.26 $X2=0 $Y2=0
cc_97 N_A_117_413#_c_87_n N_VPWR_c_283_n 0.00448433f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_98 N_A_117_413#_c_90_n N_VPWR_c_283_n 0.0317087f $X=0.73 $Y=2.26 $X2=0 $Y2=0
cc_99 N_A_117_413#_c_87_n N_VPWR_c_299_n 0.00436781f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_100 N_A_117_413#_M1002_d N_VPWR_c_280_n 0.00549204f $X=0.585 $Y=2.065 $X2=0
+ $Y2=0
cc_101 N_A_117_413#_c_90_n N_VPWR_c_280_n 0.00646998f $X=0.73 $Y=2.26 $X2=0
+ $Y2=0
cc_102 N_A_117_413#_c_87_n N_VPWR_c_289_n 0.0109006f $X=1.485 $Y=1.48 $X2=0
+ $Y2=0
cc_103 N_A_117_413#_c_89_n N_VGND_c_352_n 0.032547f $X=0.73 $Y=1.245 $X2=0 $Y2=0
cc_104 N_A_117_413#_M1000_g N_VGND_c_354_n 0.00344034f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_105 N_A_117_413#_c_89_n N_VGND_c_354_n 0.00967825f $X=0.73 $Y=1.245 $X2=0
+ $Y2=0
cc_106 N_A_117_413#_M1000_g N_VGND_c_356_n 0.00614431f $X=1.51 $Y=0.475 $X2=0
+ $Y2=0
cc_107 N_A_117_413#_c_89_n N_VGND_c_356_n 0.012569f $X=0.73 $Y=1.245 $X2=0 $Y2=0
cc_108 N_B_M1007_g N_C_M1009_g 0.0285811f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_109 N_B_c_128_n N_C_c_168_n 0.03459f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_110 N_B_M1003_g N_C_c_168_n 0.00685146f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_111 B N_C_c_168_n 0.00319465f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_112 N_B_M1007_g C 0.00509517f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_113 N_B_M1007_g N_A_225_311#_c_201_n 0.0078714f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_114 N_B_c_128_n N_A_225_311#_c_202_n 0.00805911f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_115 N_B_M1007_g N_A_225_311#_c_202_n 0.0159249f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_116 N_B_c_131_n N_A_225_311#_c_210_n 2.4825e-19 $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_117 B N_A_225_311#_c_210_n 0.0193859f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_118 N_B_c_128_n N_A_225_311#_c_231_n 0.00121429f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_119 N_B_M1003_g N_A_225_311#_c_231_n 0.00501962f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_120 B N_A_225_311#_c_231_n 7.85933e-19 $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_121 N_B_c_128_n N_A_225_311#_c_212_n 0.00622928f $X=1.955 $Y=1.48 $X2=0 $Y2=0
cc_122 N_B_c_131_n N_A_225_311#_c_212_n 3.74322e-19 $X=1.955 $Y=2.105 $X2=0
+ $Y2=0
cc_123 N_B_M1003_g N_A_225_311#_c_212_n 0.00456287f $X=1.955 $Y=1.765 $X2=0
+ $Y2=0
cc_124 B N_A_225_311#_c_212_n 0.00565787f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_125 N_B_c_131_n N_VPWR_c_284_n 0.00187778f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_126 B N_VPWR_c_284_n 0.0187455f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_127 N_B_M1003_g N_VPWR_c_299_n 0.00356134f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_128 N_B_c_131_n N_VPWR_c_285_n 0.00705703f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_129 B N_VPWR_c_285_n 0.0380394f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_130 N_B_c_131_n N_VPWR_c_280_n 0.00988926f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_131 B N_VPWR_c_280_n 0.020518f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_132 N_B_c_131_n N_VPWR_c_289_n 0.0104622f $X=1.955 $Y=2.105 $X2=0 $Y2=0
cc_133 N_B_M1003_g N_VPWR_c_289_n 0.0035201f $X=1.955 $Y=1.765 $X2=0 $Y2=0
cc_134 B N_VPWR_c_289_n 0.0295126f $X=2.165 $Y=2.125 $X2=0 $Y2=0
cc_135 N_B_M1007_g N_VGND_c_354_n 0.00498872f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_136 N_B_M1007_g N_VGND_c_356_n 0.00912581f $X=1.98 $Y=0.475 $X2=0 $Y2=0
cc_137 N_C_c_168_n N_A_225_311#_c_199_n 0.0264116f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_138 C N_A_225_311#_c_199_n 0.00190122f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_139 N_C_M1009_g N_A_225_311#_c_200_n 0.00857445f $X=2.385 $Y=0.475 $X2=0
+ $Y2=0
cc_140 C N_A_225_311#_c_200_n 0.00567069f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_141 N_C_M1009_g N_A_225_311#_c_201_n 3.55938e-19 $X=2.385 $Y=0.475 $X2=0
+ $Y2=0
cc_142 N_C_M1009_g N_A_225_311#_c_202_n 7.41404e-19 $X=2.385 $Y=0.475 $X2=0
+ $Y2=0
cc_143 N_C_c_168_n N_A_225_311#_c_202_n 8.80303e-19 $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_144 C N_A_225_311#_c_202_n 0.0297402f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_145 N_C_c_168_n N_A_225_311#_c_209_n 0.0228144f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_146 N_C_c_168_n N_A_225_311#_c_210_n 0.00236013f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_147 C N_A_225_311#_c_210_n 0.0307873f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_148 N_C_c_168_n N_A_225_311#_c_203_n 0.00255391f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_149 C N_A_225_311#_c_203_n 0.0136635f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_150 N_C_c_168_n N_VPWR_c_299_n 2.59092e-19 $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_151 N_C_c_168_n N_VPWR_c_285_n 0.00170065f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_152 N_C_c_168_n N_VPWR_c_280_n 0.00208744f $X=2.48 $Y=1.41 $X2=0 $Y2=0
cc_153 C N_VGND_M1009_d 0.00551998f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_154 N_C_M1009_g N_VGND_c_353_n 0.0036983f $X=2.385 $Y=0.475 $X2=0 $Y2=0
cc_155 C N_VGND_c_353_n 0.0256165f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_156 N_C_M1009_g N_VGND_c_354_n 0.0034758f $X=2.385 $Y=0.475 $X2=0 $Y2=0
cc_157 C N_VGND_c_354_n 0.0167959f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_158 N_C_M1009_g N_VGND_c_356_n 0.00550276f $X=2.385 $Y=0.475 $X2=0 $Y2=0
cc_159 C N_VGND_c_356_n 0.0129231f $X=2.365 $Y=0.425 $X2=0 $Y2=0
cc_160 N_A_225_311#_c_206_n N_VPWR_M1005_d 6.07398e-19 $X=1.69 $Y=1.51 $X2=0
+ $Y2=0
cc_161 N_A_225_311#_c_231_n N_VPWR_M1005_d 0.00130903f $X=1.817 $Y=1.51 $X2=0
+ $Y2=0
cc_162 N_A_225_311#_c_209_n N_VPWR_M1004_d 0.00847106f $X=2.965 $Y=1.657 $X2=0
+ $Y2=0
cc_163 N_A_225_311#_c_205_n N_VPWR_c_283_n 0.0198637f $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_164 N_A_225_311#_c_206_n N_VPWR_c_283_n 0.00498695f $X=1.69 $Y=1.51 $X2=0
+ $Y2=0
cc_165 N_A_225_311#_c_199_n N_VPWR_c_284_n 0.00574443f $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_225_311#_c_209_n N_VPWR_c_284_n 0.0143599f $X=2.965 $Y=1.657 $X2=0
+ $Y2=0
cc_167 N_A_225_311#_c_205_n N_VPWR_c_299_n 0.0134323f $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_168 N_A_225_311#_c_206_n N_VPWR_c_299_n 0.00896295f $X=1.69 $Y=1.51 $X2=0
+ $Y2=0
cc_169 N_A_225_311#_c_210_n N_VPWR_c_299_n 0.00721061f $X=2.387 $Y=1.657 $X2=0
+ $Y2=0
cc_170 N_A_225_311#_c_231_n N_VPWR_c_299_n 0.0111733f $X=1.817 $Y=1.51 $X2=0
+ $Y2=0
cc_171 N_A_225_311#_c_199_n N_VPWR_c_287_n 0.00702461f $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_225_311#_c_199_n N_VPWR_c_280_n 0.0146143f $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_225_311#_c_205_n N_VPWR_c_280_n 0.00100788f $X=1.25 $Y=1.76 $X2=0
+ $Y2=0
cc_174 N_A_225_311#_c_209_n N_VPWR_c_280_n 0.0023291f $X=2.965 $Y=1.657 $X2=0
+ $Y2=0
cc_175 N_A_225_311#_c_210_n N_VPWR_c_280_n 0.0119011f $X=2.387 $Y=1.657 $X2=0
+ $Y2=0
cc_176 N_A_225_311#_c_199_n N_X_c_335_n 0.00706371f $X=3.135 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_225_311#_c_200_n N_X_c_335_n 0.0182486f $X=3.16 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_225_311#_c_209_n N_X_c_335_n 0.0206009f $X=2.965 $Y=1.657 $X2=0 $Y2=0
cc_179 N_A_225_311#_c_203_n N_X_c_335_n 0.0313192f $X=3.1 $Y=1.16 $X2=0 $Y2=0
cc_180 N_A_225_311#_c_199_n N_VGND_c_353_n 5.93726e-19 $X=3.135 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_225_311#_c_200_n N_VGND_c_353_n 0.0106612f $X=3.16 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_225_311#_c_203_n N_VGND_c_353_n 0.00586441f $X=3.1 $Y=1.16 $X2=0
+ $Y2=0
cc_183 N_A_225_311#_c_201_n N_VGND_c_354_n 0.042298f $X=1.69 $Y=0.417 $X2=0
+ $Y2=0
cc_184 N_A_225_311#_c_200_n N_VGND_c_355_n 0.00505556f $X=3.16 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_225_311#_c_200_n N_VGND_c_356_n 0.00961922f $X=3.16 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_225_311#_c_201_n N_VGND_c_356_n 0.0304061f $X=1.69 $Y=0.417 $X2=0
+ $Y2=0
cc_187 N_A_225_311#_c_201_n A_317_53# 0.00401931f $X=1.69 $Y=0.417 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_225_311#_c_202_n A_317_53# 0.00157362f $X=1.817 $Y=1.425 $X2=-0.19
+ $Y2=-0.24
cc_189 N_VPWR_c_280_n N_X_M1008_d 0.00378012f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_190 N_VPWR_c_287_n N_X_c_340_n 0.0181772f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_191 N_VPWR_c_280_n N_X_c_340_n 0.0101314f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_192 X N_VGND_c_355_n 0.0175109f $X=3.3 $Y=0.425 $X2=0 $Y2=0
cc_193 N_X_M1001_d N_VGND_c_356_n 0.00352456f $X=3.235 $Y=0.235 $X2=0 $Y2=0
cc_194 X N_VGND_c_356_n 0.00990557f $X=3.3 $Y=0.425 $X2=0 $Y2=0
