* NGSPICE file created from sky130_fd_sc_hdll__o21ba_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VPWR a_197_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.43e+12p pd=1.286e+07u as=5.8e+11p ps=5.16e+06u
M1001 a_823_297# A2 a_197_21# VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=5.8e+11p ps=5.16e+06u
M1002 VGND A2 a_635_47# VNB nshort w=650000u l=150000u
+  ad=1.0335e+12p pd=9.68e+06u as=7.345e+11p ps=7.46e+06u
M1003 a_635_47# a_27_297# a_197_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1004 VPWR B1_N a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3.9e+11p ps=2.78e+06u
M1005 a_635_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 X a_197_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_197_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=0p ps=0u
M1008 a_197_21# A2 a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_197_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_197_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_197_21# a_27_297# a_635_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND A1 a_635_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_197_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_197_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_823_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_297# a_197_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND B1_N a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.3075e+11p ps=2.01e+06u
M1018 VPWR A1 a_823_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_635_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_197_21# a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_197_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

