# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.740000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.180000 1.075000 2.025000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 4.470000 1.285000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.695000 1.075000 6.305000 1.285000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.475000 1.075000 8.045000 1.285000 ;
    END
  END D
  PIN Y
    ANTENNADIFFAREA  2.374000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 8.630000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 4.815000 0.255000 5.195000 0.725000 ;
        RECT 5.755000 0.255000 6.135000 0.725000 ;
        RECT 6.695000 0.255000 7.075000 0.725000 ;
        RECT 6.785000 1.455000 8.630000 1.625000 ;
        RECT 6.785000 1.625000 7.035000 2.125000 ;
        RECT 7.635000 0.255000 8.015000 0.725000 ;
        RECT 7.725000 1.625000 7.975000 2.125000 ;
        RECT 8.360000 0.905000 8.630000 1.455000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 2.285000 1.625000 ;
      RECT 0.090000  1.625000 0.405000 2.465000 ;
      RECT 0.625000  1.795000 0.875000 2.635000 ;
      RECT 1.095000  1.625000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.795000 1.815000 2.635000 ;
      RECT 2.035000  1.625000 2.285000 2.295000 ;
      RECT 2.035000  2.295000 4.220000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.505000  1.455000 6.095000 1.625000 ;
      RECT 2.505000  1.625000 2.755000 2.125000 ;
      RECT 2.975000  1.795000 3.225000 2.295000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.445000  1.625000 3.695000 2.125000 ;
      RECT 3.915000  1.795000 4.220000 2.295000 ;
      RECT 3.955000  0.085000 4.645000 0.555000 ;
      RECT 4.405000  1.795000 4.685000 2.295000 ;
      RECT 4.405000  2.295000 8.445000 2.465000 ;
      RECT 4.905000  1.625000 5.155000 2.125000 ;
      RECT 5.375000  1.795000 5.625000 2.295000 ;
      RECT 5.415000  0.085000 5.585000 0.555000 ;
      RECT 5.845000  1.625000 6.095000 2.125000 ;
      RECT 6.315000  1.795000 6.565000 2.295000 ;
      RECT 6.355000  0.085000 6.525000 0.555000 ;
      RECT 7.255000  1.795000 7.505000 2.295000 ;
      RECT 7.295000  0.085000 7.465000 0.555000 ;
      RECT 8.195000  1.795000 8.445000 2.295000 ;
      RECT 8.235000  0.085000 8.405000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4_4
END LIBRARY
