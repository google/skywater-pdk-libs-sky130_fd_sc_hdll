# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor2_8
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  8.280000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.360000 1.075000 3.930000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.200000 1.075000 7.290000 1.275000 ;
    END
  END B
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.889000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.915000 0.725000 ;
        RECT 0.535000 0.725000 8.025000 0.905000 ;
        RECT 1.475000 0.255000 1.855000 0.725000 ;
        RECT 2.415000 0.255000 2.795000 0.725000 ;
        RECT 3.355000 0.255000 3.735000 0.725000 ;
        RECT 4.295000 0.255000 4.675000 0.725000 ;
        RECT 4.385000 1.445000 8.025000 1.615000 ;
        RECT 4.385000 1.615000 4.635000 2.125000 ;
        RECT 5.235000 0.255000 5.615000 0.725000 ;
        RECT 5.325000 1.615000 5.575000 2.125000 ;
        RECT 6.175000 0.255000 6.555000 0.725000 ;
        RECT 6.265000 1.615000 6.515000 2.125000 ;
        RECT 7.115000 0.255000 7.495000 0.725000 ;
        RECT 7.205000 1.615000 7.455000 2.125000 ;
        RECT 7.460000 0.905000 8.025000 1.445000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.280000 0.085000 ;
      RECT 0.000000  2.635000 8.280000 2.805000 ;
      RECT 0.090000  0.085000 0.365000 0.905000 ;
      RECT 0.090000  1.455000 4.165000 1.665000 ;
      RECT 0.090000  1.665000 0.405000 2.465000 ;
      RECT 0.625000  1.835000 0.875000 2.635000 ;
      RECT 1.095000  1.665000 1.345000 2.465000 ;
      RECT 1.135000  0.085000 1.305000 0.555000 ;
      RECT 1.565000  1.835000 1.815000 2.635000 ;
      RECT 2.035000  1.665000 2.285000 2.465000 ;
      RECT 2.075000  0.085000 2.245000 0.555000 ;
      RECT 2.505000  1.835000 2.755000 2.635000 ;
      RECT 2.975000  1.665000 3.225000 2.465000 ;
      RECT 3.015000  0.085000 3.185000 0.555000 ;
      RECT 3.445000  1.835000 3.695000 2.635000 ;
      RECT 3.915000  1.665000 4.165000 2.295000 ;
      RECT 3.915000  2.295000 7.925000 2.465000 ;
      RECT 3.955000  0.085000 4.125000 0.555000 ;
      RECT 4.855000  1.785000 5.105000 2.295000 ;
      RECT 4.895000  0.085000 5.065000 0.555000 ;
      RECT 5.795000  1.785000 6.045000 2.295000 ;
      RECT 5.835000  0.085000 6.005000 0.555000 ;
      RECT 6.735000  1.785000 6.985000 2.295000 ;
      RECT 6.775000  0.085000 6.945000 0.555000 ;
      RECT 7.675000  1.785000 7.925000 2.295000 ;
      RECT 7.715000  0.085000 8.005000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor2_8
