* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__dlrtp_4 D GATE RESET_B VGND VNB VPB VPWR Q
X0 a_702_413# a_750_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 Q a_750_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_27_363# GATE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X3 VPWR a_604_47# a_750_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_981_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_319_369# D VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_503_369# a_27_363# a_604_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X7 a_604_47# a_27_363# a_708_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VPWR a_750_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND a_319_369# a_500_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 Q a_750_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_750_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VGND a_27_363# a_203_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR a_319_369# a_503_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X14 a_27_363# GATE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 Q a_750_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR a_27_363# a_203_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X17 Q a_750_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR a_750_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_708_47# a_750_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 VGND a_750_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_750_21# a_604_47# a_981_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_500_47# a_203_47# a_604_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 a_319_369# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X24 a_604_47# a_203_47# a_702_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X25 VGND a_750_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
