* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfstp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 VGND a_693_369# a_877_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X2 a_1467_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_119_47# SCE a_201_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 VPWR a_2381_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_1075_413# a_877_369# a_1177_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VPWR SET_B a_1725_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X7 a_2381_47# a_1725_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X8 VGND a_1725_329# a_1921_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_201_47# a_349_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 a_211_369# D a_201_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X11 a_349_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X12 a_1075_413# a_693_369# a_1169_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 a_693_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_2027_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 a_1841_413# a_1921_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X16 a_201_47# a_877_369# a_1075_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X17 a_349_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1229_21# a_1075_413# a_1467_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1169_413# a_1229_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X20 a_201_47# a_693_369# a_1075_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR SCE a_211_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X22 VGND SCD a_119_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 a_1725_329# a_693_369# a_1955_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X24 VPWR a_693_369# a_877_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X25 VPWR a_1075_413# a_1229_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X26 a_295_47# a_349_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_1177_47# a_1229_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_1955_47# a_1921_295# a_2027_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_1075_413# a_1643_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X30 a_1725_329# a_877_369# a_1841_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X31 a_693_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X32 VGND a_1075_413# a_1645_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X33 a_201_47# D a_295_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 a_1229_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X35 a_2381_47# a_1725_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 VGND a_2381_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR a_1725_329# a_1921_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X38 a_1645_47# a_877_369# a_1725_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X39 a_1643_329# a_693_369# a_1725_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
.ends
