* File: sky130_fd_sc_hdll__nand3_2.pex.spice
* Created: Thu Aug 27 19:13:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%A 1 3 4 6 7 9 10 12 13 20
r44 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r45 19 20 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r46 18 19 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r47 16 18 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.495 $Y2=1.202
r48 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r49 10 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r51 7 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r53 4 19 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r54 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r55 1 18 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%B 1 3 6 8 10 13 15 16 17 24 31 35 38
c49 6 0 8.62605e-20 $X=1.46 $Y=0.56
c50 1 0 1.55098e-19 $X=1.435 $Y=1.41
r51 27 31 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=1.97 $Y=1.175
+ $X2=1.615 $Y2=1.175
r52 26 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r53 24 26 5.7381 $w=3.36e-07 $l=4e-08 $layer=POLY_cond $X=1.93 $Y=1.212 $X2=1.97
+ $Y2=1.212
r54 23 24 3.58631 $w=3.36e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.212
+ $X2=1.93 $Y2=1.212
r55 22 23 63.8363 $w=3.36e-07 $l=4.45e-07 $layer=POLY_cond $X=1.46 $Y=1.212
+ $X2=1.905 $Y2=1.212
r56 21 22 3.58631 $w=3.36e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.212
+ $X2=1.46 $Y2=1.212
r57 17 38 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=2.485 $Y=1.175
+ $X2=2.505 $Y2=1.175
r58 17 35 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=2.485 $Y=1.175
+ $X2=2.075 $Y2=1.175
r59 16 35 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=2.065 $Y=1.175
+ $X2=2.075 $Y2=1.175
r60 16 27 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=2.065 $Y=1.175
+ $X2=1.97 $Y2=1.175
r61 15 31 1.10909 $w=1.98e-07 $l=2e-08 $layer=LI1_cond $X=1.595 $Y=1.175
+ $X2=1.615 $Y2=1.175
r62 11 24 21.6522 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.93 $Y=1.015
+ $X2=1.93 $Y2=1.212
r63 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.93 $Y=1.015
+ $X2=1.93 $Y2=0.56
r64 8 23 17.3521 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.212
r65 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r66 4 22 21.6522 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.46 $Y=1.015
+ $X2=1.46 $Y2=1.212
r67 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.46 $Y=1.015
+ $X2=1.46 $Y2=0.56
r68 1 21 17.3521 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r69 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%C 3 5 7 8 10 11 13 14 15 16 23 30 33
r41 23 25 9.13411 $w=3.43e-07 $l=6.5e-08 $layer=POLY_cond $X=3.365 $Y=1.21
+ $X2=3.43 $Y2=1.21
r42 22 23 3.51312 $w=3.43e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.21
+ $X2=3.365 $Y2=1.21
r43 21 22 62.5335 $w=3.43e-07 $l=4.45e-07 $layer=POLY_cond $X=2.895 $Y=1.21
+ $X2=3.34 $Y2=1.21
r44 20 21 3.51312 $w=3.43e-07 $l=2.5e-08 $layer=POLY_cond $X=2.87 $Y=1.21
+ $X2=2.895 $Y2=1.21
r45 16 33 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.47 $Y2=1.175
r46 15 33 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=3.43 $Y=1.175 $X2=3.47
+ $Y2=1.175
r47 15 30 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=3.43 $Y=1.175
+ $X2=3.015 $Y2=1.175
r48 15 25 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.43
+ $Y=1.16 $X2=3.43 $Y2=1.16
r49 14 30 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.01 $Y=1.175
+ $X2=3.015 $Y2=1.175
r50 11 23 17.8339 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.21
r51 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r52 8 22 22.1447 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.34 $Y=1.01 $X2=3.34
+ $Y2=1.21
r53 8 10 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=3.34 $Y=1.01 $X2=3.34
+ $Y2=0.56
r54 5 21 17.8339 $w=1.8e-07 $l=2e-07 $layer=POLY_cond $X=2.895 $Y=1.41 $X2=2.895
+ $Y2=1.21
r55 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r56 1 20 22.1447 $w=1.5e-07 $l=1.95e-07 $layer=POLY_cond $X=2.87 $Y=1.015
+ $X2=2.87 $Y2=1.21
r57 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.87 $Y=1.015
+ $X2=2.87 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%VPWR 1 2 3 4 5 16 18 22 26 28 32 35 37 41
+ 43 52 55 61
r57 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 56 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 55 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r61 53 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r63 47 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 47 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r65 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 44 55 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.4 $Y2=2.72
r67 44 46 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 43 60 4.92749 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.827 $Y2=2.72
r69 43 46 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r70 41 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r71 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 37 40 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.705 $Y=1.66
+ $X2=3.705 $Y2=2.34
r73 35 60 3.2692 $w=3.8e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.705 $Y=2.635
+ $X2=3.827 $Y2=2.72
r74 35 40 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.705 $Y=2.635
+ $X2=3.705 $Y2=2.34
r75 30 55 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.4 $Y=2.635 $X2=2.4
+ $Y2=2.72
r76 30 32 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=2.4 $Y=2.635
+ $X2=2.4 $Y2=2
r77 29 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r78 28 55 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.4 $Y2=2.72
r79 28 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r80 24 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r81 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r82 23 49 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r83 22 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72 $X2=1.2
+ $Y2=2.72
r84 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r85 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r86 16 49 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r87 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r88 5 40 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.63 $Y2=2.34
r89 5 37 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.63 $Y2=1.66
r90 4 32 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=2
r91 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r92 2 26 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r93 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r94 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%Y 1 2 3 4 15 17 21 23 25 27 30 33 34 35 42
c70 42 0 2.41359e-19 $X=0.73 $Y=0.72
r71 34 35 6.69888 $w=5.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.705 $Y=1.19
+ $X2=0.705 $Y2=1.445
r72 33 34 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=0.705 $Y=0.85
+ $X2=0.705 $Y2=1.19
r73 33 42 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=0.705 $Y=0.85
+ $X2=0.705 $Y2=0.72
r74 25 32 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=3.105 $Y=1.665
+ $X2=3.105 $Y2=1.555
r75 25 27 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.105 $Y=1.665
+ $X2=3.105 $Y2=2.34
r76 24 30 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.645 $Y2=1.555
r77 23 32 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.915 $Y=1.555
+ $X2=3.105 $Y2=1.555
r78 23 24 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=2.915 $Y=1.555
+ $X2=1.835 $Y2=1.555
r79 19 30 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.555
r80 19 21 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r81 18 35 3.36699 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.555
+ $X2=0.705 $Y2=1.555
r82 17 30 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=1.645 $Y2=1.555
r83 17 18 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=0.895 $Y2=1.555
r84 13 35 3.21057 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.555
r85 13 15 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r86 4 32 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.66
r87 4 27 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.34
r88 3 30 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r89 3 21 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r90 2 35 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r91 2 15 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r92 1 42 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%A_27_47# 1 2 3 10 13 17
r27 15 17 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=0.38 $X2=2.14
+ $Y2=0.38
r28 13 15 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=0.38
+ $X2=1.2 $Y2=0.38
r29 10 13 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.345 $Y2=0.38
r30 10 12 2.15294 $w=2.55e-07 $l=4.5e-08 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.51
r31 3 17 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r32 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r33 1 12 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%A_307_47# 1 2 11
r23 8 11 62.3173 $w=2.68e-07 $l=1.46e-06 $layer=LI1_cond $X=1.67 $Y=0.77
+ $X2=3.13 $Y2=0.77
r24 2 11 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.13 $Y2=0.72
r25 1 8 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_2%VGND 1 2 9 11 13 15 17 22 28 32
r42 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r43 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r44 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r45 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r46 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r47 23 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=2.66
+ $Y2=0
r48 23 25 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.825 $Y=0 $X2=3.45
+ $Y2=0
r49 22 31 4.92749 $w=1.7e-07 $l=3.12e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.827
+ $Y2=0
r50 22 25 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.45
+ $Y2=0
r51 17 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.495 $Y=0 $X2=2.66
+ $Y2=0
r52 17 19 147.77 $w=1.68e-07 $l=2.265e-06 $layer=LI1_cond $X=2.495 $Y=0 $X2=0.23
+ $Y2=0
r53 15 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r54 15 19 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r55 11 31 3.2692 $w=3.8e-07 $l=1.58915e-07 $layer=LI1_cond $X=3.705 $Y=0.085
+ $X2=3.827 $Y2=0
r56 11 13 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.705 $Y=0.085
+ $X2=3.705 $Y2=0.38
r57 7 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085 $X2=2.66
+ $Y2=0
r58 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.38
r59 2 13 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.235 $X2=3.63 $Y2=0.38
r60 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.66 $Y2=0.38
.ends

