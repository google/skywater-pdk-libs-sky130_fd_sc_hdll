# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o31ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.930000 1.425000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.055000 4.005000 1.425000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.055000 6.590000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.165000 1.055000 8.585000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.851000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.175000 1.445000 8.625000 1.695000 ;
        RECT 6.420000 1.695000 6.590000 2.465000 ;
        RECT 6.760000 0.645000 8.080000 0.885000 ;
        RECT 6.760000 0.885000 6.995000 1.445000 ;
        RECT 7.360000 1.695000 7.530000 2.465000 ;
        RECT 8.300000 1.695000 8.625000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.090000  0.255000 0.445000 0.715000 ;
      RECT 0.090000  0.715000 6.590000 0.885000 ;
      RECT 0.090000  1.595000 2.325000 1.895000 ;
      RECT 0.090000  1.895000 0.445000 2.465000 ;
      RECT 0.665000  0.085000 0.835000 0.545000 ;
      RECT 0.665000  2.065000 0.835000 2.635000 ;
      RECT 1.005000  0.255000 1.385000 0.715000 ;
      RECT 1.005000  1.895000 1.385000 2.465000 ;
      RECT 1.605000  0.085000 1.775000 0.545000 ;
      RECT 1.605000  2.065000 1.775000 2.635000 ;
      RECT 1.945000  0.255000 2.325000 0.715000 ;
      RECT 1.945000  1.895000 2.325000 2.205000 ;
      RECT 1.945000  2.205000 4.285000 2.465000 ;
      RECT 2.545000  0.085000 2.715000 0.545000 ;
      RECT 2.545000  1.595000 4.005000 1.765000 ;
      RECT 2.545000  1.765000 2.715000 2.035000 ;
      RECT 2.885000  0.255000 3.265000 0.715000 ;
      RECT 2.885000  1.935000 3.265000 2.205000 ;
      RECT 3.485000  0.085000 3.655000 0.545000 ;
      RECT 3.485000  1.765000 4.005000 1.865000 ;
      RECT 3.485000  1.865000 6.200000 2.035000 ;
      RECT 3.825000  0.255000 4.205000 0.715000 ;
      RECT 4.445000  0.085000 5.140000 0.545000 ;
      RECT 4.530000  2.035000 6.200000 2.465000 ;
      RECT 5.360000  0.395000 5.530000 0.715000 ;
      RECT 5.790000  0.085000 6.160000 0.545000 ;
      RECT 6.420000  0.255000 8.585000 0.475000 ;
      RECT 6.420000  0.475000 6.590000 0.715000 ;
      RECT 6.760000  1.890000 7.140000 2.635000 ;
      RECT 7.700000  1.890000 8.080000 2.635000 ;
      RECT 8.300000  0.475000 8.585000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o31ai_4
