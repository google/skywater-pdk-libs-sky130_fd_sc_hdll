* File: sky130_fd_sc_hdll__muxb8to1_1.pex.spice
* Created: Thu Aug 27 19:12:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[0] 1 3 4 6 8 13 15
c28 4 0 5.33021e-20 $X=0.495 $Y=1.41
r29 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=0.51
+ $X2=0.645 $Y2=0.51
r30 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.5 $Y=1.19
+ $X2=0.645 $Y2=1.19
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=1.16 $X2=0.5 $Y2=1.16
r32 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.645 $Y=1.055
+ $X2=0.645 $Y2=1.19
r33 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=0.51
r34 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=1.055
r35 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.5 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r37 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.5 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_184_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=1.545 $Y=1.405
+ $X2=1.775 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=1.325 $Y=1.34
+ $X2=1.02 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=1.325 $Y=1.405
+ $X2=1.545 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.34 $X2=1.325 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.775 $Y=2.31
+ $X2=1.775 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.545 $Y=1.175
+ $X2=1.545 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.775 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.545 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.02 $Y=1.475
+ $X2=1.02 $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.02 $Y=1.475 $X2=1.02
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.235 $X2=1.775 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[0] 1 3 4 5 6 8 9 11 12 17
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.03 $X2=1.975 $Y2=1.03
r48 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=1.975 $Y=0.905
+ $X2=1.975 $Y2=1.03
r49 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.005 $Y=1.19
+ $X2=2.005 $Y2=1.03
r50 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=1.975 $Y2=0.905
r51 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=2.01 $Y2=0.495
r52 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.01 $Y=1.41
+ $X2=1.975 $Y2=1.03
r53 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=1.41 $X2=2.01
+ $Y2=1.985
r54 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.84 $Y=0.905
+ $X2=1.975 $Y2=0.905
r55 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.84 $Y=0.905 $X2=1.02
+ $Y2=0.905
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=1.02 $Y2=0.905
r57 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=0.945 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[1] 1 3 4 6 7 9 11 12 17
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.03 $X2=2.625 $Y2=1.03
r45 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=2.625 $Y=0.905
+ $X2=2.625 $Y2=1.03
r46 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=2.595 $Y=1.19
+ $X2=2.595 $Y2=1.03
r47 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.655 $Y=0.83
+ $X2=3.655 $Y2=0.495
r48 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=0.905
+ $X2=2.625 $Y2=0.905
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.58 $Y=0.905
+ $X2=3.655 $Y2=0.83
r50 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.58 $Y=0.905 $X2=2.76
+ $Y2=0.905
r51 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.59 $Y=0.83
+ $X2=2.625 $Y2=0.905
r52 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.59 $Y=0.83 $X2=2.59
+ $Y2=0.495
r53 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.59 $Y=1.41
+ $X2=2.625 $Y2=1.03
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.59 $Y=1.41 $X2=2.59
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_533_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=3.275 $Y=1.34
+ $X2=3.58 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.275
+ $Y=1.34 $X2=3.275 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=3.055 $Y=1.405
+ $X2=3.275 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=2.825 $Y=1.63
+ $X2=3.055 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.055 $Y=1.175
+ $X2=3.055 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=2.825 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=3.055 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.825 $Y=2.31
+ $X2=2.825 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=3.58 $Y=1.475
+ $X2=3.58 $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=3.58 $Y=1.475 $X2=3.58
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.825 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[1] 1 3 4 6 8 12 15 21
c37 8 0 1.78369e-19 $X=3.955 $Y=1.055
c38 1 0 2.31671e-19 $X=4.105 $Y=1.41
r39 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.91 $Y=0.51
+ $X2=3.955 $Y2=0.51
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.16 $X2=4.1 $Y2=1.16
r41 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.955 $Y=1.19
+ $X2=4.1 $Y2=1.19
r42 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=1.055
+ $X2=3.955 $Y2=1.19
r43 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=1.055
r45 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.13 $Y=0.995
+ $X2=4.1 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.995 $X2=4.13
+ $Y2=0.56
r47 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.1 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.105 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[2] 1 3 4 6 8 13 15
c37 8 0 1.78369e-19 $X=4.785 $Y=1.055
c38 4 0 2.31671e-19 $X=4.635 $Y=1.41
r39 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.83 $Y=0.51
+ $X2=4.785 $Y2=0.51
r40 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.64 $Y=1.19
+ $X2=4.785 $Y2=1.19
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.16 $X2=4.64 $Y2=1.16
r42 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.785 $Y=1.055
+ $X2=4.785 $Y2=1.19
r43 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=1.055
r45 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.64 $Y2=1.16
r46 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.635 $Y2=1.985
r47 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.61 $Y=0.995
+ $X2=4.64 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.61 $Y=0.995 $X2=4.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1012_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=5.685 $Y=1.405
+ $X2=5.915 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=5.465 $Y=1.34
+ $X2=5.16 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=5.465 $Y=1.405
+ $X2=5.685 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=1.34 $X2=5.465 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.915 $Y=2.31
+ $X2=5.915 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=1.175
+ $X2=5.685 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.915 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.685 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.16 $Y=1.475
+ $X2=5.16 $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=5.16 $Y=1.475 $X2=5.16
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.235 $X2=5.915 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[2] 1 3 4 5 6 8 9 11 12 17
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=1.03 $X2=6.115 $Y2=1.03
r48 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.115 $Y=0.905
+ $X2=6.115 $Y2=1.03
r49 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.145 $Y=1.19
+ $X2=6.145 $Y2=1.03
r50 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.115 $Y2=0.905
r51 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.15 $Y2=0.495
r52 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.15 $Y=1.41
+ $X2=6.115 $Y2=1.03
r53 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.15 $Y=1.41 $X2=6.15
+ $Y2=1.985
r54 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.98 $Y=0.905
+ $X2=6.115 $Y2=0.905
r55 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.98 $Y=0.905 $X2=5.16
+ $Y2=0.905
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.16 $Y2=0.905
r57 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.085 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[3] 1 3 4 6 7 9 11 12 17
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.765
+ $Y=1.03 $X2=6.765 $Y2=1.03
r45 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.765 $Y=0.905
+ $X2=6.765 $Y2=1.03
r46 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=6.735 $Y=1.19
+ $X2=6.735 $Y2=1.03
r47 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.795 $Y=0.83
+ $X2=7.795 $Y2=0.495
r48 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.9 $Y=0.905
+ $X2=6.765 $Y2=0.905
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=0.905
+ $X2=7.795 $Y2=0.83
r50 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.72 $Y=0.905 $X2=6.9
+ $Y2=0.905
r51 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.73 $Y=0.83
+ $X2=6.765 $Y2=0.905
r52 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.73 $Y=0.83 $X2=6.73
+ $Y2=0.495
r53 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.73 $Y=1.41
+ $X2=6.765 $Y2=1.03
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=1.41 $X2=6.73
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1361_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=7.415 $Y=1.34
+ $X2=7.72 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=1.34 $X2=7.415 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=7.195 $Y=1.405
+ $X2=7.415 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=6.965 $Y=1.63
+ $X2=7.195 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.195 $Y=1.175
+ $X2=7.195 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=6.965 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=7.195 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.965 $Y=2.31
+ $X2=6.965 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.72 $Y=1.475
+ $X2=7.72 $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.72 $Y=1.475 $X2=7.72
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.235 $X2=6.965 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[3] 1 3 4 6 8 12 15 21
c37 8 0 1.78369e-19 $X=8.095 $Y=1.055
c38 1 0 2.31671e-19 $X=8.245 $Y=1.41
r39 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.05 $Y=0.51
+ $X2=8.095 $Y2=0.51
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.24
+ $Y=1.16 $X2=8.24 $Y2=1.16
r41 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.095 $Y=1.19
+ $X2=8.24 $Y2=1.19
r42 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.095 $Y=1.055
+ $X2=8.095 $Y2=1.19
r43 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=1.055
r45 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.27 $Y=0.995
+ $X2=8.24 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.27 $Y=0.995 $X2=8.27
+ $Y2=0.56
r47 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.24 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.245 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[4] 1 3 4 6 8 13 15
c37 8 0 1.78369e-19 $X=8.925 $Y=1.055
c38 4 0 2.31671e-19 $X=8.775 $Y=1.41
r39 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.97 $Y=0.51
+ $X2=8.925 $Y2=0.51
r40 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.78 $Y=1.19
+ $X2=8.925 $Y2=1.19
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.78
+ $Y=1.16 $X2=8.78 $Y2=1.16
r42 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.925 $Y=1.055
+ $X2=8.925 $Y2=1.19
r43 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.925 $Y=0.625
+ $X2=8.925 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.925 $Y=0.625
+ $X2=8.925 $Y2=1.055
r45 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.775 $Y=1.41
+ $X2=8.78 $Y2=1.16
r46 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.775 $Y=1.41
+ $X2=8.775 $Y2=1.985
r47 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.75 $Y=0.995
+ $X2=8.78 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.75 $Y=0.995 $X2=8.75
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1840_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=9.825 $Y=1.405
+ $X2=10.055 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=9.605 $Y=1.34
+ $X2=9.3 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=9.605 $Y=1.405
+ $X2=9.825 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.605
+ $Y=1.34 $X2=9.605 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.055 $Y=2.31
+ $X2=10.055 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=9.825 $Y=1.175
+ $X2=9.825 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=9.825 $Y=0.755
+ $X2=10.055 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=9.825 $Y=0.755
+ $X2=9.825 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=9.3 $Y=1.475 $X2=9.3
+ $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=9.3 $Y=1.475 $X2=9.3
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.485 $X2=10.055 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=9.93
+ $Y=1.485 $X2=10.055 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.93
+ $Y=0.235 $X2=10.055 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[4] 1 3 4 5 6 8 9 11 12 17
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.255
+ $Y=1.03 $X2=10.255 $Y2=1.03
r48 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.255 $Y=0.905
+ $X2=10.255 $Y2=1.03
r49 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.285 $Y=1.19
+ $X2=10.285 $Y2=1.03
r50 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.29 $Y=0.83
+ $X2=10.255 $Y2=0.905
r51 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.29 $Y=0.83
+ $X2=10.29 $Y2=0.495
r52 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.29 $Y=1.41
+ $X2=10.255 $Y2=1.03
r53 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.29 $Y=1.41
+ $X2=10.29 $Y2=1.985
r54 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.12 $Y=0.905
+ $X2=10.255 $Y2=0.905
r55 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=10.12 $Y=0.905 $X2=9.3
+ $Y2=0.905
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=9.225 $Y=0.83
+ $X2=9.3 $Y2=0.905
r57 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.225 $Y=0.83
+ $X2=9.225 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[5] 1 3 4 6 7 9 11 12 17
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.905
+ $Y=1.03 $X2=10.905 $Y2=1.03
r45 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=10.905 $Y=0.905
+ $X2=10.905 $Y2=1.03
r46 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=10.875 $Y=1.19
+ $X2=10.875 $Y2=1.03
r47 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.935 $Y=0.83
+ $X2=11.935 $Y2=0.495
r48 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.04 $Y=0.905
+ $X2=10.905 $Y2=0.905
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.86 $Y=0.905
+ $X2=11.935 $Y2=0.83
r50 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=11.86 $Y=0.905
+ $X2=11.04 $Y2=0.905
r51 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=10.87 $Y=0.83
+ $X2=10.905 $Y2=0.905
r52 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.87 $Y=0.83
+ $X2=10.87 $Y2=0.495
r53 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=10.87 $Y=1.41
+ $X2=10.905 $Y2=1.03
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.87 $Y=1.41
+ $X2=10.87 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2189_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=11.555 $Y=1.34
+ $X2=11.86 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.555
+ $Y=1.34 $X2=11.555 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=11.335 $Y=1.405
+ $X2=11.555 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=11.105 $Y=1.63
+ $X2=11.335 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=11.335 $Y=1.175
+ $X2=11.335 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=11.335 $Y=0.755
+ $X2=11.105 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=11.335 $Y=0.755
+ $X2=11.335 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.105 $Y=2.31
+ $X2=11.105 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.86 $Y=1.475
+ $X2=11.86 $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.86 $Y=1.475 $X2=11.86
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=1.485 $X2=11.105 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.96
+ $Y=1.485 $X2=11.105 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=10.945
+ $Y=0.235 $X2=11.105 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[5] 1 3 4 6 8 12 15 21
c37 8 0 1.78369e-19 $X=12.235 $Y=1.055
c38 1 0 2.31671e-19 $X=12.385 $Y=1.41
r39 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=12.19 $Y=0.51
+ $X2=12.235 $Y2=0.51
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.38
+ $Y=1.16 $X2=12.38 $Y2=1.16
r41 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.235 $Y=1.19
+ $X2=12.38 $Y2=1.19
r42 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.235 $Y=1.055
+ $X2=12.235 $Y2=1.19
r43 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=12.235 $Y=0.625
+ $X2=12.235 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=12.235 $Y=0.625
+ $X2=12.235 $Y2=1.055
r45 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.38 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.41 $Y=0.995
+ $X2=12.41 $Y2=0.56
r47 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.385 $Y=1.41
+ $X2=12.38 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.385 $Y=1.41
+ $X2=12.385 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[6] 1 3 4 6 8 13 15
c37 8 0 1.78369e-19 $X=13.065 $Y=1.055
c38 4 0 2.31671e-19 $X=12.915 $Y=1.41
r39 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=13.11 $Y=0.51
+ $X2=13.065 $Y2=0.51
r40 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=12.92 $Y=1.19
+ $X2=13.065 $Y2=1.19
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.92
+ $Y=1.16 $X2=12.92 $Y2=1.16
r42 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.065 $Y=1.055
+ $X2=13.065 $Y2=1.19
r43 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.065 $Y=0.625
+ $X2=13.065 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=13.065 $Y=0.625
+ $X2=13.065 $Y2=1.055
r45 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.92 $Y2=1.16
r46 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.915 $Y=1.41
+ $X2=12.915 $Y2=1.985
r47 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=12.89 $Y=0.995
+ $X2=12.92 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.89 $Y=0.995
+ $X2=12.89 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2668_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=13.965 $Y=1.405
+ $X2=14.195 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=13.745 $Y=1.34
+ $X2=13.44 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=13.745 $Y=1.405
+ $X2=13.965 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.745
+ $Y=1.34 $X2=13.745 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.195 $Y=2.31
+ $X2=14.195 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=13.965 $Y=1.175
+ $X2=13.965 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=13.965 $Y=0.755
+ $X2=14.195 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.965 $Y=0.755
+ $X2=13.965 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.44 $Y=1.475
+ $X2=13.44 $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=13.44 $Y=1.475 $X2=13.44
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.485 $X2=14.195 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=14.07
+ $Y=1.485 $X2=14.195 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=14.07
+ $Y=0.235 $X2=14.195 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[6] 1 3 4 5 6 8 9 11 12 17
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.395
+ $Y=1.03 $X2=14.395 $Y2=1.03
r48 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=14.395 $Y=0.905
+ $X2=14.395 $Y2=1.03
r49 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=14.425 $Y=1.19
+ $X2=14.425 $Y2=1.03
r50 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=14.43 $Y=0.83
+ $X2=14.395 $Y2=0.905
r51 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=14.43 $Y=0.83
+ $X2=14.43 $Y2=0.495
r52 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=14.43 $Y=1.41
+ $X2=14.395 $Y2=1.03
r53 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.43 $Y=1.41
+ $X2=14.43 $Y2=1.985
r54 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=14.26 $Y=0.905
+ $X2=14.395 $Y2=0.905
r55 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=14.26 $Y=0.905
+ $X2=13.44 $Y2=0.905
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.365 $Y=0.83
+ $X2=13.44 $Y2=0.905
r57 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=13.365 $Y=0.83
+ $X2=13.365 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[7] 1 3 4 6 7 9 11 12 17
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.045
+ $Y=1.03 $X2=15.045 $Y2=1.03
r45 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=15.045 $Y=0.905
+ $X2=15.045 $Y2=1.03
r46 12 17 4.60977 $w=3.98e-07 $l=1.6e-07 $layer=LI1_cond $X=15.015 $Y=1.19
+ $X2=15.015 $Y2=1.03
r47 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.075 $Y=0.83
+ $X2=16.075 $Y2=0.495
r48 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.18 $Y=0.905
+ $X2=15.045 $Y2=0.905
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16 $Y=0.905
+ $X2=16.075 $Y2=0.83
r50 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=16 $Y=0.905 $X2=15.18
+ $Y2=0.905
r51 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=15.01 $Y=0.83
+ $X2=15.045 $Y2=0.905
r52 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.01 $Y=0.83
+ $X2=15.01 $Y2=0.495
r53 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=15.01 $Y=1.41
+ $X2=15.045 $Y2=1.03
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.01 $Y=1.41
+ $X2=15.01 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_3017_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=15.695 $Y=1.34
+ $X2=16 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.695
+ $Y=1.34 $X2=15.695 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=15.475 $Y=1.405
+ $X2=15.695 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=15.245 $Y=1.63
+ $X2=15.475 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=15.475 $Y=1.175
+ $X2=15.475 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=15.475 $Y=0.755
+ $X2=15.245 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=15.475 $Y=0.755
+ $X2=15.475 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.245 $Y=2.31
+ $X2=15.245 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=16 $Y=1.475 $X2=16
+ $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=16 $Y=1.475 $X2=16
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=1.485 $X2=15.245 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=15.1
+ $Y=1.485 $X2=15.245 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=15.085
+ $Y=0.235 $X2=15.245 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[7] 1 3 4 6 8 12 15 21
c28 1 0 5.33021e-20 $X=16.525 $Y=1.41
r29 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=16.33 $Y=0.51
+ $X2=16.375 $Y2=0.51
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.52
+ $Y=1.16 $X2=16.52 $Y2=1.16
r31 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=16.375 $Y=1.19
+ $X2=16.52 $Y2=1.19
r32 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.375 $Y=1.055
+ $X2=16.375 $Y2=1.19
r33 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.375 $Y=0.625
+ $X2=16.375 $Y2=0.51
r34 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=16.375 $Y=0.625
+ $X2=16.375 $Y2=1.055
r35 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=16.55 $Y=0.995
+ $X2=16.52 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.55 $Y=0.995
+ $X2=16.55 $Y2=0.56
r37 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.525 $Y=1.41
+ $X2=16.52 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.525 $Y=1.41
+ $X2=16.525 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VPWR 1 2 3 4 5 6 7 8 9 28 30 36 42 48
+ 54 60 66 72 76 78 83 84 86 87 89 90 92 93 94 95 96 97 98 111 125 139 153 164
+ 167 170
r265 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r266 156 159 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=14.95 $Y=2.72
+ $X2=16.33 $Y2=2.72
r267 155 158 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=14.95 $Y=2.72
+ $X2=16.33 $Y2=2.72
r268 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r269 153 173 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=16.595 $Y=2.72
+ $X2=16.807 $Y2=2.72
r270 153 158 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=16.595 $Y=2.72
+ $X2=16.33 $Y2=2.72
r271 152 156 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r272 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r273 149 152 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=14.49 $Y2=2.72
r274 148 151 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=13.11 $Y=2.72
+ $X2=14.49 $Y2=2.72
r275 148 149 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r276 146 170 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.845 $Y=2.72
+ $X2=12.65 $Y2=2.72
r277 146 148 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.845 $Y=2.72
+ $X2=13.11 $Y2=2.72
r278 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r279 142 145 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=12.19 $Y2=2.72
r280 141 144 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=2.72
+ $X2=12.19 $Y2=2.72
r281 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r282 139 170 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=12.455 $Y=2.72
+ $X2=12.65 $Y2=2.72
r283 139 144 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=12.455 $Y=2.72
+ $X2=12.19 $Y2=2.72
r284 138 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r285 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r286 135 138 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=10.35 $Y2=2.72
r287 134 137 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=10.35 $Y2=2.72
r288 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r289 132 167 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.705 $Y=2.72
+ $X2=8.51 $Y2=2.72
r290 132 134 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.705 $Y=2.72
+ $X2=8.97 $Y2=2.72
r291 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r292 128 131 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r293 127 130 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r294 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r295 125 167 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.51 $Y2=2.72
r296 125 130 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.05 $Y2=2.72
r297 124 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r298 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r299 121 124 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r300 120 123 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r301 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r302 118 164 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.37 $Y2=2.72
r303 118 120 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.83 $Y2=2.72
r304 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r305 114 117 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r306 113 116 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r307 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r308 111 164 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=4.37 $Y2=2.72
r309 111 116 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=3.91 $Y2=2.72
r310 110 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r311 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r312 107 110 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r313 106 109 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r314 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r315 104 161 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r316 104 106 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r317 98 159 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.79 $Y=2.72
+ $X2=16.33 $Y2=2.72
r318 98 173 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.79 $Y=2.72
+ $X2=16.79 $Y2=2.72
r319 97 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r320 97 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r321 97 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r322 96 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r323 96 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r324 96 167 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r325 95 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r326 95 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r327 95 164 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r328 94 107 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r329 94 161 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r330 92 151 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.555 $Y=2.72
+ $X2=14.49 $Y2=2.72
r331 92 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.555 $Y=2.72
+ $X2=14.72 $Y2=2.72
r332 91 155 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=14.95 $Y2=2.72
r333 91 93 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.885 $Y=2.72
+ $X2=14.72 $Y2=2.72
r334 89 137 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.35 $Y2=2.72
r335 89 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.58 $Y2=2.72
r336 88 141 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.745 $Y=2.72
+ $X2=10.81 $Y2=2.72
r337 88 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=2.72
+ $X2=10.58 $Y2=2.72
r338 86 123 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.21 $Y2=2.72
r339 86 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.44 $Y2=2.72
r340 85 127 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.67 $Y2=2.72
r341 85 87 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.44 $Y2=2.72
r342 83 109 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.07 $Y2=2.72
r343 83 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=2.72
+ $X2=2.3 $Y2=2.72
r344 82 113 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.53 $Y2=2.72
r345 82 84 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.3 $Y2=2.72
r346 78 81 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.76 $Y=1.66
+ $X2=16.76 $Y2=2.34
r347 76 173 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=16.76 $Y=2.635
+ $X2=16.807 $Y2=2.72
r348 76 81 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=16.76 $Y=2.635
+ $X2=16.76 $Y2=2.34
r349 72 75 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=14.72 $Y=1.63
+ $X2=14.72 $Y2=2.31
r350 70 93 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=2.635
+ $X2=14.72 $Y2=2.72
r351 70 75 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=14.72 $Y=2.635
+ $X2=14.72 $Y2=2.31
r352 66 69 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=12.65 $Y=1.66
+ $X2=12.65 $Y2=2.34
r353 64 170 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=2.635
+ $X2=12.65 $Y2=2.72
r354 64 69 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=12.65 $Y=2.635
+ $X2=12.65 $Y2=2.34
r355 60 63 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=10.58 $Y=1.63
+ $X2=10.58 $Y2=2.31
r356 58 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=2.635
+ $X2=10.58 $Y2=2.72
r357 58 63 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=10.58 $Y=2.635
+ $X2=10.58 $Y2=2.31
r358 54 57 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=8.51 $Y=1.66
+ $X2=8.51 $Y2=2.34
r359 52 167 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=2.635
+ $X2=8.51 $Y2=2.72
r360 52 57 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=8.51 $Y=2.635
+ $X2=8.51 $Y2=2.34
r361 48 51 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.44 $Y=1.63
+ $X2=6.44 $Y2=2.31
r362 46 87 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2.72
r363 46 51 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=6.44 $Y=2.635
+ $X2=6.44 $Y2=2.31
r364 42 45 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=4.37 $Y=1.66
+ $X2=4.37 $Y2=2.34
r365 40 164 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.72
r366 40 45 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.34
r367 36 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=2.3 $Y=1.63 $X2=2.3
+ $Y2=2.31
r368 34 84 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=2.635 $X2=2.3
+ $Y2=2.72
r369 34 39 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=2.3 $Y=2.635
+ $X2=2.3 $Y2=2.31
r370 30 33 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r371 28 161 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r372 28 33 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r373 9 81 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=1.485 $X2=16.76 $Y2=2.34
r374 9 78 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=16.615
+ $Y=1.485 $X2=16.76 $Y2=1.66
r375 8 75 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.485 $X2=14.72 $Y2=2.31
r376 8 72 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=14.52
+ $Y=1.485 $X2=14.72 $Y2=1.63
r377 7 69 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.65 $Y2=2.34
r378 7 66 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.65 $Y2=1.66
r379 6 63 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=1.485 $X2=10.58 $Y2=2.31
r380 6 60 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=10.38
+ $Y=1.485 $X2=10.58 $Y2=1.63
r381 5 57 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.51 $Y2=2.34
r382 5 54 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.51 $Y2=1.66
r383 4 51 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=2.31
r384 4 48 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=1.63
r385 3 45 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=2.34
r386 3 42 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=1.66
r387 2 39 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=2.31
r388 2 36 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=1.63
r389 1 33 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r390 1 30 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 50 51 53 57 61 65 68 70 71 73 77 81 85 88 90 91 93 97 101 105 108 110 111
+ 113 117 121 125 128 135 143 151 159 161 162 163 164 165 166 167 168 169 170
+ 171 172 173 174 175 176 177 178 179 180 181 182 193 198 203 208 213 218 223
+ 228
c472 159 0 5.33021e-20 $X=16.035 $Y=0.92
c473 151 0 5.33021e-20 $X=11.895 $Y=0.92
c474 143 0 5.33021e-20 $X=7.755 $Y=0.92
c475 135 0 5.33021e-20 $X=3.615 $Y=0.92
c476 111 0 5.33021e-20 $X=13.587 $Y=0.835
c477 91 0 5.33021e-20 $X=9.447 $Y=0.835
c478 71 0 5.33021e-20 $X=5.307 $Y=0.835
c479 51 0 5.33021e-20 $X=1.167 $Y=0.835
r480 228 230 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=15.87 $Y=1.87
+ $X2=16.035 $Y2=1.87
r481 221 223 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=1.87
+ $X2=13.57 $Y2=1.87
r482 218 220 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=11.73 $Y=1.87
+ $X2=11.895 $Y2=1.87
r483 211 213 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=9.265 $Y=1.87
+ $X2=9.43 $Y2=1.87
r484 208 210 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=1.87
+ $X2=7.755 $Y2=1.87
r485 201 203 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=1.87
+ $X2=5.29 $Y2=1.87
r486 198 200 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=1.87
+ $X2=3.615 $Y2=1.87
r487 191 193 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=1.87
+ $X2=1.15 $Y2=1.87
r488 182 228 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=1.87
+ $X2=15.87 $Y2=1.87
r489 181 223 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=1.87
+ $X2=13.57 $Y2=1.87
r490 180 218 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=1.87
+ $X2=11.73 $Y2=1.87
r491 179 213 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=1.87
+ $X2=9.43 $Y2=1.87
r492 178 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=1.87
+ $X2=7.59 $Y2=1.87
r493 177 203 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r494 176 198 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=1.87
+ $X2=3.45 $Y2=1.87
r495 175 193 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r496 174 181 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.715 $Y=1.87
+ $X2=13.57 $Y2=1.87
r497 173 182 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.725 $Y=1.87
+ $X2=15.87 $Y2=1.87
r498 173 174 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=15.725 $Y=1.87
+ $X2=13.715 $Y2=1.87
r499 172 180 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.875 $Y=1.87
+ $X2=11.73 $Y2=1.87
r500 171 181 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=13.425 $Y=1.87
+ $X2=13.57 $Y2=1.87
r501 171 172 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=13.425 $Y=1.87
+ $X2=11.875 $Y2=1.87
r502 170 179 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.575 $Y=1.87
+ $X2=9.43 $Y2=1.87
r503 169 180 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.585 $Y=1.87
+ $X2=11.73 $Y2=1.87
r504 169 170 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=11.585 $Y=1.87
+ $X2=9.575 $Y2=1.87
r505 168 178 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.735 $Y=1.87
+ $X2=7.59 $Y2=1.87
r506 167 179 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.285 $Y=1.87
+ $X2=9.43 $Y2=1.87
r507 167 168 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=9.285 $Y=1.87
+ $X2=7.735 $Y2=1.87
r508 166 177 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r509 165 178 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=7.59 $Y2=1.87
r510 165 166 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=5.435 $Y2=1.87
r511 164 176 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=1.87
+ $X2=3.45 $Y2=1.87
r512 163 177 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r513 163 164 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=3.595 $Y2=1.87
r514 162 175 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r515 161 176 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=3.45 $Y2=1.87
r516 161 162 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=1.295 $Y2=1.87
r517 128 230 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=16.035 $Y=1.755
+ $X2=16.035 $Y2=1.87
r518 127 159 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.035 $Y=1.005
+ $X2=16.035 $Y2=0.92
r519 127 128 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=16.035 $Y=1.005
+ $X2=16.035 $Y2=1.755
r520 123 159 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=15.852 $Y=0.92
+ $X2=16.035 $Y2=0.92
r521 123 125 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=15.852 $Y=0.835
+ $X2=15.852 $Y2=0.495
r522 119 228 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=15.765 $Y=1.87
+ $X2=15.87 $Y2=1.87
r523 119 121 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=15.765 $Y=1.985
+ $X2=15.765 $Y2=2
r524 115 223 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=13.675 $Y=1.87
+ $X2=13.57 $Y2=1.87
r525 115 117 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=13.675 $Y=1.985
+ $X2=13.675 $Y2=2
r526 111 153 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=13.587 $Y=0.92
+ $X2=13.405 $Y2=0.92
r527 111 113 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=13.587 $Y=0.835
+ $X2=13.587 $Y2=0.495
r528 110 221 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=13.405 $Y=1.755
+ $X2=13.405 $Y2=1.87
r529 109 153 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.405 $Y=1.005
+ $X2=13.405 $Y2=0.92
r530 109 110 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=13.405 $Y=1.005
+ $X2=13.405 $Y2=1.755
r531 108 220 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=11.895 $Y=1.755
+ $X2=11.895 $Y2=1.87
r532 107 151 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.895 $Y=1.005
+ $X2=11.895 $Y2=0.92
r533 107 108 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=11.895 $Y=1.005
+ $X2=11.895 $Y2=1.755
r534 103 151 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=11.712 $Y=0.92
+ $X2=11.895 $Y2=0.92
r535 103 105 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=11.712 $Y=0.835
+ $X2=11.712 $Y2=0.495
r536 99 218 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=11.625 $Y=1.87
+ $X2=11.73 $Y2=1.87
r537 99 101 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=11.625 $Y=1.985
+ $X2=11.625 $Y2=2
r538 95 213 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=1.87
+ $X2=9.43 $Y2=1.87
r539 95 97 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=9.535 $Y=1.985
+ $X2=9.535 $Y2=2
r540 91 145 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=9.447 $Y=0.92
+ $X2=9.265 $Y2=0.92
r541 91 93 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=9.447 $Y=0.835
+ $X2=9.447 $Y2=0.495
r542 90 211 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.265 $Y=1.755
+ $X2=9.265 $Y2=1.87
r543 89 145 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.265 $Y=1.005
+ $X2=9.265 $Y2=0.92
r544 89 90 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=9.265 $Y=1.005
+ $X2=9.265 $Y2=1.755
r545 88 210 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.755 $Y=1.755
+ $X2=7.755 $Y2=1.87
r546 87 143 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=0.92
r547 87 88 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=1.755
r548 83 143 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.572 $Y=0.92
+ $X2=7.755 $Y2=0.92
r549 83 85 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=7.572 $Y=0.835
+ $X2=7.572 $Y2=0.495
r550 79 208 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=1.87
+ $X2=7.59 $Y2=1.87
r551 79 81 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.485 $Y=1.985
+ $X2=7.485 $Y2=2
r552 75 203 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=1.87
+ $X2=5.29 $Y2=1.87
r553 75 77 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.395 $Y=1.985
+ $X2=5.395 $Y2=2
r554 71 137 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=5.307 $Y=0.92
+ $X2=5.125 $Y2=0.92
r555 71 73 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.307 $Y=0.835
+ $X2=5.307 $Y2=0.495
r556 70 201 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.125 $Y=1.755
+ $X2=5.125 $Y2=1.87
r557 69 137 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=0.92
r558 69 70 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=1.755
r559 68 200 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.615 $Y=1.755
+ $X2=3.615 $Y2=1.87
r560 67 135 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=0.92
r561 67 68 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=1.755
r562 63 135 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=3.432 $Y=0.92
+ $X2=3.615 $Y2=0.92
r563 63 65 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.432 $Y=0.835
+ $X2=3.432 $Y2=0.495
r564 59 198 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=1.87
+ $X2=3.45 $Y2=1.87
r565 59 61 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.345 $Y=1.985
+ $X2=3.345 $Y2=2
r566 55 193 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=1.87
+ $X2=1.15 $Y2=1.87
r567 55 57 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.255 $Y=1.985
+ $X2=1.255 $Y2=2
r568 51 129 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=1.167 $Y=0.92
+ $X2=0.985 $Y2=0.92
r569 51 53 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=0.835
+ $X2=1.167 $Y2=0.495
r570 50 191 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=1.755
+ $X2=0.985 $Y2=1.87
r571 49 129 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=0.92
r572 49 50 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=1.755
r573 16 121 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=15.64
+ $Y=1.665 $X2=15.765 $Y2=2
r574 15 117 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=13.53
+ $Y=1.665 $X2=13.675 $Y2=2
r575 14 101 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=11.5
+ $Y=1.665 $X2=11.625 $Y2=2
r576 13 97 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=9.39
+ $Y=1.665 $X2=9.535 $Y2=2
r577 12 81 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=1.665 $X2=7.485 $Y2=2
r578 11 77 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=1.665 $X2=5.395 $Y2=2
r579 10 61 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.665 $X2=3.345 $Y2=2
r580 9 57 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.665 $X2=1.255 $Y2=2
r581 8 125 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.74
+ $Y=0.235 $X2=15.865 $Y2=0.495
r582 7 113 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=13.44
+ $Y=0.235 $X2=13.575 $Y2=0.495
r583 6 105 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=11.6
+ $Y=0.235 $X2=11.725 $Y2=0.495
r584 5 93 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.3
+ $Y=0.235 $X2=9.435 $Y2=0.495
r585 4 85 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.585 $Y2=0.495
r586 3 73 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=5.16
+ $Y=0.235 $X2=5.295 $Y2=0.495
r587 2 65 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.445 $Y2=0.495
r588 1 53 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 38 42
+ 46 50 54 58 60 62 65 66 68 69 71 72 74 75 76 77 78 79 80 93 107 121 135 146
+ 149 152
r208 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r209 138 141 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=14.95 $Y=0
+ $X2=16.33 $Y2=0
r210 137 140 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=14.95 $Y=0
+ $X2=16.33 $Y2=0
r211 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r212 135 155 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=16.63 $Y=0
+ $X2=16.825 $Y2=0
r213 135 140 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=16.63 $Y=0
+ $X2=16.33 $Y2=0
r214 134 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r215 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r216 131 134 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=14.49 $Y2=0
r217 130 133 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=13.11 $Y=0
+ $X2=14.49 $Y2=0
r218 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r219 128 152 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.81 $Y=0
+ $X2=12.65 $Y2=0
r220 128 130 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.81 $Y=0
+ $X2=13.11 $Y2=0
r221 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r222 124 127 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=12.19 $Y2=0
r223 123 126 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=10.81 $Y=0
+ $X2=12.19 $Y2=0
r224 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r225 121 152 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=12.49 $Y=0
+ $X2=12.65 $Y2=0
r226 121 126 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=12.49 $Y=0
+ $X2=12.19 $Y2=0
r227 120 124 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r228 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r229 117 120 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r230 116 119 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=10.35 $Y2=0
r231 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r232 114 149 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.51
+ $Y2=0
r233 114 116 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.67 $Y=0 $X2=8.97
+ $Y2=0
r234 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r235 110 113 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r236 109 112 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r237 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r238 107 149 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.51
+ $Y2=0
r239 107 112 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.05
+ $Y2=0
r240 106 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r241 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r242 103 106 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r243 102 105 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r244 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r245 100 146 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.37
+ $Y2=0
r246 100 102 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.83
+ $Y2=0
r247 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r248 96 99 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r249 95 98 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r250 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r251 93 146 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.37
+ $Y2=0
r252 93 98 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=3.91
+ $Y2=0
r253 92 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r254 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r255 89 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r256 88 91 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r257 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r258 86 143 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0
+ $X2=0.195 $Y2=0
r259 86 88 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r260 80 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=16.79 $Y=0
+ $X2=16.33 $Y2=0
r261 80 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.79 $Y=0
+ $X2=16.79 $Y2=0
r262 79 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r263 79 127 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r264 79 152 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r265 78 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.97 $Y2=0
r266 78 113 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r267 78 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r268 77 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=4.83 $Y2=0
r269 77 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r270 77 146 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r271 76 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r272 76 143 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r273 74 133 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.555 $Y=0
+ $X2=14.49 $Y2=0
r274 74 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.555 $Y=0
+ $X2=14.72 $Y2=0
r275 73 137 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.95 $Y2=0
r276 73 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.885 $Y=0
+ $X2=14.72 $Y2=0
r277 71 119 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.35 $Y2=0
r278 71 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.58 $Y2=0
r279 70 123 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=10.745 $Y=0
+ $X2=10.81 $Y2=0
r280 70 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.745 $Y=0
+ $X2=10.58 $Y2=0
r281 68 105 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=0
+ $X2=6.21 $Y2=0
r282 68 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.44
+ $Y2=0
r283 67 109 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=0
+ $X2=6.67 $Y2=0
r284 67 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.44
+ $Y2=0
r285 65 91 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.07
+ $Y2=0
r286 65 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.3
+ $Y2=0
r287 64 95 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.53
+ $Y2=0
r288 64 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.3
+ $Y2=0
r289 60 155 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=16.76 $Y=0.085
+ $X2=16.825 $Y2=0
r290 60 62 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=16.76 $Y=0.085
+ $X2=16.76 $Y2=0.38
r291 56 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.72 $Y=0.085
+ $X2=14.72 $Y2=0
r292 56 58 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=14.72 $Y=0.085
+ $X2=14.72 $Y2=0.495
r293 52 152 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=12.65 $Y=0.085
+ $X2=12.65 $Y2=0
r294 52 54 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=12.65 $Y=0.085
+ $X2=12.65 $Y2=0.38
r295 48 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.58 $Y=0.085
+ $X2=10.58 $Y2=0
r296 48 50 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=10.58 $Y=0.085
+ $X2=10.58 $Y2=0.495
r297 44 149 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.51 $Y=0.085
+ $X2=8.51 $Y2=0
r298 44 46 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=8.51 $Y=0.085
+ $X2=8.51 $Y2=0.38
r299 40 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0
r300 40 42 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.495
r301 36 146 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0
r302 36 38 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0.38
r303 32 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.085 $X2=2.3
+ $Y2=0
r304 32 34 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.3 $Y=0.085
+ $X2=2.3 $Y2=0.495
r305 28 143 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.195 $Y2=0
r306 28 30 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r307 9 62 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=16.625
+ $Y=0.235 $X2=16.76 $Y2=0.38
r308 8 58 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=14.505
+ $Y=0.235 $X2=14.72 $Y2=0.495
r309 7 54 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=12.485
+ $Y=0.235 $X2=12.65 $Y2=0.38
r310 6 50 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=10.365
+ $Y=0.235 $X2=10.58 $Y2=0.495
r311 5 46 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=8.345
+ $Y=0.235 $X2=8.51 $Y2=0.38
r312 4 42 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=0.235 $X2=6.44 $Y2=0.495
r313 3 38 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.235 $X2=4.37 $Y2=0.38
r314 2 34 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.3 $Y2=0.495
r315 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

