* File: sky130_fd_sc_hdll__nand4_1.pex.spice
* Created: Wed Sep  2 08:38:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%D 1 3 4 6 7 12
r25 12 13 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r26 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r28 4 13 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r29 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r30 1 12 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r31 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%C 1 3 4 6 7 8 9 15 21
r36 21 23 1.11752 $w=3.28e-07 $l=3.2e-08 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.727 $Y2=1.16
r37 16 23 2.04284 $w=2.65e-07 $l=1.65e-07 $layer=LI1_cond $X=0.727 $Y=0.995
+ $X2=0.727 $Y2=1.16
r38 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r39 9 15 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.745 $Y=1.16
+ $X2=0.94 $Y2=1.16
r40 9 23 0.628605 $w=3.28e-07 $l=1.8e-08 $layer=LI1_cond $X=0.745 $Y=1.16
+ $X2=0.727 $Y2=1.16
r41 8 16 6.30582 $w=2.63e-07 $l=1.45e-07 $layer=LI1_cond $X=0.727 $Y=0.85
+ $X2=0.727 $Y2=0.995
r42 7 8 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.727 $Y=0.51
+ $X2=0.727 $Y2=0.85
r43 4 14 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.965 $Y2=1.16
r44 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.56
r45 1 14 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.16
r46 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%B 1 3 4 6 8 12 15
r42 15 22 13.079 $w=3.83e-07 $l=3.15e-07 $layer=LI1_cond $X=1.222 $Y=0.51
+ $X2=1.222 $Y2=0.825
r43 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.47
+ $Y=1.16 $X2=1.47 $Y2=1.16
r44 9 12 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.33 $Y=1.16 $X2=1.47
+ $Y2=1.16
r45 8 9 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.33 $Y=0.995 $X2=1.33
+ $Y2=1.16
r46 8 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.33 $Y=0.995
+ $X2=1.33 $Y2=0.825
r47 4 13 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.495 $Y2=1.16
r48 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r49 1 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.495 $Y2=1.16
r50 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%A 1 3 4 6 7 8 12 15
r28 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r29 12 14 39.279 $w=3.62e-07 $l=2.95e-07 $layer=POLY_cond $X=1.965 $Y=1.202
+ $X2=2.26 $Y2=1.202
r30 11 12 3.32873 $w=3.62e-07 $l=2.5e-08 $layer=POLY_cond $X=1.94 $Y=1.202
+ $X2=1.965 $Y2=1.202
r31 7 8 8.74552 $w=4.63e-07 $l=3.4e-07 $layer=LI1_cond $X=2.407 $Y=1.19
+ $X2=2.407 $Y2=1.53
r32 7 15 0.771663 $w=4.63e-07 $l=3e-08 $layer=LI1_cond $X=2.407 $Y=1.19
+ $X2=2.407 $Y2=1.16
r33 4 12 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.202
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
r35 1 11 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.94 $Y=0.995
+ $X2=1.94 $Y2=1.202
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.94 $Y=0.995 $X2=1.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%VPWR 1 2 3 10 12 16 20 24 27 28 29 36 37
+ 43
r40 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r42 34 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 34 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 31 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72 $X2=1.2
+ $Y2=2.72
r46 31 33 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 29 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 29 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 27 33 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 27 28 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.255 $Y2=2.72
r51 26 36 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.53 $Y2=2.72
r52 26 28 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.255 $Y2=2.72
r53 22 28 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2.72
r54 22 24 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2
r55 18 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r56 18 20 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r57 17 40 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r58 16 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72 $X2=1.2
+ $Y2=2.72
r59 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r60 12 15 30.1408 $w=2.58e-07 $l=6.8e-07 $layer=LI1_cond $X=0.215 $Y=1.66
+ $X2=0.215 $Y2=2.34
r61 10 40 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r62 10 15 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2.34
r63 3 24 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=1.485 $X2=2.2 $Y2=2
r64 2 20 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r65 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r66 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%Y 1 2 3 10 12 14 18 21 25 26 29
c46 21 0 1.19981e-19 $X=1.86 $Y=1.495
r47 26 33 13.4997 $w=7.43e-07 $l=3.15e-07 $layer=LI1_cond $X=2.042 $Y=0.51
+ $X2=2.042 $Y2=0.825
r48 26 29 2.08712 $w=7.43e-07 $l=1.3e-07 $layer=LI1_cond $X=2.042 $Y=0.51
+ $X2=2.042 $Y2=0.38
r49 21 25 3.70735 $w=2.5e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.86 $Y=1.495
+ $X2=1.74 $Y2=1.58
r50 21 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.86 $Y=1.495
+ $X2=1.86 $Y2=0.825
r51 16 25 3.70735 $w=2.5e-07 $l=1.03078e-07 $layer=LI1_cond $X=1.7 $Y=1.665
+ $X2=1.74 $Y2=1.58
r52 16 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.7 $Y=1.665
+ $X2=1.7 $Y2=2.34
r53 15 23 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r54 14 25 2.76166 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=1.74 $Y2=1.58
r55 14 15 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.535 $Y=1.58
+ $X2=0.895 $Y2=1.58
r56 10 23 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.58
r57 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r58 3 25 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.7 $Y2=1.66
r59 3 18 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.7 $Y2=2.34
r60 2 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r61 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r62 1 29 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.015
+ $Y=0.235 $X2=2.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_1%VGND 1 4 6 8 15 16
r26 15 16 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r27 13 16 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r28 12 15 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r29 12 13 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r30 10 19 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r31 10 12 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r32 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r33 8 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r34 4 19 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r35 4 6 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r36 1 6 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

