* File: sky130_fd_sc_hdll__or3_1.spice
* Created: Thu Aug 27 19:24:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3_1.pex.spice"
.subckt sky130_fd_sc_hdll__or3_1  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_C_M1001_g N_A_29_53#_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1007 N_A_29_53#_M1007_d N_B_M1007_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_29_53#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.0777 PD=0.816449 PS=0.79 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_29_53#_M1004_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.31525 AS=0.143516 PD=2.27 PS=1.26355 NRD=36.912 NRS=11.988 M=1 R=4.33333
+ SA=75001.2 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1002 A_119_297# N_C_M1002_g N_A_29_53#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0504 AS=0.1134 PD=0.66 PS=1.38 NRD=30.4759 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1006 A_203_297# N_B_M1006_g A_119_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0714
+ AS=0.0504 PD=0.76 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333 SA=90000.6
+ SB=90001.5 A=0.0756 P=1.2 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g A_203_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0714 PD=0.804507 PS=0.76 NRD=76.83 NRS=53.9386 M=1 R=2.33333
+ SA=90001.1 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1000 N_X_M1000_d N_A_29_53#_M1000_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.495 AS=0.218803 PD=2.99 PS=1.91549 NRD=41.3503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.8 SB=90000.4 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_12 A A PROBETYPE=1
c_52 VPB 0 1.10794e-19 $X=0.14 $Y=2.635
*
.include "sky130_fd_sc_hdll__or3_1.pxi.spice"
*
.ends
*
*
