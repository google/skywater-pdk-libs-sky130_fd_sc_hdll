* File: sky130_fd_sc_hdll__or3b_2.pxi.spice
* Created: Wed Sep  2 08:48:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3B_2%C_N N_C_N_c_77_n N_C_N_c_78_n N_C_N_M1006_g
+ N_C_N_M1009_g C_N C_N N_C_N_c_76_n PM_SKY130_FD_SC_HDLL__OR3B_2%C_N
x_PM_SKY130_FD_SC_HDLL__OR3B_2%A_186_21# N_A_186_21#_M1005_d N_A_186_21#_M1003_d
+ N_A_186_21#_M1008_d N_A_186_21#_c_106_n N_A_186_21#_M1001_g
+ N_A_186_21#_c_118_n N_A_186_21#_M1007_g N_A_186_21#_c_107_n
+ N_A_186_21#_c_108_n N_A_186_21#_M1010_g N_A_186_21#_c_109_n
+ N_A_186_21#_M1011_g N_A_186_21#_c_110_n N_A_186_21#_c_111_n
+ N_A_186_21#_c_112_n N_A_186_21#_c_172_p N_A_186_21#_c_198_p
+ N_A_186_21#_c_113_n N_A_186_21#_c_114_n N_A_186_21#_c_115_n
+ N_A_186_21#_c_116_n N_A_186_21#_c_117_n N_A_186_21#_c_124_n
+ PM_SKY130_FD_SC_HDLL__OR3B_2%A_186_21#
x_PM_SKY130_FD_SC_HDLL__OR3B_2%A N_A_c_209_n N_A_M1000_g N_A_M1005_g A A
+ PM_SKY130_FD_SC_HDLL__OR3B_2%A
x_PM_SKY130_FD_SC_HDLL__OR3B_2%B N_B_c_245_n N_B_c_248_n N_B_M1004_g N_B_M1002_g
+ B B B PM_SKY130_FD_SC_HDLL__OR3B_2%B
x_PM_SKY130_FD_SC_HDLL__OR3B_2%A_27_47# N_A_27_47#_M1009_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_282_n N_A_27_47#_M1008_g N_A_27_47#_M1003_g N_A_27_47#_c_284_n
+ N_A_27_47#_c_285_n N_A_27_47#_c_286_n N_A_27_47#_c_302_n N_A_27_47#_c_287_n
+ N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n N_A_27_47#_c_322_n
+ N_A_27_47#_c_323_n N_A_27_47#_c_294_n N_A_27_47#_c_288_n
+ PM_SKY130_FD_SC_HDLL__OR3B_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__OR3B_2%VPWR N_VPWR_M1006_d N_VPWR_M1010_d N_VPWR_c_385_n
+ N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n VPWR N_VPWR_c_389_n
+ N_VPWR_c_390_n N_VPWR_c_384_n N_VPWR_c_392_n PM_SKY130_FD_SC_HDLL__OR3B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3B_2%X N_X_M1001_d N_X_M1007_s N_X_c_432_n N_X_c_444_n
+ X X PM_SKY130_FD_SC_HDLL__OR3B_2%X
x_PM_SKY130_FD_SC_HDLL__OR3B_2%VGND N_VGND_M1009_d N_VGND_M1011_s N_VGND_M1002_d
+ N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n N_VGND_c_472_n
+ N_VGND_c_473_n N_VGND_c_474_n VGND N_VGND_c_475_n N_VGND_c_476_n
+ N_VGND_c_477_n PM_SKY130_FD_SC_HDLL__OR3B_2%VGND
cc_1 VNB N_C_N_M1009_g 0.0359511f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB C_N 0.00882738f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_76_n 0.0413107f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_186_21#_c_106_n 0.0182627f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_186_21#_c_107_n 0.0243741f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_A_186_21#_c_108_n 0.0138012f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_7 VNB N_A_186_21#_c_109_n 0.0191863f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_8 VNB N_A_186_21#_c_110_n 0.0133151f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.53
cc_9 VNB N_A_186_21#_c_111_n 6.89322e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_186_21#_c_112_n 0.0115527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_186_21#_c_113_n 0.00618952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_186_21#_c_114_n 0.0148426f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_186_21#_c_115_n 0.0228353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_186_21#_c_116_n 0.00295969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_186_21#_c_117_n 0.00991116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_c_209_n 0.0228992f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_17 VNB N_A_M1005_g 0.0276939f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_18 VNB A 0.00622854f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_19 VNB N_B_c_245_n 0.0120398f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_20 VNB N_B_M1002_g 0.032254f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_21 VNB N_A_27_47#_c_282_n 0.0239752f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_22 VNB N_A_27_47#_M1003_g 0.031502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_284_n 0.0183883f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_24 VNB N_A_27_47#_c_285_n 0.0048216f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_25 VNB N_A_27_47#_c_286_n 0.00960394f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_26 VNB N_A_27_47#_c_287_n 0.00683215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_288_n 0.00340078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_384_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_432_n 8.40947e-19 $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_30 VNB N_VGND_c_468_n 0.00467885f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_31 VNB N_VGND_c_469_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_32 VNB N_VGND_c_470_n 0.00363363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_471_n 0.0282822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_472_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_473_n 0.0188435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_474_n 0.0053059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_475_n 0.017386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_476_n 0.207769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_477_n 0.022544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_C_N_c_77_n 0.0211251f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.625
cc_41 VPB N_C_N_c_78_n 0.0324447f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.725
cc_42 VPB C_N 0.0160532f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_43 VPB N_C_N_c_76_n 0.0101485f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_44 VPB N_A_186_21#_c_118_n 0.0187325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_186_21#_c_107_n 0.0109069f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_46 VPB N_A_186_21#_c_108_n 0.0276002f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_47 VPB N_A_186_21#_c_110_n 0.0064913f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.53
cc_48 VPB N_A_186_21#_c_111_n 3.57415e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_186_21#_c_115_n 0.009285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_186_21#_c_124_n 0.0206732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_c_209_n 0.0263137f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_52 VPB A 0.00365798f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_53 VPB N_B_c_245_n 0.0066082f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_54 VPB N_B_c_248_n 0.0552099f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.625
cc_55 VPB N_B_M1004_g 0.0111506f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.01
cc_56 VPB B 0.0378463f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_57 VPB N_A_27_47#_c_282_n 0.0298363f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_58 VPB N_A_27_47#_c_287_n 0.00580119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_291_n 0.00547057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_47#_c_292_n 0.00143286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_293_n 0.0187914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_294_n 9.09856e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_288_n 4.20723e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_385_n 0.00995243f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_386_n 0.00794364f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_387_n 0.0179768f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_67 VPB N_VPWR_c_388_n 0.0051631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_389_n 0.0186913f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_390_n 0.0446991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_384_n 0.0643326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_392_n 0.00571014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_432_n 0.00175689f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_73 N_C_N_M1009_g N_A_186_21#_c_106_n 0.0181019f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_74 N_C_N_c_77_n N_A_186_21#_c_118_n 0.00844727f $X=0.495 $Y=1.625 $X2=0 $Y2=0
cc_75 N_C_N_c_78_n N_A_186_21#_c_118_n 0.015879f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_76 N_C_N_c_76_n N_A_186_21#_c_110_n 0.0181019f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_N_M1009_g N_A_27_47#_c_284_n 0.00429752f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_78 N_C_N_M1009_g N_A_27_47#_c_285_n 0.0180861f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_79 C_N N_A_27_47#_c_285_n 0.00618246f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_80 N_C_N_c_76_n N_A_27_47#_c_285_n 0.00301897f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_81 C_N N_A_27_47#_c_286_n 0.0227094f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_82 N_C_N_c_76_n N_A_27_47#_c_286_n 0.00599978f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_N_c_78_n N_A_27_47#_c_302_n 0.0183148f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_84 C_N N_A_27_47#_c_302_n 0.00421277f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_85 N_C_N_c_78_n N_A_27_47#_c_287_n 0.00209021f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_86 N_C_N_M1009_g N_A_27_47#_c_287_n 0.0117652f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_87 C_N N_A_27_47#_c_287_n 0.0350078f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_88 N_C_N_c_78_n N_A_27_47#_c_293_n 0.00472318f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_89 C_N N_A_27_47#_c_293_n 0.0226231f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_90 N_C_N_c_76_n N_A_27_47#_c_293_n 8.96314e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_91 N_C_N_c_78_n N_VPWR_c_385_n 0.00396865f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_92 N_C_N_c_78_n N_VPWR_c_389_n 0.00453698f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_93 N_C_N_c_78_n N_VPWR_c_384_n 0.00602858f $X=0.495 $Y=1.725 $X2=0 $Y2=0
cc_94 N_C_N_M1009_g N_X_c_432_n 8.22714e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_95 N_C_N_M1009_g N_VGND_c_468_n 0.00278284f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_96 N_C_N_M1009_g N_VGND_c_476_n 0.00717203f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_97 N_C_N_M1009_g N_VGND_c_477_n 0.00439206f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_98 N_A_186_21#_c_108_n N_A_c_209_n 0.042659f $X=1.61 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_186_21#_c_111_n N_A_c_209_n 7.16423e-19 $X=1.57 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_100 N_A_186_21#_c_112_n N_A_c_209_n 0.00462931f $X=2.365 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_186_21#_c_109_n N_A_M1005_g 0.0191177f $X=1.68 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_186_21#_c_111_n N_A_M1005_g 4.28033e-19 $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_186_21#_c_112_n N_A_M1005_g 0.0125796f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_104 N_A_186_21#_c_116_n N_A_M1005_g 0.0016391f $X=2.45 $Y=0.78 $X2=0 $Y2=0
cc_105 N_A_186_21#_c_108_n A 0.0075852f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_186_21#_c_111_n A 0.0130223f $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_186_21#_c_112_n A 0.0318837f $X=2.365 $Y=0.82 $X2=0 $Y2=0
cc_108 N_A_186_21#_c_116_n A 0.0155105f $X=2.45 $Y=0.78 $X2=0 $Y2=0
cc_109 N_A_186_21#_c_113_n N_B_c_245_n 0.00179638f $X=3.24 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_186_21#_c_113_n N_B_M1002_g 0.0161971f $X=3.24 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_186_21#_c_116_n N_B_M1002_g 0.00253148f $X=2.45 $Y=0.78 $X2=0 $Y2=0
cc_112 N_A_186_21#_c_124_n B 0.0214764f $X=3.46 $Y=1.71 $X2=0 $Y2=0
cc_113 N_A_186_21#_c_113_n N_A_27_47#_c_282_n 0.00389582f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_114 N_A_186_21#_c_115_n N_A_27_47#_c_282_n 0.0112574f $X=3.46 $Y=1.495 $X2=0
+ $Y2=0
cc_115 N_A_186_21#_c_117_n N_A_27_47#_c_282_n 2.9537e-19 $X=3.392 $Y=0.74 $X2=0
+ $Y2=0
cc_116 N_A_186_21#_c_124_n N_A_27_47#_c_282_n 0.00286266f $X=3.46 $Y=1.71 $X2=0
+ $Y2=0
cc_117 N_A_186_21#_c_113_n N_A_27_47#_M1003_g 0.0129827f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_118 N_A_186_21#_c_115_n N_A_27_47#_M1003_g 0.00569309f $X=3.46 $Y=1.495 $X2=0
+ $Y2=0
cc_119 N_A_186_21#_c_106_n N_A_27_47#_c_285_n 0.00132151f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_120 N_A_186_21#_c_106_n N_A_27_47#_c_287_n 0.00407679f $X=1.005 $Y=0.995
+ $X2=0 $Y2=0
cc_121 N_A_186_21#_c_118_n N_A_27_47#_c_287_n 0.00454336f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_122 N_A_186_21#_c_124_n N_A_27_47#_c_291_n 0.009394f $X=3.46 $Y=1.71 $X2=0
+ $Y2=0
cc_123 N_A_186_21#_c_115_n N_A_27_47#_c_292_n 0.0069946f $X=3.46 $Y=1.495 $X2=0
+ $Y2=0
cc_124 N_A_186_21#_c_124_n N_A_27_47#_c_292_n 0.0174776f $X=3.46 $Y=1.71 $X2=0
+ $Y2=0
cc_125 N_A_186_21#_c_118_n N_A_27_47#_c_322_n 0.00166683f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_186_21#_c_118_n N_A_27_47#_c_323_n 0.0158037f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_186_21#_c_107_n N_A_27_47#_c_323_n 0.00136921f $X=1.51 $Y=1.16 $X2=0
+ $Y2=0
cc_128 N_A_186_21#_c_108_n N_A_27_47#_c_323_n 0.0173115f $X=1.61 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_186_21#_c_111_n N_A_27_47#_c_323_n 0.0043879f $X=1.57 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_186_21#_c_108_n N_A_27_47#_c_294_n 0.00258004f $X=1.61 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_186_21#_c_113_n N_A_27_47#_c_288_n 0.0261561f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_132 N_A_186_21#_c_115_n N_A_27_47#_c_288_n 0.024341f $X=3.46 $Y=1.495 $X2=0
+ $Y2=0
cc_133 N_A_186_21#_c_118_n N_VPWR_c_385_n 0.0117335f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_186_21#_c_108_n N_VPWR_c_385_n 0.00203704f $X=1.61 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_186_21#_c_118_n N_VPWR_c_386_n 0.0020155f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_186_21#_c_108_n N_VPWR_c_386_n 0.0113201f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_186_21#_c_118_n N_VPWR_c_387_n 0.00459627f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_186_21#_c_108_n N_VPWR_c_387_n 0.00474014f $X=1.61 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_186_21#_c_118_n N_VPWR_c_384_n 0.00556431f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_186_21#_c_108_n N_VPWR_c_384_n 0.00571062f $X=1.61 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_186_21#_c_172_p N_X_M1001_d 0.00293374f $X=1.655 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_142 N_A_186_21#_c_106_n N_X_c_432_n 0.0122433f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_186_21#_c_118_n N_X_c_432_n 0.00262165f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_186_21#_c_107_n N_X_c_432_n 0.0120528f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_186_21#_c_108_n N_X_c_432_n 0.00351153f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_186_21#_c_109_n N_X_c_432_n 0.00353939f $X=1.68 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_186_21#_c_110_n N_X_c_432_n 0.0090241f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A_186_21#_c_111_n N_X_c_432_n 0.0222449f $X=1.57 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_186_21#_c_172_p N_X_c_432_n 0.0107392f $X=1.655 $Y=0.82 $X2=0 $Y2=0
cc_150 N_A_186_21#_c_118_n N_X_c_444_n 0.00598531f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_186_21#_c_107_n N_X_c_444_n 0.00801141f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_186_21#_c_108_n N_X_c_444_n 0.00413504f $X=1.61 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_186_21#_c_106_n X 0.00629929f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_186_21#_c_107_n X 0.00496114f $X=1.51 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_186_21#_c_109_n X 0.00411015f $X=1.68 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_186_21#_c_112_n N_VGND_M1011_s 0.00284211f $X=2.365 $Y=0.82 $X2=0
+ $Y2=0
cc_157 N_A_186_21#_c_113_n N_VGND_M1002_d 0.00190907f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_A_186_21#_c_106_n N_VGND_c_468_n 0.00514031f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_186_21#_c_109_n N_VGND_c_469_n 0.00523783f $X=1.68 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_186_21#_c_112_n N_VGND_c_469_n 0.0132189f $X=2.365 $Y=0.82 $X2=0
+ $Y2=0
cc_161 N_A_186_21#_c_113_n N_VGND_c_470_n 0.0163215f $X=3.24 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_186_21#_c_106_n N_VGND_c_471_n 0.00442618f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_186_21#_c_109_n N_VGND_c_471_n 0.00439161f $X=1.68 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_186_21#_c_112_n N_VGND_c_471_n 0.00248062f $X=2.365 $Y=0.82 $X2=0
+ $Y2=0
cc_165 N_A_186_21#_c_172_p N_VGND_c_471_n 0.00212913f $X=1.655 $Y=0.82 $X2=0
+ $Y2=0
cc_166 N_A_186_21#_c_112_n N_VGND_c_473_n 0.00464236f $X=2.365 $Y=0.82 $X2=0
+ $Y2=0
cc_167 N_A_186_21#_c_198_p N_VGND_c_473_n 0.00879995f $X=2.45 $Y=0.47 $X2=0
+ $Y2=0
cc_168 N_A_186_21#_c_113_n N_VGND_c_473_n 0.00283921f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_169 N_A_186_21#_c_113_n N_VGND_c_475_n 0.00232396f $X=3.24 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_186_21#_c_114_n N_VGND_c_475_n 0.0159441f $X=3.325 $Y=0.47 $X2=0
+ $Y2=0
cc_171 N_A_186_21#_c_106_n N_VGND_c_476_n 0.00797423f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A_186_21#_c_109_n N_VGND_c_476_n 0.00719016f $X=1.68 $Y=0.995 $X2=0
+ $Y2=0
cc_173 N_A_186_21#_c_112_n N_VGND_c_476_n 0.0135716f $X=2.365 $Y=0.82 $X2=0
+ $Y2=0
cc_174 N_A_186_21#_c_172_p N_VGND_c_476_n 0.00446193f $X=1.655 $Y=0.82 $X2=0
+ $Y2=0
cc_175 N_A_186_21#_c_198_p N_VGND_c_476_n 0.00627241f $X=2.45 $Y=0.47 $X2=0
+ $Y2=0
cc_176 N_A_186_21#_c_113_n N_VGND_c_476_n 0.0105277f $X=3.24 $Y=0.74 $X2=0 $Y2=0
cc_177 N_A_186_21#_c_114_n N_VGND_c_476_n 0.0113365f $X=3.325 $Y=0.47 $X2=0
+ $Y2=0
cc_178 N_A_c_209_n N_B_c_245_n 0.0146796f $X=2.15 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_179 A N_B_c_245_n 0.00349176f $X=2.3 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_180 N_A_c_209_n N_B_M1004_g 0.0248172f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_181 A N_B_M1004_g 0.00158693f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_182 N_A_M1005_g N_B_M1002_g 0.0267048f $X=2.235 $Y=0.475 $X2=0 $Y2=0
cc_183 A N_B_M1002_g 3.66953e-19 $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_184 N_A_c_209_n B 0.00131215f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_209_n N_A_27_47#_c_291_n 0.0128282f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_186 A N_A_27_47#_c_292_n 0.011742f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A_c_209_n N_A_27_47#_c_294_n 0.00255026f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_188 A N_A_27_47#_c_294_n 0.032872f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_189 A N_A_27_47#_c_288_n 0.0143501f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_190 A N_VPWR_M1010_d 0.00240272f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_191 N_A_c_209_n N_VPWR_c_390_n 0.00299159f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_c_209_n N_VPWR_c_384_n 0.0037574f $X=2.15 $Y=1.41 $X2=0 $Y2=0
cc_193 A N_X_c_444_n 0.00440295f $X=2.3 $Y=1.105 $X2=0 $Y2=0
cc_194 A A_448_297# 0.00245184f $X=2.3 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_195 N_A_M1005_g N_VGND_c_469_n 0.00593299f $X=2.235 $Y=0.475 $X2=0 $Y2=0
cc_196 N_A_M1005_g N_VGND_c_473_n 0.00413798f $X=2.235 $Y=0.475 $X2=0 $Y2=0
cc_197 N_A_M1005_g N_VGND_c_476_n 0.00610822f $X=2.235 $Y=0.475 $X2=0 $Y2=0
cc_198 N_B_c_245_n N_A_27_47#_c_282_n 0.00405288f $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_M1004_g N_A_27_47#_c_282_n 0.0283372f $X=2.64 $Y=1.695 $X2=0 $Y2=0
cc_200 N_B_M1002_g N_A_27_47#_c_282_n 0.0196008f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_201 B N_A_27_47#_c_282_n 0.00807787f $X=3.32 $Y=2.125 $X2=0 $Y2=0
cc_202 N_B_M1002_g N_A_27_47#_M1003_g 0.0219808f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_203 N_B_c_248_n N_A_27_47#_c_291_n 0.00144871f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_204 N_B_M1004_g N_A_27_47#_c_291_n 0.0172513f $X=2.64 $Y=1.695 $X2=0 $Y2=0
cc_205 B N_A_27_47#_c_291_n 0.0613864f $X=3.32 $Y=2.125 $X2=0 $Y2=0
cc_206 N_B_c_245_n N_A_27_47#_c_292_n 6.69515e-19 $X=2.64 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_M1004_g N_A_27_47#_c_292_n 0.00533878f $X=2.64 $Y=1.695 $X2=0 $Y2=0
cc_208 N_B_M1002_g N_A_27_47#_c_288_n 0.00397268f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_209 N_B_c_248_n N_VPWR_c_386_n 0.00228645f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_210 B N_VPWR_c_386_n 0.0130814f $X=3.32 $Y=2.125 $X2=0 $Y2=0
cc_211 N_B_c_248_n N_VPWR_c_390_n 0.00868974f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_212 B N_VPWR_c_390_n 0.0537216f $X=3.32 $Y=2.125 $X2=0 $Y2=0
cc_213 N_B_c_248_n N_VPWR_c_384_n 0.0122906f $X=2.64 $Y=2.035 $X2=0 $Y2=0
cc_214 B N_VPWR_c_384_n 0.0473029f $X=3.32 $Y=2.125 $X2=0 $Y2=0
cc_215 N_B_M1002_g N_VGND_c_470_n 0.00327287f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_216 N_B_M1002_g N_VGND_c_473_n 0.00402675f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_217 N_B_M1002_g N_VGND_c_476_n 0.00548116f $X=2.665 $Y=0.475 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_287_n N_VPWR_M1006_d 0.00431942f $X=0.73 $Y=1.81 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_27_47#_c_322_n N_VPWR_M1006_d 0.00255548f $X=0.73 $Y=1.925 $X2=-0.19
+ $Y2=-0.24
cc_220 N_A_27_47#_c_323_n N_VPWR_M1006_d 0.00324693f $X=1.81 $Y=1.912 $X2=-0.19
+ $Y2=-0.24
cc_221 N_A_27_47#_c_291_n N_VPWR_M1010_d 2.16905e-19 $X=2.85 $Y=1.87 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_323_n N_VPWR_M1010_d 0.00252001f $X=1.81 $Y=1.912 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_294_n N_VPWR_M1010_d 0.00894338f $X=1.98 $Y=1.912 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_322_n N_VPWR_c_385_n 0.0144404f $X=0.73 $Y=1.925 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_323_n N_VPWR_c_385_n 0.00655922f $X=1.81 $Y=1.912 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_291_n N_VPWR_c_386_n 0.00196088f $X=2.85 $Y=1.87 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_323_n N_VPWR_c_386_n 0.0185534f $X=1.81 $Y=1.912 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_323_n N_VPWR_c_387_n 0.0103188f $X=1.81 $Y=1.912 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_302_n N_VPWR_c_389_n 0.00337107f $X=0.645 $Y=1.925 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_293_n N_VPWR_c_389_n 0.00669761f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_302_n N_VPWR_c_384_n 0.00706969f $X=0.645 $Y=1.925 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_291_n N_VPWR_c_384_n 0.00727421f $X=2.85 $Y=1.87 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_293_n N_VPWR_c_384_n 0.00838075f $X=0.26 $Y=1.975 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_322_n N_VPWR_c_384_n 7.87123e-19 $X=0.73 $Y=1.925 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_323_n N_VPWR_c_384_n 0.0200852f $X=1.81 $Y=1.912 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_323_n N_X_M1007_s 0.00857304f $X=1.81 $Y=1.912 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_284_n N_X_c_432_n 0.00375501f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_285_n N_X_c_432_n 0.0138065f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_287_n N_X_c_432_n 0.0432945f $X=0.73 $Y=1.81 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_287_n N_X_c_444_n 0.0154212f $X=0.73 $Y=1.81 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_323_n N_X_c_444_n 0.027852f $X=1.81 $Y=1.912 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_284_n X 7.83518e-19 $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_291_n A_448_297# 0.00206656f $X=2.85 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_291_n A_546_297# 0.00236564f $X=2.85 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_245 N_A_27_47#_c_292_n A_546_297# 0.00327094f $X=2.935 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_246 N_A_27_47#_c_285_n N_VGND_M1009_d 0.00309755f $X=0.645 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_247 N_A_27_47#_c_285_n N_VGND_c_468_n 0.0143363f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_248 N_A_27_47#_M1003_g N_VGND_c_470_n 0.00947382f $X=3.115 $Y=0.475 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1003_g N_VGND_c_475_n 0.00322006f $X=3.115 $Y=0.475 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_M1009_s N_VGND_c_476_n 0.00302988f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1003_g N_VGND_c_476_n 0.0047132f $X=3.115 $Y=0.475 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_284_n N_VGND_c_476_n 0.00973659f $X=0.26 $Y=0.455 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_285_n N_VGND_c_476_n 0.00776442f $X=0.645 $Y=0.82 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_284_n N_VGND_c_477_n 0.01476f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_285_n N_VGND_c_477_n 0.0041864f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_256 N_VPWR_c_384_n N_X_M1007_s 0.0049337f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_257 X N_VGND_c_468_n 0.0225239f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_258 X N_VGND_c_469_n 0.0107586f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_259 X N_VGND_c_471_n 0.0230768f $X=1.17 $Y=0.425 $X2=0 $Y2=0
cc_260 N_X_M1001_d N_VGND_c_476_n 0.00832391f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_261 X N_VGND_c_476_n 0.0145315f $X=1.17 $Y=0.425 $X2=0 $Y2=0
