* File: sky130_fd_sc_hdll__clkinv_16.pxi.spice
* Created: Thu Aug 27 19:02:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_16%A N_A_c_174_n N_A_M1001_g N_A_c_175_n
+ N_A_M1002_g N_A_c_176_n N_A_M1003_g N_A_c_177_n N_A_M1004_g N_A_M1000_g
+ N_A_c_178_n N_A_M1006_g N_A_M1005_g N_A_c_179_n N_A_M1007_g N_A_M1008_g
+ N_A_c_180_n N_A_M1009_g N_A_M1010_g N_A_c_181_n N_A_M1012_g N_A_M1011_g
+ N_A_c_182_n N_A_M1015_g N_A_M1013_g N_A_c_183_n N_A_M1018_g N_A_M1014_g
+ N_A_c_184_n N_A_M1019_g N_A_c_160_n N_A_c_161_n N_A_M1016_g N_A_c_187_n
+ N_A_M1020_g N_A_M1017_g N_A_c_188_n N_A_M1021_g N_A_M1028_g N_A_c_189_n
+ N_A_M1022_g N_A_M1029_g N_A_c_190_n N_A_M1023_g N_A_M1031_g N_A_c_191_n
+ N_A_M1024_g N_A_M1033_g N_A_c_192_n N_A_M1025_g N_A_M1035_g N_A_c_193_n
+ N_A_M1026_g N_A_M1036_g N_A_c_194_n N_A_M1027_g N_A_M1038_g N_A_c_195_n
+ N_A_M1030_g N_A_c_196_n N_A_M1032_g N_A_c_197_n N_A_M1034_g N_A_c_198_n
+ N_A_M1037_g N_A_c_199_n N_A_M1039_g A N_A_c_286_p N_A_c_287_p N_A_c_293_p
+ N_A_c_348_p N_A_c_359_p N_A_c_172_n N_A_c_173_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_16%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_16%VPWR N_VPWR_M1001_d N_VPWR_M1002_d
+ N_VPWR_M1004_d N_VPWR_M1007_d N_VPWR_M1012_d N_VPWR_M1018_d N_VPWR_M1020_d
+ N_VPWR_M1022_d N_VPWR_M1024_d N_VPWR_M1026_d N_VPWR_M1030_d N_VPWR_M1034_d
+ N_VPWR_M1039_d N_VPWR_c_450_n N_VPWR_c_451_n N_VPWR_c_452_n N_VPWR_c_453_n
+ N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_457_n N_VPWR_c_458_n
+ N_VPWR_c_607_p N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_467_n
+ N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n
+ N_VPWR_c_473_n N_VPWR_c_474_n N_VPWR_c_475_n N_VPWR_c_476_n N_VPWR_c_477_n
+ N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n VPWR
+ N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_449_n N_VPWR_c_485_n N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_16%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_16%Y N_Y_M1000_d N_Y_M1008_d N_Y_M1011_d
+ N_Y_M1014_d N_Y_M1017_d N_Y_M1029_d N_Y_M1033_d N_Y_M1036_d N_Y_M1001_s
+ N_Y_M1003_s N_Y_M1006_s N_Y_M1009_s N_Y_M1015_s N_Y_M1019_s N_Y_M1021_s
+ N_Y_M1023_s N_Y_M1025_s N_Y_M1027_s N_Y_M1032_s N_Y_M1037_s N_Y_c_630_n
+ N_Y_c_773_n N_Y_c_631_n N_Y_c_632_n N_Y_c_622_n N_Y_c_634_n N_Y_c_623_n
+ N_Y_c_636_n N_Y_c_624_n N_Y_c_638_n Y N_Y_c_625_n N_Y_c_626_n N_Y_c_641_n
+ N_Y_c_627_n N_Y_c_643_n N_Y_c_628_n N_Y_c_645_n N_Y_c_629_n N_Y_c_647_n
+ N_Y_c_648_n N_Y_c_649_n N_Y_c_650_n N_Y_c_799_n N_Y_c_801_n N_Y_c_651_n
+ N_Y_c_805_n N_Y_c_807_n N_Y_c_809_n N_Y_c_652_n N_Y_c_653_n N_Y_c_654_n Y
+ PM_SKY130_FD_SC_HDLL__CLKINV_16%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_16%VGND N_VGND_M1000_s N_VGND_M1005_s
+ N_VGND_M1010_s N_VGND_M1013_s N_VGND_M1016_s N_VGND_M1028_s N_VGND_M1031_s
+ N_VGND_M1035_s N_VGND_M1038_s N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n
+ N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n N_VGND_c_855_n N_VGND_c_856_n
+ N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n N_VGND_c_860_n N_VGND_c_861_n
+ N_VGND_c_862_n N_VGND_c_863_n VGND N_VGND_c_864_n N_VGND_c_865_n
+ N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n N_VGND_c_869_n N_VGND_c_870_n
+ N_VGND_c_871_n N_VGND_c_872_n PM_SKY130_FD_SC_HDLL__CLKINV_16%VGND
cc_1 VNB N_A_M1000_g 0.0392593f $X=-0.19 $Y=-0.24 $X2=2.405 $Y2=0.445
cc_2 VNB N_A_M1005_g 0.0293323f $X=-0.19 $Y=-0.24 $X2=2.885 $Y2=0.445
cc_3 VNB N_A_M1008_g 0.029332f $X=-0.19 $Y=-0.24 $X2=3.365 $Y2=0.445
cc_4 VNB N_A_M1010_g 0.0293323f $X=-0.19 $Y=-0.24 $X2=3.845 $Y2=0.445
cc_5 VNB N_A_M1011_g 0.029332f $X=-0.19 $Y=-0.24 $X2=4.325 $Y2=0.445
cc_6 VNB N_A_M1013_g 0.029939f $X=-0.19 $Y=-0.24 $X2=4.805 $Y2=0.445
cc_7 VNB N_A_M1014_g 0.0322164f $X=-0.19 $Y=-0.24 $X2=5.32 $Y2=0.445
cc_8 VNB N_A_c_160_n 0.0231934f $X=-0.19 $Y=-0.24 $X2=5.88 $Y2=1.17
cc_9 VNB N_A_c_161_n 0.259692f $X=-0.19 $Y=-0.24 $X2=5.445 $Y2=1.17
cc_10 VNB N_A_M1016_g 0.0316207f $X=-0.19 $Y=-0.24 $X2=5.955 $Y2=0.445
cc_11 VNB N_A_M1017_g 0.0293397f $X=-0.19 $Y=-0.24 $X2=6.435 $Y2=0.445
cc_12 VNB N_A_M1028_g 0.0293325f $X=-0.19 $Y=-0.24 $X2=6.915 $Y2=0.445
cc_13 VNB N_A_M1029_g 0.0293327f $X=-0.19 $Y=-0.24 $X2=7.395 $Y2=0.445
cc_14 VNB N_A_M1031_g 0.0293325f $X=-0.19 $Y=-0.24 $X2=7.875 $Y2=0.445
cc_15 VNB N_A_M1033_g 0.0293327f $X=-0.19 $Y=-0.24 $X2=8.355 $Y2=0.445
cc_16 VNB N_A_M1035_g 0.0293325f $X=-0.19 $Y=-0.24 $X2=8.835 $Y2=0.445
cc_17 VNB N_A_M1036_g 0.0293327f $X=-0.19 $Y=-0.24 $X2=9.315 $Y2=0.445
cc_18 VNB N_A_M1038_g 0.0385631f $X=-0.19 $Y=-0.24 $X2=9.795 $Y2=0.445
cc_19 VNB A 0.0843643f $X=-0.19 $Y=-0.24 $X2=1.985 $Y2=1.105
cc_20 VNB N_A_c_172_n 0.300949f $X=-0.19 $Y=-0.24 $X2=11.61 $Y2=1.16
cc_21 VNB N_A_c_173_n 0.0853868f $X=-0.19 $Y=-0.24 $X2=11.61 $Y2=1.16
cc_22 VNB N_VPWR_c_449_n 0.516438f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.2
cc_23 VNB N_Y_c_622_n 0.00728867f $X=-0.19 $Y=-0.24 $X2=6.435 $Y2=0.445
cc_24 VNB N_Y_c_623_n 0.00782183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_624_n 0.00769318f $X=-0.19 $Y=-0.24 $X2=7.42 $Y2=1.41
cc_26 VNB N_Y_c_625_n 0.00866819f $X=-0.19 $Y=-0.24 $X2=8.355 $Y2=0.445
cc_27 VNB N_Y_c_626_n 0.00777887f $X=-0.19 $Y=-0.24 $X2=8.835 $Y2=0.99
cc_28 VNB N_Y_c_627_n 0.00777887f $X=-0.19 $Y=-0.24 $X2=9.315 $Y2=0.445
cc_29 VNB N_Y_c_628_n 0.00777887f $X=-0.19 $Y=-0.24 $X2=9.795 $Y2=0.445
cc_30 VNB N_Y_c_629_n 0.00748428f $X=-0.19 $Y=-0.24 $X2=10.78 $Y2=1.41
cc_31 VNB N_VGND_c_844_n 0.0190025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_845_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=3.845 $Y2=0.99
cc_33 VNB N_VGND_c_846_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=3.87 $Y2=1.41
cc_34 VNB N_VGND_c_847_n 0.00526426f $X=-0.19 $Y=-0.24 $X2=4.325 $Y2=0.445
cc_35 VNB N_VGND_c_848_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=4.35 $Y2=1.985
cc_36 VNB N_VGND_c_849_n 0.0197796f $X=-0.19 $Y=-0.24 $X2=4.805 $Y2=0.99
cc_37 VNB N_VGND_c_850_n 0.00503993f $X=-0.19 $Y=-0.24 $X2=4.83 $Y2=1.41
cc_38 VNB N_VGND_c_851_n 0.0211037f $X=-0.19 $Y=-0.24 $X2=4.83 $Y2=1.985
cc_39 VNB N_VGND_c_852_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_853_n 0.0197796f $X=-0.19 $Y=-0.24 $X2=5.345 $Y2=1.985
cc_41 VNB N_VGND_c_854_n 0.00526389f $X=-0.19 $Y=-0.24 $X2=5.955 $Y2=0.99
cc_42 VNB N_VGND_c_855_n 0.0189592f $X=-0.19 $Y=-0.24 $X2=5.98 $Y2=1.41
cc_43 VNB N_VGND_c_856_n 0.0200035f $X=-0.19 $Y=-0.24 $X2=6.435 $Y2=0.99
cc_44 VNB N_VGND_c_857_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=6.435 $Y2=0.445
cc_45 VNB N_VGND_c_858_n 0.0197348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_859_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=6.46 $Y2=1.41
cc_47 VNB N_VGND_c_860_n 0.0206647f $X=-0.19 $Y=-0.24 $X2=6.46 $Y2=1.985
cc_48 VNB N_VGND_c_861_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=6.915 $Y2=0.99
cc_49 VNB N_VGND_c_862_n 0.0197796f $X=-0.19 $Y=-0.24 $X2=6.915 $Y2=0.445
cc_50 VNB N_VGND_c_863_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_864_n 0.0675375f $X=-0.19 $Y=-0.24 $X2=6.94 $Y2=1.985
cc_52 VNB N_VGND_c_865_n 0.0241855f $X=-0.19 $Y=-0.24 $X2=8.355 $Y2=0.99
cc_53 VNB N_VGND_c_866_n 0.0729473f $X=-0.19 $Y=-0.24 $X2=8.86 $Y2=1.985
cc_54 VNB N_VGND_c_867_n 0.730329f $X=-0.19 $Y=-0.24 $X2=8.86 $Y2=1.985
cc_55 VNB N_VGND_c_868_n 0.00516809f $X=-0.19 $Y=-0.24 $X2=9.315 $Y2=0.445
cc_56 VNB N_VGND_c_869_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=9.34 $Y2=1.985
cc_57 VNB N_VGND_c_870_n 0.00430243f $X=-0.19 $Y=-0.24 $X2=9.795 $Y2=0.445
cc_58 VNB N_VGND_c_871_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=9.82 $Y2=1.41
cc_59 VNB N_VGND_c_872_n 0.00507191f $X=-0.19 $Y=-0.24 $X2=10.3 $Y2=1.41
cc_60 VPB N_A_c_174_n 0.0211592f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_61 VPB N_A_c_175_n 0.0161387f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.41
cc_62 VPB N_A_c_176_n 0.0161387f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.41
cc_63 VPB N_A_c_177_n 0.0160458f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.41
cc_64 VPB N_A_c_178_n 0.0160328f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.41
cc_65 VPB N_A_c_179_n 0.0156214f $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.41
cc_66 VPB N_A_c_180_n 0.0156214f $X=-0.19 $Y=1.305 $X2=3.39 $Y2=1.41
cc_67 VPB N_A_c_181_n 0.0156214f $X=-0.19 $Y=1.305 $X2=3.87 $Y2=1.41
cc_68 VPB N_A_c_182_n 0.0156214f $X=-0.19 $Y=1.305 $X2=4.35 $Y2=1.41
cc_69 VPB N_A_c_183_n 0.0158872f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.41
cc_70 VPB N_A_c_184_n 0.0169197f $X=-0.19 $Y=1.305 $X2=5.345 $Y2=1.41
cc_71 VPB N_A_c_160_n 0.0140905f $X=-0.19 $Y=1.305 $X2=5.88 $Y2=1.17
cc_72 VPB N_A_c_161_n 0.142987f $X=-0.19 $Y=1.305 $X2=5.445 $Y2=1.17
cc_73 VPB N_A_c_187_n 0.016654f $X=-0.19 $Y=1.305 $X2=5.98 $Y2=1.41
cc_74 VPB N_A_c_188_n 0.0156214f $X=-0.19 $Y=1.305 $X2=6.46 $Y2=1.41
cc_75 VPB N_A_c_189_n 0.0156214f $X=-0.19 $Y=1.305 $X2=6.94 $Y2=1.41
cc_76 VPB N_A_c_190_n 0.0156214f $X=-0.19 $Y=1.305 $X2=7.42 $Y2=1.41
cc_77 VPB N_A_c_191_n 0.0156214f $X=-0.19 $Y=1.305 $X2=7.9 $Y2=1.41
cc_78 VPB N_A_c_192_n 0.0156214f $X=-0.19 $Y=1.305 $X2=8.38 $Y2=1.41
cc_79 VPB N_A_c_193_n 0.0156214f $X=-0.19 $Y=1.305 $X2=8.86 $Y2=1.41
cc_80 VPB N_A_c_194_n 0.0156214f $X=-0.19 $Y=1.305 $X2=9.34 $Y2=1.41
cc_81 VPB N_A_c_195_n 0.0160324f $X=-0.19 $Y=1.305 $X2=9.82 $Y2=1.41
cc_82 VPB N_A_c_196_n 0.0160455f $X=-0.19 $Y=1.305 $X2=10.3 $Y2=1.41
cc_83 VPB N_A_c_197_n 0.0161387f $X=-0.19 $Y=1.305 $X2=10.78 $Y2=1.41
cc_84 VPB N_A_c_198_n 0.0161387f $X=-0.19 $Y=1.305 $X2=11.26 $Y2=1.41
cc_85 VPB N_A_c_199_n 0.0211592f $X=-0.19 $Y=1.305 $X2=11.74 $Y2=1.41
cc_86 VPB N_A_c_172_n 0.16875f $X=-0.19 $Y=1.305 $X2=11.61 $Y2=1.16
cc_87 VPB N_VPWR_c_450_n 0.0117381f $X=-0.19 $Y=1.305 $X2=3.87 $Y2=1.985
cc_88 VPB N_VPWR_c_451_n 0.00526426f $X=-0.19 $Y=1.305 $X2=4.325 $Y2=0.445
cc_89 VPB N_VPWR_c_452_n 0.0196725f $X=-0.19 $Y=1.305 $X2=4.35 $Y2=1.985
cc_90 VPB N_VPWR_c_453_n 0.00522213f $X=-0.19 $Y=1.305 $X2=4.805 $Y2=0.445
cc_91 VPB N_VPWR_c_454_n 0.0200595f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.41
cc_92 VPB N_VPWR_c_455_n 0.00519417f $X=-0.19 $Y=1.305 $X2=5.32 $Y2=0.445
cc_93 VPB N_VPWR_c_456_n 0.00522213f $X=-0.19 $Y=1.305 $X2=5.345 $Y2=1.985
cc_94 VPB N_VPWR_c_457_n 0.00519417f $X=-0.19 $Y=1.305 $X2=5.955 $Y2=0.99
cc_95 VPB N_VPWR_c_458_n 0.00519546f $X=-0.19 $Y=1.305 $X2=5.98 $Y2=1.41
cc_96 VPB N_VPWR_c_459_n 0.00522213f $X=-0.19 $Y=1.305 $X2=6.46 $Y2=1.985
cc_97 VPB N_VPWR_c_460_n 0.0201052f $X=-0.19 $Y=1.305 $X2=6.915 $Y2=0.99
cc_98 VPB N_VPWR_c_461_n 0.00519417f $X=-0.19 $Y=1.305 $X2=6.94 $Y2=1.41
cc_99 VPB N_VPWR_c_462_n 0.0201052f $X=-0.19 $Y=1.305 $X2=6.94 $Y2=1.985
cc_100 VPB N_VPWR_c_463_n 0.00519417f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_464_n 0.00519417f $X=-0.19 $Y=1.305 $X2=7.875 $Y2=0.99
cc_102 VPB N_VPWR_c_465_n 0.00519417f $X=-0.19 $Y=1.305 $X2=7.9 $Y2=1.41
cc_103 VPB N_VPWR_c_466_n 0.00519417f $X=-0.19 $Y=1.305 $X2=8.355 $Y2=0.445
cc_104 VPB N_VPWR_c_467_n 0.0287427f $X=-0.19 $Y=1.305 $X2=8.38 $Y2=1.985
cc_105 VPB N_VPWR_c_468_n 0.0201139f $X=-0.19 $Y=1.305 $X2=8.835 $Y2=0.445
cc_106 VPB N_VPWR_c_469_n 0.00497514f $X=-0.19 $Y=1.305 $X2=8.835 $Y2=0.445
cc_107 VPB N_VPWR_c_470_n 0.0200595f $X=-0.19 $Y=1.305 $X2=8.86 $Y2=1.41
cc_108 VPB N_VPWR_c_471_n 0.00487897f $X=-0.19 $Y=1.305 $X2=8.86 $Y2=1.985
cc_109 VPB N_VPWR_c_472_n 0.020833f $X=-0.19 $Y=1.305 $X2=9.315 $Y2=0.99
cc_110 VPB N_VPWR_c_473_n 0.00487897f $X=-0.19 $Y=1.305 $X2=9.315 $Y2=0.445
cc_111 VPB N_VPWR_c_474_n 0.0201052f $X=-0.19 $Y=1.305 $X2=9.34 $Y2=1.41
cc_112 VPB N_VPWR_c_475_n 0.00487897f $X=-0.19 $Y=1.305 $X2=9.34 $Y2=1.985
cc_113 VPB N_VPWR_c_476_n 0.0201052f $X=-0.19 $Y=1.305 $X2=9.795 $Y2=0.99
cc_114 VPB N_VPWR_c_477_n 0.00487897f $X=-0.19 $Y=1.305 $X2=9.795 $Y2=0.445
cc_115 VPB N_VPWR_c_478_n 0.0201965f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_479_n 0.00487897f $X=-0.19 $Y=1.305 $X2=9.82 $Y2=1.41
cc_117 VPB N_VPWR_c_480_n 0.0199004f $X=-0.19 $Y=1.305 $X2=9.82 $Y2=1.985
cc_118 VPB N_VPWR_c_481_n 0.00497514f $X=-0.19 $Y=1.305 $X2=10.3 $Y2=1.41
cc_119 VPB N_VPWR_c_482_n 0.0242138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_VPWR_c_483_n 0.0120081f $X=-0.19 $Y=1.305 $X2=1.47 $Y2=1.2
cc_121 VPB N_VPWR_c_449_n 0.0549665f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.2
cc_122 VPB N_VPWR_c_485_n 0.00497514f $X=-0.19 $Y=1.305 $X2=2.885 $Y2=1.2
cc_123 VPB N_VPWR_c_486_n 0.00487897f $X=-0.19 $Y=1.305 $X2=3.39 $Y2=1.2
cc_124 VPB N_VPWR_c_487_n 0.00497514f $X=-0.19 $Y=1.305 $X2=4.325 $Y2=1.2
cc_125 VPB N_VPWR_c_488_n 0.00487897f $X=-0.19 $Y=1.305 $X2=4.83 $Y2=1.2
cc_126 VPB N_VPWR_c_489_n 0.00487897f $X=-0.19 $Y=1.305 $X2=5.955 $Y2=1.2
cc_127 VPB N_Y_c_630_n 0.00196853f $X=-0.19 $Y=1.305 $X2=5.345 $Y2=1.985
cc_128 VPB N_Y_c_631_n 0.00204866f $X=-0.19 $Y=1.305 $X2=5.955 $Y2=0.445
cc_129 VPB N_Y_c_632_n 0.00169738f $X=-0.19 $Y=1.305 $X2=5.98 $Y2=1.985
cc_130 VPB N_Y_c_622_n 0.00112285f $X=-0.19 $Y=1.305 $X2=6.435 $Y2=0.445
cc_131 VPB N_Y_c_634_n 0.00103371f $X=-0.19 $Y=1.305 $X2=6.46 $Y2=1.985
cc_132 VPB N_Y_c_623_n 0.0011378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_Y_c_636_n 0.00103371f $X=-0.19 $Y=1.305 $X2=7.395 $Y2=0.99
cc_134 VPB N_Y_c_624_n 0.00113009f $X=-0.19 $Y=1.305 $X2=7.42 $Y2=1.41
cc_135 VPB N_Y_c_638_n 0.00116948f $X=-0.19 $Y=1.305 $X2=7.875 $Y2=0.445
cc_136 VPB N_Y_c_625_n 0.0011903f $X=-0.19 $Y=1.305 $X2=8.355 $Y2=0.445
cc_137 VPB N_Y_c_626_n 0.00113521f $X=-0.19 $Y=1.305 $X2=8.835 $Y2=0.99
cc_138 VPB N_Y_c_641_n 0.00104879f $X=-0.19 $Y=1.305 $X2=8.86 $Y2=1.41
cc_139 VPB N_Y_c_627_n 0.00113521f $X=-0.19 $Y=1.305 $X2=9.315 $Y2=0.445
cc_140 VPB N_Y_c_643_n 0.00104879f $X=-0.19 $Y=1.305 $X2=9.34 $Y2=1.985
cc_141 VPB N_Y_c_628_n 0.00113521f $X=-0.19 $Y=1.305 $X2=9.795 $Y2=0.445
cc_142 VPB N_Y_c_645_n 0.00104879f $X=-0.19 $Y=1.305 $X2=9.82 $Y2=1.985
cc_143 VPB N_Y_c_629_n 0.00113521f $X=-0.19 $Y=1.305 $X2=10.78 $Y2=1.41
cc_144 VPB N_Y_c_647_n 0.00162238f $X=-0.19 $Y=1.305 $X2=11.26 $Y2=1.985
cc_145 VPB N_Y_c_648_n 0.00178555f $X=-0.19 $Y=1.305 $X2=11.74 $Y2=1.985
cc_146 VPB N_Y_c_649_n 0.00128293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_Y_c_650_n 4.30564e-19 $X=-0.19 $Y=1.305 $X2=2.415 $Y2=1.19
cc_148 VPB N_Y_c_651_n 0.00115439f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_Y_c_652_n 4.28204e-19 $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.2
cc_150 VPB N_Y_c_653_n 0.00117346f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.16
cc_151 VPB N_Y_c_654_n 0.00197374f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.2
cc_152 N_A_c_174_n N_VPWR_c_451_n 0.00485143f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_153 A N_VPWR_c_451_n 0.00276892f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_154 N_A_c_174_n N_VPWR_c_452_n 0.00702461f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_175_n N_VPWR_c_452_n 0.00702461f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_175_n N_VPWR_c_453_n 0.00303578f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_176_n N_VPWR_c_453_n 0.00303578f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_176_n N_VPWR_c_454_n 0.00702461f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_177_n N_VPWR_c_454_n 0.00702461f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_177_n N_VPWR_c_455_n 0.0030005f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_178_n N_VPWR_c_455_n 0.00302983f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_179_n N_VPWR_c_456_n 0.00303578f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_180_n N_VPWR_c_456_n 0.00303578f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_c_181_n N_VPWR_c_457_n 0.0030005f $X=3.87 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_182_n N_VPWR_c_457_n 0.00302983f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_183_n N_VPWR_c_458_n 0.00293882f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_184_n N_VPWR_c_458_n 0.00299673f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_187_n N_VPWR_c_459_n 0.00303578f $X=5.98 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_188_n N_VPWR_c_459_n 0.00303578f $X=6.46 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_188_n N_VPWR_c_460_n 0.00702461f $X=6.46 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_189_n N_VPWR_c_460_n 0.00702461f $X=6.94 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_189_n N_VPWR_c_461_n 0.0030005f $X=6.94 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_190_n N_VPWR_c_461_n 0.00302983f $X=7.42 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_190_n N_VPWR_c_462_n 0.00702461f $X=7.42 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_191_n N_VPWR_c_462_n 0.00702461f $X=7.9 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_191_n N_VPWR_c_463_n 0.0030005f $X=7.9 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_192_n N_VPWR_c_463_n 0.00302983f $X=8.38 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_193_n N_VPWR_c_464_n 0.0030005f $X=8.86 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_194_n N_VPWR_c_464_n 0.00302983f $X=9.34 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_195_n N_VPWR_c_465_n 0.0030005f $X=9.82 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_196_n N_VPWR_c_465_n 0.00302983f $X=10.3 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_197_n N_VPWR_c_466_n 0.0030005f $X=10.78 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_198_n N_VPWR_c_466_n 0.00302983f $X=11.26 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_199_n N_VPWR_c_467_n 0.00480304f $X=11.74 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_173_n N_VPWR_c_467_n 0.00152268f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_c_178_n N_VPWR_c_468_n 0.00702461f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_c_179_n N_VPWR_c_468_n 0.00702461f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_c_180_n N_VPWR_c_470_n 0.00702461f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_181_n N_VPWR_c_470_n 0.00702461f $X=3.87 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_182_n N_VPWR_c_472_n 0.00702461f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_183_n N_VPWR_c_472_n 0.00702461f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_c_192_n N_VPWR_c_474_n 0.00702461f $X=8.38 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_c_193_n N_VPWR_c_474_n 0.00702461f $X=8.86 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_c_194_n N_VPWR_c_476_n 0.00702461f $X=9.34 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_195_n N_VPWR_c_476_n 0.00702461f $X=9.82 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_196_n N_VPWR_c_478_n 0.00702461f $X=10.3 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_197_n N_VPWR_c_478_n 0.00702461f $X=10.78 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_198_n N_VPWR_c_480_n 0.00702461f $X=11.26 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_199_n N_VPWR_c_480_n 0.00702461f $X=11.74 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_184_n N_VPWR_c_482_n 0.00702461f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_c_187_n N_VPWR_c_482_n 0.00702461f $X=5.98 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_c_174_n N_VPWR_c_449_n 0.0133471f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_c_175_n N_VPWR_c_449_n 0.0124599f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_c_176_n N_VPWR_c_449_n 0.0124927f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_177_n N_VPWR_c_449_n 0.0125053f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_178_n N_VPWR_c_449_n 0.0124927f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_c_179_n N_VPWR_c_449_n 0.0124927f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_180_n N_VPWR_c_449_n 0.0124927f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_c_181_n N_VPWR_c_449_n 0.0125053f $X=3.87 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_182_n N_VPWR_c_449_n 0.0124927f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_183_n N_VPWR_c_449_n 0.0126406f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_184_n N_VPWR_c_449_n 0.0130115f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_c_187_n N_VPWR_c_449_n 0.0128427f $X=5.98 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_c_188_n N_VPWR_c_449_n 0.0124927f $X=6.46 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_189_n N_VPWR_c_449_n 0.0125053f $X=6.94 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_190_n N_VPWR_c_449_n 0.0124927f $X=7.42 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_191_n N_VPWR_c_449_n 0.0125053f $X=7.9 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_192_n N_VPWR_c_449_n 0.0124927f $X=8.38 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_c_193_n N_VPWR_c_449_n 0.0125053f $X=8.86 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_c_194_n N_VPWR_c_449_n 0.0124927f $X=9.34 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_c_195_n N_VPWR_c_449_n 0.0125053f $X=9.82 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_196_n N_VPWR_c_449_n 0.0124927f $X=10.3 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_197_n N_VPWR_c_449_n 0.0125053f $X=10.78 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_198_n N_VPWR_c_449_n 0.0124927f $X=11.26 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_199_n N_VPWR_c_449_n 0.013511f $X=11.74 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_174_n N_Y_c_630_n 9.71261e-19 $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_c_161_n N_Y_c_630_n 0.00658682f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_228 A N_Y_c_630_n 0.0207969f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_229 N_A_c_175_n N_Y_c_631_n 0.0171085f $X=0.99 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_c_176_n N_Y_c_631_n 0.0171703f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_c_161_n N_Y_c_631_n 0.00869765f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_232 A N_Y_c_631_n 0.0506585f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A_c_177_n N_Y_c_632_n 0.0170605f $X=1.95 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_c_178_n N_Y_c_632_n 0.0174782f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_161_n N_Y_c_632_n 0.0105759f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_236 A N_Y_c_632_n 0.0302581f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_237 N_A_c_286_p N_Y_c_632_n 0.0150488f $X=2.3 $Y=1.19 $X2=0 $Y2=0
cc_238 N_A_c_287_p N_Y_c_632_n 0.00621325f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_239 N_A_M1000_g N_Y_c_622_n 0.00890007f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_240 N_A_M1005_g N_Y_c_622_n 0.00922085f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_241 N_A_c_161_n N_Y_c_622_n 0.0392547f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_242 A N_Y_c_622_n 0.0212371f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_243 N_A_c_287_p N_Y_c_622_n 0.0327219f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_244 N_A_c_293_p N_Y_c_622_n 0.00323476f $X=2.415 $Y=1.19 $X2=0 $Y2=0
cc_245 N_A_c_179_n N_Y_c_634_n 0.0192572f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_180_n N_Y_c_634_n 0.0193641f $X=3.39 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_161_n N_Y_c_634_n 0.0161743f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_248 N_A_c_287_p N_Y_c_634_n 0.0297629f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_249 N_A_M1008_g N_Y_c_623_n 0.0110171f $X=3.365 $Y=0.445 $X2=0 $Y2=0
cc_250 N_A_M1010_g N_Y_c_623_n 0.00943585f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_251 N_A_c_161_n N_Y_c_623_n 0.0488567f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_252 N_A_c_287_p N_Y_c_623_n 0.0385373f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_253 N_A_c_181_n N_Y_c_636_n 0.0193641f $X=3.87 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_182_n N_Y_c_636_n 0.0193641f $X=4.35 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_161_n N_Y_c_636_n 0.0161743f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_256 N_A_c_287_p N_Y_c_636_n 0.0297629f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_257 N_A_M1011_g N_Y_c_624_n 0.0108875f $X=4.325 $Y=0.445 $X2=0 $Y2=0
cc_258 N_A_M1013_g N_Y_c_624_n 0.00915058f $X=4.805 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_c_161_n N_Y_c_624_n 0.0477626f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_260 N_A_c_287_p N_Y_c_624_n 0.0366888f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_261 N_A_c_183_n N_Y_c_638_n 0.0196521f $X=4.83 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_184_n N_Y_c_638_n 0.0230867f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_160_n N_Y_c_638_n 4.351e-19 $X=5.88 $Y=1.17 $X2=0 $Y2=0
cc_264 N_A_c_161_n N_Y_c_638_n 0.0177489f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_265 N_A_c_287_p N_Y_c_638_n 0.0317355f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_266 N_A_M1014_g N_Y_c_625_n 0.0148494f $X=5.32 $Y=0.445 $X2=0 $Y2=0
cc_267 N_A_c_160_n N_Y_c_625_n 0.0555287f $X=5.88 $Y=1.17 $X2=0 $Y2=0
cc_268 N_A_c_161_n N_Y_c_625_n 0.00189347f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_269 N_A_M1016_g N_Y_c_625_n 0.0148387f $X=5.955 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_c_287_p N_Y_c_625_n 0.0502379f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_271 N_A_c_172_n N_Y_c_625_n 0.00173946f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_M1017_g N_Y_c_626_n 0.0109746f $X=6.435 $Y=0.445 $X2=0 $Y2=0
cc_273 N_A_M1028_g N_Y_c_626_n 0.00934041f $X=6.915 $Y=0.445 $X2=0 $Y2=0
cc_274 N_A_c_287_p N_Y_c_626_n 0.0379212f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_275 N_A_c_172_n N_Y_c_626_n 0.0484929f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_c_189_n N_Y_c_641_n 0.0193641f $X=6.94 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_c_190_n N_Y_c_641_n 0.0193641f $X=7.42 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_c_287_p N_Y_c_641_n 0.0299842f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_279 N_A_c_172_n N_Y_c_641_n 0.016416f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_M1029_g N_Y_c_627_n 0.0111734f $X=7.395 $Y=0.445 $X2=0 $Y2=0
cc_281 N_A_M1031_g N_Y_c_627_n 0.00934041f $X=7.875 $Y=0.445 $X2=0 $Y2=0
cc_282 N_A_c_287_p N_Y_c_627_n 0.0379212f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_283 N_A_c_172_n N_Y_c_627_n 0.0484929f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_c_191_n N_Y_c_643_n 0.0193641f $X=7.9 $Y=1.41 $X2=0 $Y2=0
cc_285 N_A_c_192_n N_Y_c_643_n 0.0193641f $X=8.38 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A_c_287_p N_Y_c_643_n 0.0299842f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_287 N_A_c_172_n N_Y_c_643_n 0.016416f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_288 N_A_M1033_g N_Y_c_628_n 0.0109746f $X=8.355 $Y=0.445 $X2=0 $Y2=0
cc_289 N_A_M1035_g N_Y_c_628_n 0.00934041f $X=8.835 $Y=0.445 $X2=0 $Y2=0
cc_290 N_A_c_287_p N_Y_c_628_n 0.0379212f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_291 N_A_c_172_n N_Y_c_628_n 0.0484929f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_292 N_A_c_193_n N_Y_c_645_n 0.0193641f $X=8.86 $Y=1.41 $X2=0 $Y2=0
cc_293 N_A_c_194_n N_Y_c_645_n 0.0192781f $X=9.34 $Y=1.41 $X2=0 $Y2=0
cc_294 N_A_c_287_p N_Y_c_645_n 0.0299842f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_295 N_A_c_172_n N_Y_c_645_n 0.016416f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_296 N_A_M1036_g N_Y_c_629_n 0.0109746f $X=9.315 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_M1038_g N_Y_c_629_n 0.00762872f $X=9.795 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_c_287_p N_Y_c_629_n 0.035831f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_299 N_A_c_348_p N_Y_c_629_n 0.00113197f $X=10.4 $Y=1.19 $X2=0 $Y2=0
cc_300 N_A_c_172_n N_Y_c_629_n 0.041513f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A_c_173_n N_Y_c_629_n 0.022235f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_c_195_n N_Y_c_647_n 0.0175201f $X=9.82 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_c_196_n N_Y_c_647_n 0.0170678f $X=10.3 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A_c_287_p N_Y_c_647_n 0.0112915f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_305 N_A_c_348_p N_Y_c_647_n 0.00311531f $X=10.4 $Y=1.19 $X2=0 $Y2=0
cc_306 N_A_c_172_n N_Y_c_647_n 0.00966812f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A_c_173_n N_Y_c_647_n 0.0308506f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A_c_197_n N_Y_c_648_n 0.0170605f $X=10.78 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_c_198_n N_Y_c_648_n 0.0171109f $X=11.26 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_c_359_p N_Y_c_648_n 0.0116975f $X=10.99 $Y=1.19 $X2=0 $Y2=0
cc_311 N_A_c_172_n N_Y_c_648_n 0.00907131f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_c_173_n N_Y_c_648_n 0.0452103f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_c_161_n N_Y_c_649_n 0.00658682f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_314 A N_Y_c_649_n 0.0173094f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_315 N_A_c_286_p N_Y_c_649_n 0.00572568f $X=2.3 $Y=1.19 $X2=0 $Y2=0
cc_316 N_A_c_178_n N_Y_c_650_n 0.00128387f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_c_160_n N_Y_c_651_n 0.00236888f $X=5.88 $Y=1.17 $X2=0 $Y2=0
cc_318 N_A_c_187_n N_Y_c_651_n 0.0196638f $X=5.98 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_c_188_n N_Y_c_651_n 0.0193641f $X=6.46 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A_c_287_p N_Y_c_651_n 0.0315142f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_321 N_A_c_172_n N_Y_c_651_n 0.0157121f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_322 N_A_c_195_n N_Y_c_652_n 0.00133281f $X=9.82 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_c_359_p N_Y_c_653_n 0.00610739f $X=10.99 $Y=1.19 $X2=0 $Y2=0
cc_324 N_A_c_172_n N_Y_c_653_n 0.00619936f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_c_173_n N_Y_c_653_n 0.0158536f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_326 N_A_c_199_n N_Y_c_654_n 9.77394e-19 $X=11.74 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_c_172_n N_Y_c_654_n 0.00658682f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_328 N_A_c_173_n N_Y_c_654_n 0.0207969f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_c_160_n Y 0.00135631f $X=5.88 $Y=1.17 $X2=0 $Y2=0
cc_330 N_A_c_187_n Y 0.00874017f $X=5.98 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A_c_287_p Y 0.00124485f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_332 N_A_M1000_g N_VGND_c_844_n 0.00518295f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_333 N_A_c_161_n N_VGND_c_844_n 0.00147472f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_334 A N_VGND_c_844_n 0.0131993f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_335 N_A_c_286_p N_VGND_c_844_n 0.00160784f $X=2.3 $Y=1.19 $X2=0 $Y2=0
cc_336 N_A_M1005_g N_VGND_c_845_n 0.00510286f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_337 N_A_M1008_g N_VGND_c_845_n 0.00324562f $X=3.365 $Y=0.445 $X2=0 $Y2=0
cc_338 N_A_c_161_n N_VGND_c_845_n 0.00536031f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_339 N_A_c_287_p N_VGND_c_845_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_340 N_A_M1010_g N_VGND_c_846_n 0.00510286f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_341 N_A_M1011_g N_VGND_c_846_n 0.00324562f $X=4.325 $Y=0.445 $X2=0 $Y2=0
cc_342 N_A_c_161_n N_VGND_c_846_n 0.00536031f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_343 N_A_c_287_p N_VGND_c_846_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_344 N_A_M1013_g N_VGND_c_847_n 0.00691325f $X=4.805 $Y=0.445 $X2=0 $Y2=0
cc_345 N_A_M1014_g N_VGND_c_847_n 0.00324333f $X=5.32 $Y=0.445 $X2=0 $Y2=0
cc_346 N_A_c_161_n N_VGND_c_847_n 0.00661105f $X=5.445 $Y=1.17 $X2=0 $Y2=0
cc_347 N_A_c_287_p N_VGND_c_847_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_348 N_A_M1016_g N_VGND_c_848_n 0.00542997f $X=5.955 $Y=0.445 $X2=0 $Y2=0
cc_349 N_A_M1017_g N_VGND_c_848_n 0.00324562f $X=6.435 $Y=0.445 $X2=0 $Y2=0
cc_350 N_A_c_287_p N_VGND_c_848_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_351 N_A_c_172_n N_VGND_c_848_n 0.00536031f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A_M1017_g N_VGND_c_849_n 0.00585385f $X=6.435 $Y=0.445 $X2=0 $Y2=0
cc_353 N_A_M1028_g N_VGND_c_849_n 0.00585385f $X=6.915 $Y=0.445 $X2=0 $Y2=0
cc_354 N_A_M1028_g N_VGND_c_850_n 0.00500143f $X=6.915 $Y=0.445 $X2=0 $Y2=0
cc_355 N_A_M1029_g N_VGND_c_850_n 0.00295345f $X=7.395 $Y=0.445 $X2=0 $Y2=0
cc_356 N_A_c_287_p N_VGND_c_850_n 0.00775425f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_357 N_A_c_172_n N_VGND_c_850_n 0.00536031f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_358 N_A_M1029_g N_VGND_c_851_n 0.00585385f $X=7.395 $Y=0.445 $X2=0 $Y2=0
cc_359 N_A_M1031_g N_VGND_c_851_n 0.00585385f $X=7.875 $Y=0.445 $X2=0 $Y2=0
cc_360 N_A_M1031_g N_VGND_c_852_n 0.0051287f $X=7.875 $Y=0.445 $X2=0 $Y2=0
cc_361 N_A_M1033_g N_VGND_c_852_n 0.00324562f $X=8.355 $Y=0.445 $X2=0 $Y2=0
cc_362 N_A_c_287_p N_VGND_c_852_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_363 N_A_c_172_n N_VGND_c_852_n 0.00536031f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_364 N_A_M1033_g N_VGND_c_853_n 0.00585385f $X=8.355 $Y=0.445 $X2=0 $Y2=0
cc_365 N_A_M1035_g N_VGND_c_853_n 0.00585385f $X=8.835 $Y=0.445 $X2=0 $Y2=0
cc_366 N_A_M1035_g N_VGND_c_854_n 0.0051287f $X=8.835 $Y=0.445 $X2=0 $Y2=0
cc_367 N_A_M1036_g N_VGND_c_854_n 0.00324562f $X=9.315 $Y=0.445 $X2=0 $Y2=0
cc_368 N_A_c_287_p N_VGND_c_854_n 0.00914515f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_369 N_A_c_172_n N_VGND_c_854_n 0.00536031f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_370 N_A_M1038_g N_VGND_c_855_n 0.00691977f $X=9.795 $Y=0.445 $X2=0 $Y2=0
cc_371 N_A_c_287_p N_VGND_c_855_n 0.00148989f $X=10.285 $Y=1.19 $X2=0 $Y2=0
cc_372 N_A_c_172_n N_VGND_c_855_n 0.00161098f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A_c_173_n N_VGND_c_855_n 0.0143181f $X=11.61 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_M1000_g N_VGND_c_856_n 0.00585385f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_375 N_A_M1005_g N_VGND_c_856_n 0.00585385f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_376 N_A_M1008_g N_VGND_c_858_n 0.00585385f $X=3.365 $Y=0.445 $X2=0 $Y2=0
cc_377 N_A_M1010_g N_VGND_c_858_n 0.00585385f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_378 N_A_M1011_g N_VGND_c_860_n 0.00585385f $X=4.325 $Y=0.445 $X2=0 $Y2=0
cc_379 N_A_M1013_g N_VGND_c_860_n 0.00585385f $X=4.805 $Y=0.445 $X2=0 $Y2=0
cc_380 N_A_M1036_g N_VGND_c_862_n 0.00585385f $X=9.315 $Y=0.445 $X2=0 $Y2=0
cc_381 N_A_M1038_g N_VGND_c_862_n 0.00585385f $X=9.795 $Y=0.445 $X2=0 $Y2=0
cc_382 N_A_M1014_g N_VGND_c_865_n 0.00585385f $X=5.32 $Y=0.445 $X2=0 $Y2=0
cc_383 N_A_M1016_g N_VGND_c_865_n 0.00585385f $X=5.955 $Y=0.445 $X2=0 $Y2=0
cc_384 N_A_M1000_g N_VGND_c_867_n 0.0121095f $X=2.405 $Y=0.445 $X2=0 $Y2=0
cc_385 N_A_M1005_g N_VGND_c_867_n 0.0110272f $X=2.885 $Y=0.445 $X2=0 $Y2=0
cc_386 N_A_M1008_g N_VGND_c_867_n 0.0108892f $X=3.365 $Y=0.445 $X2=0 $Y2=0
cc_387 N_A_M1010_g N_VGND_c_867_n 0.0110272f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_388 N_A_M1011_g N_VGND_c_867_n 0.0108892f $X=4.325 $Y=0.445 $X2=0 $Y2=0
cc_389 N_A_M1013_g N_VGND_c_867_n 0.0111734f $X=4.805 $Y=0.445 $X2=0 $Y2=0
cc_390 N_A_M1014_g N_VGND_c_867_n 0.0113281f $X=5.32 $Y=0.445 $X2=0 $Y2=0
cc_391 N_A_M1016_g N_VGND_c_867_n 0.0113576f $X=5.955 $Y=0.445 $X2=0 $Y2=0
cc_392 N_A_M1017_g N_VGND_c_867_n 0.0108892f $X=6.435 $Y=0.445 $X2=0 $Y2=0
cc_393 N_A_M1028_g N_VGND_c_867_n 0.0110272f $X=6.915 $Y=0.445 $X2=0 $Y2=0
cc_394 N_A_M1029_g N_VGND_c_867_n 0.0109896f $X=7.395 $Y=0.445 $X2=0 $Y2=0
cc_395 N_A_M1031_g N_VGND_c_867_n 0.0110272f $X=7.875 $Y=0.445 $X2=0 $Y2=0
cc_396 N_A_M1033_g N_VGND_c_867_n 0.0108892f $X=8.355 $Y=0.445 $X2=0 $Y2=0
cc_397 N_A_M1035_g N_VGND_c_867_n 0.0110272f $X=8.835 $Y=0.445 $X2=0 $Y2=0
cc_398 N_A_M1036_g N_VGND_c_867_n 0.0108892f $X=9.315 $Y=0.445 $X2=0 $Y2=0
cc_399 N_A_M1038_g N_VGND_c_867_n 0.0122475f $X=9.795 $Y=0.445 $X2=0 $Y2=0
cc_400 N_VPWR_c_449_n N_Y_M1001_s 0.00395511f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_449_n N_Y_M1003_s 0.00396043f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_449_n N_Y_M1006_s 0.00499658f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_c_449_n N_Y_M1009_s 0.00396043f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_449_n N_Y_M1015_s 0.00448085f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_c_449_n N_Y_M1019_s 0.00648135f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_c_449_n N_Y_M1021_s 0.0041339f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_407 N_VPWR_c_449_n N_Y_M1023_s 0.0041339f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_449_n N_Y_M1025_s 0.0041339f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_c_449_n N_Y_M1027_s 0.0041339f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_449_n N_Y_M1032_s 0.00448085f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_449_n N_Y_M1037_s 0.00396043f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_452_n N_Y_c_773_n 0.0154569f $X=1.1 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_c_449_n N_Y_c_773_n 0.00974347f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_M1002_d N_Y_c_631_n 0.00199014f $X=1.08 $Y=1.485 $X2=0 $Y2=0
cc_415 N_VPWR_c_453_n N_Y_c_631_n 0.015351f $X=1.23 $Y=2 $X2=0 $Y2=0
cc_416 N_VPWR_M1004_d N_Y_c_632_n 0.00199014f $X=2.04 $Y=1.485 $X2=0 $Y2=0
cc_417 N_VPWR_c_455_n N_Y_c_632_n 0.014828f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_418 N_VPWR_M1007_d N_Y_c_634_n 0.00200085f $X=3 $Y=1.485 $X2=0 $Y2=0
cc_419 N_VPWR_c_456_n N_Y_c_634_n 0.0150942f $X=3.15 $Y=2 $X2=0 $Y2=0
cc_420 N_VPWR_M1012_d N_Y_c_636_n 0.00200085f $X=3.96 $Y=1.485 $X2=0 $Y2=0
cc_421 N_VPWR_c_457_n N_Y_c_636_n 0.0150942f $X=4.11 $Y=2 $X2=0 $Y2=0
cc_422 N_VPWR_M1018_d N_Y_c_638_n 0.00237736f $X=4.92 $Y=1.485 $X2=0 $Y2=0
cc_423 N_VPWR_c_458_n N_Y_c_638_n 0.0179346f $X=5.09 $Y=2 $X2=0 $Y2=0
cc_424 N_VPWR_M1022_d N_Y_c_641_n 0.00200085f $X=7.03 $Y=1.485 $X2=0 $Y2=0
cc_425 N_VPWR_c_461_n N_Y_c_641_n 0.0150942f $X=7.18 $Y=2 $X2=0 $Y2=0
cc_426 N_VPWR_M1024_d N_Y_c_643_n 0.00200085f $X=7.99 $Y=1.485 $X2=0 $Y2=0
cc_427 N_VPWR_c_463_n N_Y_c_643_n 0.0150942f $X=8.14 $Y=2 $X2=0 $Y2=0
cc_428 N_VPWR_M1026_d N_Y_c_645_n 0.00200085f $X=8.95 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_464_n N_Y_c_645_n 0.0150942f $X=9.1 $Y=2 $X2=0 $Y2=0
cc_430 N_VPWR_M1030_d N_Y_c_647_n 0.00199014f $X=9.91 $Y=1.485 $X2=0 $Y2=0
cc_431 N_VPWR_c_465_n N_Y_c_647_n 0.0149091f $X=10.06 $Y=2 $X2=0 $Y2=0
cc_432 N_VPWR_M1034_d N_Y_c_648_n 0.00199014f $X=10.87 $Y=1.485 $X2=0 $Y2=0
cc_433 N_VPWR_c_466_n N_Y_c_648_n 0.014828f $X=11.02 $Y=2 $X2=0 $Y2=0
cc_434 N_VPWR_c_454_n N_Y_c_649_n 0.0141142f $X=2.065 $Y=2.72 $X2=0 $Y2=0
cc_435 N_VPWR_c_449_n N_Y_c_649_n 0.00967382f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_436 N_VPWR_c_468_n N_Y_c_650_n 0.0143924f $X=3.02 $Y=2.72 $X2=0 $Y2=0
cc_437 N_VPWR_c_449_n N_Y_c_650_n 0.0085829f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_c_470_n N_Y_c_799_n 0.0141142f $X=3.985 $Y=2.72 $X2=0 $Y2=0
cc_439 N_VPWR_c_449_n N_Y_c_799_n 0.00967382f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_440 N_VPWR_c_472_n N_Y_c_801_n 0.0136252f $X=4.965 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_449_n N_Y_c_801_n 0.00910028f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_M1020_d N_Y_c_651_n 0.00200085f $X=6.07 $Y=1.485 $X2=0 $Y2=0
cc_443 N_VPWR_c_607_p N_Y_c_651_n 0.0150942f $X=6.215 $Y=2 $X2=0 $Y2=0
cc_444 N_VPWR_c_460_n N_Y_c_805_n 0.0139512f $X=7.055 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_c_449_n N_Y_c_805_n 0.00948264f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_462_n N_Y_c_807_n 0.0139512f $X=8.015 $Y=2.72 $X2=0 $Y2=0
cc_447 N_VPWR_c_449_n N_Y_c_807_n 0.00948264f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_474_n N_Y_c_809_n 0.0139512f $X=8.975 $Y=2.72 $X2=0 $Y2=0
cc_449 N_VPWR_c_449_n N_Y_c_809_n 0.00948264f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_476_n N_Y_c_652_n 0.0139512f $X=9.935 $Y=2.72 $X2=0 $Y2=0
cc_451 N_VPWR_c_449_n N_Y_c_652_n 0.00948264f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_452 N_VPWR_c_478_n N_Y_c_653_n 0.0136252f $X=10.895 $Y=2.72 $X2=0 $Y2=0
cc_453 N_VPWR_c_449_n N_Y_c_653_n 0.00910028f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_c_480_n N_Y_c_654_n 0.0141142f $X=11.85 $Y=2.72 $X2=0 $Y2=0
cc_455 N_VPWR_c_449_n N_Y_c_654_n 0.00967382f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_456 N_VPWR_c_482_n Y 0.0227887f $X=6.09 $Y=2.72 $X2=0 $Y2=0
cc_457 N_VPWR_c_449_n Y 0.0142622f $X=12.19 $Y=2.72 $X2=0 $Y2=0
cc_458 N_Y_c_625_n N_VGND_c_848_n 0.0178784f $X=5.615 $Y=0.445 $X2=0 $Y2=0
cc_459 N_Y_c_626_n N_VGND_c_849_n 0.0138079f $X=6.7 $Y=0.445 $X2=0 $Y2=0
cc_460 N_Y_c_627_n N_VGND_c_851_n 0.0138079f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_461 N_Y_c_628_n N_VGND_c_853_n 0.0138079f $X=8.62 $Y=0.445 $X2=0 $Y2=0
cc_462 N_Y_c_622_n N_VGND_c_856_n 0.0121454f $X=2.67 $Y=0.445 $X2=0 $Y2=0
cc_463 N_Y_c_623_n N_VGND_c_858_n 0.0139627f $X=3.63 $Y=0.445 $X2=0 $Y2=0
cc_464 N_Y_c_624_n N_VGND_c_860_n 0.0134985f $X=4.59 $Y=0.445 $X2=0 $Y2=0
cc_465 N_Y_c_629_n N_VGND_c_862_n 0.0138079f $X=9.58 $Y=0.445 $X2=0 $Y2=0
cc_466 N_Y_c_625_n N_VGND_c_865_n 0.0210802f $X=5.615 $Y=0.445 $X2=0 $Y2=0
cc_467 N_Y_M1000_d N_VGND_c_867_n 0.00637397f $X=2.48 $Y=0.235 $X2=0 $Y2=0
cc_468 N_Y_M1008_d N_VGND_c_867_n 0.00533378f $X=3.44 $Y=0.235 $X2=0 $Y2=0
cc_469 N_Y_M1011_d N_VGND_c_867_n 0.00585388f $X=4.4 $Y=0.235 $X2=0 $Y2=0
cc_470 N_Y_M1014_d N_VGND_c_867_n 0.00868643f $X=5.395 $Y=0.235 $X2=0 $Y2=0
cc_471 N_Y_M1017_d N_VGND_c_867_n 0.00550715f $X=6.51 $Y=0.235 $X2=0 $Y2=0
cc_472 N_Y_M1029_d N_VGND_c_867_n 0.00550715f $X=7.47 $Y=0.235 $X2=0 $Y2=0
cc_473 N_Y_M1033_d N_VGND_c_867_n 0.00550715f $X=8.43 $Y=0.235 $X2=0 $Y2=0
cc_474 N_Y_M1036_d N_VGND_c_867_n 0.00550715f $X=9.39 $Y=0.235 $X2=0 $Y2=0
cc_475 N_Y_c_622_n N_VGND_c_867_n 0.00848423f $X=2.67 $Y=0.445 $X2=0 $Y2=0
cc_476 N_Y_c_623_n N_VGND_c_867_n 0.00962561f $X=3.63 $Y=0.445 $X2=0 $Y2=0
cc_477 N_Y_c_624_n N_VGND_c_867_n 0.00905492f $X=4.59 $Y=0.445 $X2=0 $Y2=0
cc_478 N_Y_c_625_n N_VGND_c_867_n 0.01324f $X=5.615 $Y=0.445 $X2=0 $Y2=0
cc_479 N_Y_c_626_n N_VGND_c_867_n 0.00943538f $X=6.7 $Y=0.445 $X2=0 $Y2=0
cc_480 N_Y_c_627_n N_VGND_c_867_n 0.00943538f $X=7.66 $Y=0.445 $X2=0 $Y2=0
cc_481 N_Y_c_628_n N_VGND_c_867_n 0.00943538f $X=8.62 $Y=0.445 $X2=0 $Y2=0
cc_482 N_Y_c_629_n N_VGND_c_867_n 0.00943538f $X=9.58 $Y=0.445 $X2=0 $Y2=0
