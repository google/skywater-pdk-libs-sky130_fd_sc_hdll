* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkmux2_2 VGND VPWR S A1 A0 X VPB VNB
X0 VGND S a_337_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 a_337_47# A1 a_79_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 a_79_199# A1 a_691_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X4 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X5 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_691_309# a_741_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X7 VPWR S a_335_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X8 VPWR S a_741_21# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X9 a_79_199# A0 a_570_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 a_335_309# A0 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X11 a_570_47# a_741_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND S a_741_21# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_4 VPB VNB VGND VPWR Z S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] D[0]
X0 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X5 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_559_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_3135_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X10 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_3135_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 VGND S[3] a_4006_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 a_1430_325# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR S[2] a_3135_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X22 VGND S[0] a_559_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_4006_325# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_559_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X30 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X31 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 VPWR S[3] a_4006_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X35 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X39 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 VGND S[1] a_1430_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X44 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 VGND S[2] a_3135_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X46 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X49 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X52 VPWR S[1] a_1430_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X53 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X56 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X58 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 VPWR S[0] a_559_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X62 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X63 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X68 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X69 a_1430_325# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X70 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X71 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X73 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X74 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 a_4006_325# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X77 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X78 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X79 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_1 Z VGND VPWR VNB VPB D[0] S[12] S[13] S[8] S[9]
+ S[10] S[11] S[14] S[15] D[12] D[9] D[10] D[13] D[14] D[15] D[8] D[11] S[0] S[1]
+ D[1] D[2] S[2] S[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] D[3]
X0 VGND S[11] a_1361_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X1 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VPWR S[1] a_533_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_109_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 VGND D[2] a_937_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_1840_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_1012_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X7 VGND D[4] a_1765_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_3218_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND D[10] a_937_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_2402_47# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND S[7] a_3017_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X12 VPWR S[13] a_2189_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR D[4] a_1773_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR D[10] a_945_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR S[15] a_3017_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 Z S[7] a_3230_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_937_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 a_2390_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_1574_47# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1765_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_1012_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_1765_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X23 VPWR S[11] a_1361_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_109_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X26 VGND S[13] a_2189_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X27 Z a_3017_937# a_3218_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 a_2593_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X29 VGND S[9] a_533_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X30 a_117_591# a_184_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X31 Z a_533_937# a_734_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X32 VGND S[15] a_3017_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 a_1562_591# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VPWR D[2] a_945_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 VPWR S[5] a_2189_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_2668_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X37 Z S[13] a_2402_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X38 VPWR S[7] a_3017_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VGND D[8] a_109_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 a_3230_937# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 Z a_2189_937# a_2390_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X42 a_2601_591# a_2668_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 VPWR S[3] a_1361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 Z a_3017_47# a_3218_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X45 Z S[11] a_1574_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X46 a_117_297# a_184_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X47 Z a_533_47# a_734_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X48 a_184_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X49 VGND S[3] a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_1840_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X51 VGND D[14] a_2593_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 a_2593_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X53 VGND S[1] a_533_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X54 a_184_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 a_2402_937# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_2668_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_734_591# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 a_945_591# a_1012_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X59 a_2668_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 Z a_1361_937# a_1562_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 a_1562_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_1773_591# a_1840_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X63 Z a_2189_47# a_2390_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X64 VGND S[5] a_2189_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X65 a_746_937# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X66 a_2601_297# a_2668_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 a_1012_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_184_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X69 VGND D[12] a_1765_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X70 Z S[15] a_3230_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X71 Z S[5] a_2402_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X72 a_1574_937# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X73 VPWR D[14] a_2601_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X74 a_945_297# a_1012_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X75 VGND D[0] a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X76 Z a_1361_47# a_1562_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X77 a_937_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 VPWR S[9] a_533_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X79 a_3218_591# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X80 a_1773_297# a_1840_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 Z S[3] a_1574_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X82 a_2668_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X83 a_1840_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 Z S[1] a_746_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X85 VPWR D[12] a_1773_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X86 a_734_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X87 Z S[9] a_746_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X88 a_2390_591# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X89 VGND D[6] a_2593_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X90 a_1012_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X91 a_184_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X92 a_746_47# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X93 a_1840_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X94 a_3230_47# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X95 VPWR D[6] a_2601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_2 VGND VPWR Z VNB VPB S[1] S[2] S[3] D[1] D[0]
+ D[2] D[3] S[0]
X0 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X2 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X3 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X5 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X15 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X19 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X26 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X27 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X36 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X39 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_1 VGND Z VPWR VNB VPB D[0] S[0] S[1] D[1] D[2]
+ S[2] S[3] D[4] S[4] S[5] D[5] D[6] S[6] S[7] D[7] D[3]
X0 VPWR S[1] a_533_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND D[2] a_937_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1840_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_1012_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 VGND D[4] a_1765_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_3218_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_2402_47# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND S[7] a_3017_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 VPWR D[4] a_1773_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 Z S[7] a_3230_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X10 a_2390_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_1574_47# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_1765_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X13 a_1012_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_109_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X16 a_2593_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 VPWR D[2] a_945_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR S[5] a_2189_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_2668_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 VPWR S[7] a_3017_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR S[3] a_1361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 Z a_3017_47# a_3218_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X23 a_117_297# a_184_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X24 Z a_533_47# a_734_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X25 a_184_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X26 VGND S[3] a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X27 VGND S[1] a_533_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X28 a_1562_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 Z a_2189_47# a_2390_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X30 VGND S[5] a_2189_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 a_2601_297# a_2668_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X32 Z S[5] a_2402_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 a_945_297# a_1012_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X34 VGND D[0] a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 Z a_1361_47# a_1562_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X36 a_937_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X37 a_1773_297# a_1840_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 Z S[3] a_1574_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X39 a_2668_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 Z S[1] a_746_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X41 a_734_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VGND D[6] a_2593_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_184_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 a_746_47# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 a_1840_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X46 a_3230_47# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 VPWR D[6] a_2601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_4 VGND Z VPWR VNB VPB S[6] S[10] D[12] D[13]
+ D[8] D[15] D[10] D[9] D[14] S[14] D[11] S[11] S[8] S[15] S[12] S[9] S[13] D[3] D[0]
+ D[4] D[5] D[2] D[1] D[6] S[2] S[3] S[7] S[0] S[1] S[4] S[5] D[7]
X0 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Z S[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 VGND D[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_9250_599# S[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X4 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR D[7] a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_6937_918# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND D[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Z a_4006_599# a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 VPWR D[13] a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_6937_66# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z S[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X15 Z S[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X16 VGND S[8] a_559_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X18 Z a_9250_599# a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 a_7939_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 VPWR S[8] a_559_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X21 VGND D[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND D[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR D[12] a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Z a_8379_265# a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X25 VGND D[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_4269_918# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Z S[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X28 Z a_3135_793# a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X29 Z a_5803_793# a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X30 a_559_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_7939_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_117_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VPWR D[11] a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_1430_599# S[9] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_3135_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 a_7937_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 a_9463_613# a_9250_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X40 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 a_9463_311# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X44 Z a_559_793# a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X45 a_5361_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VPWR S[14] a_8379_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X47 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_559_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 a_2693_591# a_3135_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X52 VGND S[3] a_4006_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X53 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 Z S[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 a_4219_613# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X56 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_3135_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X58 Z S[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X59 VGND S[14] a_8379_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X60 a_2695_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X61 a_9463_613# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 VPWR D[6] a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X63 Z S[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 VGND S[13] a_6674_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X65 a_4269_918# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X66 Z S[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X67 Z S[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_117_591# a_559_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_1430_325# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X70 a_6887_311# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X71 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X72 a_2693_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X73 VPWR S[2] a_3135_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X74 VGND S[0] a_559_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X75 Z a_6674_599# a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X77 VGND S[12] a_5803_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X78 a_4006_599# S[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X79 VGND S[4] a_5803_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X80 a_6674_325# S[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 a_5803_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X82 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X83 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X84 Z S[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X85 VPWR D[5] a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X86 a_4006_325# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X87 VPWR D[9] a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X88 VGND D[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X89 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X90 a_5361_297# a_5803_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X91 a_4006_599# S[11] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X92 VPWR D[10] a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X93 a_8379_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X94 a_6937_66# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X95 a_9250_325# S[7] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X96 Z S[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X97 a_1643_613# a_1430_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X98 a_9513_66# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X99 VGND D[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X100 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X101 a_6937_66# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X102 VPWR S[5] a_6674_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X103 VPWR S[12] a_5803_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X104 VPWR D[14] a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X105 VPWR D[4] a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X106 Z a_8379_793# a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X107 VGND D[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X108 a_5363_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X109 Z S[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X110 a_9513_918# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X111 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X112 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X113 VPWR S[15] a_9250_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X114 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X115 a_559_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X116 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X117 VGND D[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X118 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X119 a_5361_297# a_5803_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X120 Z S[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X121 VGND S[15] a_9250_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X122 VGND D[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X123 a_4219_613# a_4006_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X124 a_7939_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 a_6887_613# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X126 Z a_3135_793# a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X127 VPWR S[3] a_4006_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X128 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X129 a_5361_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X130 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X131 VGND D[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X132 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X133 a_8379_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X134 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X135 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X136 VGND S[7] a_9250_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X137 Z S[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X138 Z a_5803_265# a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X139 a_9513_918# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 a_9463_311# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X141 a_7937_297# a_8379_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X142 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X143 VGND S[1] a_1430_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X144 a_9463_311# a_9250_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X145 a_6937_918# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X146 a_7937_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X147 a_9513_918# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X148 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X149 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 VGND S[9] a_1430_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X151 a_9250_599# S[15] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X152 VGND S[2] a_3135_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X153 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X154 a_2695_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X155 VPWR D[12] a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X156 VGND D[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X157 a_6887_311# a_6674_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X158 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X159 a_117_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X160 a_2693_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X161 VPWR D[11] a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X162 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X163 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X164 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X165 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X166 a_1693_918# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X167 a_6937_918# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X168 a_5361_591# a_5803_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X169 Z S[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X170 VPWR D[15] a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X171 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X172 a_3135_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X173 Z a_559_793# a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X174 VPWR S[1] a_1430_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X175 a_6674_325# S[5] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X176 VPWR D[6] a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X177 a_7939_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X178 a_5803_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X179 Z a_6674_325# a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X180 a_3135_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X181 VGND D[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X182 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X183 a_8379_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X184 Z S[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X185 a_1430_599# S[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X186 a_4219_613# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X187 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X188 Z a_9250_325# a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X189 a_7939_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X190 a_2695_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X191 VPWR S[10] a_3135_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X192 Z a_4006_599# a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X193 a_5361_591# a_5803_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X194 a_9250_325# S[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X195 a_6887_311# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X196 a_1643_613# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X197 a_6674_599# S[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X198 Z S[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X199 a_5363_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X200 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X201 a_6887_311# a_6674_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X202 a_9513_918# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X203 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X204 a_9513_66# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X205 Z a_1430_599# a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X206 VGND D[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X207 a_7939_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X208 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X209 a_6937_918# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X210 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X211 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X212 Z S[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X213 Z a_8379_265# a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X214 VGND D[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X215 a_4269_918# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X216 Z S[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X217 Z a_5803_793# a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X218 VPWR D[9] a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X219 VPWR S[13] a_6674_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X220 a_7937_591# a_8379_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X221 a_119_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X222 VPWR S[0] a_559_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X223 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X224 Z S[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X225 a_7937_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X226 VGND D[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X227 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X228 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X229 a_7939_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X230 a_1643_613# a_1430_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X231 VGND D[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X232 a_9463_613# a_9250_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X233 VGND S[6] a_8379_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X234 a_559_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X235 a_5361_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X236 VPWR D[13] a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X237 a_7937_297# a_8379_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X238 VPWR D[4] a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X239 a_2693_591# a_3135_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X240 a_1693_918# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X241 a_5363_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X242 a_6887_613# a_6674_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X243 Z S[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X244 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X245 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X246 VPWR S[11] a_4006_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X247 a_7939_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X248 VPWR D[15] a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X249 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X250 VPWR S[6] a_8379_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X251 a_5363_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X252 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X253 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X254 a_9513_66# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X255 VGND D[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X256 a_1430_325# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X257 VPWR D[7] a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X258 a_1693_918# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X259 a_8379_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X260 VGND D[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X261 a_9513_66# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X262 Z a_9250_325# a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X263 Z a_6674_599# a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X264 a_5363_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X265 a_5363_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X266 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X267 VGND D[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X268 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X269 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X270 Z a_5803_265# a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X271 a_119_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X272 VGND S[11] a_4006_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X273 a_6674_599# S[13] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X274 Z a_9250_599# a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X275 Z S[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X276 VPWR D[10] a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X277 VGND D[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X278 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X279 a_4006_325# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X280 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X281 a_9463_311# a_9250_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X282 a_5803_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X283 a_5803_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X284 a_7937_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X285 a_2695_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X286 a_6887_613# a_6674_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X287 a_9463_613# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X288 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X289 VGND D[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X290 Z S[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X291 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X292 VGND D[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X293 a_1693_918# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X294 VGND S[10] a_3135_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X295 a_117_591# a_559_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X296 a_6937_66# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X297 Z a_8379_793# a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X298 Z S[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X299 a_119_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X300 a_1643_613# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X301 VGND S[5] a_6674_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X302 a_4269_918# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X303 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X304 VPWR S[9] a_1430_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X305 VPWR S[4] a_5803_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X306 Z a_1430_599# a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X307 VPWR D[14] a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X308 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X309 a_5363_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X310 a_4219_613# a_4006_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X311 a_6887_613# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X312 a_119_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X313 VPWR S[7] a_9250_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X314 VPWR D[5] a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X315 a_5361_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X316 a_5363_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X317 a_7937_591# a_8379_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X318 VGND D[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X319 Z a_6674_325# a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
.subckt sky130_fd_sc_hdll__clkmux2_1 VGND VPWR S A1 A0 X VPB VNB
X0 VPWR S a_649_21# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X1 a_243_309# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X2 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VPWR S a_243_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X4 a_79_21# A1 a_599_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X5 VGND S a_649_21# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X6 a_79_21# A0 a_478_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_478_47# a_649_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND S a_245_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X10 a_245_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_599_309# a_649_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
.ends
.subckt sky130_fd_sc_hdll__muxb16to1_2 Z VGND VPWR VNB VPB D[2] D[1] S[7] S[6] S[5]
+ D[9] D[8] S[14] S[13] S[12] S[11] S[10] S[9] S[8] D[15] D[14] D[13] D[12] D[11]
+ D[10] S[15] S[4] S[3] S[2] S[1] S[0] D[7] D[6] D[5] D[4] D[3] D[0]
X0 a_27_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_3421_915# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2603_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_3891_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_4709_915# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X6 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X7 VGND S[13] a_3277_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_1566_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_3891_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X10 VPWR D[5] a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Z a_4142_793# a_3891_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 a_27_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND D[15] a_4709_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X15 VGND S[11] a_1989_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X16 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_4688_591# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND D[13] a_3421_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z S[15] a_4709_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_4142_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X22 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_1315_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR S[9] a_701_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Z a_701_937# a_824_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_3400_591# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_3891_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VPWR D[12] a_2603_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_1315_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X30 a_27_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 Z a_4142_265# a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X34 a_824_591# a_701_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X35 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VGND D[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VGND S[15] a_4565_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X38 a_27_591# a_278_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X39 a_2112_591# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 a_278_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_2603_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VPWR D[9] a_824_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 VPWR D[10] a_1315_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 VGND S[5] a_3277_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VGND S[7] a_4565_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 Z S[10] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 VPWR S[15] a_4565_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_4688_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 Z a_4565_937# a_4688_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X51 VGND D[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X53 a_824_591# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 a_1315_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 a_2603_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 a_3421_69# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 a_3891_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_2603_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X63 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 a_3891_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_3400_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 a_3891_591# a_4142_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 Z a_3277_937# a_3400_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X68 VPWR S[13] a_3277_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X69 a_2854_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X70 Z S[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X71 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 a_4142_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X73 a_4142_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X74 VPWR D[4] a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 VGND D[14] a_3891_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X76 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X77 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 VGND D[12] a_2603_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X79 Z S[9] a_845_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X80 Z a_4565_47# a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 VPWR D[8] a_27_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X82 Z S[14] a_3891_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X83 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X85 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X86 a_2603_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X87 a_2854_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X88 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X89 Z S[12] a_2603_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X90 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X91 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X92 a_2603_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X93 a_3891_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X94 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X95 VPWR S[7] a_4565_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X96 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X97 Z S[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X98 VPWR D[15] a_4688_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X99 a_845_915# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X100 Z S[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X101 a_3891_297# a_4142_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X102 Z a_3277_47# a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X103 a_2133_915# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X104 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X105 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X106 Z a_2854_793# a_2603_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X107 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X108 a_4709_69# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X109 a_4709_915# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X110 VGND S[9] a_701_937# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X111 VPWR S[5] a_3277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X112 VPWR S[11] a_1989_937# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X113 a_4142_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X114 VPWR D[14] a_3891_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X115 a_2603_591# a_2854_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X116 a_4688_591# a_4565_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X117 VGND D[9] a_845_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X118 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X119 Z a_1566_793# a_1315_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X120 a_3421_69# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X121 Z S[11] a_2133_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X122 a_4709_69# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X123 VGND D[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X124 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X126 a_2854_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X127 a_1315_591# a_1566_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X128 a_3400_591# a_3277_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X129 Z a_2854_265# a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X130 a_2133_915# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X131 a_3421_915# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X132 Z a_1989_937# a_2112_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X133 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X134 VPWR D[7] a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X135 VGND D[10] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X136 VPWR D[13] a_3400_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X137 VGND D[8] a_27_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X138 a_845_915# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X139 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 a_2603_297# a_2854_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X141 a_4688_333# a_4565_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X142 a_2112_591# a_1989_937# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X143 VGND D[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X144 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X145 Z S[8] a_27_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X146 VGND D[11] a_2133_915# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X147 VPWR D[6] a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X148 Z a_278_793# a_27_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X149 Z S[13] a_3421_915# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 VPWR D[11] a_2112_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X151 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X152 Z S[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X153 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X154 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X155 a_3400_333# a_3277_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X156 a_2854_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X157 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X158 a_1566_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X159 a_278_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
.subckt sky130_fd_sc_hdll__muxb4to1_1 S[0] D[0] D[1] S[1] S[2] D[2] D[3] S[3] VPB
+ VNB VGND VPWR Z
X0 VPWR S[1] a_533_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND D[2] a_937_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_1012_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X3 a_1574_47# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1012_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_109_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X7 VPWR D[2] a_945_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR S[3] a_1361_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_117_297# a_184_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X10 Z a_533_47# a_734_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_184_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X12 VGND S[3] a_1361_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X13 VGND S[1] a_533_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X14 a_1562_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_945_297# a_1012_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 VGND D[0] a_109_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Z a_1361_47# a_1562_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X18 a_937_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X19 Z S[3] a_1574_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 Z S[1] a_746_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X21 a_734_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_184_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_746_47# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_4 VGND Z VPWR VNB VPB S[6] D[3] D[0] D[4] D[5]
+ D[2] D[1] D[6] S[2] S[3] S[7] S[0] S[1] S[4] S[5] D[7]
X0 VGND D[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_1313_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND D[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_355_613# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_3797_297# a_4239_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X5 VPWR S[6] a_4239_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X6 a_1313_591# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VPWR D[2] a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR D[5] a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR D[1] a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_4239_793# S[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_1755_793# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 a_2839_613# a_2626_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X13 VPWR D[7] a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Z S[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X15 a_142_599# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 Z a_142_325# a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X17 a_1315_911# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND D[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z a_2626_599# a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X20 a_2626_599# S[5] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR S[3] a_1755_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X22 a_3797_591# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 Z S[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X24 Z S[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X25 a_355_311# a_142_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_1313_297# a_1755_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X27 Z a_142_325# a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 Z a_4239_793# a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X29 a_1755_793# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND S[2] a_1755_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_3799_911# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 a_142_325# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X33 a_405_66# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_3799_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 a_405_66# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_2839_311# a_2626_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X37 a_355_311# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 a_1315_911# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_355_311# a_142_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X40 a_3797_591# a_4239_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X41 a_3799_911# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VPWR S[0] a_142_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 a_2839_613# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 VGND D[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 VPWR D[4] a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 a_1313_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X47 a_355_613# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 VPWR S[5] a_2626_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X49 a_3799_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_405_66# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X51 VPWR D[0] a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X52 VPWR D[6] a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X53 a_3799_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 VGND S[0] a_142_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X56 VPWR D[1] a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 VGND D[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 Z a_4239_265# a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X59 Z S[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 Z a_142_599# a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 a_3799_911# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X62 VGND D[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X63 VPWR D[7] a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X64 VPWR D[3] a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_3797_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 Z S[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X67 VPWR S[7] a_4239_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X68 a_355_613# a_142_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_1313_591# a_1755_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X70 Z a_142_599# a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X71 Z a_2626_325# a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 VGND S[1] a_142_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X73 VGND S[5] a_2626_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X74 a_2839_613# a_2626_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X75 a_3799_911# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X76 a_2626_325# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X77 a_355_613# a_142_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X78 a_2839_311# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X79 a_1315_911# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X80 a_405_918# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X81 VGND S[3] a_1755_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X82 Z a_1755_265# a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X83 a_355_311# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 a_2626_325# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X85 a_405_918# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X86 a_2889_66# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X87 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X88 VGND D[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X89 a_142_599# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X90 a_1313_297# a_1755_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X91 VPWR D[0] a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X92 Z a_4239_793# a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X93 VPWR D[6] a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X94 VPWR D[5] a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X95 VPWR D[2] a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X96 Z S[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X97 VPWR S[1] a_142_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X98 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X99 Z a_1755_265# a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X100 Z S[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X101 a_142_325# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X102 VGND D[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X103 a_4239_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X104 a_405_918# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X105 VGND D[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X106 VGND D[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X107 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X108 a_1755_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X109 a_2839_613# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X110 a_3797_297# a_4239_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X111 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X112 VGND D[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X113 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X114 Z a_2626_599# a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X115 a_405_66# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X116 a_3797_591# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X117 a_1315_911# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X118 a_1313_591# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X119 a_405_918# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X120 VPWR S[2] a_1755_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X121 VGND S[7] a_4239_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X122 a_2889_918# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X123 Z a_1755_793# a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X124 a_2889_66# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 a_2889_918# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X126 VPWR D[3] a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X127 a_4239_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X128 a_2839_311# a_2626_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X129 a_2889_918# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X130 VGND D[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X131 VGND D[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X132 a_1755_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X133 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X134 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X135 a_1313_591# a_1755_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X136 Z S[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X137 a_2889_66# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X138 Z S[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X139 Z S[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 Z S[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X141 VGND S[4] a_2626_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X142 VPWR D[4] a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X143 Z a_2626_325# a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X144 a_4239_793# S[7] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X145 VGND D[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X146 VPWR S[4] a_2626_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X147 Z a_1755_793# a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X148 Z S[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X149 Z S[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 a_3799_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X151 a_2839_311# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X152 a_2626_599# S[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X153 VGND S[6] a_4239_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X154 Z a_4239_265# a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X155 a_2889_918# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X156 a_3797_591# a_4239_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X157 Z S[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X158 a_3797_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X159 a_2889_66# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
.subckt sky130_fd_sc_hdll__clkmux2_4 VGND VPWR S A1 A0 X VPB VNB
X0 VPWR S a_523_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X1 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 a_523_309# A0 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X3 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 a_79_199# A0 a_754_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_79_199# A1 a_875_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X7 a_754_47# a_925_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X11 VGND S a_525_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_875_309# a_925_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X13 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X14 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR S a_925_21# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X16 a_525_47# A1 a_79_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND S a_925_21# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
.subckt sky130_fd_sc_hdll__muxb8to1_2 Z VGND VPWR VNB VPB D[2] D[1] S[7] S[6] S[5]
+ S[4] S[3] S[2] S[1] S[0] D[7] D[6] D[5] D[4] D[3] D[0]
X0 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_2603_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_3891_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X4 VPWR D[5] a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_3891_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X6 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X7 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Z a_4142_265# a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND D[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VGND S[5] a_3277_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 VGND S[7] a_4565_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 a_4688_333# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 VGND D[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_3421_69# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X27 VPWR D[4] a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_3400_333# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_3891_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 Z S[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 a_2854_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 a_4142_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X36 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 Z a_4565_47# a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X39 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_2603_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X44 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 VPWR S[7] a_4565_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 a_2603_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X50 Z a_3277_47# a_3400_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X51 a_3891_297# a_4142_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X52 Z S[5] a_3421_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X53 Z S[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X54 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X55 a_4709_69# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 VPWR S[5] a_3277_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_4142_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X59 a_3421_69# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 a_4709_69# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X61 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 a_2854_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X63 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 VGND D[7] a_4709_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X65 Z a_2854_265# a_2603_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X66 VPWR D[7] a_4688_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X67 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_2603_297# a_2854_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X70 a_4688_333# a_4565_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X71 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 VGND D[4] a_2603_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X73 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X74 VPWR D[6] a_3891_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 a_3400_333# a_3277_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X77 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X78 Z S[6] a_3891_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X79 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
* Top level circuit sky130_fd_sc_hdll__muxb
Xsky130_fd_sc_hdll__clkmux2_2_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__clkmux2_1_0/VPWR
+ sky130_fd_sc_hdll__clkmux2_2_0/S sky130_fd_sc_hdll__clkmux2_2_0/A1 sky130_fd_sc_hdll__clkmux2_2_0/A0
+ sky130_fd_sc_hdll__clkmux2_2_0/X sky130_fd_sc_hdll__clkmux2_1_0/VPB SUBS sky130_fd_sc_hdll__clkmux2_2
Xsky130_fd_sc_hdll__muxb4to1_4_0 sky130_fd_sc_hdll__clkmux2_1_0/VPB SUBS sky130_fd_sc_hdll__clkmux2_1_0/VGND
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR sky130_fd_sc_hdll__muxb4to1_4_0/Z sky130_fd_sc_hdll__muxb4to1_4_0/S[0]
+ sky130_fd_sc_hdll__muxb4to1_4_0/S[1] sky130_fd_sc_hdll__muxb4to1_4_0/D[1] sky130_fd_sc_hdll__muxb4to1_4_0/D[2]
+ sky130_fd_sc_hdll__muxb4to1_4_0/S[2] sky130_fd_sc_hdll__muxb4to1_4_0/S[3] sky130_fd_sc_hdll__muxb4to1_4_0/D[3]
+ sky130_fd_sc_hdll__muxb4to1_4_0/D[0] sky130_fd_sc_hdll__muxb4to1_4
Xsky130_fd_sc_hdll__muxb16to1_1_0 sky130_fd_sc_hdll__muxb16to1_1_0/Z sky130_fd_sc_hdll__clkmux2_1_0/VGND
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb16to1_1_0/D[0]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[12] sky130_fd_sc_hdll__muxb16to1_1_0/S[13] sky130_fd_sc_hdll__muxb16to1_1_0/S[8]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[9] sky130_fd_sc_hdll__muxb16to1_1_0/S[10] sky130_fd_sc_hdll__muxb16to1_1_0/S[11]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[14] sky130_fd_sc_hdll__muxb16to1_1_0/S[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[12]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[9] sky130_fd_sc_hdll__muxb16to1_1_0/D[10] sky130_fd_sc_hdll__muxb16to1_1_0/D[13]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[14] sky130_fd_sc_hdll__muxb16to1_1_0/D[15] sky130_fd_sc_hdll__muxb16to1_1_0/D[8]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[11] sky130_fd_sc_hdll__muxb16to1_1_0/S[0] sky130_fd_sc_hdll__muxb16to1_1_0/S[1]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[1] sky130_fd_sc_hdll__muxb16to1_1_0/D[2] sky130_fd_sc_hdll__muxb16to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[3] sky130_fd_sc_hdll__muxb16to1_1_0/D[4] sky130_fd_sc_hdll__muxb16to1_1_0/S[4]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[5] sky130_fd_sc_hdll__muxb16to1_1_0/D[5] sky130_fd_sc_hdll__muxb16to1_1_0/D[6]
+ sky130_fd_sc_hdll__muxb16to1_1_0/S[6] sky130_fd_sc_hdll__muxb16to1_1_0/S[7] sky130_fd_sc_hdll__muxb16to1_1_0/D[7]
+ sky130_fd_sc_hdll__muxb16to1_1_0/D[3] sky130_fd_sc_hdll__muxb16to1_1
Xsky130_fd_sc_hdll__muxb4to1_2_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__clkmux2_1_0/VPWR
+ sky130_fd_sc_hdll__muxb4to1_2_0/Z SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb4to1_2_0/S[1]
+ sky130_fd_sc_hdll__muxb4to1_2_0/S[2] sky130_fd_sc_hdll__muxb4to1_2_0/S[3] sky130_fd_sc_hdll__muxb4to1_2_0/D[1]
+ sky130_fd_sc_hdll__muxb4to1_2_0/D[0] sky130_fd_sc_hdll__muxb4to1_2_0/D[2] sky130_fd_sc_hdll__muxb4to1_2_0/D[3]
+ sky130_fd_sc_hdll__muxb4to1_2_0/S[0] sky130_fd_sc_hdll__muxb4to1_2
Xsky130_fd_sc_hdll__muxb8to1_1_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__muxb8to1_1_0/Z
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb8to1_1_0/D[0]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[0] sky130_fd_sc_hdll__muxb8to1_1_0/S[1] sky130_fd_sc_hdll__muxb8to1_1_0/D[1]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[2] sky130_fd_sc_hdll__muxb8to1_1_0/S[2] sky130_fd_sc_hdll__muxb8to1_1_0/S[3]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[4] sky130_fd_sc_hdll__muxb8to1_1_0/S[4] sky130_fd_sc_hdll__muxb8to1_1_0/S[5]
+ sky130_fd_sc_hdll__muxb8to1_1_0/D[5] sky130_fd_sc_hdll__muxb8to1_1_0/D[6] sky130_fd_sc_hdll__muxb8to1_1_0/S[6]
+ sky130_fd_sc_hdll__muxb8to1_1_0/S[7] sky130_fd_sc_hdll__muxb8to1_1_0/D[7] sky130_fd_sc_hdll__muxb8to1_1_0/D[3]
+ sky130_fd_sc_hdll__muxb8to1_1
Xsky130_fd_sc_hdll__muxb16to1_4_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__muxb16to1_4_0/Z
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb16to1_4_0/S[6]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[10] sky130_fd_sc_hdll__muxb16to1_4_0/D[12] sky130_fd_sc_hdll__muxb16to1_4_0/D[13]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[8] sky130_fd_sc_hdll__muxb16to1_4_0/D[15] sky130_fd_sc_hdll__muxb16to1_4_0/D[10]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[9] sky130_fd_sc_hdll__muxb16to1_4_0/D[14] sky130_fd_sc_hdll__muxb16to1_4_0/S[14]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[11] sky130_fd_sc_hdll__muxb16to1_4_0/S[11] sky130_fd_sc_hdll__muxb16to1_4_0/S[8]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[15] sky130_fd_sc_hdll__muxb16to1_4_0/S[12] sky130_fd_sc_hdll__muxb16to1_4_0/S[9]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[13] sky130_fd_sc_hdll__muxb16to1_4_0/D[3] sky130_fd_sc_hdll__muxb16to1_4_0/D[0]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[4] sky130_fd_sc_hdll__muxb16to1_4_0/D[5] sky130_fd_sc_hdll__muxb16to1_4_0/D[2]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[1] sky130_fd_sc_hdll__muxb16to1_4_0/D[6] sky130_fd_sc_hdll__muxb16to1_4_0/S[2]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[3] sky130_fd_sc_hdll__muxb16to1_4_0/S[7] sky130_fd_sc_hdll__muxb16to1_4_0/S[0]
+ sky130_fd_sc_hdll__muxb16to1_4_0/S[1] sky130_fd_sc_hdll__muxb16to1_4_0/S[4] sky130_fd_sc_hdll__muxb16to1_4_0/S[5]
+ sky130_fd_sc_hdll__muxb16to1_4_0/D[7] sky130_fd_sc_hdll__muxb16to1_4
Xsky130_fd_sc_hdll__clkmux2_1_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__clkmux2_1_0/VPWR
+ sky130_fd_sc_hdll__clkmux2_1_0/S sky130_fd_sc_hdll__clkmux2_1_0/A1 sky130_fd_sc_hdll__clkmux2_1_0/A0
+ sky130_fd_sc_hdll__clkmux2_1_0/X sky130_fd_sc_hdll__clkmux2_1_0/VPB SUBS sky130_fd_sc_hdll__clkmux2_1
Xsky130_fd_sc_hdll__muxb16to1_2_0 sky130_fd_sc_hdll__muxb16to1_2_0/Z sky130_fd_sc_hdll__clkmux2_1_0/VGND
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb16to1_2_0/D[2]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[1] sky130_fd_sc_hdll__muxb16to1_2_0/S[7] sky130_fd_sc_hdll__muxb16to1_2_0/S[6]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[5] sky130_fd_sc_hdll__muxb16to1_2_0/D[9] sky130_fd_sc_hdll__muxb16to1_2_0/D[8]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[14] sky130_fd_sc_hdll__muxb16to1_2_0/S[13] sky130_fd_sc_hdll__muxb16to1_2_0/S[12]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[11] sky130_fd_sc_hdll__muxb16to1_2_0/S[10] sky130_fd_sc_hdll__muxb16to1_2_0/S[9]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[8] sky130_fd_sc_hdll__muxb16to1_2_0/D[15] sky130_fd_sc_hdll__muxb16to1_2_0/D[14]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[13] sky130_fd_sc_hdll__muxb16to1_2_0/D[12] sky130_fd_sc_hdll__muxb16to1_2_0/D[11]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[10] sky130_fd_sc_hdll__muxb16to1_2_0/S[15] sky130_fd_sc_hdll__muxb16to1_2_0/S[4]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[3] sky130_fd_sc_hdll__muxb16to1_2_0/S[2] sky130_fd_sc_hdll__muxb16to1_2_0/S[1]
+ sky130_fd_sc_hdll__muxb16to1_2_0/S[0] sky130_fd_sc_hdll__muxb16to1_2_0/D[7] sky130_fd_sc_hdll__muxb16to1_2_0/D[6]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[5] sky130_fd_sc_hdll__muxb16to1_2_0/D[4] sky130_fd_sc_hdll__muxb16to1_2_0/D[3]
+ sky130_fd_sc_hdll__muxb16to1_2_0/D[0] sky130_fd_sc_hdll__muxb16to1_2
Xsky130_fd_sc_hdll__muxb4to1_1_0 sky130_fd_sc_hdll__muxb4to1_1_0/S[0] sky130_fd_sc_hdll__muxb4to1_1_0/D[0]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[1] sky130_fd_sc_hdll__muxb4to1_1_0/S[2]
+ sky130_fd_sc_hdll__muxb4to1_1_0/D[2] sky130_fd_sc_hdll__muxb4to1_1_0/D[3] sky130_fd_sc_hdll__muxb4to1_1_0/S[3]
+ sky130_fd_sc_hdll__clkmux2_1_0/VPB SUBS sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__clkmux2_1_0/VPWR
+ sky130_fd_sc_hdll__muxb4to1_1_0/Z sky130_fd_sc_hdll__muxb4to1_1
Xsky130_fd_sc_hdll__muxb8to1_4_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__muxb8to1_4_0/Z
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb8to1_4_0/S[6]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[3] sky130_fd_sc_hdll__muxb8to1_4_0/D[0] sky130_fd_sc_hdll__muxb8to1_4_0/D[4]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[5] sky130_fd_sc_hdll__muxb8to1_4_0/D[2] sky130_fd_sc_hdll__muxb8to1_4_0/D[1]
+ sky130_fd_sc_hdll__muxb8to1_4_0/D[6] sky130_fd_sc_hdll__muxb8to1_4_0/S[2] sky130_fd_sc_hdll__muxb8to1_4_0/S[3]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[7] sky130_fd_sc_hdll__muxb8to1_4_0/S[0] sky130_fd_sc_hdll__muxb8to1_4_0/S[1]
+ sky130_fd_sc_hdll__muxb8to1_4_0/S[4] sky130_fd_sc_hdll__muxb8to1_4_0/S[5] sky130_fd_sc_hdll__muxb8to1_4_0/D[7]
+ sky130_fd_sc_hdll__muxb8to1_4
Xsky130_fd_sc_hdll__clkmux2_4_0 sky130_fd_sc_hdll__clkmux2_1_0/VGND sky130_fd_sc_hdll__clkmux2_1_0/VPWR
+ sky130_fd_sc_hdll__clkmux2_4_0/S sky130_fd_sc_hdll__clkmux2_4_0/A1 sky130_fd_sc_hdll__clkmux2_4_0/A0
+ sky130_fd_sc_hdll__clkmux2_4_0/X sky130_fd_sc_hdll__clkmux2_1_0/VPB SUBS sky130_fd_sc_hdll__clkmux2_4
Xsky130_fd_sc_hdll__muxb8to1_2_0 sky130_fd_sc_hdll__muxb8to1_2_0/Z sky130_fd_sc_hdll__clkmux2_1_0/VGND
+ sky130_fd_sc_hdll__clkmux2_1_0/VPWR SUBS sky130_fd_sc_hdll__clkmux2_1_0/VPB sky130_fd_sc_hdll__muxb8to1_2_0/D[2]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[1] sky130_fd_sc_hdll__muxb8to1_2_0/S[7] sky130_fd_sc_hdll__muxb8to1_2_0/S[6]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[5] sky130_fd_sc_hdll__muxb8to1_2_0/S[4] sky130_fd_sc_hdll__muxb8to1_2_0/S[3]
+ sky130_fd_sc_hdll__muxb8to1_2_0/S[2] sky130_fd_sc_hdll__muxb8to1_2_0/S[1] sky130_fd_sc_hdll__muxb8to1_2_0/S[0]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[7] sky130_fd_sc_hdll__muxb8to1_2_0/D[6] sky130_fd_sc_hdll__muxb8to1_2_0/D[5]
+ sky130_fd_sc_hdll__muxb8to1_2_0/D[4] sky130_fd_sc_hdll__muxb8to1_2_0/D[3] sky130_fd_sc_hdll__muxb8to1_2_0/D[0]
+ sky130_fd_sc_hdll__muxb8to1_2
.end
