* File: sky130_fd_sc_hdll__nor3_1.spice
* Created: Wed Sep  2 08:40:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor3_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor3_1  VNB VPB C B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_C_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.104
+ AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75001.5
+ A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.4225
+ AS=0.08775 PD=2.6 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1 SB=75000.6
+ A=0.0975 P=1.6 MULT=1
MM1003 A_117_297# N_C_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=17.7103 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.5 A=0.18 P=2.36 MULT=1
MM1000 A_211_297# N_B_M1000_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=17.7103 M=1 R=5.55556 SA=90000.6
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_211_297# VPB PHIGHVT L=0.18 W=1 AD=0.61
+ AS=0.145 PD=3.22 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90001.1
+ SB=90000.5 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__nor3_1.pxi.spice"
*
.ends
*
*
