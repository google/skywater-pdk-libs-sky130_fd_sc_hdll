* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfsbp_2 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
X0 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X1 VGND a_693_369# a_877_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 Q a_2739_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_1467_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_1870_413# a_1930_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 VPWR a_2739_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_1075_413# a_877_369# a_1177_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_199_47# a_349_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X8 a_211_369# D a_199_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X9 a_349_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 a_1075_413# a_693_369# a_1169_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 a_693_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_2739_47# a_1735_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X13 Q_N a_1735_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_199_47# a_877_369# a_1075_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X15 VPWR a_1075_413# a_1652_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X16 a_349_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1219_21# a_1075_413# a_1467_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_1169_413# a_1219_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X19 VPWR a_1735_329# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 Q_N a_1735_329# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_1219_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X22 a_199_47# a_693_369# a_1075_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND a_1075_413# a_1655_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 VPWR SCE a_211_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X25 a_1735_329# a_693_369# a_1977_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_693_369# a_877_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X27 a_295_47# a_349_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2739_47# a_1735_329# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 a_693_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X30 a_1652_329# a_693_369# a_1735_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X31 a_1977_47# a_1930_295# a_2049_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 VGND SCD a_109_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_199_47# D a_295_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X34 Q a_2739_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 VPWR a_1735_329# a_1930_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X36 a_1177_47# a_1219_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1655_47# a_877_369# a_1735_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X38 a_2049_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_1735_329# a_1930_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X40 VGND a_2739_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VPWR a_1075_413# a_1219_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X42 a_109_47# SCE a_199_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_1735_329# a_877_369# a_1870_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X44 VPWR SET_B a_1735_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X45 VGND a_1735_329# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
