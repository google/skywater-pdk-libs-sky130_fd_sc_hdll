* File: sky130_fd_sc_hdll__nor4b_1.spice
* Created: Thu Aug 27 19:17:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor4b_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor4b_1  VNB VPB C B A D_N Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* D_N	D_N
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_A_91_199#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2145 PD=0.97 PS=1.96 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.3
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_C_M1004_g N_Y_M1006_d VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.104 PD=1.03 PS=0.97 NRD=4.608 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.1235 PD=0.92 PS=1.03 NRD=0 NRS=13.836 M=1 R=4.33333 SA=75001.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_M1007_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.208425 AS=0.08775 PD=1.47617 PS=0.92 NRD=21.228 NRS=0 M=1 R=4.33333
+ SA=75001.7 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1008 N_A_91_199#_M1008_d N_D_N_M1008_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.134675 PD=1.46 PS=0.953832 NRD=12.852 NRS=49.284 M=1 R=2.8
+ SA=75002.4 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_169_297# N_A_91_199#_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.53 PD=1.29 PS=3.06 NRD=17.7103 NRS=52.1853 M=1 R=5.55556
+ SA=90000.4 SB=90002 A=0.18 P=2.36 MULT=1
MM1000 A_263_297# N_C_M1000_g A_169_297# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.145 PD=1.35 PS=1.29 NRD=23.6203 NRS=17.7103 M=1 R=5.55556 SA=90000.9
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1009 A_369_297# N_B_M1009_g A_263_297# VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.175 PD=1.29 PS=1.35 NRD=17.7103 NRS=23.6203 M=1 R=5.55556 SA=90001.4
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_369_297# VPB PHIGHVT L=0.18 W=1 AD=0.337958
+ AS=0.145 PD=2.16197 PS=1.29 NRD=16.7253 NRS=17.7103 M=1 R=5.55556 SA=90001.9
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_91_199#_M1002_d N_D_N_M1002_g N_VPWR_M1005_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.141942 PD=1.38 PS=0.908028 NRD=2.3443 NRS=132.719 M=1
+ R=2.33333 SA=90002.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_14 B B PROBETYPE=1
*
.include "sky130_fd_sc_hdll__nor4b_1.pxi.spice"
*
.ends
*
*
