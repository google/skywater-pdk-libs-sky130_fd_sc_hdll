* File: sky130_fd_sc_hdll__einvp_8.pxi.spice
* Created: Thu Aug 27 19:08:10 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVP_8%TE N_TE_c_131_n N_TE_M1031_g N_TE_c_132_n
+ N_TE_M1013_g N_TE_c_133_n N_TE_c_134_n N_TE_M1001_g N_TE_c_135_n N_TE_c_136_n
+ N_TE_M1002_g N_TE_c_137_n N_TE_c_138_n N_TE_M1010_g N_TE_c_139_n N_TE_c_140_n
+ N_TE_M1012_g N_TE_c_141_n N_TE_c_142_n N_TE_M1016_g N_TE_c_143_n N_TE_c_144_n
+ N_TE_M1022_g N_TE_c_145_n N_TE_c_146_n N_TE_M1023_g N_TE_c_147_n N_TE_c_148_n
+ N_TE_M1025_g N_TE_c_149_n N_TE_c_150_n N_TE_c_151_n N_TE_c_152_n N_TE_c_153_n
+ N_TE_c_154_n N_TE_c_155_n TE TE PM_SKY130_FD_SC_HDLL__EINVP_8%TE
x_PM_SKY130_FD_SC_HDLL__EINVP_8%A_27_47# N_A_27_47#_M1031_s N_A_27_47#_M1013_s
+ N_A_27_47#_c_275_n N_A_27_47#_M1003_g N_A_27_47#_c_276_n N_A_27_47#_c_277_n
+ N_A_27_47#_c_278_n N_A_27_47#_M1006_g N_A_27_47#_c_279_n N_A_27_47#_c_280_n
+ N_A_27_47#_M1009_g N_A_27_47#_c_281_n N_A_27_47#_c_282_n N_A_27_47#_M1014_g
+ N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_M1018_g N_A_27_47#_c_285_n
+ N_A_27_47#_c_286_n N_A_27_47#_M1027_g N_A_27_47#_c_287_n N_A_27_47#_c_288_n
+ N_A_27_47#_M1029_g N_A_27_47#_c_289_n N_A_27_47#_c_290_n N_A_27_47#_M1033_g
+ N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n N_A_27_47#_c_294_n
+ N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_297_n N_A_27_47#_c_270_n
+ N_A_27_47#_c_298_n N_A_27_47#_c_271_n N_A_27_47#_c_272_n N_A_27_47#_c_299_n
+ N_A_27_47#_c_273_n N_A_27_47#_c_274_n N_A_27_47#_c_343_n
+ PM_SKY130_FD_SC_HDLL__EINVP_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVP_8%A N_A_c_447_n N_A_M1007_g N_A_c_457_n
+ N_A_M1000_g N_A_c_448_n N_A_M1008_g N_A_c_458_n N_A_M1004_g N_A_M1017_g
+ N_A_c_459_n N_A_M1005_g N_A_M1019_g N_A_c_460_n N_A_M1011_g N_A_c_451_n
+ N_A_M1020_g N_A_c_461_n N_A_M1015_g N_A_c_452_n N_A_M1026_g N_A_c_462_n
+ N_A_M1021_g N_A_M1028_g N_A_c_463_n N_A_M1024_g N_A_M1032_g N_A_c_464_n
+ N_A_M1030_g A A A A A A A N_A_c_455_n A A A A A A
+ PM_SKY130_FD_SC_HDLL__EINVP_8%A
x_PM_SKY130_FD_SC_HDLL__EINVP_8%VPWR N_VPWR_M1013_d N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_M1018_d N_VPWR_M1029_d N_VPWR_c_584_n N_VPWR_c_585_n
+ N_VPWR_c_586_n N_VPWR_c_587_n N_VPWR_c_588_n N_VPWR_c_589_n N_VPWR_c_590_n
+ N_VPWR_c_591_n N_VPWR_c_592_n N_VPWR_c_593_n N_VPWR_c_594_n N_VPWR_c_595_n
+ VPWR N_VPWR_c_596_n N_VPWR_c_597_n N_VPWR_c_583_n N_VPWR_c_599_n
+ N_VPWR_c_600_n PM_SKY130_FD_SC_HDLL__EINVP_8%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVP_8%A_235_309# N_A_235_309#_M1003_s
+ N_A_235_309#_M1006_s N_A_235_309#_M1014_s N_A_235_309#_M1027_s
+ N_A_235_309#_M1033_s N_A_235_309#_M1004_s N_A_235_309#_M1011_s
+ N_A_235_309#_M1021_s N_A_235_309#_M1030_s N_A_235_309#_c_717_n
+ N_A_235_309#_c_718_n N_A_235_309#_c_714_n N_A_235_309#_c_731_n
+ N_A_235_309#_c_721_n N_A_235_309#_c_737_n N_A_235_309#_c_722_n
+ N_A_235_309#_c_743_n N_A_235_309#_c_745_n N_A_235_309#_c_749_n
+ N_A_235_309#_c_758_n N_A_235_309#_c_805_n N_A_235_309#_c_834_p
+ N_A_235_309#_c_760_n N_A_235_309#_c_826_p N_A_235_309#_c_762_n
+ N_A_235_309#_c_828_p N_A_235_309#_c_715_n N_A_235_309#_c_716_n
+ N_A_235_309#_c_750_n N_A_235_309#_c_752_n N_A_235_309#_c_754_n
+ N_A_235_309#_c_814_n N_A_235_309#_c_816_n N_A_235_309#_c_818_n
+ PM_SKY130_FD_SC_HDLL__EINVP_8%A_235_309#
x_PM_SKY130_FD_SC_HDLL__EINVP_8%Z N_Z_M1007_d N_Z_M1017_d N_Z_M1020_d
+ N_Z_M1028_d N_Z_M1000_d N_Z_M1005_d N_Z_M1015_d N_Z_M1024_d N_Z_c_846_n
+ N_Z_c_866_n Z Z Z Z Z Z Z Z Z N_Z_c_850_n Z N_Z_c_851_n Z Z N_Z_c_852_n
+ N_Z_c_906_n N_Z_c_910_n PM_SKY130_FD_SC_HDLL__EINVP_8%Z
x_PM_SKY130_FD_SC_HDLL__EINVP_8%VGND N_VGND_M1031_d N_VGND_M1002_s
+ N_VGND_M1012_s N_VGND_M1022_s N_VGND_M1025_s N_VGND_c_958_n N_VGND_c_959_n
+ N_VGND_c_960_n N_VGND_c_961_n N_VGND_c_962_n N_VGND_c_963_n VGND
+ N_VGND_c_964_n N_VGND_c_965_n N_VGND_c_966_n N_VGND_c_967_n N_VGND_c_968_n
+ N_VGND_c_969_n N_VGND_c_970_n N_VGND_c_971_n N_VGND_c_972_n N_VGND_c_973_n
+ N_VGND_c_974_n PM_SKY130_FD_SC_HDLL__EINVP_8%VGND
x_PM_SKY130_FD_SC_HDLL__EINVP_8%A_213_47# N_A_213_47#_M1001_d
+ N_A_213_47#_M1010_d N_A_213_47#_M1016_d N_A_213_47#_M1023_d
+ N_A_213_47#_M1007_s N_A_213_47#_M1008_s N_A_213_47#_M1019_s
+ N_A_213_47#_M1026_s N_A_213_47#_M1032_s N_A_213_47#_c_1092_n
+ N_A_213_47#_c_1094_n N_A_213_47#_c_1097_n N_A_213_47#_c_1099_n
+ N_A_213_47#_c_1100_n N_A_213_47#_c_1103_n N_A_213_47#_c_1104_n
+ N_A_213_47#_c_1107_n N_A_213_47#_c_1088_n N_A_213_47#_c_1089_n
+ N_A_213_47#_c_1090_n N_A_213_47#_c_1091_n N_A_213_47#_c_1111_n
+ N_A_213_47#_c_1112_n N_A_213_47#_c_1113_n
+ PM_SKY130_FD_SC_HDLL__EINVP_8%A_213_47#
cc_1 VNB N_TE_c_131_n 0.0193865f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_2 VNB N_TE_c_132_n 0.0409119f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_TE_c_133_n 0.0195237f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.035
cc_4 VNB N_TE_c_134_n 0.0155801f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.96
cc_5 VNB N_TE_c_135_n 0.0185436f $X=-0.19 $Y=-0.24 $X2=1.405 $Y2=1.035
cc_6 VNB N_TE_c_136_n 0.0143142f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.96
cc_7 VNB N_TE_c_137_n 0.00896117f $X=-0.19 $Y=-0.24 $X2=1.825 $Y2=1.035
cc_8 VNB N_TE_c_138_n 0.01444f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=0.96
cc_9 VNB N_TE_c_139_n 0.0113601f $X=-0.19 $Y=-0.24 $X2=2.295 $Y2=1.035
cc_10 VNB N_TE_c_140_n 0.01485f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.96
cc_11 VNB N_TE_c_141_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=2.765 $Y2=1.035
cc_12 VNB N_TE_c_142_n 0.01485f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.96
cc_13 VNB N_TE_c_143_n 0.0113601f $X=-0.19 $Y=-0.24 $X2=3.235 $Y2=1.035
cc_14 VNB N_TE_c_144_n 0.01485f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=0.96
cc_15 VNB N_TE_c_145_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=3.705 $Y2=1.035
cc_16 VNB N_TE_c_146_n 0.0152276f $X=-0.19 $Y=-0.24 $X2=3.78 $Y2=0.96
cc_17 VNB N_TE_c_147_n 0.0208718f $X=-0.19 $Y=-0.24 $X2=4.225 $Y2=1.035
cc_18 VNB N_TE_c_148_n 0.0187961f $X=-0.19 $Y=-0.24 $X2=4.3 $Y2=0.96
cc_19 VNB N_TE_c_149_n 0.00661167f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.035
cc_20 VNB N_TE_c_150_n 0.00446222f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.035
cc_21 VNB N_TE_c_151_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.9 $Y2=1.035
cc_22 VNB N_TE_c_152_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.035
cc_23 VNB N_TE_c_153_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.035
cc_24 VNB N_TE_c_154_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=1.035
cc_25 VNB N_TE_c_155_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=3.78 $Y2=1.035
cc_26 VNB TE 0.0134173f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_A_27_47#_c_270_n 0.0156779f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_28 VNB N_A_27_47#_c_271_n 0.00761104f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_29 VNB N_A_27_47#_c_272_n 7.52914e-19 $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_30 VNB N_A_27_47#_c_273_n 0.00767716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_274_n 0.0303505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_c_447_n 0.0219887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_33 VNB N_A_c_448_n 0.0164911f $X=-0.19 $Y=-0.24 $X2=0.915 $Y2=1.035
cc_34 VNB N_A_M1017_g 0.0184652f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.56
cc_35 VNB N_A_M1019_g 0.0184806f $X=-0.19 $Y=-0.24 $X2=2.295 $Y2=1.035
cc_36 VNB N_A_c_451_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=2.765 $Y2=1.035
cc_37 VNB N_A_c_452_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=2.915 $Y2=1.035
cc_38 VNB N_A_M1028_g 0.0184806f $X=-0.19 $Y=-0.24 $X2=3.78 $Y2=0.56
cc_39 VNB N_A_M1032_g 0.0241067f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.035
cc_40 VNB N_A_c_455_n 0.202919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB A 0.0240879f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VPWR_c_583_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Z_c_846_n 0.0108089f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.56
cc_44 VNB N_VGND_c_958_n 0.00244569f $X=-0.19 $Y=-0.24 $X2=1.555 $Y2=1.035
cc_45 VNB N_VGND_c_959_n 3.22956e-19 $X=-0.19 $Y=-0.24 $X2=2.295 $Y2=1.035
cc_46 VNB N_VGND_c_960_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.56
cc_47 VNB N_VGND_c_961_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=0.56
cc_48 VNB N_VGND_c_962_n 0.0124004f $X=-0.19 $Y=-0.24 $X2=3.235 $Y2=1.035
cc_49 VNB N_VGND_c_963_n 0.00526805f $X=-0.19 $Y=-0.24 $X2=3.31 $Y2=0.56
cc_50 VNB N_VGND_c_964_n 0.014319f $X=-0.19 $Y=-0.24 $X2=3.78 $Y2=0.56
cc_51 VNB N_VGND_c_965_n 0.0150315f $X=-0.19 $Y=-0.24 $X2=4.3 $Y2=0.56
cc_52 VNB N_VGND_c_966_n 0.0124004f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.035
cc_53 VNB N_VGND_c_967_n 0.0124004f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_54 VNB N_VGND_c_968_n 0.104157f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_55 VNB N_VGND_c_969_n 0.432569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_970_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_971_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_972_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_973_n 0.00502768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_974_n 0.00592999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_213_47#_c_1088_n 0.00668623f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=1.035
cc_62 VNB N_A_213_47#_c_1089_n 0.00339064f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_63 VNB N_A_213_47#_c_1090_n 0.00355109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_213_47#_c_1091_n 0.0102574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_TE_c_132_n 0.0384411f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_66 VPB TE 0.0127325f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_67 VPB N_A_27_47#_c_275_n 0.0195251f $X=-0.19 $Y=1.305 $X2=0.915 $Y2=1.035
cc_68 VPB N_A_27_47#_c_276_n 0.00987291f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_69 VPB N_A_27_47#_c_277_n 0.0100079f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_70 VPB N_A_27_47#_c_278_n 0.0160921f $X=-0.19 $Y=1.305 $X2=1.405 $Y2=1.035
cc_71 VPB N_A_27_47#_c_279_n 0.00987215f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.56
cc_72 VPB N_A_27_47#_c_280_n 0.0160921f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.035
cc_73 VPB N_A_27_47#_c_281_n 0.00987291f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_74 VPB N_A_27_47#_c_282_n 0.0160921f $X=-0.19 $Y=1.305 $X2=2.295 $Y2=1.035
cc_75 VPB N_A_27_47#_c_283_n 0.00987215f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=0.56
cc_76 VPB N_A_27_47#_c_284_n 0.0160921f $X=-0.19 $Y=1.305 $X2=2.765 $Y2=1.035
cc_77 VPB N_A_27_47#_c_285_n 0.00987291f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.56
cc_78 VPB N_A_27_47#_c_286_n 0.0160921f $X=-0.19 $Y=1.305 $X2=3.235 $Y2=1.035
cc_79 VPB N_A_27_47#_c_287_n 0.00987215f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=0.56
cc_80 VPB N_A_27_47#_c_288_n 0.0160921f $X=-0.19 $Y=1.305 $X2=3.705 $Y2=1.035
cc_81 VPB N_A_27_47#_c_289_n 0.00851129f $X=-0.19 $Y=1.305 $X2=3.78 $Y2=0.56
cc_82 VPB N_A_27_47#_c_290_n 0.0166808f $X=-0.19 $Y=1.305 $X2=4.225 $Y2=1.035
cc_83 VPB N_A_27_47#_c_291_n 0.0046927f $X=-0.19 $Y=1.305 $X2=4.3 $Y2=0.56
cc_84 VPB N_A_27_47#_c_292_n 0.0046927f $X=-0.19 $Y=1.305 $X2=4.3 $Y2=0.56
cc_85 VPB N_A_27_47#_c_293_n 0.0046927f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.035
cc_86 VPB N_A_27_47#_c_294_n 0.0046927f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.035
cc_87 VPB N_A_27_47#_c_295_n 0.0046927f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.035
cc_88 VPB N_A_27_47#_c_296_n 0.00597984f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=1.035
cc_89 VPB N_A_27_47#_c_297_n 0.00949374f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=1.035
cc_90 VPB N_A_27_47#_c_298_n 0.0198678f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_91 VPB N_A_27_47#_c_299_n 0.0173666f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_27_47#_c_273_n 0.0152209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_27_47#_c_274_n 0.00108677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_c_457_n 0.0164945f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_95 VPB N_A_c_458_n 0.0157312f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_96 VPB N_A_c_459_n 0.0158662f $X=-0.19 $Y=1.305 $X2=1.825 $Y2=1.035
cc_97 VPB N_A_c_460_n 0.0158869f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=0.96
cc_98 VPB N_A_c_461_n 0.0158869f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=0.56
cc_99 VPB N_A_c_462_n 0.0158869f $X=-0.19 $Y=1.305 $X2=3.31 $Y2=0.56
cc_100 VPB N_A_c_463_n 0.0158869f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.035
cc_101 VPB N_A_c_464_n 0.0198539f $X=-0.19 $Y=1.305 $X2=2.37 $Y2=1.035
cc_102 VPB N_A_c_455_n 0.0763706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_584_n 0.00773567f $X=-0.19 $Y=1.305 $X2=1.555 $Y2=1.035
cc_104 VPB N_VPWR_c_585_n 0.0185717f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=0.56
cc_105 VPB N_VPWR_c_586_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=2.37 $Y2=0.96
cc_106 VPB N_VPWR_c_587_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=2.445 $Y2=1.035
cc_107 VPB N_VPWR_c_588_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=3.235 $Y2=1.035
cc_108 VPB N_VPWR_c_589_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=3.31 $Y2=0.56
cc_109 VPB N_VPWR_c_590_n 0.0156737f $X=-0.19 $Y=1.305 $X2=3.78 $Y2=0.96
cc_110 VPB N_VPWR_c_591_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.78 $Y2=0.56
cc_111 VPB N_VPWR_c_592_n 0.0156737f $X=-0.19 $Y=1.305 $X2=4.225 $Y2=1.035
cc_112 VPB N_VPWR_c_593_n 0.00436868f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.035
cc_113 VPB N_VPWR_c_594_n 0.0156737f $X=-0.19 $Y=1.305 $X2=4.3 $Y2=0.56
cc_114 VPB N_VPWR_c_595_n 0.00436868f $X=-0.19 $Y=1.305 $X2=4.3 $Y2=0.56
cc_115 VPB N_VPWR_c_596_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.9 $Y2=1.035
cc_116 VPB N_VPWR_c_597_n 0.10271f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_583_n 0.0559277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_599_n 0.00638089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_600_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_235_309#_c_714_n 0.00147984f $X=-0.19 $Y=1.305 $X2=2.915
+ $Y2=1.035
cc_121 VPB N_A_235_309#_c_715_n 0.00821273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_235_309#_c_716_n 0.0371051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB Z 0.00172031f $X=-0.19 $Y=1.305 $X2=3.385 $Y2=1.035
cc_124 VPB Z 0.00174301f $X=-0.19 $Y=1.305 $X2=3.78 $Y2=0.56
cc_125 VPB Z 0.00176159f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.035
cc_126 VPB N_Z_c_850_n 0.00198646f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_127 VPB N_Z_c_851_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Z_c_852_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 TE N_A_27_47#_M1013_s 0.00430377f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_130 N_TE_c_137_n N_A_27_47#_c_276_n 0.015894f $X=1.825 $Y=1.035 $X2=0 $Y2=0
cc_131 N_TE_c_150_n N_A_27_47#_c_277_n 0.015894f $X=1.48 $Y=1.035 $X2=0 $Y2=0
cc_132 N_TE_c_139_n N_A_27_47#_c_279_n 0.015894f $X=2.295 $Y=1.035 $X2=0 $Y2=0
cc_133 N_TE_c_141_n N_A_27_47#_c_281_n 0.015894f $X=2.765 $Y=1.035 $X2=0 $Y2=0
cc_134 N_TE_c_143_n N_A_27_47#_c_283_n 0.015894f $X=3.235 $Y=1.035 $X2=0 $Y2=0
cc_135 N_TE_c_145_n N_A_27_47#_c_285_n 0.015894f $X=3.705 $Y=1.035 $X2=0 $Y2=0
cc_136 N_TE_c_147_n N_A_27_47#_c_287_n 0.015894f $X=4.225 $Y=1.035 $X2=0 $Y2=0
cc_137 N_TE_c_151_n N_A_27_47#_c_291_n 0.015894f $X=1.9 $Y=1.035 $X2=0 $Y2=0
cc_138 N_TE_c_152_n N_A_27_47#_c_292_n 0.015894f $X=2.37 $Y=1.035 $X2=0 $Y2=0
cc_139 N_TE_c_153_n N_A_27_47#_c_293_n 0.015894f $X=2.84 $Y=1.035 $X2=0 $Y2=0
cc_140 N_TE_c_154_n N_A_27_47#_c_294_n 0.015894f $X=3.31 $Y=1.035 $X2=0 $Y2=0
cc_141 N_TE_c_155_n N_A_27_47#_c_295_n 0.015894f $X=3.78 $Y=1.035 $X2=0 $Y2=0
cc_142 N_TE_c_132_n N_A_27_47#_c_298_n 0.00707894f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_143 N_TE_c_131_n N_A_27_47#_c_271_n 0.0155568f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_144 N_TE_c_132_n N_A_27_47#_c_271_n 0.00303485f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_145 N_TE_c_133_n N_A_27_47#_c_271_n 6.18261e-19 $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_146 N_TE_c_134_n N_A_27_47#_c_271_n 0.00177148f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_147 TE N_A_27_47#_c_271_n 0.019129f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_148 N_TE_c_131_n N_A_27_47#_c_272_n 0.00738997f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_149 N_TE_c_132_n N_A_27_47#_c_272_n 0.00164422f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_TE_c_133_n N_A_27_47#_c_272_n 0.00389967f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_151 N_TE_c_134_n N_A_27_47#_c_272_n 0.00311815f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_152 N_TE_c_132_n N_A_27_47#_c_299_n 0.0427085f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_153 N_TE_c_133_n N_A_27_47#_c_299_n 5.76168e-19 $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_154 TE N_A_27_47#_c_299_n 0.042355f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_155 N_TE_c_135_n N_A_27_47#_c_273_n 0.0157059f $X=1.405 $Y=1.035 $X2=0 $Y2=0
cc_156 N_TE_c_137_n N_A_27_47#_c_273_n 0.0083577f $X=1.825 $Y=1.035 $X2=0 $Y2=0
cc_157 N_TE_c_139_n N_A_27_47#_c_273_n 0.00963335f $X=2.295 $Y=1.035 $X2=0 $Y2=0
cc_158 N_TE_c_141_n N_A_27_47#_c_273_n 0.00963839f $X=2.765 $Y=1.035 $X2=0 $Y2=0
cc_159 N_TE_c_143_n N_A_27_47#_c_273_n 0.00963335f $X=3.235 $Y=1.035 $X2=0 $Y2=0
cc_160 N_TE_c_145_n N_A_27_47#_c_273_n 0.00963839f $X=3.705 $Y=1.035 $X2=0 $Y2=0
cc_161 N_TE_c_147_n N_A_27_47#_c_273_n 0.017158f $X=4.225 $Y=1.035 $X2=0 $Y2=0
cc_162 N_TE_c_149_n N_A_27_47#_c_273_n 0.0107224f $X=0.99 $Y=1.035 $X2=0 $Y2=0
cc_163 N_TE_c_150_n N_A_27_47#_c_273_n 0.00538458f $X=1.48 $Y=1.035 $X2=0 $Y2=0
cc_164 N_TE_c_151_n N_A_27_47#_c_273_n 0.0051004f $X=1.9 $Y=1.035 $X2=0 $Y2=0
cc_165 N_TE_c_152_n N_A_27_47#_c_273_n 0.0051004f $X=2.37 $Y=1.035 $X2=0 $Y2=0
cc_166 N_TE_c_153_n N_A_27_47#_c_273_n 0.0051004f $X=2.84 $Y=1.035 $X2=0 $Y2=0
cc_167 N_TE_c_154_n N_A_27_47#_c_273_n 0.0051004f $X=3.31 $Y=1.035 $X2=0 $Y2=0
cc_168 N_TE_c_155_n N_A_27_47#_c_273_n 0.0051004f $X=3.78 $Y=1.035 $X2=0 $Y2=0
cc_169 N_TE_c_147_n N_A_27_47#_c_274_n 0.00670692f $X=4.225 $Y=1.035 $X2=0 $Y2=0
cc_170 N_TE_c_132_n N_A_27_47#_c_343_n 0.0130827f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_171 N_TE_c_133_n N_A_27_47#_c_343_n 0.0149982f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_172 N_TE_c_149_n N_A_27_47#_c_343_n 8.40576e-19 $X=0.99 $Y=1.035 $X2=0 $Y2=0
cc_173 TE N_A_27_47#_c_343_n 0.025787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_174 N_TE_c_132_n N_VPWR_c_584_n 0.0144429f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_175 N_TE_c_132_n N_VPWR_c_596_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_176 N_TE_c_132_n N_VPWR_c_583_n 0.0049402f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_177 N_TE_c_132_n N_A_235_309#_c_717_n 0.00532598f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_TE_c_137_n N_A_235_309#_c_718_n 2.02846e-19 $X=1.825 $Y=1.035 $X2=0
+ $Y2=0
cc_179 N_TE_c_132_n N_A_235_309#_c_714_n 6.86088e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_TE_c_135_n N_A_235_309#_c_714_n 0.00104058f $X=1.405 $Y=1.035 $X2=0
+ $Y2=0
cc_181 N_TE_c_141_n N_A_235_309#_c_721_n 2.03088e-19 $X=2.765 $Y=1.035 $X2=0
+ $Y2=0
cc_182 N_TE_c_145_n N_A_235_309#_c_722_n 2.03088e-19 $X=3.705 $Y=1.035 $X2=0
+ $Y2=0
cc_183 N_TE_c_131_n N_VGND_c_958_n 0.00877186f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_184 N_TE_c_133_n N_VGND_c_958_n 0.00135012f $X=0.915 $Y=1.035 $X2=0 $Y2=0
cc_185 N_TE_c_134_n N_VGND_c_958_n 0.00173422f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_186 N_TE_c_134_n N_VGND_c_959_n 6.09064e-19 $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_187 N_TE_c_136_n N_VGND_c_959_n 0.00997405f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_188 N_TE_c_138_n N_VGND_c_959_n 0.00726222f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_189 N_TE_c_140_n N_VGND_c_959_n 5.61602e-19 $X=2.37 $Y=0.96 $X2=0 $Y2=0
cc_190 N_TE_c_138_n N_VGND_c_960_n 5.45578e-19 $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_191 N_TE_c_140_n N_VGND_c_960_n 0.00722185f $X=2.37 $Y=0.96 $X2=0 $Y2=0
cc_192 N_TE_c_142_n N_VGND_c_960_n 0.00748964f $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_193 N_TE_c_144_n N_VGND_c_960_n 5.61602e-19 $X=3.31 $Y=0.96 $X2=0 $Y2=0
cc_194 N_TE_c_142_n N_VGND_c_961_n 5.45578e-19 $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_195 N_TE_c_144_n N_VGND_c_961_n 0.00722185f $X=3.31 $Y=0.96 $X2=0 $Y2=0
cc_196 N_TE_c_146_n N_VGND_c_961_n 0.00751483f $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_197 N_TE_c_148_n N_VGND_c_961_n 5.2779e-19 $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_198 N_TE_c_146_n N_VGND_c_962_n 0.00341689f $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_199 N_TE_c_148_n N_VGND_c_962_n 0.00199015f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_200 N_TE_c_146_n N_VGND_c_963_n 5.79224e-19 $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_201 N_TE_c_148_n N_VGND_c_963_n 0.0110574f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_202 N_TE_c_131_n N_VGND_c_964_n 0.00341689f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_203 N_TE_c_134_n N_VGND_c_965_n 0.00585385f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_204 N_TE_c_136_n N_VGND_c_965_n 0.00199015f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_205 N_TE_c_138_n N_VGND_c_966_n 0.00341689f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_206 N_TE_c_140_n N_VGND_c_966_n 0.00341689f $X=2.37 $Y=0.96 $X2=0 $Y2=0
cc_207 N_TE_c_142_n N_VGND_c_967_n 0.00341689f $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_208 N_TE_c_144_n N_VGND_c_967_n 0.00341689f $X=3.31 $Y=0.96 $X2=0 $Y2=0
cc_209 N_TE_c_131_n N_VGND_c_969_n 0.0050171f $X=0.47 $Y=0.96 $X2=0 $Y2=0
cc_210 N_TE_c_134_n N_VGND_c_969_n 0.0109612f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_211 N_TE_c_136_n N_VGND_c_969_n 0.00283749f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_212 N_TE_c_138_n N_VGND_c_969_n 0.00415805f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_213 N_TE_c_140_n N_VGND_c_969_n 0.00415805f $X=2.37 $Y=0.96 $X2=0 $Y2=0
cc_214 N_TE_c_142_n N_VGND_c_969_n 0.00415805f $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_215 N_TE_c_144_n N_VGND_c_969_n 0.00415805f $X=3.31 $Y=0.96 $X2=0 $Y2=0
cc_216 N_TE_c_146_n N_VGND_c_969_n 0.00427783f $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_217 N_TE_c_148_n N_VGND_c_969_n 0.00290797f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_218 N_TE_c_134_n N_A_213_47#_c_1092_n 0.00452417f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_219 N_TE_c_136_n N_A_213_47#_c_1092_n 0.00413033f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_220 N_TE_c_136_n N_A_213_47#_c_1094_n 0.0100271f $X=1.48 $Y=0.96 $X2=0 $Y2=0
cc_221 N_TE_c_137_n N_A_213_47#_c_1094_n 0.00179137f $X=1.825 $Y=1.035 $X2=0
+ $Y2=0
cc_222 N_TE_c_138_n N_A_213_47#_c_1094_n 0.0106582f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_223 N_TE_c_134_n N_A_213_47#_c_1097_n 0.00182133f $X=0.99 $Y=0.96 $X2=0 $Y2=0
cc_224 N_TE_c_135_n N_A_213_47#_c_1097_n 0.00310054f $X=1.405 $Y=1.035 $X2=0
+ $Y2=0
cc_225 N_TE_c_138_n N_A_213_47#_c_1099_n 0.00426436f $X=1.9 $Y=0.96 $X2=0 $Y2=0
cc_226 N_TE_c_140_n N_A_213_47#_c_1100_n 0.0109985f $X=2.37 $Y=0.96 $X2=0 $Y2=0
cc_227 N_TE_c_141_n N_A_213_47#_c_1100_n 0.00278658f $X=2.765 $Y=1.035 $X2=0
+ $Y2=0
cc_228 N_TE_c_142_n N_A_213_47#_c_1100_n 0.0109985f $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_229 N_TE_c_142_n N_A_213_47#_c_1103_n 0.00426436f $X=2.84 $Y=0.96 $X2=0 $Y2=0
cc_230 N_TE_c_144_n N_A_213_47#_c_1104_n 0.0109985f $X=3.31 $Y=0.96 $X2=0 $Y2=0
cc_231 N_TE_c_145_n N_A_213_47#_c_1104_n 0.00278658f $X=3.705 $Y=1.035 $X2=0
+ $Y2=0
cc_232 N_TE_c_146_n N_A_213_47#_c_1104_n 0.0111434f $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_233 N_TE_c_146_n N_A_213_47#_c_1107_n 0.00431325f $X=3.78 $Y=0.96 $X2=0 $Y2=0
cc_234 N_TE_c_148_n N_A_213_47#_c_1107_n 0.00415942f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_235 N_TE_c_148_n N_A_213_47#_c_1088_n 0.0124528f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_236 N_TE_c_148_n N_A_213_47#_c_1089_n 0.00371f $X=4.3 $Y=0.96 $X2=0 $Y2=0
cc_237 N_TE_c_139_n N_A_213_47#_c_1111_n 0.00268716f $X=2.295 $Y=1.035 $X2=0
+ $Y2=0
cc_238 N_TE_c_143_n N_A_213_47#_c_1112_n 0.00268716f $X=3.235 $Y=1.035 $X2=0
+ $Y2=0
cc_239 N_TE_c_147_n N_A_213_47#_c_1113_n 0.00351409f $X=4.225 $Y=1.035 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_290_n N_A_c_457_n 0.0146185f $X=4.825 $Y=1.47 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_297_n N_A_c_457_n 0.00254398f $X=4.765 $Y=1.395 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_273_n N_A_c_455_n 0.00354582f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_274_n N_A_c_455_n 0.0158325f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_299_n N_VPWR_M1013_d 0.00571933f $X=0.712 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_245 N_A_27_47#_c_275_n N_VPWR_c_584_n 0.00320248f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_298_n N_VPWR_c_584_n 0.0263462f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_299_n N_VPWR_c_584_n 0.0276039f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_275_n N_VPWR_c_585_n 0.00622633f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_275_n N_VPWR_c_586_n 0.0128003f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_278_n N_VPWR_c_586_n 0.0111045f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_280_n N_VPWR_c_586_n 6.18043e-19 $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_278_n N_VPWR_c_587_n 6.18043e-19 $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_280_n N_VPWR_c_587_n 0.0111045f $X=2.475 $Y=1.47 $X2=0 $Y2=0
cc_254 N_A_27_47#_c_282_n N_VPWR_c_587_n 0.0111045f $X=2.945 $Y=1.47 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_284_n N_VPWR_c_587_n 6.18043e-19 $X=3.415 $Y=1.47 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_282_n N_VPWR_c_588_n 6.18043e-19 $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_284_n N_VPWR_c_588_n 0.0111045f $X=3.415 $Y=1.47 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_286_n N_VPWR_c_588_n 0.0111045f $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_288_n N_VPWR_c_588_n 6.18043e-19 $X=4.355 $Y=1.47 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_286_n N_VPWR_c_589_n 6.18043e-19 $X=3.885 $Y=1.47 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_288_n N_VPWR_c_589_n 0.0111045f $X=4.355 $Y=1.47 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_290_n N_VPWR_c_589_n 0.0121047f $X=4.825 $Y=1.47 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_278_n N_VPWR_c_590_n 0.00622633f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_280_n N_VPWR_c_590_n 0.00622633f $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_282_n N_VPWR_c_592_n 0.00622633f $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_284_n N_VPWR_c_592_n 0.00622633f $X=3.415 $Y=1.47 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_286_n N_VPWR_c_594_n 0.00622633f $X=3.885 $Y=1.47 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_288_n N_VPWR_c_594_n 0.00622633f $X=4.355 $Y=1.47 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_298_n N_VPWR_c_596_n 0.0178308f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_290_n N_VPWR_c_597_n 0.00622633f $X=4.825 $Y=1.47 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_M1013_s N_VPWR_c_583_n 0.00252291f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_275_n N_VPWR_c_583_n 0.0118107f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_278_n N_VPWR_c_583_n 0.0104011f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_280_n N_VPWR_c_583_n 0.0104011f $X=2.475 $Y=1.47 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_282_n N_VPWR_c_583_n 0.0104011f $X=2.945 $Y=1.47 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_284_n N_VPWR_c_583_n 0.0104011f $X=3.415 $Y=1.47 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_286_n N_VPWR_c_583_n 0.0104011f $X=3.885 $Y=1.47 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_288_n N_VPWR_c_583_n 0.0104011f $X=4.355 $Y=1.47 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_290_n N_VPWR_c_583_n 0.0105515f $X=4.825 $Y=1.47 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_298_n N_VPWR_c_583_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_299_n N_VPWR_c_583_n 0.00695765f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_275_n N_A_235_309#_c_717_n 0.0124981f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_283 N_A_27_47#_c_299_n N_A_235_309#_c_717_n 0.014384f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_275_n N_A_235_309#_c_718_n 0.018301f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_276_n N_A_235_309#_c_718_n 0.0024163f $X=1.915 $Y=1.395
+ $X2=0 $Y2=0
cc_286 N_A_27_47#_c_278_n N_A_235_309#_c_718_n 0.0170681f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_287 N_A_27_47#_c_273_n N_A_235_309#_c_718_n 0.0375096f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_c_299_n N_A_235_309#_c_714_n 0.0113703f $X=0.712 $Y=1.785
+ $X2=0 $Y2=0
cc_289 N_A_27_47#_c_273_n N_A_235_309#_c_714_n 0.0146313f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_278_n N_A_235_309#_c_731_n 0.00546277f $X=2.005 $Y=1.47
+ $X2=0 $Y2=0
cc_291 N_A_27_47#_c_280_n N_A_235_309#_c_731_n 0.00546277f $X=2.475 $Y=1.47
+ $X2=0 $Y2=0
cc_292 N_A_27_47#_c_280_n N_A_235_309#_c_721_n 0.0170681f $X=2.475 $Y=1.47 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_281_n N_A_235_309#_c_721_n 0.0024163f $X=2.855 $Y=1.395
+ $X2=0 $Y2=0
cc_294 N_A_27_47#_c_282_n N_A_235_309#_c_721_n 0.0170681f $X=2.945 $Y=1.47 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_273_n N_A_235_309#_c_721_n 0.0372681f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_282_n N_A_235_309#_c_737_n 0.00546277f $X=2.945 $Y=1.47
+ $X2=0 $Y2=0
cc_297 N_A_27_47#_c_284_n N_A_235_309#_c_737_n 0.00546277f $X=3.415 $Y=1.47
+ $X2=0 $Y2=0
cc_298 N_A_27_47#_c_284_n N_A_235_309#_c_722_n 0.0170681f $X=3.415 $Y=1.47 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_285_n N_A_235_309#_c_722_n 0.0024163f $X=3.795 $Y=1.395
+ $X2=0 $Y2=0
cc_300 N_A_27_47#_c_286_n N_A_235_309#_c_722_n 0.0170681f $X=3.885 $Y=1.47 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_273_n N_A_235_309#_c_722_n 0.0372681f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_c_286_n N_A_235_309#_c_743_n 0.00546277f $X=3.885 $Y=1.47
+ $X2=0 $Y2=0
cc_303 N_A_27_47#_c_288_n N_A_235_309#_c_743_n 0.00546277f $X=4.355 $Y=1.47
+ $X2=0 $Y2=0
cc_304 N_A_27_47#_c_288_n N_A_235_309#_c_745_n 0.0171405f $X=4.355 $Y=1.47 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_289_n N_A_235_309#_c_745_n 0.00262074f $X=4.605 $Y=1.395
+ $X2=0 $Y2=0
cc_306 N_A_27_47#_c_290_n N_A_235_309#_c_745_n 0.017123f $X=4.825 $Y=1.47 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_273_n N_A_235_309#_c_745_n 0.053186f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_290_n N_A_235_309#_c_749_n 0.00521089f $X=4.825 $Y=1.47
+ $X2=0 $Y2=0
cc_309 N_A_27_47#_c_279_n N_A_235_309#_c_750_n 0.0025662f $X=2.385 $Y=1.395
+ $X2=0 $Y2=0
cc_310 N_A_27_47#_c_273_n N_A_235_309#_c_750_n 0.0111227f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_283_n N_A_235_309#_c_752_n 0.0025662f $X=3.325 $Y=1.395
+ $X2=0 $Y2=0
cc_312 N_A_27_47#_c_273_n N_A_235_309#_c_752_n 0.0111227f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_c_287_n N_A_235_309#_c_754_n 0.0025662f $X=4.265 $Y=1.395
+ $X2=0 $Y2=0
cc_314 N_A_27_47#_c_273_n N_A_235_309#_c_754_n 0.0111227f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_290_n Z 4.61547e-19 $X=4.825 $Y=1.47 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_297_n Z 6.99971e-19 $X=4.765 $Y=1.395 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_273_n Z 0.0281682f $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_274_n Z 2.32681e-19 $X=4.74 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_27_47#_c_271_n N_VGND_M1031_d 0.00403359f $X=0.622 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_320 N_A_27_47#_c_272_n N_VGND_M1031_d 0.00114418f $X=0.622 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_321 N_A_27_47#_c_271_n N_VGND_c_958_n 0.0130205f $X=0.622 $Y=0.825 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_343_n N_VGND_c_958_n 0.00474116f $X=0.712 $Y=1.16 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_270_n N_VGND_c_964_n 0.0173297f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_271_n N_VGND_c_964_n 0.00235711f $X=0.622 $Y=0.825 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_M1031_s N_VGND_c_969_n 0.00230206f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_270_n N_VGND_c_969_n 0.00980382f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_271_n N_VGND_c_969_n 0.00520552f $X=0.622 $Y=0.825 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_277_n N_A_213_47#_c_1094_n 2.11378e-19 $X=1.625 $Y=1.395
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_273_n N_A_213_47#_c_1094_n 0.047625f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_271_n N_A_213_47#_c_1097_n 0.00815106f $X=0.622 $Y=0.825
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_273_n N_A_213_47#_c_1097_n 0.0138439f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_273_n N_A_213_47#_c_1100_n 0.0479154f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_333 N_A_27_47#_c_273_n N_A_213_47#_c_1104_n 0.0479154f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_296_n N_A_213_47#_c_1088_n 7.28392e-19 $X=4.355 $Y=1.395
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_273_n N_A_213_47#_c_1088_n 0.0796403f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_274_n N_A_213_47#_c_1088_n 0.00837424f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_273_n N_A_213_47#_c_1111_n 0.0135367f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_27_47#_c_273_n N_A_213_47#_c_1112_n 0.0135367f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_c_273_n N_A_213_47#_c_1113_n 0.0138438f $X=4.74 $Y=1.16 $X2=0
+ $Y2=0
cc_340 N_A_c_457_n N_VPWR_c_589_n 9.24125e-19 $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_c_457_n N_VPWR_c_597_n 0.00429453f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A_c_458_n N_VPWR_c_597_n 0.00429453f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_c_459_n N_VPWR_c_597_n 0.00429453f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_c_460_n N_VPWR_c_597_n 0.00429453f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A_c_461_n N_VPWR_c_597_n 0.00429453f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A_c_462_n N_VPWR_c_597_n 0.00429453f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_c_463_n N_VPWR_c_597_n 0.00429453f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A_c_464_n N_VPWR_c_597_n 0.00429453f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A_c_457_n N_VPWR_c_583_n 0.00621534f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_c_458_n N_VPWR_c_583_n 0.00606499f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_c_459_n N_VPWR_c_583_n 0.00606499f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_c_460_n N_VPWR_c_583_n 0.00606499f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A_c_461_n N_VPWR_c_583_n 0.00606499f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A_c_462_n N_VPWR_c_583_n 0.00606499f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A_c_463_n N_VPWR_c_583_n 0.00606499f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A_c_464_n N_VPWR_c_583_n 0.00703152f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A_c_457_n N_A_235_309#_c_745_n 0.00155606f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A_c_457_n N_A_235_309#_c_749_n 0.00491432f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_c_457_n N_A_235_309#_c_758_n 0.0122062f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A_c_458_n N_A_235_309#_c_758_n 0.013747f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_c_459_n N_A_235_309#_c_760_n 0.0122199f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A_c_460_n N_A_235_309#_c_760_n 0.013747f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_c_461_n N_A_235_309#_c_762_n 0.0122476f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_c_462_n N_A_235_309#_c_762_n 0.0137768f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_c_463_n N_A_235_309#_c_715_n 0.0122476f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A_c_464_n N_A_235_309#_c_715_n 0.0137768f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_c_464_n N_A_235_309#_c_716_n 0.0128337f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_c_455_n N_A_235_309#_c_716_n 0.00562759f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_369 A N_A_235_309#_c_716_n 0.0215429f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_370 N_A_c_448_n N_Z_c_846_n 0.00700139f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_371 N_A_M1017_g N_Z_c_846_n 0.00992634f $X=6.265 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_M1019_g N_Z_c_846_n 0.00992634f $X=6.735 $Y=0.56 $X2=0 $Y2=0
cc_373 N_A_c_451_n N_Z_c_846_n 0.00992634f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A_c_452_n N_Z_c_846_n 0.00992634f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_375 N_A_M1028_g N_Z_c_846_n 0.00992634f $X=8.145 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A_M1032_g N_Z_c_846_n 0.0116762f $X=8.615 $Y=0.56 $X2=0 $Y2=0
cc_377 N_A_c_455_n N_Z_c_846_n 0.0169289f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_378 A N_Z_c_846_n 0.200975f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_379 N_A_c_447_n N_Z_c_866_n 0.00369523f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A_c_448_n N_Z_c_866_n 0.00273142f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_c_447_n Z 0.00789115f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A_c_457_n Z 0.00543634f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A_c_448_n Z 0.00480247f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A_c_458_n Z 0.0053556f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A_M1017_g Z 8.97777e-19 $X=6.265 $Y=0.56 $X2=0 $Y2=0
cc_386 N_A_c_455_n Z 0.037262f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_387 A Z 0.0167546f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_388 N_A_c_459_n Z 0.00276155f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A_c_460_n Z 0.00112083f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_390 N_A_c_455_n Z 0.00721593f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_391 A Z 0.0278197f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_392 N_A_c_461_n Z 0.00258847f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A_c_462_n Z 0.00106327f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_394 N_A_c_455_n Z 0.00785193f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_395 A Z 0.031084f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_396 N_A_c_460_n Z 5.88772e-19 $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_397 N_A_c_461_n Z 0.00939814f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_398 N_A_c_462_n Z 0.00734069f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_399 N_A_c_463_n Z 5.53873e-19 $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_400 N_A_c_463_n Z 0.00258847f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_401 N_A_c_464_n Z 0.00286468f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_402 N_A_c_455_n Z 0.00746666f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_403 A Z 0.031085f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_404 N_A_c_462_n Z 5.88979e-19 $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_405 N_A_c_463_n Z 0.00940839f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_406 N_A_c_464_n Z 0.00653869f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_407 N_A_c_458_n N_Z_c_850_n 0.0115096f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_408 N_A_c_459_n N_Z_c_850_n 0.0101048f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_409 N_A_c_455_n N_Z_c_850_n 0.00771017f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_410 A N_Z_c_850_n 0.0209277f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_411 N_A_c_460_n N_Z_c_851_n 0.0137916f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_412 N_A_c_461_n N_Z_c_851_n 0.0101048f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_413 N_A_c_455_n N_Z_c_851_n 0.00720931f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_414 A N_Z_c_851_n 0.0401943f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_415 N_A_c_462_n N_Z_c_852_n 0.0137916f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_416 N_A_c_463_n N_Z_c_852_n 0.0101048f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_417 N_A_c_455_n N_Z_c_852_n 0.00720931f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_418 A N_Z_c_852_n 0.0401943f $X=8.94 $Y=1.19 $X2=0 $Y2=0
cc_419 N_A_c_457_n N_Z_c_906_n 0.00832922f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_420 N_A_c_458_n N_Z_c_906_n 0.00742278f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_421 N_A_c_459_n N_Z_c_906_n 5.51689e-19 $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_422 N_A_c_455_n N_Z_c_906_n 9.31598e-19 $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_423 N_A_c_458_n N_Z_c_910_n 5.86616e-19 $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_424 N_A_c_459_n N_Z_c_910_n 0.00963799f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_425 N_A_c_460_n N_Z_c_910_n 0.00742548f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_426 N_A_c_461_n N_Z_c_910_n 5.51873e-19 $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_427 N_A_c_447_n N_VGND_c_963_n 0.00275505f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A_c_447_n N_VGND_c_968_n 0.00357877f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_c_448_n N_VGND_c_968_n 0.00357877f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_430 N_A_M1017_g N_VGND_c_968_n 0.00357877f $X=6.265 $Y=0.56 $X2=0 $Y2=0
cc_431 N_A_M1019_g N_VGND_c_968_n 0.00357877f $X=6.735 $Y=0.56 $X2=0 $Y2=0
cc_432 N_A_c_451_n N_VGND_c_968_n 0.00357877f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A_c_452_n N_VGND_c_968_n 0.00357877f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_M1028_g N_VGND_c_968_n 0.00357877f $X=8.145 $Y=0.56 $X2=0 $Y2=0
cc_435 N_A_M1032_g N_VGND_c_968_n 0.00357877f $X=8.615 $Y=0.56 $X2=0 $Y2=0
cc_436 N_A_c_447_n N_VGND_c_969_n 0.00677297f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_437 N_A_c_448_n N_VGND_c_969_n 0.00548399f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A_M1017_g N_VGND_c_969_n 0.00548399f $X=6.265 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_M1019_g N_VGND_c_969_n 0.00548399f $X=6.735 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_c_451_n N_VGND_c_969_n 0.00548399f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A_c_452_n N_VGND_c_969_n 0.00548399f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_442 N_A_M1028_g N_VGND_c_969_n 0.00548399f $X=8.145 $Y=0.56 $X2=0 $Y2=0
cc_443 N_A_M1032_g N_VGND_c_969_n 0.00640469f $X=8.615 $Y=0.56 $X2=0 $Y2=0
cc_444 N_A_c_447_n N_A_213_47#_c_1091_n 0.014599f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_445 N_A_c_448_n N_A_213_47#_c_1091_n 0.00903041f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_446 N_A_M1017_g N_A_213_47#_c_1091_n 0.00903374f $X=6.265 $Y=0.56 $X2=0 $Y2=0
cc_447 N_A_M1019_g N_A_213_47#_c_1091_n 0.00903374f $X=6.735 $Y=0.56 $X2=0 $Y2=0
cc_448 N_A_c_451_n N_A_213_47#_c_1091_n 0.00903374f $X=7.205 $Y=0.995 $X2=0
+ $Y2=0
cc_449 N_A_c_452_n N_A_213_47#_c_1091_n 0.00903374f $X=7.675 $Y=0.995 $X2=0
+ $Y2=0
cc_450 N_A_M1028_g N_A_213_47#_c_1091_n 0.00903374f $X=8.145 $Y=0.56 $X2=0 $Y2=0
cc_451 N_A_M1032_g N_A_213_47#_c_1091_n 0.00903374f $X=8.615 $Y=0.56 $X2=0 $Y2=0
cc_452 N_A_c_455_n N_A_213_47#_c_1091_n 4.68623e-19 $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_453 N_VPWR_c_583_n N_A_235_309#_M1003_s 0.00429283f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_454 N_VPWR_c_583_n N_A_235_309#_M1006_s 0.00647849f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_583_n N_A_235_309#_M1014_s 0.00647849f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_583_n N_A_235_309#_M1027_s 0.00647849f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_583_n N_A_235_309#_M1033_s 0.00480254f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_583_n N_A_235_309#_M1004_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_583_n N_A_235_309#_M1011_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_583_n N_A_235_309#_M1021_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_c_583_n N_A_235_309#_M1030_s 0.00217523f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_584_n N_A_235_309#_c_717_n 0.0207729f $X=0.73 $Y=2.34 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_585_n N_A_235_309#_c_717_n 0.0146267f $X=1.605 $Y=2.72 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_586_n N_A_235_309#_c_717_n 0.0350594f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_583_n N_A_235_309#_c_717_n 0.00801045f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_M1003_d N_A_235_309#_c_718_n 0.00357692f $X=1.625 $Y=1.545 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_586_n N_A_235_309#_c_718_n 0.0171295f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_586_n N_A_235_309#_c_731_n 0.0345089f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_587_n N_A_235_309#_c_731_n 0.0345089f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_590_n N_A_235_309#_c_731_n 0.0118139f $X=2.545 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_583_n N_A_235_309#_c_731_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_472 N_VPWR_M1009_d N_A_235_309#_c_721_n 0.00357692f $X=2.565 $Y=1.545 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_587_n N_A_235_309#_c_721_n 0.0171295f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_587_n N_A_235_309#_c_737_n 0.0345089f $X=2.71 $Y=2.02 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_588_n N_A_235_309#_c_737_n 0.0345089f $X=3.65 $Y=2.02 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_592_n N_A_235_309#_c_737_n 0.0118139f $X=3.485 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_583_n N_A_235_309#_c_737_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_M1018_d N_A_235_309#_c_722_n 0.00357692f $X=3.505 $Y=1.545 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_588_n N_A_235_309#_c_722_n 0.0171295f $X=3.65 $Y=2.02 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_588_n N_A_235_309#_c_743_n 0.0345089f $X=3.65 $Y=2.02 $X2=0
+ $Y2=0
cc_481 N_VPWR_c_589_n N_A_235_309#_c_743_n 0.0345089f $X=4.59 $Y=2.02 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_594_n N_A_235_309#_c_743_n 0.0118139f $X=4.425 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_583_n N_A_235_309#_c_743_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_M1029_d N_A_235_309#_c_745_n 0.0036863f $X=4.445 $Y=1.545 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_589_n N_A_235_309#_c_745_n 0.0171295f $X=4.59 $Y=2.02 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_589_n N_A_235_309#_c_749_n 0.0247004f $X=4.59 $Y=2.02 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_597_n N_A_235_309#_c_758_n 0.0415032f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_583_n N_A_235_309#_c_758_n 0.0268781f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_589_n N_A_235_309#_c_805_n 0.0115076f $X=4.59 $Y=2.02 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_597_n N_A_235_309#_c_805_n 0.0158221f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_583_n N_A_235_309#_c_805_n 0.00866514f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_597_n N_A_235_309#_c_760_n 0.0415032f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_583_n N_A_235_309#_c_760_n 0.0268781f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_597_n N_A_235_309#_c_762_n 0.0415032f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_583_n N_A_235_309#_c_762_n 0.0268781f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_597_n N_A_235_309#_c_715_n 0.0630468f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_583_n N_A_235_309#_c_715_n 0.0386189f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_597_n N_A_235_309#_c_814_n 0.0119545f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_583_n N_A_235_309#_c_814_n 0.006547f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_c_597_n N_A_235_309#_c_816_n 0.0119545f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_501 N_VPWR_c_583_n N_A_235_309#_c_816_n 0.006547f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_502 N_VPWR_c_597_n N_A_235_309#_c_818_n 0.0119545f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_503 N_VPWR_c_583_n N_A_235_309#_c_818_n 0.006547f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_504 N_VPWR_c_583_n N_Z_M1000_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_505 N_VPWR_c_583_n N_Z_M1005_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_506 N_VPWR_c_583_n N_Z_M1015_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_507 N_VPWR_c_583_n N_Z_M1024_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_508 N_A_235_309#_c_758_n N_Z_M1000_d 0.00352848f $X=5.97 $Y=2.38 $X2=0 $Y2=0
cc_509 N_A_235_309#_c_760_n N_Z_M1005_d 0.00352848f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_510 N_A_235_309#_c_762_n N_Z_M1015_d 0.00352392f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_511 N_A_235_309#_c_715_n N_Z_M1024_d 0.00352392f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_512 N_A_235_309#_c_716_n N_Z_c_846_n 0.00157651f $X=8.942 $Y=2.295 $X2=0
+ $Y2=0
cc_513 N_A_235_309#_c_745_n Z 0.00524418f $X=4.975 $Y=1.64 $X2=0 $Y2=0
cc_514 N_A_235_309#_c_826_p Z 0.0253827f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_515 N_A_235_309#_c_762_n Z 0.0196128f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_516 N_A_235_309#_c_828_p Z 0.0208108f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_517 N_A_235_309#_c_716_n Z 0.0114695f $X=8.942 $Y=2.295 $X2=0 $Y2=0
cc_518 N_A_235_309#_c_828_p Z 0.0253827f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_519 N_A_235_309#_c_715_n Z 0.0196128f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_520 N_A_235_309#_c_716_n Z 0.0325841f $X=8.942 $Y=2.295 $X2=0 $Y2=0
cc_521 N_A_235_309#_M1004_s N_Z_c_850_n 0.00178587f $X=5.91 $Y=1.485 $X2=0 $Y2=0
cc_522 N_A_235_309#_c_834_p N_Z_c_850_n 0.0136682f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_523 N_A_235_309#_M1011_s N_Z_c_851_n 0.00178587f $X=6.85 $Y=1.485 $X2=0 $Y2=0
cc_524 N_A_235_309#_c_826_p N_Z_c_851_n 0.0136682f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_525 N_A_235_309#_M1021_s N_Z_c_852_n 0.00178587f $X=7.79 $Y=1.485 $X2=0 $Y2=0
cc_526 N_A_235_309#_c_828_p N_Z_c_852_n 0.0136682f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_527 N_A_235_309#_c_745_n N_Z_c_906_n 0.00913595f $X=4.975 $Y=1.64 $X2=0 $Y2=0
cc_528 N_A_235_309#_c_749_n N_Z_c_906_n 0.0305225f $X=5.09 $Y=1.96 $X2=0 $Y2=0
cc_529 N_A_235_309#_c_758_n N_Z_c_906_n 0.0191829f $X=5.97 $Y=2.38 $X2=0 $Y2=0
cc_530 N_A_235_309#_c_834_p N_Z_c_906_n 0.0208308f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_531 N_A_235_309#_c_834_p N_Z_c_910_n 0.0254345f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_532 N_A_235_309#_c_760_n N_Z_c_910_n 0.0192183f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_533 N_A_235_309#_c_826_p N_Z_c_910_n 0.0208308f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_534 N_Z_M1007_d N_VGND_c_969_n 0.00256987f $X=5.4 $Y=0.235 $X2=0 $Y2=0
cc_535 N_Z_M1017_d N_VGND_c_969_n 0.00256987f $X=6.34 $Y=0.235 $X2=0 $Y2=0
cc_536 N_Z_M1020_d N_VGND_c_969_n 0.00256987f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_537 N_Z_M1028_d N_VGND_c_969_n 0.00256987f $X=8.22 $Y=0.235 $X2=0 $Y2=0
cc_538 N_Z_c_846_n N_A_213_47#_M1008_s 0.00456735f $X=8.405 $Y=0.76 $X2=0 $Y2=0
cc_539 N_Z_c_846_n N_A_213_47#_M1019_s 0.00401761f $X=8.405 $Y=0.76 $X2=0 $Y2=0
cc_540 N_Z_c_846_n N_A_213_47#_M1026_s 0.00401761f $X=8.405 $Y=0.76 $X2=0 $Y2=0
cc_541 N_Z_c_846_n N_A_213_47#_M1032_s 0.00681836f $X=8.405 $Y=0.76 $X2=0 $Y2=0
cc_542 N_Z_M1007_d N_A_213_47#_c_1091_n 0.00399738f $X=5.4 $Y=0.235 $X2=0 $Y2=0
cc_543 N_Z_M1017_d N_A_213_47#_c_1091_n 0.00401386f $X=6.34 $Y=0.235 $X2=0 $Y2=0
cc_544 N_Z_M1020_d N_A_213_47#_c_1091_n 0.00400219f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_545 N_Z_M1028_d N_A_213_47#_c_1091_n 0.00401386f $X=8.22 $Y=0.235 $X2=0 $Y2=0
cc_546 N_Z_c_846_n N_A_213_47#_c_1091_n 0.177184f $X=8.405 $Y=0.76 $X2=0 $Y2=0
cc_547 N_Z_c_866_n N_A_213_47#_c_1091_n 0.0240274f $X=5.585 $Y=0.85 $X2=0 $Y2=0
cc_548 N_VGND_c_969_n N_A_213_47#_M1001_d 0.00560278f $X=8.97 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_549 N_VGND_c_969_n N_A_213_47#_M1010_d 0.00314422f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_969_n N_A_213_47#_M1016_d 0.00314422f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_969_n N_A_213_47#_M1023_d 0.00376968f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_969_n N_A_213_47#_M1007_s 0.00210127f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_553 N_VGND_c_969_n N_A_213_47#_M1008_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_554 N_VGND_c_969_n N_A_213_47#_M1019_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_969_n N_A_213_47#_M1026_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_969_n N_A_213_47#_M1032_s 0.00266737f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_959_n N_A_213_47#_c_1092_n 0.0171708f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_558 N_VGND_c_965_n N_A_213_47#_c_1092_n 0.0116627f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_969_n N_A_213_47#_c_1092_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_M1002_s N_A_213_47#_c_1094_n 0.00297022f $X=1.555 $Y=0.235 $X2=0
+ $Y2=0
cc_561 N_VGND_c_959_n N_A_213_47#_c_1094_n 0.0196541f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_562 N_VGND_c_965_n N_A_213_47#_c_1094_n 0.0023206f $X=1.475 $Y=0 $X2=0 $Y2=0
cc_563 N_VGND_c_966_n N_A_213_47#_c_1094_n 0.00310196f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_c_969_n N_A_213_47#_c_1094_n 0.0115456f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_c_959_n N_A_213_47#_c_1099_n 0.0140781f $X=1.69 $Y=0.36 $X2=0
+ $Y2=0
cc_566 N_VGND_c_966_n N_A_213_47#_c_1099_n 0.011459f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_969_n N_A_213_47#_c_1099_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_M1012_s N_A_213_47#_c_1100_n 0.0038973f $X=2.445 $Y=0.235 $X2=0
+ $Y2=0
cc_569 N_VGND_c_960_n N_A_213_47#_c_1100_n 0.0198997f $X=2.63 $Y=0.36 $X2=0
+ $Y2=0
cc_570 N_VGND_c_966_n N_A_213_47#_c_1100_n 0.00232396f $X=2.415 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_967_n N_A_213_47#_c_1100_n 0.00310196f $X=3.355 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_969_n N_A_213_47#_c_1100_n 0.0113143f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_960_n N_A_213_47#_c_1103_n 0.0140781f $X=2.63 $Y=0.36 $X2=0
+ $Y2=0
cc_574 N_VGND_c_967_n N_A_213_47#_c_1103_n 0.011459f $X=3.355 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_c_969_n N_A_213_47#_c_1103_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_M1022_s N_A_213_47#_c_1104_n 0.0038973f $X=3.385 $Y=0.235 $X2=0
+ $Y2=0
cc_577 N_VGND_c_961_n N_A_213_47#_c_1104_n 0.0198997f $X=3.57 $Y=0.36 $X2=0
+ $Y2=0
cc_578 N_VGND_c_962_n N_A_213_47#_c_1104_n 0.00310196f $X=4.295 $Y=0 $X2=0 $Y2=0
cc_579 N_VGND_c_967_n N_A_213_47#_c_1104_n 0.00232396f $X=3.355 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_969_n N_A_213_47#_c_1104_n 0.0113143f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_c_961_n N_A_213_47#_c_1107_n 0.0140781f $X=3.57 $Y=0.36 $X2=0
+ $Y2=0
cc_582 N_VGND_c_962_n N_A_213_47#_c_1107_n 0.0116627f $X=4.295 $Y=0 $X2=0 $Y2=0
cc_583 N_VGND_c_963_n N_A_213_47#_c_1107_n 0.0172059f $X=4.51 $Y=0.36 $X2=0
+ $Y2=0
cc_584 N_VGND_c_969_n N_A_213_47#_c_1107_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_M1025_s N_A_213_47#_c_1088_n 0.00522868f $X=4.375 $Y=0.235 $X2=0
+ $Y2=0
cc_586 N_VGND_c_962_n N_A_213_47#_c_1088_n 0.0023206f $X=4.295 $Y=0 $X2=0 $Y2=0
cc_587 N_VGND_c_963_n N_A_213_47#_c_1088_n 0.0250655f $X=4.51 $Y=0.36 $X2=0
+ $Y2=0
cc_588 N_VGND_c_968_n N_A_213_47#_c_1088_n 0.00296166f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_c_969_n N_A_213_47#_c_1088_n 0.0108207f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_590 N_VGND_c_963_n N_A_213_47#_c_1089_n 0.00165038f $X=4.51 $Y=0.36 $X2=0
+ $Y2=0
cc_591 N_VGND_c_963_n N_A_213_47#_c_1090_n 0.0188013f $X=4.51 $Y=0.36 $X2=0
+ $Y2=0
cc_592 N_VGND_c_968_n N_A_213_47#_c_1090_n 0.0238916f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_969_n N_A_213_47#_c_1090_n 0.0132257f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_968_n N_A_213_47#_c_1091_n 0.221762f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_969_n N_A_213_47#_c_1091_n 0.13977f $X=8.97 $Y=0 $X2=0 $Y2=0
