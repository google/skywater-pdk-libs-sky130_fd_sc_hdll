* File: sky130_fd_sc_hdll__o211ai_4.pxi.spice
* Created: Wed Sep  2 08:42:54 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211AI_4%A1 N_A1_c_98_n N_A1_M1007_g N_A1_c_106_n
+ N_A1_M1011_g N_A1_c_99_n N_A1_M1015_g N_A1_c_107_n N_A1_M1014_g N_A1_c_108_n
+ N_A1_M1017_g N_A1_c_100_n N_A1_M1016_g N_A1_c_101_n N_A1_M1024_g N_A1_c_102_n
+ N_A1_M1022_g N_A1_c_103_n N_A1_c_116_p N_A1_c_104_n A1 N_A1_c_112_n
+ N_A1_c_105_n PM_SKY130_FD_SC_HDLL__O211AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O211AI_4%A2 N_A2_c_214_n N_A2_M1000_g N_A2_c_220_n
+ N_A2_M1002_g N_A2_c_215_n N_A2_M1003_g N_A2_c_221_n N_A2_M1021_g N_A2_c_216_n
+ N_A2_M1026_g N_A2_c_222_n N_A2_M1027_g N_A2_c_223_n N_A2_M1029_g N_A2_c_217_n
+ N_A2_M1030_g A2 N_A2_c_218_n N_A2_c_219_n A2 PM_SKY130_FD_SC_HDLL__O211AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O211AI_4%B1 N_B1_c_290_n N_B1_M1008_g N_B1_c_299_n
+ N_B1_M1006_g N_B1_c_291_n N_B1_M1013_g N_B1_c_300_n N_B1_M1009_g N_B1_c_301_n
+ N_B1_M1012_g N_B1_c_292_n N_B1_M1010_g N_B1_c_293_n N_B1_M1025_g N_B1_c_294_n
+ N_B1_M1018_g N_B1_c_318_p N_B1_c_295_n B1 N_B1_c_296_n B1 N_B1_c_297_n
+ N_B1_c_298_n PM_SKY130_FD_SC_HDLL__O211AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O211AI_4%C1 N_C1_c_403_n N_C1_M1005_g N_C1_c_408_n
+ N_C1_M1001_g N_C1_c_404_n N_C1_M1004_g N_C1_c_409_n N_C1_M1019_g N_C1_c_405_n
+ N_C1_M1028_g N_C1_c_410_n N_C1_M1023_g N_C1_c_411_n N_C1_M1031_g N_C1_c_406_n
+ N_C1_M1020_g C1 N_C1_c_412_n N_C1_c_407_n C1 PM_SKY130_FD_SC_HDLL__O211AI_4%C1
x_PM_SKY130_FD_SC_HDLL__O211AI_4%VPWR N_VPWR_M1011_s N_VPWR_M1014_s
+ N_VPWR_M1024_s N_VPWR_M1009_s N_VPWR_M1001_d N_VPWR_M1023_d N_VPWR_M1025_s
+ N_VPWR_c_484_n N_VPWR_c_485_n N_VPWR_c_486_n N_VPWR_c_487_n N_VPWR_c_488_n
+ N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n N_VPWR_c_493_n
+ N_VPWR_c_494_n VPWR N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_483_n
+ PM_SKY130_FD_SC_HDLL__O211AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O211AI_4%A_118_297# N_A_118_297#_M1011_d
+ N_A_118_297#_M1017_d N_A_118_297#_M1021_s N_A_118_297#_M1029_s
+ N_A_118_297#_c_607_n N_A_118_297#_c_631_n N_A_118_297#_c_613_n
+ N_A_118_297#_c_615_n PM_SKY130_FD_SC_HDLL__O211AI_4%A_118_297#
x_PM_SKY130_FD_SC_HDLL__O211AI_4%Y N_Y_M1005_s N_Y_M1028_s N_Y_M1002_d
+ N_Y_M1027_d N_Y_M1006_d N_Y_M1012_d N_Y_M1019_s N_Y_M1031_s N_Y_c_652_n
+ N_Y_c_666_n N_Y_c_667_n N_Y_c_668_n N_Y_c_693_n N_Y_c_654_n N_Y_c_646_n
+ N_Y_c_645_n Y N_Y_c_649_n N_Y_c_656_n Y PM_SKY130_FD_SC_HDLL__O211AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O211AI_4%A_27_47# N_A_27_47#_M1007_s N_A_27_47#_M1015_s
+ N_A_27_47#_M1000_d N_A_27_47#_M1026_d N_A_27_47#_M1022_s N_A_27_47#_M1013_d
+ N_A_27_47#_M1018_d N_A_27_47#_c_760_n N_A_27_47#_c_772_n N_A_27_47#_c_761_n
+ N_A_27_47#_c_781_n N_A_27_47#_c_798_n N_A_27_47#_c_762_n N_A_27_47#_c_763_n
+ N_A_27_47#_c_764_n N_A_27_47#_c_784_n N_A_27_47#_c_765_n N_A_27_47#_c_766_n
+ PM_SKY130_FD_SC_HDLL__O211AI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O211AI_4%VGND N_VGND_M1007_d N_VGND_M1016_d
+ N_VGND_M1003_s N_VGND_M1030_s N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n
+ VGND N_VGND_c_891_n N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n
+ N_VGND_c_895_n N_VGND_c_896_n N_VGND_c_897_n N_VGND_c_898_n
+ PM_SKY130_FD_SC_HDLL__O211AI_4%VGND
x_PM_SKY130_FD_SC_HDLL__O211AI_4%A_886_47# N_A_886_47#_M1008_s
+ N_A_886_47#_M1004_d N_A_886_47#_c_1007_n
+ PM_SKY130_FD_SC_HDLL__O211AI_4%A_886_47#
cc_1 VNB N_A1_c_98_n 0.0218629f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A1_c_99_n 0.0171779f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_A1_c_100_n 0.016863f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_4 VNB N_A1_c_101_n 0.0291732f $X=-0.19 $Y=-0.24 $X2=3.86 $Y2=1.41
cc_5 VNB N_A1_c_102_n 0.0174867f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_6 VNB N_A1_c_103_n 0.00921322f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.202
cc_7 VNB N_A1_c_104_n 0.00158596f $X=-0.19 $Y=-0.24 $X2=3.855 $Y2=1.16
cc_8 VNB N_A1_c_105_n 0.0635045f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.202
cc_9 VNB N_A2_c_214_n 0.0164314f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_10 VNB N_A2_c_215_n 0.0167376f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_11 VNB N_A2_c_216_n 0.0171693f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_12 VNB N_A2_c_217_n 0.017118f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_13 VNB N_A2_c_218_n 0.00191239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_219_n 0.0756404f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.202
cc_15 VNB N_B1_c_290_n 0.0171932f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_16 VNB N_B1_c_291_n 0.017593f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_17 VNB N_B1_c_292_n 0.0172615f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.995
cc_18 VNB N_B1_c_293_n 0.0276436f $X=-0.19 $Y=-0.24 $X2=3.86 $Y2=1.41
cc_19 VNB N_B1_c_294_n 0.0204299f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_20 VNB N_B1_c_295_n 0.0010116f $X=-0.19 $Y=-0.24 $X2=3.855 $Y2=1.16
cc_21 VNB N_B1_c_296_n 0.0537902f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_22 VNB N_B1_c_297_n 0.00276098f $X=-0.19 $Y=-0.24 $X2=1.287 $Y2=1.53
cc_23 VNB N_B1_c_298_n 0.00365784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C1_c_403_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_25 VNB N_C1_c_404_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_26 VNB N_C1_c_405_n 0.0174167f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_27 VNB N_C1_c_406_n 0.0181302f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_28 VNB N_C1_c_407_n 0.0770371f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_29 VNB N_VPWR_c_483_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_645_n 0.0199827f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_31 VNB N_A_27_47#_c_760_n 0.00498999f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.995
cc_32 VNB N_A_27_47#_c_761_n 0.0146992f $X=-0.19 $Y=-0.24 $X2=1.015 $Y2=1.202
cc_33 VNB N_A_27_47#_c_762_n 0.00224113f $X=-0.19 $Y=-0.24 $X2=3.855 $Y2=1.16
cc_34 VNB N_A_27_47#_c_763_n 0.00837836f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.202
cc_35 VNB N_A_27_47#_c_764_n 4.96561e-19 $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_36 VNB N_A_27_47#_c_765_n 0.0208627f $X=-0.19 $Y=-0.24 $X2=1.287 $Y2=1.16
cc_37 VNB N_A_27_47#_c_766_n 0.0124137f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_888_n 0.0145889f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.41
cc_39 VNB N_VGND_c_889_n 3.34065e-19 $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=0.56
cc_40 VNB N_VGND_c_890_n 0.0137175f $X=-0.19 $Y=-0.24 $X2=3.86 $Y2=1.41
cc_41 VNB N_VGND_c_891_n 0.0159706f $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.56
cc_42 VNB N_VGND_c_892_n 0.0136961f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.16
cc_43 VNB N_VGND_c_893_n 0.120506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_894_n 0.416701f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=1.202
cc_45 VNB N_VGND_c_895_n 0.00547466f $X=-0.19 $Y=-0.24 $X2=1.345 $Y2=1.202
cc_46 VNB N_VGND_c_896_n 0.00436092f $X=-0.19 $Y=-0.24 $X2=1.287 $Y2=1.16
cc_47 VNB N_VGND_c_897_n 0.00537617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_898_n 0.00855845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VPB N_A1_c_106_n 0.0211647f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_50 VPB N_A1_c_107_n 0.0156758f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_51 VPB N_A1_c_108_n 0.0156704f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.41
cc_52 VPB N_A1_c_101_n 0.0275851f $X=-0.19 $Y=1.305 $X2=3.86 $Y2=1.41
cc_53 VPB N_A1_c_103_n 0.00534617f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.202
cc_54 VPB N_A1_c_104_n 0.00301589f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.16
cc_55 VPB N_A1_c_112_n 9.021e-19 $X=-0.19 $Y=1.305 $X2=1.345 $Y2=1.16
cc_56 VPB N_A1_c_105_n 0.0377353f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.202
cc_57 VPB N_A2_c_220_n 0.0165923f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_58 VPB N_A2_c_221_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_59 VPB N_A2_c_222_n 0.0164285f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=0.995
cc_60 VPB N_A2_c_223_n 0.0165879f $X=-0.19 $Y=1.305 $X2=3.86 $Y2=1.41
cc_61 VPB N_A2_c_218_n 7.05409e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A2_c_219_n 0.0454748f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=1.202
cc_63 VPB N_B1_c_299_n 0.0168695f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_64 VPB N_B1_c_300_n 0.0153391f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_65 VPB N_B1_c_301_n 0.0155911f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.41
cc_66 VPB N_B1_c_293_n 0.030195f $X=-0.19 $Y=1.305 $X2=3.86 $Y2=1.41
cc_67 VPB N_B1_c_295_n 0.00315868f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.16
cc_68 VPB N_B1_c_296_n 0.0329278f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.202
cc_69 VPB N_B1_c_297_n 0.00496449f $X=-0.19 $Y=1.305 $X2=1.287 $Y2=1.53
cc_70 VPB N_B1_c_298_n 0.00286634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_C1_c_408_n 0.015975f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_72 VPB N_C1_c_409_n 0.0160912f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_73 VPB N_C1_c_410_n 0.0158129f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=0.995
cc_74 VPB N_C1_c_411_n 0.0162318f $X=-0.19 $Y=1.305 $X2=3.86 $Y2=1.41
cc_75 VPB N_C1_c_412_n 0.00710388f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.202
cc_76 VPB N_C1_c_407_n 0.0478432f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_77 VPB N_VPWR_c_484_n 0.0107202f $X=-0.19 $Y=1.305 $X2=3.895 $Y2=0.995
cc_78 VPB N_VPWR_c_485_n 0.0379999f $X=-0.19 $Y=1.305 $X2=3.895 $Y2=0.56
cc_79 VPB N_VPWR_c_486_n 0.00468573f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.16
cc_80 VPB N_VPWR_c_487_n 0.0166095f $X=-0.19 $Y=1.305 $X2=3.7 $Y2=1.6
cc_81 VPB N_VPWR_c_488_n 0.0136265f $X=-0.19 $Y=1.305 $X2=3.865 $Y2=1.515
cc_82 VPB N_VPWR_c_489_n 0.0595126f $X=-0.19 $Y=1.305 $X2=3.855 $Y2=1.16
cc_83 VPB N_VPWR_c_490_n 0.0051645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_491_n 0.00537679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_492_n 0.0153463f $X=-0.19 $Y=1.305 $X2=0.955 $Y2=1.202
cc_86 VPB N_VPWR_c_493_n 0.00537832f $X=-0.19 $Y=1.305 $X2=1.345 $Y2=1.16
cc_87 VPB N_VPWR_c_494_n 0.013262f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.16
cc_88 VPB N_VPWR_c_495_n 0.0166052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_496_n 0.013126f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_497_n 0.026119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_498_n 0.00547308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_499_n 0.00553786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_483_n 0.0503528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_646_n 0.0260018f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.202
cc_95 VPB N_Y_c_645_n 0.00160692f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.202
cc_96 VPB Y 0.0105287f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.16
cc_97 VPB N_Y_c_649_n 0.0104015f $X=-0.19 $Y=1.305 $X2=1.287 $Y2=1.202
cc_98 N_A1_c_100_n N_A2_c_214_n 0.0238053f $X=1.485 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_99 N_A1_c_108_n N_A2_c_220_n 0.0350071f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A1_c_116_p N_A2_c_220_n 0.0131725f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_101 N_A1_c_112_n N_A2_c_220_n 0.0017846f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_c_116_p N_A2_c_221_n 0.0120284f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_103 N_A1_c_116_p N_A2_c_222_n 0.0120284f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_104 N_A1_c_101_n N_A2_c_223_n 0.0386994f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A1_c_116_p N_A2_c_223_n 0.0119833f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_106 N_A1_c_104_n N_A2_c_223_n 0.00231257f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_c_102_n N_A2_c_217_n 0.0259747f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A1_c_101_n N_A2_c_218_n 0.00164951f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_116_p N_A2_c_218_n 0.105751f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_110 N_A1_c_104_n N_A2_c_218_n 0.0226789f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A1_c_112_n N_A2_c_218_n 0.0142578f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_c_105_n N_A2_c_218_n 0.00116297f $X=1.46 $Y=1.202 $X2=0 $Y2=0
cc_113 N_A1_c_101_n N_A2_c_219_n 0.0253824f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A1_c_116_p N_A2_c_219_n 0.0205773f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_115 N_A1_c_104_n N_A2_c_219_n 0.00245023f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_c_112_n N_A2_c_219_n 0.00167732f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A1_c_105_n N_A2_c_219_n 0.0238053f $X=1.46 $Y=1.202 $X2=0 $Y2=0
cc_118 N_A1_c_102_n N_B1_c_290_n 0.0210315f $X=3.895 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A1_c_101_n N_B1_c_299_n 0.0328714f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A1_c_116_p N_B1_c_299_n 0.00205823f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_121 N_A1_c_104_n N_B1_c_299_n 0.00226989f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A1_c_101_n N_B1_c_296_n 0.024061f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A1_c_104_n N_B1_c_296_n 5.74505e-19 $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A1_c_101_n N_B1_c_297_n 0.00251603f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_104_n N_B1_c_297_n 0.035173f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A1_c_116_p N_B1_c_298_n 0.00528583f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_127 N_A1_c_112_n N_VPWR_M1014_s 0.00244652f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A1_c_116_p N_VPWR_M1024_s 0.00299168f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_129 N_A1_c_104_n N_VPWR_M1024_s 3.90316e-19 $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_130 N_A1_c_106_n N_VPWR_c_485_n 0.00586821f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_c_101_n N_VPWR_c_486_n 0.005745f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A1_c_108_n N_VPWR_c_489_n 0.00464324f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A1_c_101_n N_VPWR_c_489_n 0.00510168f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_106_n N_VPWR_c_495_n 0.00702461f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_107_n N_VPWR_c_495_n 0.0032362f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_106_n N_VPWR_c_498_n 0.00114359f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_107_n N_VPWR_c_498_n 0.0107306f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_108_n N_VPWR_c_498_n 0.00735595f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A1_c_106_n N_VPWR_c_483_n 0.013442f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A1_c_107_n N_VPWR_c_483_n 0.00388795f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A1_c_108_n N_VPWR_c_483_n 0.00532287f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_101_n N_VPWR_c_483_n 0.00691261f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A1_c_116_p N_A_118_297#_M1017_d 0.00613866f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_144 N_A1_c_116_p N_A_118_297#_M1021_s 0.00352397f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_145 N_A1_c_116_p N_A_118_297#_M1029_s 0.00817675f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_146 N_A1_c_104_n N_A_118_297#_M1029_s 3.80829e-19 $X=3.855 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A1_c_107_n N_A_118_297#_c_607_n 0.0126212f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A1_c_108_n N_A_118_297#_c_607_n 0.0120623f $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A1_c_103_n N_A_118_297#_c_607_n 0.00419569f $X=1.015 $Y=1.202 $X2=0
+ $Y2=0
cc_150 N_A1_c_116_p N_A_118_297#_c_607_n 0.010665f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_151 N_A1_c_112_n N_A_118_297#_c_607_n 0.0242314f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A1_c_105_n N_A_118_297#_c_607_n 9.19106e-19 $X=1.46 $Y=1.202 $X2=0
+ $Y2=0
cc_153 N_A1_c_101_n N_A_118_297#_c_613_n 0.002515f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A1_c_116_p N_A_118_297#_c_613_n 0.00277337f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_155 N_A1_c_103_n N_A_118_297#_c_615_n 0.00703433f $X=1.015 $Y=1.202 $X2=0
+ $Y2=0
cc_156 N_A1_c_105_n N_A_118_297#_c_615_n 0.00111457f $X=1.46 $Y=1.202 $X2=0
+ $Y2=0
cc_157 N_A1_c_116_p N_Y_M1002_d 0.00352397f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_158 N_A1_c_116_p N_Y_M1027_d 0.00352397f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_159 N_A1_c_108_n N_Y_c_652_n 4.63455e-19 $X=1.46 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A1_c_116_p N_Y_c_652_n 0.0974125f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_161 N_A1_c_101_n N_Y_c_654_n 0.00747676f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A1_c_116_p N_Y_c_654_n 0.016669f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_163 N_A1_c_101_n N_Y_c_656_n 0.0104857f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_c_98_n N_A_27_47#_c_760_n 0.0132853f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_99_n N_A_27_47#_c_760_n 0.0131977f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_103_n N_A_27_47#_c_760_n 0.0460086f $X=1.015 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A1_c_112_n N_A_27_47#_c_760_n 0.00881237f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A1_c_105_n N_A_27_47#_c_760_n 0.00386608f $X=1.46 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A1_c_101_n N_A_27_47#_c_772_n 0.00288519f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_102_n N_A_27_47#_c_772_n 0.0110591f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_104_n N_A_27_47#_c_772_n 0.0170843f $X=3.855 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A1_c_99_n N_A_27_47#_c_761_n 0.00340518f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_100_n N_A_27_47#_c_761_n 0.0157917f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A1_c_102_n N_A_27_47#_c_761_n 6.5376e-19 $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A1_c_116_p N_A_27_47#_c_761_n 0.00753594f $X=3.7 $Y=1.6 $X2=0 $Y2=0
cc_176 N_A1_c_112_n N_A_27_47#_c_761_n 0.0345931f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A1_c_105_n N_A_27_47#_c_761_n 0.00494155f $X=1.46 $Y=1.202 $X2=0 $Y2=0
cc_178 N_A1_c_102_n N_A_27_47#_c_781_n 3.29317e-19 $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A1_c_100_n N_A_27_47#_c_764_n 0.00272001f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_102_n N_A_27_47#_c_764_n 0.00352307f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A1_c_99_n N_A_27_47#_c_784_n 0.00419048f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A1_c_100_n N_A_27_47#_c_784_n 8.07403e-19 $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A1_c_112_n N_A_27_47#_c_784_n 0.00117031f $X=1.345 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A1_c_99_n N_VGND_c_888_n 0.00353009f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A1_c_100_n N_VGND_c_888_n 0.00352186f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A1_c_99_n N_VGND_c_889_n 0.00101018f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_100_n N_VGND_c_889_n 0.00789494f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_98_n N_VGND_c_891_n 0.00353009f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_102_n N_VGND_c_893_n 0.0042361f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A1_c_98_n N_VGND_c_894_n 0.00510538f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A1_c_99_n N_VGND_c_894_n 0.00438375f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_100_n N_VGND_c_894_n 0.00366404f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A1_c_102_n N_VGND_c_894_n 0.00516079f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A1_c_98_n N_VGND_c_895_n 0.0144723f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A1_c_99_n N_VGND_c_895_n 0.00828763f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A1_c_100_n N_VGND_c_895_n 0.0010058f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A1_c_102_n N_VGND_c_898_n 0.00420474f $X=3.895 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_220_n N_VPWR_c_489_n 0.00429453f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A2_c_221_n N_VPWR_c_489_n 0.00429453f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A2_c_222_n N_VPWR_c_489_n 0.00429453f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A2_c_223_n N_VPWR_c_489_n 0.00429453f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A2_c_220_n N_VPWR_c_498_n 0.00112655f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_220_n N_VPWR_c_483_n 0.00618304f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_c_221_n N_VPWR_c_483_n 0.00611674f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A2_c_222_n N_VPWR_c_483_n 0.00611674f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_223_n N_VPWR_c_483_n 0.00614026f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_220_n N_A_118_297#_c_607_n 7.99602e-19 $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_220_n N_A_118_297#_c_613_n 0.01205f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_221_n N_A_118_297#_c_613_n 0.00955231f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_222_n N_A_118_297#_c_613_n 0.00955231f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_223_n N_A_118_297#_c_613_n 0.00955231f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A2_c_220_n N_Y_c_652_n 0.00638895f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A2_c_221_n N_Y_c_652_n 0.0122704f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A2_c_222_n N_Y_c_652_n 0.0122704f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A2_c_223_n N_Y_c_652_n 0.0122038f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A2_c_214_n N_A_27_47#_c_761_n 0.0126072f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A2_c_215_n N_A_27_47#_c_761_n 0.0129944f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_c_216_n N_A_27_47#_c_761_n 0.0130229f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A2_c_217_n N_A_27_47#_c_761_n 0.011746f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A2_c_218_n N_A_27_47#_c_761_n 0.119169f $X=3.19 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_c_219_n N_A_27_47#_c_761_n 0.0128516f $X=3.38 $Y=1.202 $X2=0 $Y2=0
cc_222 N_A2_c_214_n N_A_27_47#_c_764_n 0.00307664f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A2_c_215_n N_A_27_47#_c_764_n 0.00315083f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_224 N_A2_c_216_n N_A_27_47#_c_764_n 0.00321611f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A2_c_217_n N_A_27_47#_c_764_n 0.00275293f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A2_c_214_n N_VGND_c_889_n 0.00796693f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A2_c_215_n N_VGND_c_889_n 0.00113111f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A2_c_216_n N_VGND_c_890_n 0.00352884f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A2_c_217_n N_VGND_c_890_n 0.00211731f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A2_c_214_n N_VGND_c_892_n 0.00352186f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A2_c_215_n N_VGND_c_892_n 0.00352884f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_214_n N_VGND_c_894_n 0.00354654f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_215_n N_VGND_c_894_n 0.00354658f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_216_n N_VGND_c_894_n 0.00366408f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_217_n N_VGND_c_894_n 0.00259142f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A2_c_214_n N_VGND_c_897_n 0.00106158f $X=1.915 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_215_n N_VGND_c_897_n 0.00802029f $X=2.395 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_216_n N_VGND_c_897_n 0.00807014f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A2_c_217_n N_VGND_c_897_n 0.00103793f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_216_n N_VGND_c_898_n 0.00115166f $X=2.875 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_217_n N_VGND_c_898_n 0.0102967f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B1_c_292_n N_C1_c_403_n 0.0317774f $X=5.365 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_243 N_B1_c_301_n N_C1_c_408_n 0.0363576f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B1_c_318_p N_C1_c_408_n 0.0173644f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_245 N_B1_c_298_n N_C1_c_408_n 0.00282927f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_246 N_B1_c_318_p N_C1_c_409_n 0.01191f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_247 N_B1_c_318_p N_C1_c_410_n 0.01191f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_248 N_B1_c_293_n N_C1_c_411_n 0.0373375f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B1_c_318_p N_C1_c_411_n 0.017059f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_250 N_B1_c_295_n N_C1_c_411_n 0.00153214f $X=7.665 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B1_c_294_n N_C1_c_406_n 0.0280119f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_293_n N_C1_c_412_n 6.9292e-19 $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B1_c_318_p N_C1_c_412_n 0.076816f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_254 N_B1_c_295_n N_C1_c_412_n 0.00967173f $X=7.665 $Y=1.16 $X2=0 $Y2=0
cc_255 N_B1_c_298_n N_C1_c_412_n 0.011651f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_256 N_B1_c_293_n N_C1_c_407_n 0.0263368f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B1_c_318_p N_C1_c_407_n 0.00604008f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_258 N_B1_c_295_n N_C1_c_407_n 0.00301923f $X=7.665 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B1_c_296_n N_C1_c_407_n 0.0317774f $X=5.34 $Y=1.202 $X2=0 $Y2=0
cc_260 N_B1_c_298_n N_C1_c_407_n 0.00710365f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_261 N_B1_c_298_n N_VPWR_M1009_s 0.00206918f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_262 N_B1_c_318_p N_VPWR_M1001_d 0.00340201f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_263 N_B1_c_318_p N_VPWR_M1023_d 0.0033587f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_264 N_B1_c_299_n N_VPWR_c_486_n 0.0017535f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B1_c_293_n N_VPWR_c_488_n 0.00892439f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B1_c_299_n N_VPWR_c_491_n 0.00113168f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B1_c_300_n N_VPWR_c_491_n 0.01063f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B1_c_301_n N_VPWR_c_491_n 0.00762757f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B1_c_299_n N_VPWR_c_492_n 0.0052046f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B1_c_300_n N_VPWR_c_492_n 0.0032362f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B1_c_301_n N_VPWR_c_493_n 0.00112575f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_301_n N_VPWR_c_494_n 0.00464324f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_293_n N_VPWR_c_497_n 0.00506535f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_293_n N_VPWR_c_499_n 0.00194382f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B1_c_299_n N_VPWR_c_483_n 0.00690188f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_300_n N_VPWR_c_483_n 0.00388795f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_301_n N_VPWR_c_483_n 0.00529826f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B1_c_293_n N_VPWR_c_483_n 0.00814165f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B1_c_298_n N_Y_M1006_d 0.00315346f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_280 N_B1_c_318_p N_Y_M1012_d 0.0066872f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_281 N_B1_c_298_n N_Y_M1012_d 8.41019e-19 $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_282 N_B1_c_318_p N_Y_M1019_s 0.0033587f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_283 N_B1_c_318_p N_Y_M1031_s 0.0082477f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_284 N_B1_c_294_n N_Y_c_666_n 0.00218558f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B1_c_294_n N_Y_c_667_n 0.00337628f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_286 N_B1_c_293_n N_Y_c_668_n 0.0026207f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B1_c_294_n N_Y_c_668_n 0.0139653f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B1_c_295_n N_Y_c_668_n 0.0139672f $X=7.665 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B1_c_299_n N_Y_c_654_n 2.52786e-19 $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_290 N_B1_c_293_n N_Y_c_646_n 0.00200441f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B1_c_293_n N_Y_c_645_n 6.23164e-19 $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B1_c_294_n N_Y_c_645_n 0.0138429f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B1_c_295_n N_Y_c_645_n 0.0370345f $X=7.665 $Y=1.16 $X2=0 $Y2=0
cc_294 N_B1_c_293_n Y 0.00655601f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_295 N_B1_c_300_n N_Y_c_649_n 0.0132286f $X=4.86 $Y=1.41 $X2=0 $Y2=0
cc_296 N_B1_c_301_n N_Y_c_649_n 0.0136581f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_297 N_B1_c_293_n N_Y_c_649_n 0.0176f $X=7.69 $Y=1.41 $X2=0 $Y2=0
cc_298 N_B1_c_318_p N_Y_c_649_n 0.0140665f $X=7.58 $Y=1.6 $X2=0 $Y2=0
cc_299 N_B1_c_296_n N_Y_c_649_n 0.00199669f $X=5.34 $Y=1.202 $X2=0 $Y2=0
cc_300 N_B1_c_298_n N_Y_c_649_n 0.159976f $X=5.525 $Y=1.34 $X2=0 $Y2=0
cc_301 N_B1_c_299_n N_Y_c_656_n 0.0136821f $X=4.38 $Y=1.41 $X2=0 $Y2=0
cc_302 N_B1_c_297_n N_Y_c_656_n 0.0172505f $X=4.71 $Y=1.34 $X2=0 $Y2=0
cc_303 N_B1_c_297_n N_A_27_47#_c_772_n 0.00205362f $X=4.71 $Y=1.34 $X2=0 $Y2=0
cc_304 N_B1_c_290_n N_A_27_47#_c_798_n 0.00972566f $X=4.355 $Y=0.995 $X2=0 $Y2=0
cc_305 N_B1_c_291_n N_A_27_47#_c_798_n 0.00796047f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_306 N_B1_c_292_n N_A_27_47#_c_798_n 0.0059805f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_307 N_B1_c_297_n N_A_27_47#_c_798_n 0.00251253f $X=4.71 $Y=1.34 $X2=0 $Y2=0
cc_308 N_B1_c_294_n N_A_27_47#_c_762_n 0.00514577f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_309 N_B1_c_290_n N_A_27_47#_c_764_n 0.00235806f $X=4.355 $Y=0.995 $X2=0 $Y2=0
cc_310 N_B1_c_291_n N_A_27_47#_c_764_n 0.0021112f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_311 N_B1_c_292_n N_A_27_47#_c_764_n 0.00232103f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_312 N_B1_c_294_n N_A_27_47#_c_764_n 0.00256483f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_313 N_B1_c_297_n N_A_27_47#_c_764_n 0.00602013f $X=4.71 $Y=1.34 $X2=0 $Y2=0
cc_314 N_B1_c_294_n N_A_27_47#_c_765_n 8.38249e-19 $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B1_c_294_n N_A_27_47#_c_766_n 9.94574e-19 $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B1_c_290_n N_VGND_c_893_n 0.00357877f $X=4.355 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_291_n N_VGND_c_893_n 0.00357877f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_292_n N_VGND_c_893_n 0.00357877f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_319 N_B1_c_294_n N_VGND_c_893_n 0.00380901f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_320 N_B1_c_290_n N_VGND_c_894_n 0.00504961f $X=4.355 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B1_c_291_n N_VGND_c_894_n 0.00515079f $X=4.835 $Y=0.995 $X2=0 $Y2=0
cc_322 N_B1_c_292_n N_VGND_c_894_n 0.0050223f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B1_c_294_n N_VGND_c_894_n 0.00640034f $X=7.775 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B1_c_290_n N_A_886_47#_c_1007_n 0.00265506f $X=4.355 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_B1_c_291_n N_A_886_47#_c_1007_n 0.00929367f $X=4.835 $Y=0.995 $X2=0
+ $Y2=0
cc_326 N_B1_c_292_n N_A_886_47#_c_1007_n 0.011351f $X=5.365 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B1_c_296_n N_A_886_47#_c_1007_n 0.00780733f $X=5.34 $Y=1.202 $X2=0
+ $Y2=0
cc_328 N_B1_c_297_n N_A_886_47#_c_1007_n 0.0680068f $X=4.71 $Y=1.34 $X2=0 $Y2=0
cc_329 N_C1_c_408_n N_VPWR_c_491_n 9.99588e-19 $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_330 N_C1_c_408_n N_VPWR_c_493_n 0.0106707f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_331 N_C1_c_409_n N_VPWR_c_493_n 0.00783855f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_332 N_C1_c_410_n N_VPWR_c_493_n 0.00100747f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_333 N_C1_c_408_n N_VPWR_c_494_n 0.00309549f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_334 N_C1_c_409_n N_VPWR_c_496_n 0.00450253f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_335 N_C1_c_410_n N_VPWR_c_496_n 0.00309549f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_336 N_C1_c_411_n N_VPWR_c_497_n 0.00436183f $X=7.22 $Y=1.41 $X2=0 $Y2=0
cc_337 N_C1_c_409_n N_VPWR_c_499_n 0.00112282f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_338 N_C1_c_410_n N_VPWR_c_499_n 0.010644f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_339 N_C1_c_411_n N_VPWR_c_499_n 0.00928909f $X=7.22 $Y=1.41 $X2=0 $Y2=0
cc_340 N_C1_c_408_n N_VPWR_c_483_n 0.00374672f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_341 N_C1_c_409_n N_VPWR_c_483_n 0.00513103f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_342 N_C1_c_410_n N_VPWR_c_483_n 0.00372054f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_343 N_C1_c_411_n N_VPWR_c_483_n 0.00501617f $X=7.22 $Y=1.41 $X2=0 $Y2=0
cc_344 N_C1_c_403_n N_Y_c_666_n 0.00307758f $X=5.785 $Y=0.995 $X2=0 $Y2=0
cc_345 N_C1_c_404_n N_Y_c_666_n 0.00748475f $X=6.255 $Y=0.995 $X2=0 $Y2=0
cc_346 N_C1_c_405_n N_Y_c_666_n 0.00748475f $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_347 N_C1_c_406_n N_Y_c_666_n 0.0078804f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_348 N_C1_c_412_n N_Y_c_666_n 0.00345838f $X=6.975 $Y=1.16 $X2=0 $Y2=0
cc_349 N_C1_c_407_n N_Y_c_666_n 0.00300671f $X=7.22 $Y=1.202 $X2=0 $Y2=0
cc_350 N_C1_c_405_n N_Y_c_667_n 0.00102729f $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_351 N_C1_c_406_n N_Y_c_667_n 0.00657128f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_352 N_C1_c_405_n N_Y_c_693_n 2.14776e-19 $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_353 N_C1_c_406_n N_Y_c_693_n 0.00831067f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_354 N_C1_c_408_n N_Y_c_649_n 0.0130983f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_355 N_C1_c_409_n N_Y_c_649_n 0.0135278f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_356 N_C1_c_410_n N_Y_c_649_n 0.0130983f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_357 N_C1_c_411_n N_Y_c_649_n 0.0134848f $X=7.22 $Y=1.41 $X2=0 $Y2=0
cc_358 N_C1_c_403_n N_A_27_47#_c_798_n 6.02163e-19 $X=5.785 $Y=0.995 $X2=0 $Y2=0
cc_359 N_C1_c_403_n N_A_27_47#_c_764_n 0.00336823f $X=5.785 $Y=0.995 $X2=0 $Y2=0
cc_360 N_C1_c_404_n N_A_27_47#_c_764_n 0.0021087f $X=6.255 $Y=0.995 $X2=0 $Y2=0
cc_361 N_C1_c_405_n N_A_27_47#_c_764_n 0.00212645f $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_362 N_C1_c_406_n N_A_27_47#_c_764_n 0.00410005f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_363 N_C1_c_412_n N_A_27_47#_c_764_n 0.00760746f $X=6.975 $Y=1.16 $X2=0 $Y2=0
cc_364 N_C1_c_407_n N_A_27_47#_c_764_n 0.00397112f $X=7.22 $Y=1.202 $X2=0 $Y2=0
cc_365 N_C1_c_403_n N_VGND_c_893_n 0.00412276f $X=5.785 $Y=0.995 $X2=0 $Y2=0
cc_366 N_C1_c_404_n N_VGND_c_893_n 0.00361001f $X=6.255 $Y=0.995 $X2=0 $Y2=0
cc_367 N_C1_c_405_n N_VGND_c_893_n 0.00361001f $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_368 N_C1_c_406_n N_VGND_c_893_n 0.00360925f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_369 N_C1_c_403_n N_VGND_c_894_n 0.00507704f $X=5.785 $Y=0.995 $X2=0 $Y2=0
cc_370 N_C1_c_404_n N_VGND_c_894_n 0.00499047f $X=6.255 $Y=0.995 $X2=0 $Y2=0
cc_371 N_C1_c_405_n N_VGND_c_894_n 0.00510581f $X=6.725 $Y=0.995 $X2=0 $Y2=0
cc_372 N_C1_c_406_n N_VGND_c_894_n 0.00525824f $X=7.245 $Y=0.995 $X2=0 $Y2=0
cc_373 N_C1_c_403_n N_A_886_47#_c_1007_n 0.0164769f $X=5.785 $Y=0.995 $X2=0
+ $Y2=0
cc_374 N_C1_c_404_n N_A_886_47#_c_1007_n 0.00945706f $X=6.255 $Y=0.995 $X2=0
+ $Y2=0
cc_375 N_C1_c_405_n N_A_886_47#_c_1007_n 0.00835265f $X=6.725 $Y=0.995 $X2=0
+ $Y2=0
cc_376 N_C1_c_406_n N_A_886_47#_c_1007_n 0.00150053f $X=7.245 $Y=0.995 $X2=0
+ $Y2=0
cc_377 N_C1_c_412_n N_A_886_47#_c_1007_n 0.0363925f $X=6.975 $Y=1.16 $X2=0 $Y2=0
cc_378 N_C1_c_407_n N_A_886_47#_c_1007_n 0.00678446f $X=7.22 $Y=1.202 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_483_n N_A_118_297#_M1011_d 0.00365219f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_380 N_VPWR_c_483_n N_A_118_297#_M1017_d 0.00259393f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_483_n N_A_118_297#_M1021_s 0.00239319f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_483_n N_A_118_297#_M1029_s 0.00239319f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_M1014_s N_A_118_297#_c_607_n 0.00402698f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_384 N_VPWR_c_489_n N_A_118_297#_c_607_n 0.0033904f $X=4.015 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_495_n N_A_118_297#_c_607_n 0.00269991f $X=1.005 $Y=2.72 $X2=0
+ $Y2=0
cc_386 N_VPWR_c_498_n N_A_118_297#_c_607_n 0.019553f $X=1.22 $Y=2.36 $X2=0 $Y2=0
cc_387 N_VPWR_c_483_n N_A_118_297#_c_607_n 0.011867f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_c_489_n N_A_118_297#_c_631_n 0.012363f $X=4.015 $Y=2.72 $X2=0
+ $Y2=0
cc_389 N_VPWR_c_483_n N_A_118_297#_c_631_n 0.00687765f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_390 N_VPWR_c_486_n N_A_118_297#_c_613_n 0.0120827f $X=4.12 $Y=2.36 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_489_n N_A_118_297#_c_613_n 0.111532f $X=4.015 $Y=2.72 $X2=0
+ $Y2=0
cc_392 N_VPWR_c_483_n N_A_118_297#_c_613_n 0.0710383f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_495_n N_A_118_297#_c_615_n 0.00469289f $X=1.005 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_VPWR_c_483_n N_A_118_297#_c_615_n 0.00686953f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_395 N_VPWR_c_483_n N_Y_M1002_d 0.00240926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_396 N_VPWR_c_483_n N_Y_M1027_d 0.00240926f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_483_n N_Y_M1006_d 0.00344662f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_483_n N_Y_M1012_d 0.00330361f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_483_n N_Y_M1019_s 0.00330361f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_483_n N_Y_M1031_s 0.00330361f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_483_n N_Y_c_652_n 0.00455889f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_489_n N_Y_c_654_n 6.14891e-19 $X=4.015 $Y=2.72 $X2=0 $Y2=0
cc_403 N_VPWR_M1025_s N_Y_c_646_n 0.00374076f $X=7.78 $Y=1.485 $X2=0 $Y2=0
cc_404 N_VPWR_M1025_s Y 0.0116145f $X=7.78 $Y=1.485 $X2=0 $Y2=0
cc_405 N_VPWR_M1009_s N_Y_c_649_n 0.00371648f $X=4.95 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_M1001_d N_Y_c_649_n 0.00351667f $X=5.9 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_M1023_d N_Y_c_649_n 0.00351667f $X=6.84 $Y=1.485 $X2=0 $Y2=0
cc_408 N_VPWR_M1025_s N_Y_c_649_n 0.0224909f $X=7.78 $Y=1.485 $X2=0 $Y2=0
cc_409 N_VPWR_c_488_n N_Y_c_649_n 0.0252336f $X=8.32 $Y=2.36 $X2=0 $Y2=0
cc_410 N_VPWR_c_491_n N_Y_c_649_n 0.0200578f $X=5.1 $Y=2.36 $X2=0 $Y2=0
cc_411 N_VPWR_c_492_n N_Y_c_649_n 0.00642399f $X=4.885 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_493_n N_Y_c_649_n 0.0200084f $X=6.045 $Y=2.36 $X2=0 $Y2=0
cc_413 N_VPWR_c_494_n N_Y_c_649_n 0.00929776f $X=5.83 $Y=2.72 $X2=0 $Y2=0
cc_414 N_VPWR_c_496_n N_Y_c_649_n 0.00920992f $X=6.77 $Y=2.72 $X2=0 $Y2=0
cc_415 N_VPWR_c_497_n N_Y_c_649_n 0.0169011f $X=8.155 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_499_n N_Y_c_649_n 0.0203724f $X=6.985 $Y=2.36 $X2=0 $Y2=0
cc_417 N_VPWR_c_483_n N_Y_c_649_n 0.0755095f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_418 N_VPWR_M1024_s N_Y_c_656_n 0.00875315f $X=3.95 $Y=1.485 $X2=0 $Y2=0
cc_419 N_VPWR_c_486_n N_Y_c_656_n 0.0168509f $X=4.12 $Y=2.36 $X2=0 $Y2=0
cc_420 N_VPWR_c_489_n N_Y_c_656_n 0.00244379f $X=4.015 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_c_492_n N_Y_c_656_n 0.00280903f $X=4.885 $Y=2.72 $X2=0 $Y2=0
cc_422 N_VPWR_c_483_n N_Y_c_656_n 0.0104153f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_423 N_A_118_297#_c_613_n N_Y_M1002_d 0.00374179f $X=3.62 $Y=2.36 $X2=0.475
+ $Y2=0.56
cc_424 N_A_118_297#_c_613_n N_Y_M1027_d 0.00374179f $X=3.62 $Y=2.36 $X2=0.5
+ $Y2=1.41
cc_425 N_A_118_297#_M1021_s N_Y_c_652_n 0.00369302f $X=2.51 $Y=1.485 $X2=1.015
+ $Y2=1.202
cc_426 N_A_118_297#_M1029_s N_Y_c_652_n 0.00345095f $X=3.47 $Y=1.485 $X2=1.015
+ $Y2=1.202
cc_427 N_A_118_297#_c_607_n N_Y_c_652_n 0.0147711f $X=1.605 $Y=2.02 $X2=1.015
+ $Y2=1.202
cc_428 N_A_118_297#_c_613_n N_Y_c_652_n 0.0945885f $X=3.62 $Y=2.36 $X2=1.015
+ $Y2=1.202
cc_429 N_A_118_297#_M1029_s N_Y_c_654_n 3.50153e-19 $X=3.47 $Y=1.485 $X2=1.345
+ $Y2=1.16
cc_430 N_Y_c_668_n N_A_27_47#_M1018_d 0.0141187f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_431 N_Y_c_645_n N_A_27_47#_M1018_d 0.0033607f $X=8.23 $Y=1.34 $X2=0 $Y2=0
cc_432 N_Y_c_666_n N_A_27_47#_c_798_n 0.004097f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_433 N_Y_c_666_n N_A_27_47#_c_762_n 0.00887123f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_434 N_Y_c_667_n N_A_27_47#_c_762_n 0.00130172f $X=7.375 $Y=0.655 $X2=0 $Y2=0
cc_435 N_Y_c_668_n N_A_27_47#_c_762_n 0.0244243f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_436 N_Y_M1005_s N_A_27_47#_c_764_n 0.00231205f $X=5.86 $Y=0.235 $X2=0 $Y2=0
cc_437 N_Y_M1028_s N_A_27_47#_c_764_n 0.00499996f $X=6.8 $Y=0.235 $X2=0 $Y2=0
cc_438 N_Y_c_666_n N_A_27_47#_c_764_n 0.0329018f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_439 N_Y_c_667_n N_A_27_47#_c_764_n 0.0201476f $X=7.375 $Y=0.655 $X2=0 $Y2=0
cc_440 N_Y_c_668_n N_A_27_47#_c_764_n 0.0200613f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_441 N_Y_c_666_n N_VGND_c_893_n 0.085761f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_442 N_Y_c_668_n N_VGND_c_893_n 0.00326381f $X=7.98 $Y=0.74 $X2=0 $Y2=0
cc_443 N_Y_M1005_s N_VGND_c_894_n 0.00144449f $X=5.86 $Y=0.235 $X2=0 $Y2=0
cc_444 N_Y_M1028_s N_VGND_c_894_n 0.00167161f $X=6.8 $Y=0.235 $X2=0 $Y2=0
cc_445 N_Y_c_666_n N_VGND_c_894_n 0.0155663f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_446 N_Y_c_666_n N_A_886_47#_M1004_d 0.00306559f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_447 N_Y_M1005_s N_A_886_47#_c_1007_n 0.00513447f $X=5.86 $Y=0.235 $X2=0 $Y2=0
cc_448 N_Y_M1028_s N_A_886_47#_c_1007_n 0.00262923f $X=6.8 $Y=0.235 $X2=0 $Y2=0
cc_449 N_Y_c_666_n N_A_886_47#_c_1007_n 0.0466828f $X=7.265 $Y=0.36 $X2=0 $Y2=0
cc_450 N_Y_c_667_n N_A_886_47#_c_1007_n 7.79711e-19 $X=7.375 $Y=0.655 $X2=0
+ $Y2=0
cc_451 N_Y_c_693_n N_A_886_47#_c_1007_n 0.00722787f $X=7.485 $Y=0.74 $X2=0 $Y2=0
cc_452 N_Y_c_666_n A_1464_47# 0.00305272f $X=7.265 $Y=0.36 $X2=-0.19 $Y2=-0.24
cc_453 N_Y_c_667_n A_1464_47# 0.0028236f $X=7.375 $Y=0.655 $X2=-0.19 $Y2=-0.24
cc_454 N_Y_c_668_n A_1464_47# 0.00541918f $X=7.98 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_455 N_Y_c_693_n A_1464_47# 0.00475485f $X=7.485 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_456 N_A_27_47#_c_760_n N_VGND_M1007_d 0.0022909f $X=1.125 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_457 N_A_27_47#_c_761_n N_VGND_M1016_d 0.00158f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_764_n N_VGND_M1016_d 0.00201451f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_459 N_A_27_47#_c_761_n N_VGND_M1003_s 0.00210124f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_764_n N_VGND_M1003_s 0.00237425f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_772_n N_VGND_M1030_s 0.00869456f $X=4.005 $Y=0.71 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_764_n N_VGND_M1030_s 0.0026406f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_463 N_A_27_47#_c_760_n N_VGND_c_888_n 0.00338958f $X=1.125 $Y=0.765 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_761_n N_VGND_c_888_n 0.0104158f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_465 N_A_27_47#_c_764_n N_VGND_c_888_n 3.74208e-19 $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_466 N_A_27_47#_c_784_n N_VGND_c_888_n 8.52016e-19 $X=1.4 $Y=0.51 $X2=0 $Y2=0
cc_467 N_A_27_47#_c_761_n N_VGND_c_889_n 0.0178786f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_468 N_A_27_47#_c_764_n N_VGND_c_889_n 0.00817983f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_469 N_A_27_47#_c_784_n N_VGND_c_889_n 0.0015315f $X=1.4 $Y=0.51 $X2=0 $Y2=0
cc_470 N_A_27_47#_c_761_n N_VGND_c_890_n 0.00858711f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_471 N_A_27_47#_c_764_n N_VGND_c_890_n 0.00177014f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_472 N_A_27_47#_c_760_n N_VGND_c_891_n 0.0026054f $X=1.125 $Y=0.765 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_763_n N_VGND_c_891_n 0.00453599f $X=0.355 $Y=0.72 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_761_n N_VGND_c_892_n 0.00853161f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_475 N_A_27_47#_c_764_n N_VGND_c_892_n 0.00174721f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_772_n N_VGND_c_893_n 0.00295179f $X=4.005 $Y=0.71 $X2=0
+ $Y2=0
cc_477 N_A_27_47#_c_781_n N_VGND_c_893_n 0.0147597f $X=4.235 $Y=0.355 $X2=0
+ $Y2=0
cc_478 N_A_27_47#_c_798_n N_VGND_c_893_n 0.0695034f $X=5.1 $Y=0.365 $X2=0 $Y2=0
cc_479 N_A_27_47#_c_762_n N_VGND_c_893_n 0.0264198f $X=8.32 $Y=0.395 $X2=0 $Y2=0
cc_480 N_A_27_47#_c_764_n N_VGND_c_893_n 0.00510596f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_481 N_A_27_47#_c_765_n N_VGND_c_893_n 5.08791e-19 $X=8.405 $Y=0.51 $X2=0
+ $Y2=0
cc_482 N_A_27_47#_c_766_n N_VGND_c_893_n 0.00838914f $X=8.405 $Y=0.395 $X2=0
+ $Y2=0
cc_483 N_A_27_47#_M1007_s N_VGND_c_894_n 0.00344766f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_27_47#_M1015_s N_VGND_c_894_n 0.00237391f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_485 N_A_27_47#_M1000_d N_VGND_c_894_n 0.00194336f $X=1.99 $Y=0.235 $X2=0
+ $Y2=0
cc_486 N_A_27_47#_M1026_d N_VGND_c_894_n 0.0022674f $X=2.95 $Y=0.235 $X2=0 $Y2=0
cc_487 N_A_27_47#_M1022_s N_VGND_c_894_n 0.00145272f $X=3.97 $Y=0.235 $X2=0
+ $Y2=0
cc_488 N_A_27_47#_M1013_d N_VGND_c_894_n 0.00171342f $X=4.91 $Y=0.235 $X2=0
+ $Y2=0
cc_489 N_A_27_47#_M1018_d N_VGND_c_894_n 0.00184732f $X=7.85 $Y=0.235 $X2=0
+ $Y2=0
cc_490 N_A_27_47#_c_760_n N_VGND_c_894_n 0.0115485f $X=1.125 $Y=0.765 $X2=0
+ $Y2=0
cc_491 N_A_27_47#_c_761_n N_VGND_c_894_n 0.00107448f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_492 N_A_27_47#_c_781_n N_VGND_c_894_n 0.00244609f $X=4.235 $Y=0.355 $X2=0
+ $Y2=0
cc_493 N_A_27_47#_c_798_n N_VGND_c_894_n 0.011443f $X=5.1 $Y=0.365 $X2=0 $Y2=0
cc_494 N_A_27_47#_c_762_n N_VGND_c_894_n 0.00543455f $X=8.32 $Y=0.395 $X2=0
+ $Y2=0
cc_495 N_A_27_47#_c_763_n N_VGND_c_894_n 0.00630153f $X=0.355 $Y=0.72 $X2=0
+ $Y2=0
cc_496 N_A_27_47#_c_764_n N_VGND_c_894_n 0.581415f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_497 N_A_27_47#_c_784_n N_VGND_c_894_n 0.0298383f $X=1.4 $Y=0.51 $X2=0 $Y2=0
cc_498 N_A_27_47#_c_765_n N_VGND_c_894_n 0.0288358f $X=8.405 $Y=0.51 $X2=0 $Y2=0
cc_499 N_A_27_47#_c_766_n N_VGND_c_894_n 0.00152175f $X=8.405 $Y=0.395 $X2=0
+ $Y2=0
cc_500 N_A_27_47#_c_760_n N_VGND_c_895_n 0.0193953f $X=1.125 $Y=0.765 $X2=0
+ $Y2=0
cc_501 N_A_27_47#_c_761_n N_VGND_c_895_n 9.97233e-19 $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_502 N_A_27_47#_c_784_n N_VGND_c_895_n 0.00158555f $X=1.4 $Y=0.51 $X2=0 $Y2=0
cc_503 N_A_27_47#_c_761_n N_VGND_c_897_n 0.018283f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_504 N_A_27_47#_c_764_n N_VGND_c_897_n 0.00883914f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_505 N_A_27_47#_c_772_n N_VGND_c_898_n 0.0149026f $X=4.005 $Y=0.71 $X2=0 $Y2=0
cc_506 N_A_27_47#_c_761_n N_VGND_c_898_n 0.00429609f $X=3.48 $Y=0.71 $X2=0 $Y2=0
cc_507 N_A_27_47#_c_764_n N_VGND_c_898_n 0.00881372f $X=8.26 $Y=0.51 $X2=0 $Y2=0
cc_508 N_A_27_47#_c_798_n N_A_886_47#_M1008_s 0.0031236f $X=5.1 $Y=0.365
+ $X2=-0.19 $Y2=-0.24
cc_509 N_A_27_47#_c_764_n N_A_886_47#_M1008_s 0.00236985f $X=8.26 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_510 N_A_27_47#_c_764_n N_A_886_47#_M1004_d 0.0022976f $X=8.26 $Y=0.51 $X2=0
+ $Y2=0
cc_511 N_A_27_47#_M1013_d N_A_886_47#_c_1007_n 0.00520425f $X=4.91 $Y=0.235
+ $X2=0 $Y2=0
cc_512 N_A_27_47#_c_798_n N_A_886_47#_c_1007_n 0.0508149f $X=5.1 $Y=0.365 $X2=0
+ $Y2=0
cc_513 N_A_27_47#_c_764_n N_A_886_47#_c_1007_n 0.0701774f $X=8.26 $Y=0.51 $X2=0
+ $Y2=0
cc_514 N_A_27_47#_c_764_n A_1088_47# 0.00331135f $X=8.26 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_515 N_A_27_47#_c_764_n A_1464_47# 0.00279275f $X=8.26 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_516 N_VGND_c_894_n N_A_886_47#_M1008_s 0.00149584f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_517 N_VGND_c_894_n N_A_886_47#_M1004_d 0.00145358f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_893_n N_A_886_47#_c_1007_n 0.00500307f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_519 N_VGND_c_894_n A_1088_47# 0.00156226f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_520 N_VGND_c_894_n A_1464_47# 0.00204794f $X=8.51 $Y=0 $X2=-0.19 $Y2=-0.24
cc_521 N_A_886_47#_c_1007_n A_1088_47# 0.00762341f $X=6.515 $Y=0.725 $X2=0.475
+ $Y2=0.995
