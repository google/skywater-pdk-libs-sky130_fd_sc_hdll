* File: sky130_fd_sc_hdll__mux2_12.spice
* Created: Wed Sep  2 08:34:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2_12.pex.spice"
.subckt sky130_fd_sc_hdll__mux2_12  VNB VPB A1 S A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* S	S
* A1	A1
* VPB	VPB
* VNB	VNB
MM1016 N_A_27_47#_M1016_d N_A1_M1016_g N_A_119_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1040 N_A_27_47#_M1040_d N_A1_M1040_g N_A_119_47#_M1016_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1051 N_A_27_47#_M1040_d N_A1_M1051_g N_A_119_47#_M1051_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1058 N_A_27_47#_M1058_d N_A1_M1058_g N_A_119_47#_M1051_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_119_47#_M1000_d N_S_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1020 N_A_119_47#_M1000_d N_S_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1023 N_A_119_47#_M1023_d N_S_M1023_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1054 N_A_119_47#_M1023_d N_S_M1054_g N_VGND_M1054_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1038 N_A_973_297#_M1038_d N_S_M1038_g N_VGND_M1054_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1039 N_A_973_297#_M1038_d N_S_M1039_g N_VGND_M1039_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1039_s N_A_973_297#_M1001_g N_A_1163_47#_M1001_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75003.1 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_973_297#_M1009_g N_A_1163_47#_M1001_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75003.5 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1009_d N_A_973_297#_M1024_g N_A_1163_47#_M1024_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75004 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1044 N_VGND_M1044_d N_A_973_297#_M1044_g N_A_1163_47#_M1024_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1
+ R=4.33333 SA=75004.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_27_47#_M1004_d N_A0_M1004_g N_A_1163_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1011_d N_A0_M1011_g N_A_1163_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1041 N_A_27_47#_M1011_d N_A0_M1041_g N_A_1163_47#_M1041_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1046 N_A_27_47#_M1046_d N_A0_M1046_g N_A_1163_47#_M1041_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_X_M1014_d N_A_27_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1017 N_X_M1014_d N_A_27_47#_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1021_d N_A_27_47#_M1021_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1025 N_X_M1021_d N_A_27_47#_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1027 N_X_M1027_d N_A_27_47#_M1027_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1033 N_X_M1027_d N_A_27_47#_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1034 N_X_M1034_d N_A_27_47#_M1034_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.1
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1043 N_X_M1034_d N_A_27_47#_M1043_g N_VGND_M1043_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1047 N_X_M1047_d N_A_27_47#_M1047_g N_VGND_M1043_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1052 N_X_M1047_d N_A_27_47#_M1052_g N_VGND_M1052_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1055 N_X_M1055_d N_A_27_47#_M1055_g N_VGND_M1052_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1059 N_X_M1055_d N_A_27_47#_M1059_g N_VGND_M1059_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1002_d N_A1_M1002_g N_A_117_297#_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1026 N_A_27_47#_M1026_d N_A1_M1026_g N_A_117_297#_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1035 N_A_27_47#_M1026_d N_A1_M1035_g N_A_117_297#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1048 N_A_27_47#_M1048_d N_A1_M1048_g N_A_117_297#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_S_M1006_g N_A_597_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_S_M1015_g N_A_597_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1042 N_VPWR_M1015_d N_S_M1042_g N_A_597_297#_M1042_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1056 N_VPWR_M1056_d N_S_M1056_g N_A_597_297#_M1042_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1056_d N_S_M1012_g N_A_973_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1032 N_VPWR_M1032_d N_S_M1032_g N_A_973_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1005 N_A_117_297#_M1005_d N_A_973_297#_M1005_g N_VPWR_M1032_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1029 N_A_117_297#_M1005_d N_A_973_297#_M1029_g N_VPWR_M1029_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1036 N_A_117_297#_M1036_d N_A_973_297#_M1036_g N_VPWR_M1029_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1049 N_A_117_297#_M1036_d N_A_973_297#_M1049_g N_VPWR_M1049_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90004.4 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_597_297#_M1008_d N_A0_M1008_g N_A_27_47#_M1008_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1010 N_A_597_297#_M1008_d N_A0_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1018 N_A_597_297#_M1018_d N_A0_M1018_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1030 N_A_597_297#_M1018_d N_A0_M1030_g N_A_27_47#_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_27_47#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90005.3 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_47#_M1007_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1007_d N_A_27_47#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A_27_47#_M1019_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1019_d N_A_27_47#_M1022_g N_X_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_A_27_47#_M1028_g N_X_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1031 N_VPWR_M1028_d N_A_27_47#_M1031_g N_X_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1037 N_VPWR_M1037_d N_A_27_47#_M1037_g N_X_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1045 N_VPWR_M1037_d N_A_27_47#_M1045_g N_X_M1045_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1050 N_VPWR_M1050_d N_A_27_47#_M1050_g N_X_M1045_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1053 N_VPWR_M1050_d N_A_27_47#_M1053_g N_X_M1053_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1057 N_VPWR_M1057_d N_A_27_47#_M1057_g N_X_M1053_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX60_noxref VNB VPB NWDIODE A=27.1887 P=37.09
*
.include "sky130_fd_sc_hdll__mux2_12.pxi.spice"
*
.ends
*
*
