* File: sky130_fd_sc_hdll__clkbuf_1.pxi.spice
* Created: Thu Aug 27 19:01:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_1%A_75_212# N_A_75_212#_M1001_d
+ N_A_75_212#_M1002_d N_A_75_212#_c_33_n N_A_75_212#_M1000_g N_A_75_212#_M1003_g
+ N_A_75_212#_c_35_n N_A_75_212#_c_39_n N_A_75_212#_c_36_n N_A_75_212#_c_59_p
+ N_A_75_212#_c_40_n N_A_75_212#_c_61_p N_A_75_212#_c_85_p N_A_75_212#_c_49_p
+ N_A_75_212#_c_37_n PM_SKY130_FD_SC_HDLL__CLKBUF_1%A_75_212#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_1%A N_A_M1001_g N_A_c_101_n N_A_c_102_n
+ N_A_M1002_g A N_A_c_99_n A PM_SKY130_FD_SC_HDLL__CLKBUF_1%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_1%X N_X_M1003_s N_X_M1000_s N_X_c_128_n
+ N_X_c_131_n N_X_c_129_n X X X PM_SKY130_FD_SC_HDLL__CLKBUF_1%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_1%VPWR N_VPWR_M1000_d N_VPWR_c_153_n VPWR
+ N_VPWR_c_154_n N_VPWR_c_155_n N_VPWR_c_152_n N_VPWR_c_157_n VPWR
+ PM_SKY130_FD_SC_HDLL__CLKBUF_1%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_1%VGND N_VGND_M1003_d VGND N_VGND_c_176_n
+ N_VGND_c_177_n N_VGND_c_178_n N_VGND_c_179_n VGND
+ PM_SKY130_FD_SC_HDLL__CLKBUF_1%VGND
cc_1 VNB N_A_75_212#_c_33_n 0.0258937f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.62
cc_2 VNB N_A_75_212#_M1003_g 0.0328054f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.495
cc_3 VNB N_A_75_212#_c_35_n 0.00338912f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.06
cc_4 VNB N_A_75_212#_c_36_n 0.020701f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.72
cc_5 VNB N_A_75_212#_c_37_n 0.00302584f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.225
cc_6 VNB N_A_M1001_g 0.0350981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_c_99_n 0.0424504f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.39
cc_8 VNB A 0.0188192f $X=-0.19 $Y=-0.24 $X2=1.54 $Y2=0.635
cc_9 VNB N_X_c_128_n 0.00850613f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.06
cc_10 VNB N_X_c_129_n 0.0255134f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.495
cc_11 VNB X 0.0145716f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_152_n 0.079965f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=0.72
cc_13 VNB N_VGND_c_176_n 0.0166815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_VGND_c_177_n 0.126858f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=0.805
cc_15 VNB N_VGND_c_178_n 0.01537f $X=-0.19 $Y=-0.24 $X2=0.76 $Y2=0.72
cc_16 VNB N_VGND_c_179_n 0.0137863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VPB N_A_75_212#_c_33_n 0.0470586f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.62
cc_18 VPB N_A_75_212#_c_39_n 0.00206391f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.535
cc_19 VPB N_A_75_212#_c_40_n 0.0263515f $X=-0.19 $Y=1.305 $X2=1.495 $Y2=1.62
cc_20 VPB N_A_75_212#_c_37_n 0.00123503f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.225
cc_21 VPB N_A_c_101_n 0.0185466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_22 VPB N_A_c_102_n 0.0293303f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.62
cc_23 VPB N_A_c_99_n 0.00985919f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.39
cc_24 VPB A 0.00696807f $X=-0.19 $Y=1.305 $X2=1.54 $Y2=0.635
cc_25 VPB N_X_c_131_n 0.0110422f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.495
cc_26 VPB N_X_c_129_n 0.0119024f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.495
cc_27 VPB X 0.0297138f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=0.805
cc_28 VPB N_VPWR_c_153_n 0.0022004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_154_n 0.0152818f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.06
cc_30 VPB N_VPWR_c_155_n 0.0174954f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.535
cc_31 VPB N_VPWR_c_152_n 0.0449489f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=0.72
cc_32 VPB N_VPWR_c_157_n 0.0117963f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=1.62
cc_33 N_A_75_212#_M1003_g N_A_M1001_g 0.00793399f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_34 N_A_75_212#_c_35_n N_A_M1001_g 0.00375164f $X=0.65 $Y=1.06 $X2=0 $Y2=0
cc_35 N_A_75_212#_c_36_n N_A_M1001_g 0.0177047f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_36 N_A_75_212#_c_33_n N_A_c_101_n 0.0027433f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_37 N_A_75_212#_c_39_n N_A_c_101_n 0.0025074f $X=0.65 $Y=1.535 $X2=0 $Y2=0
cc_38 N_A_75_212#_c_33_n N_A_c_102_n 0.00369035f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_39 N_A_75_212#_c_40_n N_A_c_102_n 0.0236505f $X=1.495 $Y=1.62 $X2=0 $Y2=0
cc_40 N_A_75_212#_c_49_p N_A_c_102_n 0.00654464f $X=1.58 $Y=1.96 $X2=0 $Y2=0
cc_41 N_A_75_212#_c_33_n N_A_c_99_n 0.00578119f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_42 N_A_75_212#_c_36_n N_A_c_99_n 0.00167163f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_43 N_A_75_212#_c_40_n N_A_c_99_n 0.00155496f $X=1.495 $Y=1.62 $X2=0 $Y2=0
cc_44 N_A_75_212#_c_37_n N_A_c_99_n 0.00321913f $X=0.65 $Y=1.225 $X2=0 $Y2=0
cc_45 N_A_75_212#_c_33_n A 2.65858e-19 $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_46 N_A_75_212#_c_35_n A 0.00217834f $X=0.65 $Y=1.06 $X2=0 $Y2=0
cc_47 N_A_75_212#_c_36_n A 0.0209602f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_48 N_A_75_212#_c_40_n A 0.0238708f $X=1.495 $Y=1.62 $X2=0 $Y2=0
cc_49 N_A_75_212#_c_37_n A 0.00899296f $X=0.65 $Y=1.225 $X2=0 $Y2=0
cc_50 N_A_75_212#_c_59_p N_X_c_128_n 0.00910805f $X=0.76 $Y=0.72 $X2=0 $Y2=0
cc_51 N_A_75_212#_c_33_n N_X_c_131_n 0.00358938f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_52 N_A_75_212#_c_61_p N_X_c_131_n 0.0107806f $X=0.76 $Y=1.62 $X2=0 $Y2=0
cc_53 N_A_75_212#_c_33_n N_X_c_129_n 0.0116224f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_54 N_A_75_212#_M1003_g N_X_c_129_n 0.0059516f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_55 N_A_75_212#_c_35_n N_X_c_129_n 0.0126005f $X=0.65 $Y=1.06 $X2=0 $Y2=0
cc_56 N_A_75_212#_c_39_n N_X_c_129_n 0.00716662f $X=0.65 $Y=1.535 $X2=0 $Y2=0
cc_57 N_A_75_212#_c_59_p N_X_c_129_n 0.00241035f $X=0.76 $Y=0.72 $X2=0 $Y2=0
cc_58 N_A_75_212#_c_61_p N_X_c_129_n 0.00132712f $X=0.76 $Y=1.62 $X2=0 $Y2=0
cc_59 N_A_75_212#_c_37_n N_X_c_129_n 0.0247996f $X=0.65 $Y=1.225 $X2=0 $Y2=0
cc_60 N_A_75_212#_M1003_g X 0.00660891f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_61 N_A_75_212#_c_40_n N_VPWR_M1000_d 0.00478986f $X=1.495 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A_75_212#_c_61_p N_VPWR_M1000_d 0.00126472f $X=0.76 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_63 N_A_75_212#_c_33_n N_VPWR_c_153_n 0.0172722f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_64 N_A_75_212#_c_40_n N_VPWR_c_153_n 0.0370038f $X=1.495 $Y=1.62 $X2=0 $Y2=0
cc_65 N_A_75_212#_c_61_p N_VPWR_c_153_n 0.0136314f $X=0.76 $Y=1.62 $X2=0 $Y2=0
cc_66 N_A_75_212#_c_49_p N_VPWR_c_153_n 0.0378335f $X=1.58 $Y=1.96 $X2=0 $Y2=0
cc_67 N_A_75_212#_c_37_n N_VPWR_c_153_n 5.10987e-19 $X=0.65 $Y=1.225 $X2=0 $Y2=0
cc_68 N_A_75_212#_c_33_n N_VPWR_c_154_n 0.0046653f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_69 N_A_75_212#_c_49_p N_VPWR_c_155_n 0.0118139f $X=1.58 $Y=1.96 $X2=0 $Y2=0
cc_70 N_A_75_212#_M1002_d N_VPWR_c_152_n 0.00568146f $X=1.435 $Y=1.695 $X2=0
+ $Y2=0
cc_71 N_A_75_212#_c_33_n N_VPWR_c_152_n 0.00885548f $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_72 N_A_75_212#_c_49_p N_VPWR_c_152_n 0.00646998f $X=1.58 $Y=1.96 $X2=0 $Y2=0
cc_73 N_A_75_212#_c_36_n N_VGND_M1003_d 0.00628718f $X=1.455 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_75_212#_c_59_p N_VGND_M1003_d 0.00112549f $X=0.76 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_75_212#_c_36_n N_VGND_c_176_n 0.00253436f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_76 N_A_75_212#_c_85_p N_VGND_c_176_n 0.0116326f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_77 N_A_75_212#_M1001_d N_VGND_c_177_n 0.00381741f $X=1.395 $Y=0.235 $X2=0
+ $Y2=0
cc_78 N_A_75_212#_M1003_g N_VGND_c_177_n 0.0065495f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_79 N_A_75_212#_c_36_n N_VGND_c_177_n 0.00675301f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_80 N_A_75_212#_c_59_p N_VGND_c_177_n 0.00104135f $X=0.76 $Y=0.72 $X2=0 $Y2=0
cc_81 N_A_75_212#_c_85_p N_VGND_c_177_n 0.00643448f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_82 N_A_75_212#_M1003_g N_VGND_c_178_n 0.00310428f $X=0.52 $Y=0.495 $X2=0
+ $Y2=0
cc_83 N_A_75_212#_c_33_n N_VGND_c_179_n 2.5127e-19 $X=0.495 $Y=1.62 $X2=0 $Y2=0
cc_84 N_A_75_212#_M1003_g N_VGND_c_179_n 0.0121205f $X=0.52 $Y=0.495 $X2=0 $Y2=0
cc_85 N_A_75_212#_c_36_n N_VGND_c_179_n 0.0345378f $X=1.455 $Y=0.72 $X2=0 $Y2=0
cc_86 N_A_75_212#_c_59_p N_VGND_c_179_n 0.0129045f $X=0.76 $Y=0.72 $X2=0 $Y2=0
cc_87 N_A_75_212#_c_85_p N_VGND_c_179_n 0.0157111f $X=1.54 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_75_212#_c_37_n N_VGND_c_179_n 4.4673e-19 $X=0.65 $Y=1.225 $X2=0 $Y2=0
cc_89 N_A_c_102_n N_VPWR_c_153_n 0.0141428f $X=1.345 $Y=1.62 $X2=0 $Y2=0
cc_90 N_A_c_102_n N_VPWR_c_155_n 0.00622633f $X=1.345 $Y=1.62 $X2=0 $Y2=0
cc_91 N_A_c_102_n N_VPWR_c_152_n 0.0113126f $X=1.345 $Y=1.62 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_VGND_c_176_n 0.00339367f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_93 N_A_M1001_g N_VGND_c_177_n 0.00500869f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_94 N_A_M1001_g N_VGND_c_179_n 0.00959243f $X=1.32 $Y=0.495 $X2=0 $Y2=0
cc_95 X N_VPWR_c_154_n 0.0187043f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_96 N_X_M1000_s N_VPWR_c_152_n 0.00391095f $X=0.135 $Y=1.695 $X2=0 $Y2=0
cc_97 X N_VPWR_c_152_n 0.0103212f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_98 N_X_M1003_s N_VGND_c_177_n 0.0060443f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_99 X N_VGND_c_177_n 0.00990988f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_100 X N_VGND_c_178_n 0.0180762f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_101 X N_VGND_c_179_n 0.016191f $X=0.145 $Y=0.425 $X2=0 $Y2=0
