* File: sky130_fd_sc_hdll__o221ai_4.pex.spice
* Created: Wed Sep  2 08:45:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%C1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 45
r61 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r62 38 45 28.0045 $w=1.98e-07 $l=5.05e-07 $layer=LI1_cond $X=1.66 $Y=1.175
+ $X2=1.155 $Y2=1.175
r63 37 39 34.5216 $w=3.7e-07 $l=2.65e-07 $layer=POLY_cond $X=1.66 $Y=1.202
+ $X2=1.925 $Y2=1.202
r64 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.66
+ $Y=1.16 $X2=1.66 $Y2=1.16
r65 35 37 23.4486 $w=3.7e-07 $l=1.8e-07 $layer=POLY_cond $X=1.48 $Y=1.202
+ $X2=1.66 $Y2=1.202
r66 34 35 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r67 33 34 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=1.01 $Y=1.202
+ $X2=1.455 $Y2=1.202
r68 32 33 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r69 31 32 57.9703 $w=3.7e-07 $l=4.45e-07 $layer=POLY_cond $X=0.54 $Y=1.202
+ $X2=0.985 $Y2=1.202
r70 30 31 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r71 28 30 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r72 28 29 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r73 25 45 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.14 $Y=1.175
+ $X2=1.155 $Y2=1.175
r74 25 29 36.0455 $w=1.98e-07 $l=6.5e-07 $layer=LI1_cond $X=1.14 $Y=1.175
+ $X2=0.49 $Y2=1.175
r75 22 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r76 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r77 19 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r78 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r79 16 35 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r80 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r81 13 34 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r82 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r83 10 33 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r84 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r85 7 32 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r86 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r87 4 31 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r88 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r89 1 30 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r90 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 26 27 28 29 31 36 48 53
c99 28 0 1.6089e-19 $X=4.925 $Y=1.53
r100 48 49 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.855 $Y=1.202
+ $X2=3.88 $Y2=1.202
r101 46 48 18.0912 $w=3.73e-07 $l=1.4e-07 $layer=POLY_cond $X=3.715 $Y=1.202
+ $X2=3.855 $Y2=1.202
r102 46 47 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.715
+ $Y=1.16 $X2=3.715 $Y2=1.16
r103 44 46 39.4129 $w=3.73e-07 $l=3.05e-07 $layer=POLY_cond $X=3.41 $Y=1.202
+ $X2=3.715 $Y2=1.202
r104 43 44 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.385 $Y=1.202
+ $X2=3.41 $Y2=1.202
r105 42 43 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=2.94 $Y=1.202
+ $X2=3.385 $Y2=1.202
r106 40 42 0.646113 $w=3.73e-07 $l=5e-09 $layer=POLY_cond $X=2.935 $Y=1.202
+ $X2=2.94 $Y2=1.202
r107 40 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r108 38 40 2.58445 $w=3.73e-07 $l=2e-08 $layer=POLY_cond $X=2.915 $Y=1.202
+ $X2=2.935 $Y2=1.202
r109 36 47 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=3.265 $Y=1.175
+ $X2=3.715 $Y2=1.175
r110 36 53 18.3 $w=1.98e-07 $l=3.3e-07 $layer=LI1_cond $X=3.265 $Y=1.175
+ $X2=2.935 $Y2=1.175
r111 31 34 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.205 $Y=1.16
+ $X2=6.205 $Y2=1.53
r112 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=1.16 $X2=6.18 $Y2=1.16
r113 29 47 56.5636 $w=1.98e-07 $l=1.02e-06 $layer=LI1_cond $X=4.735 $Y=1.175
+ $X2=3.715 $Y2=1.175
r114 27 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.015 $Y=1.53
+ $X2=6.205 $Y2=1.53
r115 27 28 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=6.015 $Y=1.53
+ $X2=4.925 $Y2=1.53
r116 26 28 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=4.83 $Y=1.445
+ $X2=4.925 $Y2=1.53
r117 25 29 6.82232 $w=2e-07 $l=1.39642e-07 $layer=LI1_cond $X=4.83 $Y=1.275
+ $X2=4.735 $Y2=1.175
r118 25 26 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=4.83 $Y=1.275
+ $X2=4.83 $Y2=1.445
r119 22 32 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.205 $Y2=1.16
r120 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.23 $Y2=0.56
r121 19 32 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.16
r122 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.985
r123 16 49 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=1.202
r124 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.88 $Y=0.995
+ $X2=3.88 $Y2=0.56
r125 13 48 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.202
r126 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.985
r127 10 44 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=1.202
r128 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r129 7 43 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.202
r130 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.985
r131 4 42 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=1.202
r132 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.94 $Y=0.995
+ $X2=2.94 $Y2=0.56
r133 1 38 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.202
r134 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.915 $Y=1.41
+ $X2=2.915 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 35 36 41
c72 4 0 1.6089e-19 $X=4.325 $Y=1.41
r73 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.735 $Y=1.202
+ $X2=5.76 $Y2=1.202
r74 35 41 8.02594 $w=2.78e-07 $l=1.95e-07 $layer=LI1_cond $X=5.65 $Y=1.135
+ $X2=5.455 $Y2=1.135
r75 34 36 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=5.65 $Y=1.202
+ $X2=5.735 $Y2=1.202
r76 34 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.65
+ $Y=1.16 $X2=5.65 $Y2=1.16
r77 32 34 49.8844 $w=3.72e-07 $l=3.85e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.65 $Y2=1.202
r78 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.265 $Y2=1.202
r79 30 31 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=5.24 $Y2=1.202
r80 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.77 $Y=1.202
+ $X2=4.795 $Y2=1.202
r81 28 29 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=4.325 $Y=1.202
+ $X2=4.77 $Y2=1.202
r82 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.3 $Y=1.202
+ $X2=4.325 $Y2=1.202
r83 25 41 6.1738 $w=2.78e-07 $l=1.5e-07 $layer=LI1_cond $X=5.305 $Y=1.135
+ $X2=5.455 $Y2=1.135
r84 22 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=1.202
r85 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.76 $Y=0.995
+ $X2=5.76 $Y2=0.56
r86 19 36 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.202
r87 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.985
r88 16 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.202
r89 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.985
r90 13 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r91 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r92 10 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.202
r93 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.985
r94 7 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.202
r95 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995 $X2=4.77
+ $Y2=0.56
r96 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.202
r97 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.985
r98 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=0.995 $X2=4.3
+ $Y2=1.202
r99 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.3 $Y=0.995 $X2=4.3
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 39 49 50 54
c114 4 0 2.98607e-20 $X=6.78 $Y=0.995
r115 50 51 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=10.02 $Y=1.202
+ $X2=10.045 $Y2=1.202
r116 49 54 25.7864 $w=1.98e-07 $l=4.65e-07 $layer=LI1_cond $X=9.95 $Y=1.175
+ $X2=9.485 $Y2=1.175
r117 48 50 9.04558 $w=3.73e-07 $l=7e-08 $layer=POLY_cond $X=9.95 $Y=1.202
+ $X2=10.02 $Y2=1.202
r118 48 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.95
+ $Y=1.16 $X2=9.95 $Y2=1.16
r119 46 48 48.4584 $w=3.73e-07 $l=3.75e-07 $layer=POLY_cond $X=9.575 $Y=1.202
+ $X2=9.95 $Y2=1.202
r120 45 46 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=9.55 $Y=1.202
+ $X2=9.575 $Y2=1.202
r121 42 43 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=9.08 $Y=1.202
+ $X2=9.105 $Y2=1.202
r122 39 54 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=9.435 $Y=1.175
+ $X2=9.485 $Y2=1.175
r123 38 45 49.1046 $w=3.73e-07 $l=3.8e-07 $layer=POLY_cond $X=9.17 $Y=1.202
+ $X2=9.55 $Y2=1.202
r124 38 43 8.39946 $w=3.73e-07 $l=6.5e-08 $layer=POLY_cond $X=9.17 $Y=1.202
+ $X2=9.105 $Y2=1.202
r125 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.17
+ $Y=1.16 $X2=9.17 $Y2=1.16
r126 35 39 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=9.32 $Y=1.175
+ $X2=9.435 $Y2=1.175
r127 35 37 4.45102 $w=2e-07 $l=1.58e-07 $layer=LI1_cond $X=9.32 $Y=1.175
+ $X2=9.162 $Y2=1.175
r128 30 33 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=6.755 $Y=1.16
+ $X2=6.755 $Y2=1.53
r129 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.73
+ $Y=1.16 $X2=6.73 $Y2=1.16
r130 27 37 2.8171 $w=3.15e-07 $l=1e-07 $layer=LI1_cond $X=9.162 $Y=1.275
+ $X2=9.162 $Y2=1.175
r131 27 28 6.21953 $w=3.13e-07 $l=1.7e-07 $layer=LI1_cond $X=9.162 $Y=1.275
+ $X2=9.162 $Y2=1.445
r132 26 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.945 $Y=1.53
+ $X2=6.755 $Y2=1.53
r133 25 28 7.64049 $w=1.7e-07 $l=1.94921e-07 $layer=LI1_cond $X=9.005 $Y=1.53
+ $X2=9.162 $Y2=1.445
r134 25 26 134.396 $w=1.68e-07 $l=2.06e-06 $layer=LI1_cond $X=9.005 $Y=1.53
+ $X2=6.945 $Y2=1.53
r135 22 51 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.045 $Y=1.41
+ $X2=10.045 $Y2=1.202
r136 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.045 $Y=1.41
+ $X2=10.045 $Y2=1.985
r137 19 50 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.02 $Y=0.995
+ $X2=10.02 $Y2=1.202
r138 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.02 $Y=0.995
+ $X2=10.02 $Y2=0.56
r139 16 46 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.575 $Y=1.41
+ $X2=9.575 $Y2=1.202
r140 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.575 $Y=1.41
+ $X2=9.575 $Y2=1.985
r141 13 45 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.55 $Y=0.995
+ $X2=9.55 $Y2=1.202
r142 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.55 $Y=0.995
+ $X2=9.55 $Y2=0.56
r143 10 43 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.105 $Y=1.41
+ $X2=9.105 $Y2=1.202
r144 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.105 $Y=1.41
+ $X2=9.105 $Y2=1.985
r145 7 42 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=1.202
r146 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=0.56
r147 4 31 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.755 $Y2=1.16
r148 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.78 $Y2=0.56
r149 1 31 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.755 $Y=1.41
+ $X2=6.755 $Y2=1.16
r150 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.755 $Y=1.41
+ $X2=6.755 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39 44
c81 22 0 2.98607e-20 $X=8.66 $Y=0.995
r82 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.635 $Y=1.202
+ $X2=8.66 $Y2=1.202
r83 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=8.46 $Y=1.202
+ $X2=8.635 $Y2=1.202
r84 37 38 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.46
+ $Y=1.16 $X2=8.46 $Y2=1.16
r85 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=8.165 $Y=1.202
+ $X2=8.46 $Y2=1.202
r86 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.14 $Y=1.202
+ $X2=8.165 $Y2=1.202
r87 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.695 $Y=1.202
+ $X2=8.14 $Y2=1.202
r88 32 44 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=7.68 $Y=1.175 $X2=7.9
+ $Y2=1.175
r89 31 33 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=7.68 $Y=1.202
+ $X2=7.695 $Y2=1.202
r90 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.68
+ $Y=1.16 $X2=7.68 $Y2=1.16
r91 29 31 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=7.67 $Y=1.202 $X2=7.68
+ $Y2=1.202
r92 28 29 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.225 $Y=1.202
+ $X2=7.67 $Y2=1.202
r93 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.2 $Y=1.202
+ $X2=7.225 $Y2=1.202
r94 25 38 30.7773 $w=1.98e-07 $l=5.55e-07 $layer=LI1_cond $X=7.905 $Y=1.175
+ $X2=8.46 $Y2=1.175
r95 25 44 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=7.905 $Y=1.175
+ $X2=7.9 $Y2=1.175
r96 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.66 $Y2=1.202
r97 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.66 $Y2=0.56
r98 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.635 $Y=1.41
+ $X2=8.635 $Y2=1.202
r99 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.635 $Y=1.41
+ $X2=8.635 $Y2=1.985
r100 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.165 $Y=1.41
+ $X2=8.165 $Y2=1.202
r101 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.165 $Y=1.41
+ $X2=8.165 $Y2=1.985
r102 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=1.202
r103 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=0.56
r104 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.695 $Y=1.41
+ $X2=7.695 $Y2=1.202
r105 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.695 $Y=1.41
+ $X2=7.695 $Y2=1.985
r106 7 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=1.202
r107 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.67 $Y=0.995
+ $X2=7.67 $Y2=0.56
r108 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.225 $Y=1.41
+ $X2=7.225 $Y2=1.202
r109 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.225 $Y=1.41
+ $X2=7.225 $Y2=1.985
r110 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.2 $Y=0.995
+ $X2=7.2 $Y2=1.202
r111 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.2 $Y=0.995 $X2=7.2
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 38 42 46
+ 48 50 55 56 58 59 61 62 63 81 89 94 100 103
r130 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r131 99 100 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.68 $Y=2.465
+ $X2=2.805 $Y2=2.465
r132 96 99 2.63841 $w=6.78e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=2.465
+ $X2=2.68 $Y2=2.465
r133 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 93 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r135 92 96 8.09112 $w=6.78e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=2.465
+ $X2=2.53 $Y2=2.465
r136 92 94 8.38974 $w=6.78e-07 $l=3.5e-08 $layer=LI1_cond $X=2.07 $Y=2.465
+ $X2=2.035 $Y2=2.465
r137 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r138 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r139 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 84 103 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r141 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r142 81 102 3.94362 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=10.367 $Y2=2.72
r143 81 83 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=10.155 $Y=2.72
+ $X2=9.89 $Y2=2.72
r144 80 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r145 79 80 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r146 77 80 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.97 $Y2=2.72
r147 76 79 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.97 $Y2=2.72
r148 76 77 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r149 74 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r150 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r151 71 74 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=6.21 $Y2=2.72
r152 70 73 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=6.21 $Y2=2.72
r153 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r154 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r155 68 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r156 67 100 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.805 $Y2=2.72
r157 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r158 63 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r159 63 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r160 61 79 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.215 $Y=2.72
+ $X2=8.97 $Y2=2.72
r161 61 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.215 $Y=2.72
+ $X2=9.34 $Y2=2.72
r162 60 83 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=9.465 $Y=2.72
+ $X2=9.89 $Y2=2.72
r163 60 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.465 $Y=2.72
+ $X2=9.34 $Y2=2.72
r164 58 73 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.21 $Y2=2.72
r165 58 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.355 $Y=2.72
+ $X2=6.48 $Y2=2.72
r166 57 76 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.67 $Y2=2.72
r167 57 59 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.48 $Y2=2.72
r168 55 67 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.495 $Y=2.72
+ $X2=3.45 $Y2=2.72
r169 55 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.495 $Y=2.72
+ $X2=3.62 $Y2=2.72
r170 54 70 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.745 $Y=2.72
+ $X2=3.91 $Y2=2.72
r171 54 56 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.745 $Y=2.72
+ $X2=3.62 $Y2=2.72
r172 50 53 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=10.28 $Y=1.62
+ $X2=10.28 $Y2=2.3
r173 48 102 3.19954 $w=2.5e-07 $l=1.22327e-07 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.367 $Y2=2.72
r174 48 53 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.28 $Y2=2.3
r175 44 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.34 $Y=2.635
+ $X2=9.34 $Y2=2.72
r176 44 46 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.34 $Y=2.635
+ $X2=9.34 $Y2=2.3
r177 40 59 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=2.635
+ $X2=6.48 $Y2=2.72
r178 40 42 13.1378 $w=2.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.48 $Y=2.635
+ $X2=6.48 $Y2=2.35
r179 36 56 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.72
r180 36 38 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.62 $Y=2.635
+ $X2=3.62 $Y2=2.3
r181 35 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.22 $Y2=2.72
r182 35 94 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=2.035 $Y2=2.72
r183 30 89 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r184 30 32 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=1.99
r185 29 86 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r186 28 89 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=1.22 $Y2=2.72
r187 28 29 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.405 $Y2=2.72
r188 24 27 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.28 $Y=1.65
+ $X2=0.28 $Y2=2.33
r189 22 86 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.202 $Y2=2.72
r190 22 27 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=2.33
r191 7 53 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.485 $X2=10.28 $Y2=2.3
r192 7 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.485 $X2=10.28 $Y2=1.62
r193 6 46 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.195
+ $Y=1.485 $X2=9.34 $Y2=2.3
r194 5 42 600 $w=1.7e-07 $l=9.53021e-07 $layer=licon1_PDIFF $count=1 $X=6.295
+ $Y=1.485 $X2=6.48 $Y2=2.35
r195 4 38 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.62 $Y2=2.3
r196 3 99 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.68 $Y2=2.3
r197 2 32 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.99
r198 1 27 400 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.33
r199 1 24 400 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%Y 1 2 3 4 5 6 7 8 25 33 38 41 44 45 48 51
+ 53 57 66
r115 64 66 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=7.46 $Y=1.895
+ $X2=8.4 $Y2=1.895
r116 57 64 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=6.67 $Y=1.895
+ $X2=7.46 $Y2=1.895
r117 57 60 61.289 $w=2.18e-07 $l=1.17e-06 $layer=LI1_cond $X=6.67 $Y=1.895
+ $X2=5.5 $Y2=1.895
r118 54 60 48.9788 $w=2.18e-07 $l=9.35e-07 $layer=LI1_cond $X=4.565 $Y=1.895
+ $X2=5.5 $Y2=1.895
r119 54 56 3.40825 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.565 $Y=1.895
+ $X2=4.455 $Y2=1.895
r120 52 53 8.12479 $w=5.08e-07 $l=1.03e-07 $layer=LI1_cond $X=2.222 $Y=1.7
+ $X2=2.325 $Y2=1.7
r121 50 52 12.4767 $w=5.08e-07 $l=5.32e-07 $layer=LI1_cond $X=1.69 $Y=1.7
+ $X2=2.222 $Y2=1.7
r122 50 51 8.64074 $w=5.08e-07 $l=1.25e-07 $layer=LI1_cond $X=1.69 $Y=1.7
+ $X2=1.565 $Y2=1.7
r123 48 56 3.40825 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=4.455 $Y=1.785
+ $X2=4.455 $Y2=1.895
r124 47 48 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=4.455 $Y=1.615
+ $X2=4.455 $Y2=1.785
r125 45 47 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.345 $Y=1.53
+ $X2=4.455 $Y2=1.615
r126 45 53 131.786 $w=1.68e-07 $l=2.02e-06 $layer=LI1_cond $X=4.345 $Y=1.53
+ $X2=2.325 $Y2=1.53
r127 44 52 6.13047 $w=2.05e-07 $l=2.55e-07 $layer=LI1_cond $X=2.222 $Y=1.445
+ $X2=2.222 $Y2=1.7
r128 43 44 31.3792 $w=2.03e-07 $l=5.8e-07 $layer=LI1_cond $X=2.222 $Y=0.865
+ $X2=2.222 $Y2=1.445
r129 39 50 4.91917 $w=2.5e-07 $l=2.55e-07 $layer=LI1_cond $X=1.69 $Y=1.955
+ $X2=1.69 $Y2=1.7
r130 39 41 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.69 $Y=1.955
+ $X2=1.69 $Y2=1.96
r131 38 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.875 $Y=1.53
+ $X2=1.565 $Y2=1.53
r132 33 35 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.75 $Y=1.62
+ $X2=0.75 $Y2=2.3
r133 31 38 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.75 $Y=1.615
+ $X2=0.875 $Y2=1.53
r134 31 33 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.75 $Y=1.615
+ $X2=0.75 $Y2=1.62
r135 27 30 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=0.75 $Y=0.755
+ $X2=1.69 $Y2=0.755
r136 25 43 6.82754 $w=2.2e-07 $l=1.52709e-07 $layer=LI1_cond $X=2.12 $Y=0.755
+ $X2=2.222 $Y2=0.865
r137 25 30 22.525 $w=2.18e-07 $l=4.3e-07 $layer=LI1_cond $X=2.12 $Y=0.755
+ $X2=1.69 $Y2=0.755
r138 8 66 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=8.255
+ $Y=1.485 $X2=8.4 $Y2=1.92
r139 7 64 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=7.315
+ $Y=1.485 $X2=7.46 $Y2=1.92
r140 6 60 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=5.355
+ $Y=1.485 $X2=5.5 $Y2=1.92
r141 5 56 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.485 $X2=4.56 $Y2=1.92
r142 4 50 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r143 4 41 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
r144 3 35 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.3
r145 3 33 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.62
r146 2 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.73
r147 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A_601_297# 1 2 3 4 15 17 18 22 23 27
r37 25 27 52.1273 $w=1.98e-07 $l=9.4e-07 $layer=LI1_cond $X=5.03 $Y=2.365
+ $X2=5.97 $Y2=2.365
r38 23 25 47.4136 $w=1.98e-07 $l=8.55e-07 $layer=LI1_cond $X=4.175 $Y=2.365
+ $X2=5.03 $Y2=2.365
r39 20 23 6.82177 $w=2e-07 $l=1.46714e-07 $layer=LI1_cond $X=4.07 $Y=2.265
+ $X2=4.175 $Y2=2.365
r40 20 22 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=4.07 $Y=2.265
+ $X2=4.07 $Y2=1.96
r41 19 22 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=4.07 $Y=1.955
+ $X2=4.07 $Y2=1.96
r42 17 19 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.965 $Y=1.87
+ $X2=4.07 $Y2=1.955
r43 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.965 $Y=1.87
+ $X2=3.275 $Y2=1.87
r44 13 18 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.15 $Y=1.955
+ $X2=3.275 $Y2=1.87
r45 13 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.15 $Y=1.955
+ $X2=3.15 $Y2=1.96
r46 4 27 600 $w=1.7e-07 $l=9.34692e-07 $layer=licon1_PDIFF $count=1 $X=5.825
+ $Y=1.485 $X2=5.97 $Y2=2.35
r47 3 25 600 $w=1.7e-07 $l=9.34692e-07 $layer=licon1_PDIFF $count=1 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=2.35
r48 2 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=1.96
r49 1 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.005
+ $Y=1.485 $X2=3.15 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A_1369_297# 1 2 3 4 13 22 23 24 27 31
r42 29 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=1.955
+ $X2=9.81 $Y2=1.87
r43 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=9.81 $Y=1.955
+ $X2=9.81 $Y2=1.96
r44 25 33 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=1.785
+ $X2=9.81 $Y2=1.87
r45 25 27 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=9.81 $Y=1.785
+ $X2=9.81 $Y2=1.62
r46 23 33 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.685 $Y=1.87
+ $X2=9.81 $Y2=1.87
r47 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.685 $Y=1.87
+ $X2=8.995 $Y2=1.87
r48 20 22 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=8.89 $Y=2.265
+ $X2=8.89 $Y2=1.96
r49 19 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.89 $Y=1.955
+ $X2=8.995 $Y2=1.87
r50 19 22 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=8.89 $Y=1.955
+ $X2=8.89 $Y2=1.96
r51 15 18 52.1273 $w=1.98e-07 $l=9.4e-07 $layer=LI1_cond $X=6.99 $Y=2.365
+ $X2=7.93 $Y2=2.365
r52 13 20 6.82177 $w=2e-07 $l=1.46714e-07 $layer=LI1_cond $X=8.785 $Y=2.365
+ $X2=8.89 $Y2=2.265
r53 13 18 47.4136 $w=1.98e-07 $l=8.55e-07 $layer=LI1_cond $X=8.785 $Y=2.365
+ $X2=7.93 $Y2=2.365
r54 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.665
+ $Y=1.485 $X2=9.81 $Y2=1.96
r55 4 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.665
+ $Y=1.485 $X2=9.81 $Y2=1.62
r56 3 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.725
+ $Y=1.485 $X2=8.87 $Y2=1.96
r57 2 18 600 $w=1.7e-07 $l=9.34692e-07 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=1.485 $X2=7.93 $Y2=2.35
r58 1 15 600 $w=1.7e-07 $l=9.34692e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.485 $X2=6.99 $Y2=2.35
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A_27_47# 1 2 3 4 5 6 7 22 24 38
r47 36 38 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=5.03 $Y=0.365
+ $X2=5.97 $Y2=0.365
r48 34 36 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=4.09 $Y=0.365
+ $X2=5.03 $Y2=0.365
r49 32 34 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=3.15 $Y=0.365
+ $X2=4.09 $Y2=0.365
r50 30 32 51.8599 $w=2.18e-07 $l=9.9e-07 $layer=LI1_cond $X=2.16 $Y=0.365
+ $X2=3.15 $Y2=0.365
r51 28 30 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=1.22 $Y=0.365
+ $X2=2.16 $Y2=0.365
r52 26 41 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.365 $Y=0.365
+ $X2=0.24 $Y2=0.365
r53 26 28 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=0.365 $Y=0.365
+ $X2=1.22 $Y2=0.365
r54 22 41 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.24 $Y=0.475
+ $X2=0.24 $Y2=0.365
r55 22 24 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=0.475
+ $X2=0.24 $Y2=0.73
r56 7 38 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.835
+ $Y=0.235 $X2=5.97 $Y2=0.39
r57 6 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=5.03 $Y2=0.39
r58 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.39
r59 4 32 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.015
+ $Y=0.235 $X2=3.15 $Y2=0.39
r60 3 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r61 2 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r62 1 41 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
r63 1 24 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%A_511_47# 1 2 3 4 5 6 7 8 9 40 42 46 48
+ 52 54 58 60 64 67 69 70 71 72
c127 72 0 2.98607e-20 $X=9.315 $Y=0.815
c128 70 0 2.98607e-20 $X=7.435 $Y=0.815
r129 62 64 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.255 $Y=0.725
+ $X2=10.255 $Y2=0.39
r130 61 72 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=9.505 $Y=0.815
+ $X2=9.315 $Y2=0.815
r131 60 62 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=10.065 $Y=0.815
+ $X2=10.255 $Y2=0.725
r132 60 61 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=10.065 $Y=0.815
+ $X2=9.505 $Y2=0.815
r133 56 72 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=9.315 $Y=0.725
+ $X2=9.315 $Y2=0.815
r134 56 58 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.315 $Y=0.725
+ $X2=9.315 $Y2=0.39
r135 55 71 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=8.565 $Y=0.82
+ $X2=8.375 $Y2=0.815
r136 54 72 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=9.125 $Y=0.82
+ $X2=9.315 $Y2=0.815
r137 54 55 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.125 $Y=0.82
+ $X2=8.565 $Y2=0.82
r138 50 71 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=8.375 $Y=0.725
+ $X2=8.375 $Y2=0.815
r139 50 52 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.375 $Y=0.725
+ $X2=8.375 $Y2=0.39
r140 49 70 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=7.625 $Y=0.815
+ $X2=7.435 $Y2=0.815
r141 48 71 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=8.185 $Y=0.815
+ $X2=8.375 $Y2=0.815
r142 48 49 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.185 $Y=0.815
+ $X2=7.625 $Y2=0.815
r143 44 70 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.435 $Y=0.725
+ $X2=7.435 $Y2=0.815
r144 44 46 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.435 $Y=0.725
+ $X2=7.435 $Y2=0.39
r145 42 70 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=7.245 $Y=0.82
+ $X2=7.435 $Y2=0.815
r146 42 69 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.245 $Y=0.82
+ $X2=6.685 $Y2=0.82
r147 38 69 8.69362 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=6.52 $Y=0.775
+ $X2=6.685 $Y2=0.775
r148 38 67 23.6207 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=6.52 $Y=0.775
+ $X2=6.015 $Y2=0.775
r149 38 40 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.52 $Y=0.645
+ $X2=6.52 $Y2=0.39
r150 37 67 32.639 $w=1.73e-07 $l=5.15e-07 $layer=LI1_cond $X=5.5 $Y=0.732
+ $X2=6.015 $Y2=0.732
r151 35 37 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=4.56 $Y=0.732
+ $X2=5.5 $Y2=0.732
r152 33 35 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=3.62 $Y=0.732
+ $X2=4.56 $Y2=0.732
r153 30 33 59.574 $w=1.73e-07 $l=9.4e-07 $layer=LI1_cond $X=2.68 $Y=0.732
+ $X2=3.62 $Y2=0.732
r154 9 64 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=10.095
+ $Y=0.235 $X2=10.28 $Y2=0.39
r155 8 58 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.155
+ $Y=0.235 $X2=9.34 $Y2=0.39
r156 7 52 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.215
+ $Y=0.235 $X2=8.4 $Y2=0.39
r157 6 46 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.275
+ $Y=0.235 $X2=7.46 $Y2=0.39
r158 5 38 182 $w=1.7e-07 $l=5.92832e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.235 $X2=6.52 $Y2=0.73
r159 5 40 182 $w=1.7e-07 $l=2.82046e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.235 $X2=6.52 $Y2=0.39
r160 4 37 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.73
r161 3 35 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.375
+ $Y=0.235 $X2=4.56 $Y2=0.73
r162 2 33 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.73
r163 1 30 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.68 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_4%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36
+ 37 39 40 41 60 61
r118 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r119 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r120 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r121 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r122 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r123 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r124 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r125 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r126 48 49 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r127 44 48 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=6.67
+ $Y2=0
r128 41 49 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=6.67
+ $Y2=0
r129 41 44 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r130 39 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.725 $Y=0 $X2=9.43
+ $Y2=0
r131 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.725 $Y=0 $X2=9.81
+ $Y2=0
r132 38 60 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=9.895 $Y=0
+ $X2=10.35 $Y2=0
r133 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.895 $Y=0 $X2=9.81
+ $Y2=0
r134 36 54 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.785 $Y=0
+ $X2=8.51 $Y2=0
r135 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.785 $Y=0 $X2=8.87
+ $Y2=0
r136 35 57 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=8.955 $Y=0
+ $X2=9.43 $Y2=0
r137 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.955 $Y=0 $X2=8.87
+ $Y2=0
r138 33 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.845 $Y=0
+ $X2=7.59 $Y2=0
r139 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=0 $X2=7.93
+ $Y2=0
r140 32 54 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.015 $Y=0
+ $X2=8.51 $Y2=0
r141 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.015 $Y=0 $X2=7.93
+ $Y2=0
r142 30 48 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.905 $Y=0
+ $X2=6.67 $Y2=0
r143 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0 $X2=6.99
+ $Y2=0
r144 29 51 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.075 $Y=0
+ $X2=7.59 $Y2=0
r145 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.075 $Y=0 $X2=6.99
+ $Y2=0
r146 25 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.81 $Y=0.085
+ $X2=9.81 $Y2=0
r147 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.81 $Y=0.085
+ $X2=9.81 $Y2=0.39
r148 21 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0
r149 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.87 $Y=0.085
+ $X2=8.87 $Y2=0.39
r150 17 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r151 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.39
r152 13 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0
r153 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.99 $Y=0.085
+ $X2=6.99 $Y2=0.39
r154 4 27 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.625
+ $Y=0.235 $X2=9.81 $Y2=0.39
r155 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=8.735
+ $Y=0.235 $X2=8.87 $Y2=0.39
r156 2 19 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.93 $Y2=0.39
r157 1 15 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.855
+ $Y=0.235 $X2=6.99 $Y2=0.39
.ends

