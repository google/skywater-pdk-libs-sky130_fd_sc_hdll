* File: sky130_fd_sc_hdll__a21bo_1.pex.spice
* Created: Wed Sep  2 08:16:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%B1_N 1 2 3 5 6 8 11 13 14 15 16 22
r37 15 16 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16
+ $X2=0.22 $Y2=1.53
r38 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r39 14 15 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=0.22 $Y=0.85
+ $X2=0.22 $Y2=1.16
r40 13 14 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=0.51
+ $X2=0.22 $Y2=0.85
r41 11 22 145.524 $w=2.7e-07 $l=6.55e-07 $layer=POLY_cond $X=0.24 $Y=1.815
+ $X2=0.24 $Y2=1.16
r42 9 22 56.6543 $w=2.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=0.905
+ $X2=0.24 $Y2=1.16
r43 6 8 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.865 $Y=0.755
+ $X2=0.865 $Y2=0.445
r44 3 11 76.8187 $w=1.6e-07 $l=2.55e-07 $layer=POLY_cond $X=0.495 $Y=1.902
+ $X2=0.24 $Y2=1.902
r45 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r46 2 9 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.375 $Y=0.83
+ $X2=0.24 $Y2=0.905
r47 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.79 $Y=0.83
+ $X2=0.865 $Y2=0.755
r48 1 2 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.79 $Y=0.83
+ $X2=0.375 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%A_27_413# 1 2 7 9 11 14 16 19 23 26 32 35
c67 16 0 1.55807e-19 $X=1.54 $Y=1.297
r68 33 35 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=0.85 $Y=1.35
+ $X2=0.85 $Y2=1.285
r69 32 34 6.61431 $w=4.48e-07 $l=1.85e-07 $layer=LI1_cond $X=0.74 $Y=1.35
+ $X2=0.74 $Y2=1.165
r70 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.85
+ $Y=1.35 $X2=0.85 $Y2=1.35
r71 25 32 1.06318 $w=4.48e-07 $l=4e-08 $layer=LI1_cond $X=0.74 $Y=1.39 $X2=0.74
+ $Y2=1.35
r72 25 26 12.0937 $w=4.48e-07 $l=4.55e-07 $layer=LI1_cond $X=0.74 $Y=1.39
+ $X2=0.74 $Y2=1.845
r73 23 34 29.4285 $w=2.78e-07 $l=7.15e-07 $layer=LI1_cond $X=0.655 $Y=0.45
+ $X2=0.655 $Y2=1.165
r74 17 26 28.5591 $w=1.98e-07 $l=5.15e-07 $layer=LI1_cond $X=0.225 $Y=1.945
+ $X2=0.74 $Y2=1.945
r75 17 19 10.8042 $w=2.38e-07 $l=2.25e-07 $layer=LI1_cond $X=0.225 $Y=2.045
+ $X2=0.225 $Y2=2.27
r76 12 16 23.8791 $w=1.65e-07 $l=1.23871e-07 $layer=POLY_cond $X=1.565 $Y=1.185
+ $X2=1.54 $Y2=1.297
r77 12 14 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.565 $Y=1.185
+ $X2=1.565 $Y2=0.56
r78 9 16 23.8791 $w=1.65e-07 $l=1.13e-07 $layer=POLY_cond $X=1.54 $Y=1.41
+ $X2=1.54 $Y2=1.297
r79 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.54 $Y=1.41
+ $X2=1.54 $Y2=1.985
r80 8 35 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.985 $Y=1.285
+ $X2=0.85 $Y2=1.285
r81 7 16 2.60714 $w=2e-07 $l=1.0583e-07 $layer=POLY_cond $X=1.44 $Y=1.285
+ $X2=1.54 $Y2=1.297
r82 7 8 150.868 $w=2e-07 $l=4.55e-07 $layer=POLY_cond $X=1.44 $Y=1.285 $X2=0.985
+ $Y2=1.285
r83 2 19 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.27
r84 1 23 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.475
+ $Y=0.235 $X2=0.6 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%A1 1 3 4 6 7 8
c35 4 0 1.64481e-19 $X=2.01 $Y=1.41
r36 7 8 11.3708 $w=3.73e-07 $l=3.7e-07 $layer=LI1_cond $X=2.087 $Y=1.16
+ $X2=2.087 $Y2=1.53
r37 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.045
+ $Y=1.16 $X2=2.045 $Y2=1.16
r38 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.01 $Y=1.41
+ $X2=2.045 $Y2=1.16
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=1.41 $X2=2.01
+ $Y2=1.985
r40 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=2.045 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%A2 1 3 4 6 7 8
c30 4 0 1.04739e-19 $X=2.49 $Y=1.41
r31 7 8 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=2.575 $Y=1.16
+ $X2=2.575 $Y2=1.53
r32 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.16 $X2=2.53 $Y2=1.16
r33 4 12 51.0578 $w=2.59e-07 $l=2.67862e-07 $layer=POLY_cond $X=2.49 $Y=1.41
+ $X2=2.527 $Y2=1.16
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.49 $Y=1.41 $X2=2.49
+ $Y2=1.985
r35 1 12 39.1718 $w=2.59e-07 $l=1.93533e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.527 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.465 $Y=0.995
+ $X2=2.465 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%A_235_297# 1 2 7 9 10 12 15 20 21 25 30 33
c72 20 0 3.20288e-19 $X=1.595 $Y=1.045
c73 7 0 1.25047e-19 $X=3.485 $Y=1.41
r74 35 36 4.63806 $w=4.78e-07 $l=9.5e-08 $layer=LI1_cond $X=1.7 $Y=0.72 $X2=1.7
+ $Y2=0.815
r75 33 35 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.7 $Y=0.38 $X2=1.7
+ $Y2=0.72
r76 28 30 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=1.3 $Y=1.195
+ $X2=1.595 $Y2=1.195
r77 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.16 $X2=3.45 $Y2=1.16
r78 23 25 15.292 $w=2.58e-07 $l=3.45e-07 $layer=LI1_cond $X=3.415 $Y=0.815
+ $X2=3.415 $Y2=1.16
r79 22 35 6.21271 $w=1.9e-07 $l=2.4e-07 $layer=LI1_cond $X=1.94 $Y=0.72 $X2=1.7
+ $Y2=0.72
r80 21 23 7.03324 $w=1.9e-07 $l=1.71026e-07 $layer=LI1_cond $X=3.285 $Y=0.72
+ $X2=3.415 $Y2=0.815
r81 21 22 78.512 $w=1.88e-07 $l=1.345e-06 $layer=LI1_cond $X=3.285 $Y=0.72
+ $X2=1.94 $Y2=0.72
r82 20 30 1.35108 $w=2.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.595 $Y=1.045
+ $X2=1.595 $Y2=1.195
r83 20 36 9.81711 $w=2.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.595 $Y=1.045
+ $X2=1.595 $Y2=0.815
r84 15 17 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.3 $Y=1.63 $X2=1.3
+ $Y2=2.31
r85 13 28 0.126616 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=1.3 $Y=1.345 $X2=1.3
+ $Y2=1.195
r86 13 15 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=1.3 $Y=1.345
+ $X2=1.3 $Y2=1.63
r87 10 26 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.45 $Y2=1.16
r88 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r89 7 26 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.45 $Y2=1.16
r90 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.985
r91 2 17 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.485 $X2=1.3 $Y2=2.31
r92 2 15 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.485 $X2=1.3 $Y2=1.63
r93 1 33 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.64
+ $Y=0.235 $X2=1.775 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%VPWR 1 2 3 12 16 20 25 26 27 29 34 44 45
+ 48 51
r61 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r63 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r64 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r65 42 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r67 39 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.225 $Y2=2.72
r68 39 41 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.415 $Y=2.72
+ $X2=2.99 $Y2=2.72
r69 38 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r70 38 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 37 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 35 48 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.915 $Y=2.72 $X2=0.715
+ $Y2=2.72
r73 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 34 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=2.225 $Y2=2.72
r75 34 37 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 29 48 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.515 $Y=2.72 $X2=0.715
+ $Y2=2.72
r77 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 27 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 25 41 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 25 26 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.075 $Y=2.72
+ $X2=3.217 $Y2=2.72
r82 24 44 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.36 $Y=2.72
+ $X2=3.91 $Y2=2.72
r83 24 26 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.36 $Y=2.72
+ $X2=3.217 $Y2=2.72
r84 20 23 27.4969 $w=2.83e-07 $l=6.8e-07 $layer=LI1_cond $X=3.217 $Y=1.66
+ $X2=3.217 $Y2=2.34
r85 18 26 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.217 $Y=2.635
+ $X2=3.217 $Y2=2.72
r86 18 23 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=3.217 $Y=2.635
+ $X2=3.217 $Y2=2.34
r87 14 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.72
r88 14 16 11.9793 $w=3.78e-07 $l=3.95e-07 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.24
r89 10 48 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r90 10 12 8.49927 $w=3.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.34
r91 3 23 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=1.485 $X2=3.25 $Y2=2.34
r92 3 20 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=3.125
+ $Y=1.485 $X2=3.25 $Y2=1.66
r93 2 16 600 $w=1.7e-07 $l=8.26604e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.25 $Y2=2.24
r94 1 12 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%A_326_297# 1 2 9 14 16
c20 16 0 1.04739e-19 $X=2.725 $Y=1.95
r21 10 14 3.24051 $w=2e-07 $l=9e-08 $layer=LI1_cond $X=1.865 $Y=1.885 $X2=1.775
+ $Y2=1.885
r22 9 16 3.15876 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=1.885 $X2=2.725
+ $Y2=1.885
r23 9 10 42.9773 $w=1.98e-07 $l=7.75e-07 $layer=LI1_cond $X=2.64 $Y=1.885
+ $X2=1.865 $Y2=1.885
r24 2 16 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.485 $X2=2.725 $Y2=1.95
r25 1 14 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.63
+ $Y=1.485 $X2=1.775 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%X 1 2 7 8 9 10 11 12
r13 11 12 16.8751 $w=2.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.855 $Y=1.8
+ $X2=3.855 $Y2=2.21
r14 10 11 11.1128 $w=2.78e-07 $l=2.7e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=3.855 $Y2=1.8
r15 9 10 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.855 $Y=1.19
+ $X2=3.855 $Y2=1.53
r16 8 9 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.855 $Y=0.85 $X2=3.855
+ $Y2=1.19
r17 7 8 13.994 $w=2.78e-07 $l=3.4e-07 $layer=LI1_cond $X=3.855 $Y=0.51 $X2=3.855
+ $Y2=0.85
r18 2 11 300 $w=1.7e-07 $l=4.25588e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.485 $X2=3.835 $Y2=1.8
r19 1 7 182 $w=1.7e-07 $l=4.42691e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.835 $Y2=0.57
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_1%VGND 1 2 9 13 15 30 31 34 39 42
c46 42 0 1.25047e-19 $X=3.35 $Y=0.185
r47 41 42 10.3217 $w=5.38e-07 $l=1.9e-07 $layer=LI1_cond $X=3.16 $Y=0.185
+ $X2=3.35 $Y2=0.185
r48 37 41 3.76543 $w=5.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.99 $Y=0.185
+ $X2=3.16 $Y2=0.185
r49 37 39 14.3086 $w=5.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.99 $Y=0.185
+ $X2=2.62 $Y2=0.185
r50 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r51 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 31 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r53 30 42 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=3.35
+ $Y2=0
r54 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r55 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r56 26 39 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.62
+ $Y2=0
r57 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r58 24 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r59 24 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r60 23 26 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r61 23 24 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r62 21 34 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.167
+ $Y2=0
r63 21 23 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.29 $Y=0 $X2=1.61
+ $Y2=0
r64 18 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r65 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r66 15 34 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.167
+ $Y2=0
r67 15 17 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.69
+ $Y2=0
r68 13 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 9 11 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=0.36
+ $X2=1.167 $Y2=0.7
r70 7 34 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=1.167 $Y=0.085
+ $X2=1.167 $Y2=0
r71 7 9 12.9356 $w=2.43e-07 $l=2.75e-07 $layer=LI1_cond $X=1.167 $Y=0.085
+ $X2=1.167 $Y2=0.36
r72 2 41 91 $w=1.7e-07 $l=6.79632e-07 $layer=licon1_NDIFF $count=2 $X=2.54
+ $Y=0.235 $X2=3.16 $Y2=0.36
r73 1 11 182 $w=1.7e-07 $l=5.82623e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.235 $X2=1.205 $Y2=0.7
r74 1 9 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.94
+ $Y=0.235 $X2=1.205 $Y2=0.36
.ends

