* File: sky130_fd_sc_hdll__a31o_2.pex.spice
* Created: Thu Aug 27 18:55:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A31O_2%A_79_21# 1 2 7 9 10 12 13 15 16 18 20 21 22
+ 25 27 31 35 38 42
c90 35 0 1.01582e-19 $X=0.68 $Y=1.16
c91 25 0 1.11805e-19 $X=2.87 $Y=0.42
c92 20 0 1.51137e-19 $X=0.6 $Y=1.495
r93 42 43 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r94 39 40 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r95 36 42 36.15 $w=3.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.68 $Y=1.202
+ $X2=0.965 $Y2=1.202
r96 36 40 23.4658 $w=3.8e-07 $l=1.85e-07 $layer=POLY_cond $X=0.68 $Y=1.202
+ $X2=0.495 $Y2=1.202
r97 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.68
+ $Y=1.16 $X2=0.68 $Y2=1.16
r98 29 31 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.26 $Y=1.665
+ $X2=3.26 $Y2=1.96
r99 28 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.955 $Y=1.58
+ $X2=2.87 $Y2=1.58
r100 27 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.175 $Y=1.58
+ $X2=3.26 $Y2=1.665
r101 27 28 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.175 $Y=1.58
+ $X2=2.955 $Y2=1.58
r102 23 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.87 $Y=1.495
+ $X2=2.87 $Y2=1.58
r103 23 25 70.1337 $w=1.68e-07 $l=1.075e-06 $layer=LI1_cond $X=2.87 $Y=1.495
+ $X2=2.87 $Y2=0.42
r104 21 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.785 $Y=1.58
+ $X2=2.87 $Y2=1.58
r105 21 22 137.005 $w=1.68e-07 $l=2.1e-06 $layer=LI1_cond $X=2.785 $Y=1.58
+ $X2=0.685 $Y2=1.58
r106 20 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=1.495
+ $X2=0.685 $Y2=1.58
r107 19 35 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.6 $Y=1.245
+ $X2=0.6 $Y2=1.16
r108 19 20 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.6 $Y=1.245
+ $X2=0.6 $Y2=1.495
r109 16 43 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r110 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r111 13 42 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r112 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r113 10 40 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r114 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r115 7 39 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r116 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
r117 2 31 300 $w=1.7e-07 $l=5.68331e-07 $layer=licon1_PDIFF $count=2 $X=3.055
+ $Y=1.485 $X2=3.26 $Y2=1.96
r118 1 25 182 $w=1.7e-07 $l=4.68455e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.87 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%A3 1 3 4 6 7 8
c34 1 0 1.46885e-19 $X=1.435 $Y=1.41
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r36 8 13 0.828054 $w=4.42e-07 $l=3e-08 $layer=LI1_cond $X=1.287 $Y=1.19
+ $X2=1.287 $Y2=1.16
r37 7 13 8.55656 $w=4.42e-07 $l=3.1e-07 $layer=LI1_cond $X=1.287 $Y=0.85
+ $X2=1.287 $Y2=1.16
r38 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.435 $Y2=1.16
r39 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995 $X2=1.46
+ $Y2=0.56
r40 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.16
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%A2 1 3 4 6 7
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.16 $X2=1.99 $Y2=1.16
r31 7 11 29.9635 $w=2.48e-07 $l=6.5e-07 $layer=LI1_cond $X=2.03 $Y=0.51 $X2=2.03
+ $Y2=1.16
r32 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.965 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r34 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.965 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995 $X2=1.88
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%A1 1 3 4 6 7
r30 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.16 $X2=2.47 $Y2=1.16
r31 7 11 32.569 $w=2.28e-07 $l=6.5e-07 $layer=LI1_cond $X=2.5 $Y=0.51 $X2=2.5
+ $Y2=1.16
r32 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.495 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.435 $Y=1.41
+ $X2=2.435 $Y2=1.985
r34 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.41 $Y=0.995
+ $X2=2.495 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.41 $Y=0.995 $X2=2.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%B1 1 3 4 6 7 8 12
r31 12 14 26.7778 $w=3.6e-07 $l=2e-07 $layer=POLY_cond $X=3.08 $Y=1.202 $X2=3.28
+ $Y2=1.202
r32 11 12 15.3972 $w=3.6e-07 $l=1.15e-07 $layer=POLY_cond $X=2.965 $Y=1.202
+ $X2=3.08 $Y2=1.202
r33 7 8 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=3.365 $Y=1.16
+ $X2=3.365 $Y2=0.85
r34 7 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.28
+ $Y=1.16 $X2=3.28 $Y2=1.16
r35 4 12 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.08 $Y=0.995
+ $X2=3.08 $Y2=1.202
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.08 $Y=0.995 $X2=3.08
+ $Y2=0.56
r37 1 11 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.202
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%VPWR 1 2 3 10 12 16 18 22 24 26 36 37 43 46
r61 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r62 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 33 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 31 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.18 $Y2=2.72
r70 31 33 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 30 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 27 40 3.98448 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.192 $Y2=2.72
r74 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.385 $Y=2.72
+ $X2=0.69 $Y2=2.72
r75 26 43 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=1.135 $Y2=2.72
r76 26 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=2.72
+ $X2=0.69 $Y2=2.72
r77 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 24 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r79 20 46 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.635
+ $X2=2.18 $Y2=2.72
r80 20 22 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=2.18 $Y=2.635
+ $X2=2.18 $Y2=2.26
r81 19 43 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.135 $Y2=2.72
r82 18 46 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.18 $Y2=2.72
r83 18 19 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.285 $Y2=2.72
r84 14 43 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=2.635
+ $X2=1.135 $Y2=2.72
r85 14 16 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=1.135 $Y=2.635
+ $X2=1.135 $Y2=2
r86 10 40 3.15868 $w=2.5e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.192 $Y2=2.72
r87 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r88 3 22 600 $w=1.7e-07 $l=8.62554e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.18 $Y2=2.26
r89 2 16 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r90 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%X 1 2 7 9 13 17 19 20 21 22 29 30
c49 2 0 1.05833e-19 $X=0.585 $Y=1.485
r50 22 30 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.92
+ $X2=0.217 $Y2=1.835
r51 22 30 1.12985 $w=2.53e-07 $l=2.5e-08 $layer=LI1_cond $X=0.217 $Y=1.81
+ $X2=0.217 $Y2=1.835
r52 21 22 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=0.217 $Y=1.53
+ $X2=0.217 $Y2=1.81
r53 20 21 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=1.19
+ $X2=0.217 $Y2=1.53
r54 19 29 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=0.8
+ $X2=0.217 $Y2=0.885
r55 19 20 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=0.217 $Y=0.91
+ $X2=0.217 $Y2=1.19
r56 19 29 1.12985 $w=2.53e-07 $l=2.5e-08 $layer=LI1_cond $X=0.217 $Y=0.91
+ $X2=0.217 $Y2=0.885
r57 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=2.005
+ $X2=0.73 $Y2=2.3
r58 11 13 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.715
+ $X2=0.73 $Y2=0.42
r59 10 22 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.92
+ $X2=0.217 $Y2=1.92
r60 9 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=1.92
+ $X2=0.73 $Y2=2.005
r61 9 10 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=1.92 $X2=0.345
+ $Y2=1.92
r62 8 19 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.8
+ $X2=0.217 $Y2=0.8
r63 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.645 $Y=0.8
+ $X2=0.73 $Y2=0.715
r64 7 8 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=0.8 $X2=0.345
+ $Y2=0.8
r65 2 17 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
r66 1 13 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%A_305_297# 1 2 7 9 11 13 15
c30 2 0 1.11805e-19 $X=2.525 $Y=1.485
r31 13 20 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=2.005
+ $X2=2.74 $Y2=1.92
r32 13 15 9.47977 $w=3.08e-07 $l=2.55e-07 $layer=LI1_cond $X=2.74 $Y=2.005
+ $X2=2.74 $Y2=2.26
r33 12 18 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.755 $Y=1.92
+ $X2=1.605 $Y2=1.92
r34 11 20 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=2.585 $Y=1.92
+ $X2=2.74 $Y2=1.92
r35 11 12 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=2.585 $Y=1.92
+ $X2=1.755 $Y2=1.92
r36 7 18 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.005 $X2=1.605
+ $Y2=1.92
r37 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.605 $Y=2.005
+ $X2=1.605 $Y2=2.26
r38 2 20 600 $w=1.7e-07 $l=5.27636e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.73 $Y2=1.92
r39 2 15 600 $w=1.7e-07 $l=8.71493e-07 $layer=licon1_PDIFF $count=1 $X=2.525
+ $Y=1.485 $X2=2.73 $Y2=2.26
r40 1 18 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.92
r41 1 9 600 $w=1.7e-07 $l=8.44393e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.26
.ends

.subckt PM_SKY130_FD_SC_HDLL__A31O_2%VGND 1 2 3 10 12 14 16 18 20 25 38 45
r56 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r57 38 41 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.195 $Y=0 $X2=1.195
+ $Y2=0.38
r58 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r59 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r60 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r61 29 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r62 29 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r63 28 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r64 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r65 26 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.195
+ $Y2=0
r66 26 28 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.61
+ $Y2=0
r67 25 44 4.22148 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=3.427
+ $Y2=0
r68 25 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.175 $Y=0 $X2=2.99
+ $Y2=0
r69 24 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r70 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r71 21 34 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r72 21 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r73 20 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.195
+ $Y2=0
r74 20 23 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.69
+ $Y2=0
r75 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r76 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r77 14 44 3.21636 $w=2.9e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.32 $Y=0.085
+ $X2=3.427 $Y2=0
r78 14 16 12.5179 $w=2.88e-07 $l=3.15e-07 $layer=LI1_cond $X=3.32 $Y=0.085
+ $X2=3.32 $Y2=0.4
r79 10 34 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r80 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r81 3 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.235 $X2=3.29 $Y2=0.4
r82 2 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r83 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

