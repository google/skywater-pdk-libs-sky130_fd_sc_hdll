* File: sky130_fd_sc_hdll__o2bb2ai_2.pxi.spice
* Created: Wed Sep  2 08:46:28 2020
* 
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A1_N N_A1_N_c_88_n N_A1_N_M1000_g
+ N_A1_N_c_89_n N_A1_N_M1004_g N_A1_N_c_90_n N_A1_N_M1006_g N_A1_N_c_91_n
+ N_A1_N_M1003_g N_A1_N_c_96_n N_A1_N_c_92_n A1_N A1_N N_A1_N_c_93_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A1_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A2_N N_A2_N_c_158_n N_A2_N_M1001_g
+ N_A2_N_c_162_n N_A2_N_M1007_g N_A2_N_c_163_n N_A2_N_M1015_g N_A2_N_c_159_n
+ N_A2_N_M1011_g A2_N N_A2_N_c_161_n PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A2_N
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_121_297# N_A_121_297#_M1001_d
+ N_A_121_297#_M1000_d N_A_121_297#_M1015_d N_A_121_297#_c_208_n
+ N_A_121_297#_M1009_g N_A_121_297#_c_202_n N_A_121_297#_M1010_g
+ N_A_121_297#_c_209_n N_A_121_297#_M1016_g N_A_121_297#_c_203_n
+ N_A_121_297#_M1012_g N_A_121_297#_c_216_n N_A_121_297#_c_204_n
+ N_A_121_297#_c_205_n N_A_121_297#_c_211_n N_A_121_297#_c_228_n
+ N_A_121_297#_c_206_n N_A_121_297#_c_207_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_121_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B1 N_B1_c_297_n N_B1_M1014_g N_B1_c_298_n
+ N_B1_M1013_g N_B1_c_299_n N_B1_M1018_g N_B1_c_300_n N_B1_M1019_g N_B1_c_305_n
+ N_B1_c_301_n B1 PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B2 N_B2_c_371_n N_B2_M1002_g N_B2_c_375_n
+ N_B2_M1005_g N_B2_c_376_n N_B2_M1008_g N_B2_c_372_n N_B2_M1017_g B2
+ N_B2_c_374_n B2 PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B2
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VPWR N_VPWR_M1000_s N_VPWR_M1007_s
+ N_VPWR_M1003_s N_VPWR_M1016_d N_VPWR_M1019_s N_VPWR_c_419_n N_VPWR_c_420_n
+ N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n
+ N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n VPWR N_VPWR_c_429_n
+ N_VPWR_c_418_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%Y N_Y_M1010_s N_Y_M1009_s N_Y_M1005_s
+ N_Y_c_496_n N_Y_c_504_n N_Y_c_516_n N_Y_c_497_n N_Y_c_508_n N_Y_c_521_n Y
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_788_297# N_A_788_297#_M1014_d
+ N_A_788_297#_M1008_d N_A_788_297#_c_547_n N_A_788_297#_c_546_n
+ N_A_788_297#_c_553_n PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_788_297#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_M1013_s N_VGND_M1017_s N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n
+ N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n N_VGND_c_567_n
+ N_VGND_c_568_n VGND N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n
+ N_VGND_c_572_n PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VGND
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_123_47# N_A_123_47#_M1004_s
+ N_A_123_47#_M1011_s N_A_123_47#_c_643_n N_A_123_47#_c_642_n
+ N_A_123_47#_c_647_n PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_123_47#
x_PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_503_47# N_A_503_47#_M1010_d
+ N_A_503_47#_M1012_d N_A_503_47#_M1002_d N_A_503_47#_M1018_d
+ N_A_503_47#_c_670_n N_A_503_47#_c_704_n N_A_503_47#_c_664_n
+ N_A_503_47#_c_665_n N_A_503_47#_c_681_n N_A_503_47#_c_666_n
+ N_A_503_47#_c_667_n N_A_503_47#_c_668_n N_A_503_47#_c_669_n
+ PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_503_47#
cc_1 VNB N_A1_N_c_88_n 0.0297694f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_2 VNB N_A1_N_c_89_n 0.0218895f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_3 VNB N_A1_N_c_90_n 0.0197773f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.995
cc_4 VNB N_A1_N_c_91_n 0.021967f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.41
cc_5 VNB N_A1_N_c_92_n 0.00429224f $X=-0.19 $Y=-0.24 $X2=1.97 $Y2=1.16
cc_6 VNB N_A1_N_c_93_n 0.0175715f $X=-0.19 $Y=-0.24 $X2=0.675 $Y2=1.345
cc_7 VNB N_A2_N_c_158_n 0.0170715f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_8 VNB N_A2_N_c_159_n 0.0170327f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.41
cc_9 VNB A2_N 0.00225501f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.53
cc_10 VNB N_A2_N_c_161_n 0.037357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_121_297#_c_202_n 0.0195832f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.53
cc_12 VNB N_A_121_297#_c_203_n 0.0174298f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.53
cc_13 VNB N_A_121_297#_c_204_n 0.0123094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_121_297#_c_205_n 0.0120923f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.19
cc_15 VNB N_A_121_297#_c_206_n 0.00259728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_121_297#_c_207_n 0.0554826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B1_c_297_n 0.0202739f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_18 VNB N_B1_c_298_n 0.0169765f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_19 VNB N_B1_c_299_n 0.021688f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.995
cc_20 VNB N_B1_c_300_n 0.0348333f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.41
cc_21 VNB N_B1_c_301_n 0.00421058f $X=-0.19 $Y=-0.24 $X2=1.97 $Y2=1.16
cc_22 VNB B1 0.00198218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B2_c_371_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_24 VNB N_B2_c_372_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.41
cc_25 VNB B2 0.00158585f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.53
cc_26 VNB N_B2_c_374_n 0.0372287f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_418_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_496_n 0.00101052f $X=-0.19 $Y=-0.24 $X2=1.935 $Y2=1.985
cc_29 VNB N_Y_c_497_n 0.0017908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_560_n 0.0116911f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.53
cc_31 VNB N_VGND_c_561_n 0.00670844f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.16
cc_32 VNB N_VGND_c_562_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.53
cc_33 VNB N_VGND_c_563_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_34 VNB N_VGND_c_564_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.345
cc_35 VNB N_VGND_c_565_n 0.0427121f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.19
cc_36 VNB N_VGND_c_566_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_567_n 0.0193035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_568_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_569_n 0.0411697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_570_n 0.0255062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_571_n 0.309249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_572_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_123_47#_c_642_n 0.00311909f $X=-0.19 $Y=-0.24 $X2=1.91 $Y2=0.56
cc_44 VNB N_A_503_47#_c_664_n 0.00363741f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.53
cc_45 VNB N_A_503_47#_c_665_n 0.00735292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_503_47#_c_666_n 0.0200032f $X=-0.19 $Y=-0.24 $X2=0.48 $Y2=1.16
cc_47 VNB N_A_503_47#_c_667_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.345
cc_48 VNB N_A_503_47#_c_668_n 0.0036207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_503_47#_c_669_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_A1_N_c_88_n 0.0286525f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_51 VPB N_A1_N_c_91_n 0.0285361f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.41
cc_52 VPB N_A1_N_c_96_n 0.00823075f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.53
cc_53 VPB N_A1_N_c_92_n 0.00298462f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.16
cc_54 VPB N_A1_N_c_93_n 0.0165886f $X=-0.19 $Y=1.305 $X2=0.675 $Y2=1.345
cc_55 VPB N_A2_N_c_162_n 0.0159776f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_56 VPB N_A2_N_c_163_n 0.0160572f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.995
cc_57 VPB N_A2_N_c_161_n 0.0194393f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_121_297#_c_208_n 0.0190428f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.41
cc_59 VPB N_A_121_297#_c_209_n 0.0159231f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.16
cc_60 VPB N_A_121_297#_c_205_n 0.00907516f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.19
cc_61 VPB N_A_121_297#_c_211_n 0.00240692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_121_297#_c_207_n 0.0304684f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B1_c_297_n 0.0237318f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_64 VPB N_B1_c_300_n 0.0306194f $X=-0.19 $Y=1.305 $X2=1.935 $Y2=1.41
cc_65 VPB N_B1_c_305_n 0.0098044f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.53
cc_66 VPB N_B1_c_301_n 0.00273476f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.16
cc_67 VPB B1 0.00596434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_B2_c_375_n 0.0159964f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_69 VPB N_B2_c_376_n 0.0159786f $X=-0.19 $Y=1.305 $X2=1.91 $Y2=0.995
cc_70 VPB N_B2_c_374_n 0.0193751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_419_n 0.0117686f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.16
cc_72 VPB N_VPWR_c_420_n 0.00518019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_421_n 0.018941f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_422_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.48 $Y2=1.16
cc_75 VPB N_VPWR_c_423_n 0.0053627f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.19
cc_76 VPB N_VPWR_c_424_n 0.0049401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_425_n 0.0198475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_426_n 0.00545601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_427_n 0.0417635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_428_n 0.00391723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_429_n 0.0135992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_418_n 0.0549979f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_431_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_432_n 0.0194879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_433_n 0.0208899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Y_c_497_n 3.62521e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB Y 8.24654e-19 $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.345
cc_88 N_A1_N_c_89_n N_A2_N_c_158_n 0.0164857f $X=0.54 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A1_N_c_88_n N_A2_N_c_162_n 0.022609f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A1_N_c_96_n N_A2_N_c_162_n 0.0118239f $X=1.765 $Y=1.53 $X2=0 $Y2=0
cc_91 N_A1_N_c_93_n N_A2_N_c_162_n 8.76396e-19 $X=0.675 $Y=1.345 $X2=0 $Y2=0
cc_92 N_A1_N_c_91_n N_A2_N_c_163_n 0.0346822f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A1_N_c_96_n N_A2_N_c_163_n 0.0119735f $X=1.765 $Y=1.53 $X2=0 $Y2=0
cc_94 N_A1_N_c_92_n N_A2_N_c_163_n 9.75029e-19 $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A1_N_c_90_n N_A2_N_c_159_n 0.0228293f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A1_N_c_88_n A2_N 6.68904e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A1_N_c_91_n A2_N 2.09039e-19 $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A1_N_c_96_n A2_N 0.0463839f $X=1.765 $Y=1.53 $X2=0 $Y2=0
cc_99 N_A1_N_c_92_n A2_N 0.012001f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A1_N_c_93_n A2_N 0.0182871f $X=0.675 $Y=1.345 $X2=0 $Y2=0
cc_101 N_A1_N_c_88_n N_A2_N_c_161_n 0.0164857f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A1_N_c_91_n N_A2_N_c_161_n 0.0228293f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A1_N_c_96_n N_A2_N_c_161_n 0.00803891f $X=1.765 $Y=1.53 $X2=0 $Y2=0
cc_104 N_A1_N_c_92_n N_A2_N_c_161_n 0.00482702f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A1_N_c_93_n N_A2_N_c_161_n 0.00417633f $X=0.675 $Y=1.345 $X2=0 $Y2=0
cc_106 N_A1_N_c_96_n N_A_121_297#_M1000_d 0.00172209f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_107 N_A1_N_c_96_n N_A_121_297#_M1015_d 0.00204196f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_108 N_A1_N_c_92_n N_A_121_297#_M1015_d 5.59275e-19 $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_109 N_A1_N_c_91_n N_A_121_297#_c_216_n 0.0142628f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_110 N_A1_N_c_96_n N_A_121_297#_c_216_n 0.0491691f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_111 N_A1_N_c_92_n N_A_121_297#_c_216_n 0.0202038f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A1_N_c_90_n N_A_121_297#_c_204_n 0.0142809f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_113 N_A1_N_c_91_n N_A_121_297#_c_204_n 0.00314385f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_114 N_A1_N_c_96_n N_A_121_297#_c_204_n 0.00861691f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_115 N_A1_N_c_92_n N_A_121_297#_c_204_n 0.0296937f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A1_N_c_90_n N_A_121_297#_c_205_n 0.00259035f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_117 N_A1_N_c_91_n N_A_121_297#_c_205_n 0.00287586f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A1_N_c_92_n N_A_121_297#_c_205_n 0.0214817f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A1_N_c_91_n N_A_121_297#_c_211_n 0.00674247f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A1_N_c_92_n N_A_121_297#_c_211_n 0.0228362f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A1_N_c_93_n N_A_121_297#_c_228_n 0.014372f $X=0.675 $Y=1.345 $X2=0
+ $Y2=0
cc_122 N_A1_N_c_91_n N_A_121_297#_c_207_n 0.0101735f $X=1.935 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A1_N_c_92_n N_A_121_297#_c_207_n 6.55835e-19 $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A1_N_c_93_n N_VPWR_M1000_s 0.00380009f $X=0.675 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_125 N_A1_N_c_96_n N_VPWR_M1007_s 0.00187547f $X=1.765 $Y=1.53 $X2=0 $Y2=0
cc_126 N_A1_N_c_92_n N_VPWR_M1003_s 0.001994f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A1_N_c_88_n N_VPWR_c_420_n 0.00492139f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A1_N_c_93_n N_VPWR_c_420_n 0.0183449f $X=0.675 $Y=1.345 $X2=0 $Y2=0
cc_129 N_A1_N_c_88_n N_VPWR_c_421_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A1_N_c_88_n N_VPWR_c_418_n 0.0133765f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_N_c_91_n N_VPWR_c_418_n 0.00825746f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A1_N_c_91_n N_VPWR_c_432_n 0.0053025f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A1_N_c_91_n N_VPWR_c_433_n 0.0052211f $X=1.935 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_N_c_88_n N_VGND_c_561_n 4.85489e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_N_c_89_n N_VGND_c_561_n 0.00695086f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A1_N_c_93_n N_VGND_c_561_n 0.0147074f $X=0.675 $Y=1.345 $X2=0 $Y2=0
cc_137 N_A1_N_c_90_n N_VGND_c_562_n 0.00438629f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A1_N_c_89_n N_VGND_c_569_n 0.00469405f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_N_c_90_n N_VGND_c_569_n 0.00428555f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_N_c_89_n N_VGND_c_571_n 0.00879116f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_N_c_90_n N_VGND_c_571_n 0.00716151f $X=1.91 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_N_c_89_n N_A_123_47#_c_643_n 0.00328522f $X=0.54 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A1_N_c_89_n N_A_123_47#_c_642_n 0.00725592f $X=0.54 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A1_N_c_96_n N_A_123_47#_c_642_n 0.00584717f $X=1.765 $Y=1.53 $X2=0
+ $Y2=0
cc_145 N_A1_N_c_93_n N_A_123_47#_c_642_n 0.0114026f $X=0.675 $Y=1.345 $X2=0
+ $Y2=0
cc_146 N_A1_N_c_90_n N_A_123_47#_c_647_n 0.00230812f $X=1.91 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A2_N_c_162_n N_A_121_297#_c_216_n 0.0123176f $X=0.985 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A2_N_c_163_n N_A_121_297#_c_216_n 0.0123176f $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A2_N_c_159_n N_A_121_297#_c_204_n 0.0100355f $X=1.48 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A2_N_c_158_n N_A_121_297#_c_206_n 0.00387597f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_151 A2_N N_A_121_297#_c_206_n 0.0363061f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A2_N_c_161_n N_A_121_297#_c_206_n 0.0047334f $X=1.455 $Y=1.202 $X2=0
+ $Y2=0
cc_153 N_A2_N_c_162_n N_VPWR_c_421_n 0.0053025f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_N_c_162_n N_VPWR_c_422_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A2_N_c_163_n N_VPWR_c_422_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A2_N_c_162_n N_VPWR_c_418_n 0.00693014f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A2_N_c_163_n N_VPWR_c_418_n 0.00700267f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_N_c_163_n N_VPWR_c_432_n 0.0053025f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A2_N_c_158_n N_VGND_c_569_n 0.00368123f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_N_c_159_n N_VGND_c_569_n 0.00368123f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_N_c_158_n N_VGND_c_571_n 0.00552518f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_N_c_159_n N_VGND_c_571_n 0.00554968f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_N_c_158_n N_A_123_47#_c_647_n 0.0101308f $X=0.96 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A2_N_c_159_n N_A_123_47#_c_647_n 0.00897812f $X=1.48 $Y=0.995 $X2=0
+ $Y2=0
cc_165 A2_N N_A_123_47#_c_647_n 0.00353291f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_166 N_A_121_297#_c_209_n N_B1_c_297_n 0.0315042f $X=3.345 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_121_297#_c_207_n N_B1_c_297_n 0.0228211f $X=3.345 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_121_297#_c_203_n N_B1_c_298_n 0.017558f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_121_297#_c_209_n N_B1_c_301_n 7.28691e-19 $X=3.345 $Y=1.41 $X2=0
+ $Y2=0
cc_170 N_A_121_297#_c_207_n N_B1_c_301_n 0.00115234f $X=3.345 $Y=1.202 $X2=0
+ $Y2=0
cc_171 N_A_121_297#_c_216_n N_VPWR_M1007_s 0.00348321f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_172 N_A_121_297#_c_216_n N_VPWR_M1003_s 0.0165797f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_173 N_A_121_297#_c_211_n N_VPWR_M1003_s 0.00969652f $X=2.4 $Y=1.785 $X2=0
+ $Y2=0
cc_174 N_A_121_297#_c_216_n N_VPWR_c_421_n 0.00254499f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_175 N_A_121_297#_c_228_n N_VPWR_c_421_n 0.0149311f $X=0.75 $Y=1.96 $X2=0
+ $Y2=0
cc_176 N_A_121_297#_c_216_n N_VPWR_c_422_n 0.0139299f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_177 N_A_121_297#_c_209_n N_VPWR_c_423_n 0.0031043f $X=3.345 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A_121_297#_c_208_n N_VPWR_c_425_n 0.00597712f $X=2.875 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_121_297#_c_209_n N_VPWR_c_425_n 0.00702461f $X=3.345 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_121_297#_M1000_d N_VPWR_c_418_n 0.00310186f $X=0.605 $Y=1.485 $X2=0
+ $Y2=0
cc_181 N_A_121_297#_M1015_d N_VPWR_c_418_n 0.00403478f $X=1.545 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_A_121_297#_c_208_n N_VPWR_c_418_n 0.0112745f $X=2.875 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_121_297#_c_209_n N_VPWR_c_418_n 0.00703789f $X=3.345 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_121_297#_c_216_n N_VPWR_c_418_n 0.0232697f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_185 N_A_121_297#_c_228_n N_VPWR_c_418_n 0.00955092f $X=0.75 $Y=1.96 $X2=0
+ $Y2=0
cc_186 N_A_121_297#_c_216_n N_VPWR_c_432_n 0.00809105f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_187 N_A_121_297#_c_208_n N_VPWR_c_433_n 0.0064896f $X=2.875 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_121_297#_c_216_n N_VPWR_c_433_n 0.0329633f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_189 N_A_121_297#_c_202_n N_Y_c_496_n 0.0117243f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_121_297#_c_203_n N_Y_c_496_n 0.00285271f $X=3.37 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_121_297#_c_205_n N_Y_c_496_n 0.0376426f $X=2.4 $Y=1.325 $X2=0 $Y2=0
cc_192 N_A_121_297#_c_207_n N_Y_c_496_n 0.00815911f $X=3.345 $Y=1.202 $X2=0
+ $Y2=0
cc_193 N_A_121_297#_c_208_n N_Y_c_504_n 0.0136564f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_121_297#_c_216_n N_Y_c_504_n 4.01087e-19 $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_195 N_A_121_297#_c_211_n N_Y_c_497_n 0.0180917f $X=2.4 $Y=1.785 $X2=0 $Y2=0
cc_196 N_A_121_297#_c_207_n N_Y_c_497_n 0.0311337f $X=3.345 $Y=1.202 $X2=0 $Y2=0
cc_197 N_A_121_297#_c_208_n N_Y_c_508_n 0.00350666f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_121_297#_c_209_n N_Y_c_508_n 0.00967792f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_121_297#_c_216_n N_Y_c_508_n 0.00750299f $X=2.315 $Y=1.875 $X2=0
+ $Y2=0
cc_200 N_A_121_297#_c_208_n Y 0.00857296f $X=2.875 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_121_297#_c_209_n Y 0.00900172f $X=3.345 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_121_297#_c_207_n Y 0.00402829f $X=3.345 $Y=1.202 $X2=0 $Y2=0
cc_203 N_A_121_297#_c_204_n N_VGND_M1006_d 0.00315681f $X=2.315 $Y=0.815 $X2=0
+ $Y2=0
cc_204 N_A_121_297#_c_202_n N_VGND_c_562_n 0.00179926f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_121_297#_c_204_n N_VGND_c_562_n 0.0127273f $X=2.315 $Y=0.815 $X2=0
+ $Y2=0
cc_206 N_A_121_297#_c_202_n N_VGND_c_565_n 0.00357877f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_121_297#_c_203_n N_VGND_c_565_n 0.00357877f $X=3.37 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A_121_297#_c_204_n N_VGND_c_565_n 0.00163764f $X=2.315 $Y=0.815 $X2=0
+ $Y2=0
cc_209 N_A_121_297#_c_205_n N_VGND_c_565_n 0.0027238f $X=2.4 $Y=1.325 $X2=0
+ $Y2=0
cc_210 N_A_121_297#_c_204_n N_VGND_c_569_n 0.00212702f $X=2.315 $Y=0.815 $X2=0
+ $Y2=0
cc_211 N_A_121_297#_M1001_d N_VGND_c_571_n 0.00301822f $X=1.035 $Y=0.235 $X2=0
+ $Y2=0
cc_212 N_A_121_297#_c_202_n N_VGND_c_571_n 0.00668309f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_121_297#_c_203_n N_VGND_c_571_n 0.00557903f $X=3.37 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_121_297#_c_204_n N_VGND_c_571_n 0.00871706f $X=2.315 $Y=0.815 $X2=0
+ $Y2=0
cc_215 N_A_121_297#_c_205_n N_VGND_c_571_n 0.00452669f $X=2.4 $Y=1.325 $X2=0
+ $Y2=0
cc_216 N_A_121_297#_c_204_n N_A_123_47#_M1011_s 0.00204044f $X=2.315 $Y=0.815
+ $X2=0 $Y2=0
cc_217 N_A_121_297#_c_206_n N_A_123_47#_c_642_n 0.0105775f $X=1.385 $Y=0.775
+ $X2=0 $Y2=0
cc_218 N_A_121_297#_M1001_d N_A_123_47#_c_647_n 0.00527949f $X=1.035 $Y=0.235
+ $X2=0 $Y2=0
cc_219 N_A_121_297#_c_204_n N_A_123_47#_c_647_n 0.0160411f $X=2.315 $Y=0.815
+ $X2=0 $Y2=0
cc_220 N_A_121_297#_c_206_n N_A_123_47#_c_647_n 0.0201898f $X=1.385 $Y=0.775
+ $X2=0 $Y2=0
cc_221 N_A_121_297#_c_202_n N_A_503_47#_c_670_n 0.0115292f $X=2.9 $Y=0.995 $X2=0
+ $Y2=0
cc_222 N_A_121_297#_c_203_n N_A_503_47#_c_670_n 0.0113611f $X=3.37 $Y=0.995
+ $X2=0 $Y2=0
cc_223 N_A_121_297#_c_207_n N_A_503_47#_c_670_n 0.00253348f $X=3.345 $Y=1.202
+ $X2=0 $Y2=0
cc_224 N_A_121_297#_c_205_n N_A_503_47#_c_668_n 0.00978984f $X=2.4 $Y=1.325
+ $X2=0 $Y2=0
cc_225 N_A_121_297#_c_207_n N_A_503_47#_c_668_n 0.00150611f $X=3.345 $Y=1.202
+ $X2=0 $Y2=0
cc_226 N_B1_c_298_n N_B2_c_371_n 0.0232181f $X=3.875 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_227 N_B1_c_297_n N_B2_c_375_n 0.0378352f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_228 N_B1_c_305_n N_B2_c_375_n 0.0116479f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_229 N_B1_c_301_n N_B2_c_375_n 0.00101886f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B1_c_300_n N_B2_c_376_n 0.0226184f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B1_c_305_n N_B2_c_376_n 0.0173214f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_232 B1 N_B2_c_376_n 7.35049e-19 $X=5.195 $Y=1.105 $X2=0 $Y2=0
cc_233 N_B1_c_299_n N_B2_c_372_n 0.0233179f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B1_c_297_n B2 2.04595e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B1_c_300_n B2 7.83557e-19 $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_236 N_B1_c_305_n B2 0.0451262f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_237 N_B1_c_301_n B2 0.0137935f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_238 B1 B2 0.0140899f $X=5.195 $Y=1.105 $X2=0 $Y2=0
cc_239 N_B1_c_297_n N_B2_c_374_n 0.0232181f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B1_c_300_n N_B2_c_374_n 0.0233179f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B1_c_305_n N_B2_c_374_n 0.00803891f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B1_c_301_n N_B2_c_374_n 0.00489731f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_243 B1 N_B2_c_374_n 0.00372544f $X=5.195 $Y=1.105 $X2=0 $Y2=0
cc_244 N_B1_c_301_n N_VPWR_M1016_d 0.00174439f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B1_c_305_n N_VPWR_M1019_s 0.00674339f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_246 N_B1_c_297_n N_VPWR_c_423_n 0.0031043f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B1_c_300_n N_VPWR_c_424_n 0.00840787f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B1_c_305_n N_VPWR_c_424_n 0.00373767f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_249 N_B1_c_297_n N_VPWR_c_427_n 0.00702461f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B1_c_300_n N_VPWR_c_427_n 0.00702461f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B1_c_297_n N_VPWR_c_418_n 0.00706607f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B1_c_300_n N_VPWR_c_418_n 0.013611f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B1_c_305_n N_Y_M1005_s 0.00187091f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_254 N_B1_c_297_n N_Y_c_496_n 3.82e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B1_c_297_n N_Y_c_516_n 0.0136916f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B1_c_305_n N_Y_c_516_n 0.0218268f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_257 N_B1_c_301_n N_Y_c_516_n 0.0209561f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_297_n N_Y_c_497_n 0.00115808f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B1_c_301_n N_Y_c_497_n 0.0388852f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_260 N_B1_c_305_n N_Y_c_521_n 0.0135474f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_261 N_B1_c_297_n Y 3.26911e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B1_c_305_n N_A_788_297#_M1014_d 0.00172342f $X=5.13 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_263 N_B1_c_301_n N_A_788_297#_M1014_d 7.76441e-19 $X=3.815 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_264 N_B1_c_305_n N_A_788_297#_M1008_d 0.00187091f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_265 N_B1_c_305_n N_A_788_297#_c_546_n 0.0143191f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_266 N_B1_c_298_n N_VGND_c_563_n 0.00268723f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B1_c_299_n N_VGND_c_564_n 0.00268723f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B1_c_298_n N_VGND_c_565_n 0.00439206f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_269 N_B1_c_299_n N_VGND_c_570_n 0.00423334f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B1_c_298_n N_VGND_c_571_n 0.00621366f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B1_c_299_n N_VGND_c_571_n 0.00687714f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_272 N_B1_c_297_n N_A_503_47#_c_664_n 5.76059e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_298_n N_A_503_47#_c_664_n 0.0121961f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B1_c_305_n N_A_503_47#_c_664_n 0.00717126f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_275 N_B1_c_301_n N_A_503_47#_c_664_n 0.0201153f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B1_c_297_n N_A_503_47#_c_665_n 0.00265533f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_301_n N_A_503_47#_c_665_n 0.0113987f $X=3.815 $Y=1.16 $X2=0 $Y2=0
cc_278 N_B1_c_298_n N_A_503_47#_c_681_n 5.32212e-19 $X=3.875 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_B1_c_299_n N_A_503_47#_c_666_n 0.00995989f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_B1_c_300_n N_A_503_47#_c_666_n 0.00499986f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B1_c_305_n N_A_503_47#_c_666_n 0.00779194f $X=5.13 $Y=1.53 $X2=0 $Y2=0
cc_282 B1 N_A_503_47#_c_666_n 0.0268868f $X=5.195 $Y=1.105 $X2=0 $Y2=0
cc_283 N_B1_c_299_n N_A_503_47#_c_667_n 0.00644736f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_B2_c_375_n N_VPWR_c_427_n 0.00429453f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_285 N_B2_c_376_n N_VPWR_c_427_n 0.00429453f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B2_c_375_n N_VPWR_c_418_n 0.00609021f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B2_c_376_n N_VPWR_c_418_n 0.00609021f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_288 N_B2_c_375_n N_Y_c_516_n 0.0108425f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_289 N_B2_c_375_n N_A_788_297#_c_547_n 0.0100164f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_290 N_B2_c_376_n N_A_788_297#_c_547_n 0.0143148f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B2_c_371_n N_VGND_c_563_n 0.00268723f $X=4.295 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_372_n N_VGND_c_564_n 0.00268723f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B2_c_371_n N_VGND_c_567_n 0.00424416f $X=4.295 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B2_c_372_n N_VGND_c_567_n 0.00437852f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_295 N_B2_c_371_n N_VGND_c_571_n 0.00600559f $X=4.295 $Y=0.995 $X2=0 $Y2=0
cc_296 N_B2_c_372_n N_VGND_c_571_n 0.00615622f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_297 N_B2_c_371_n N_A_503_47#_c_664_n 0.00891961f $X=4.295 $Y=0.995 $X2=0
+ $Y2=0
cc_298 B2 N_A_503_47#_c_664_n 0.00545718f $X=4.66 $Y=1.105 $X2=0 $Y2=0
cc_299 N_B2_c_371_n N_A_503_47#_c_681_n 0.00644736f $X=4.295 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_B2_c_372_n N_A_503_47#_c_666_n 0.0106151f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_301 B2 N_A_503_47#_c_666_n 0.012523f $X=4.66 $Y=1.105 $X2=0 $Y2=0
cc_302 N_B2_c_372_n N_A_503_47#_c_667_n 5.32212e-19 $X=4.815 $Y=0.995 $X2=0
+ $Y2=0
cc_303 N_B2_c_371_n N_A_503_47#_c_669_n 0.00135102f $X=4.295 $Y=0.995 $X2=0
+ $Y2=0
cc_304 B2 N_A_503_47#_c_669_n 0.0307352f $X=4.66 $Y=1.105 $X2=0 $Y2=0
cc_305 N_B2_c_374_n N_A_503_47#_c_669_n 0.00486271f $X=4.79 $Y=1.202 $X2=0 $Y2=0
cc_306 N_VPWR_c_418_n N_Y_M1009_s 0.0024101f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_307 N_VPWR_c_418_n N_Y_M1005_s 0.00232092f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_308 N_VPWR_c_425_n N_Y_c_504_n 0.0203479f $X=3.455 $Y=2.72 $X2=0 $Y2=0
cc_309 N_VPWR_c_418_n N_Y_c_504_n 0.012629f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_310 N_VPWR_c_433_n N_Y_c_504_n 0.0272573f $X=2.725 $Y=2.47 $X2=0 $Y2=0
cc_311 N_VPWR_M1016_d N_Y_c_516_n 0.00878823f $X=3.435 $Y=1.485 $X2=0 $Y2=0
cc_312 N_VPWR_c_423_n N_Y_c_516_n 0.0166773f $X=3.58 $Y=2.3 $X2=0 $Y2=0
cc_313 N_VPWR_c_418_n N_Y_c_516_n 0.00865823f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_418_n N_Y_c_508_n 0.00773108f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_418_n N_A_788_297#_M1014_d 0.00241598f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_316 N_VPWR_c_418_n N_A_788_297#_M1008_d 0.00297222f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_427_n N_A_788_297#_c_547_n 0.0536835f $X=5.415 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_418_n N_A_788_297#_c_547_n 0.0335464f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_427_n N_A_788_297#_c_553_n 0.0143006f $X=5.415 $Y=2.72 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_418_n N_A_788_297#_c_553_n 0.00938288f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_Y_c_516_n N_A_788_297#_M1014_d 0.00368732f $X=4.43 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_322 N_Y_M1005_s N_A_788_297#_c_547_n 0.00352392f $X=4.41 $Y=1.485 $X2=0 $Y2=0
cc_323 N_Y_c_516_n N_A_788_297#_c_547_n 0.00608347f $X=4.43 $Y=1.87 $X2=0 $Y2=0
cc_324 N_Y_c_521_n N_A_788_297#_c_547_n 0.0127274f $X=4.555 $Y=1.87 $X2=0 $Y2=0
cc_325 N_Y_c_516_n N_A_788_297#_c_553_n 0.0130645f $X=4.43 $Y=1.87 $X2=0 $Y2=0
cc_326 N_Y_M1010_s N_VGND_c_571_n 0.00256987f $X=2.975 $Y=0.235 $X2=0 $Y2=0
cc_327 N_Y_M1010_s N_A_503_47#_c_670_n 0.00399909f $X=2.975 $Y=0.235 $X2=0 $Y2=0
cc_328 N_Y_c_496_n N_A_503_47#_c_670_n 0.0219167f $X=3.11 $Y=0.73 $X2=0 $Y2=0
cc_329 N_Y_c_497_n N_A_503_47#_c_670_n 0.00473744f $X=3.18 $Y=1.36 $X2=0 $Y2=0
cc_330 N_Y_c_496_n N_A_503_47#_c_665_n 0.00141443f $X=3.11 $Y=0.73 $X2=0 $Y2=0
cc_331 N_VGND_c_571_n N_A_123_47#_M1004_s 0.00218529f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_332 N_VGND_c_571_n N_A_123_47#_M1011_s 0.00226774f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_561_n N_A_123_47#_c_643_n 0.0133617f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_334 N_VGND_c_569_n N_A_123_47#_c_643_n 0.0140015f $X=2.035 $Y=0 $X2=0 $Y2=0
cc_335 N_VGND_c_571_n N_A_123_47#_c_643_n 0.0107693f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_336 N_VGND_c_561_n N_A_123_47#_c_642_n 0.0307592f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_337 N_VGND_c_569_n N_A_123_47#_c_647_n 0.0427166f $X=2.035 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_c_571_n N_A_123_47#_c_647_n 0.0351264f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_571_n N_A_503_47#_M1010_d 0.00250339f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_340 N_VGND_c_571_n N_A_503_47#_M1012_d 0.00294504f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_571_n N_A_503_47#_M1002_d 0.00304143f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_571_n N_A_503_47#_M1018_d 0.00250309f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_565_n N_A_503_47#_c_704_n 0.0184525f $X=4 $Y=0 $X2=0 $Y2=0
cc_344 N_VGND_c_571_n N_A_503_47#_c_704_n 0.0109628f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_345 N_VGND_M1013_s N_A_503_47#_c_664_n 0.00165819f $X=3.95 $Y=0.235 $X2=0
+ $Y2=0
cc_346 N_VGND_c_563_n N_A_503_47#_c_664_n 0.0116529f $X=4.085 $Y=0.39 $X2=0
+ $Y2=0
cc_347 N_VGND_c_565_n N_A_503_47#_c_664_n 0.00248756f $X=4 $Y=0 $X2=0 $Y2=0
cc_348 N_VGND_c_567_n N_A_503_47#_c_664_n 0.00193763f $X=4.94 $Y=0 $X2=0 $Y2=0
cc_349 N_VGND_c_571_n N_A_503_47#_c_664_n 0.00943347f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_350 N_VGND_c_567_n N_A_503_47#_c_681_n 0.0231806f $X=4.94 $Y=0 $X2=0 $Y2=0
cc_351 N_VGND_c_571_n N_A_503_47#_c_681_n 0.0143352f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_M1017_s N_A_503_47#_c_666_n 0.00162089f $X=4.89 $Y=0.235 $X2=0
+ $Y2=0
cc_353 N_VGND_c_564_n N_A_503_47#_c_666_n 0.0122559f $X=5.025 $Y=0.39 $X2=0
+ $Y2=0
cc_354 N_VGND_c_567_n N_A_503_47#_c_666_n 0.00254521f $X=4.94 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_570_n N_A_503_47#_c_666_n 0.00198695f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_571_n N_A_503_47#_c_666_n 0.0094839f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_c_570_n N_A_503_47#_c_667_n 0.0244796f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_358 N_VGND_c_571_n N_A_503_47#_c_667_n 0.0143352f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_359 N_VGND_c_562_n N_A_503_47#_c_668_n 0.0174095f $X=2.12 $Y=0.39 $X2=0 $Y2=0
cc_360 N_VGND_c_565_n N_A_503_47#_c_668_n 0.0590629f $X=4 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_571_n N_A_503_47#_c_668_n 0.0367524f $X=5.75 $Y=0 $X2=0 $Y2=0
