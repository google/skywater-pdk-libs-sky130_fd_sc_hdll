* File: sky130_fd_sc_hdll__inv_4.pex.spice
* Created: Wed Sep  2 08:33:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 27 28 33 46 47 54 57 60
c78 7 0 6.33157e-20 $X=1.015 $Y=1.41
r79 47 48 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.202
+ $X2=1.98 $Y2=1.202
r80 46 60 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=1.72 $Y=1.2 $X2=1.61
+ $Y2=1.2
r81 45 47 30.4489 $w=3.72e-07 $l=2.35e-07 $layer=POLY_cond $X=1.72 $Y=1.202
+ $X2=1.955 $Y2=1.202
r82 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.72
+ $Y=1.16 $X2=1.72 $Y2=1.16
r83 43 45 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.72 $Y2=1.202
r84 42 43 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r85 41 42 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.04 $Y=1.202
+ $X2=1.485 $Y2=1.202
r86 40 41 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.015 $Y=1.202
+ $X2=1.04 $Y2=1.202
r87 39 40 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.57 $Y=1.202
+ $X2=1.015 $Y2=1.202
r88 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.545 $Y=1.202
+ $X2=0.57 $Y2=1.202
r89 33 38 13.6879 $w=3.72e-07 $l=1.19164e-07 $layer=POLY_cond $X=0.445 $Y=1.16
+ $X2=0.545 $Y2=1.202
r90 33 35 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=0.445 $Y=1.16
+ $X2=0.27 $Y2=1.16
r91 28 60 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.605 $Y=1.2 $X2=1.61
+ $Y2=1.2
r92 28 57 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=1.605 $Y=1.2
+ $X2=1.15 $Y2=1.2
r93 27 57 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=1.14 $Y=1.2 $X2=1.15
+ $Y2=1.2
r94 27 54 20.744 $w=2.48e-07 $l=4.5e-07 $layer=LI1_cond $X=1.14 $Y=1.2 $X2=0.69
+ $Y2=1.2
r95 26 54 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=0.675 $Y=1.2
+ $X2=0.69 $Y2=1.2
r96 25 26 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=0.23 $Y=1.2
+ $X2=0.675 $Y2=1.2
r97 25 35 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r98 22 48 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.98 $Y2=1.202
r99 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.98 $Y2=0.56
r100 19 47 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.202
r101 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r102 16 43 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r103 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r104 13 42 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r105 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r106 10 41 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.04 $Y=0.995
+ $X2=1.04 $Y2=1.202
r107 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.04 $Y=0.995
+ $X2=1.04 $Y2=0.56
r108 7 40 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.202
r109 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.985
r110 4 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.57 $Y=0.995
+ $X2=0.57 $Y2=1.202
r111 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.57 $Y=0.995
+ $X2=0.57 $Y2=0.56
r112 1 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.545 $Y=1.41
+ $X2=0.545 $Y2=1.202
r113 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.545 $Y=1.41
+ $X2=0.545 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_4%VPWR 1 2 3 10 12 18 22 25 26 28 29 30 40 41
r42 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r43 38 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r44 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 32 44 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r48 32 34 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 30 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r50 30 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r51 28 37 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 28 29 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.21 $Y2=2.72
r53 27 40 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.53 $Y2=2.72
r54 27 29 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.21 $Y2=2.72
r55 25 34 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.25 $Y2=2.72
r57 24 37 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.25 $Y2=2.72
r59 20 29 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.21 $Y=2.635
+ $X2=2.21 $Y2=2.72
r60 20 22 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.21 $Y=2.635
+ $X2=2.21 $Y2=2.34
r61 16 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=2.635
+ $X2=1.25 $Y2=2.72
r62 16 18 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.25 $Y=2.635
+ $X2=1.25 $Y2=2
r63 12 15 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=0.262 $Y=1.66
+ $X2=0.262 $Y2=2.34
r64 10 44 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.197 $Y2=2.72
r65 10 15 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.262 $Y2=2.34
r66 3 22 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2.34
r67 2 18 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=2
r68 1 15 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=2.34
r69 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_4%Y 1 2 3 4 15 17 19 21 22 23 27 31 33 35 39
+ 41 42 43 44 50 51
c82 41 0 6.33157e-20 $X=1.72 $Y=1.66
r83 44 51 2.9277 $w=2.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.53 $Y=1.59 $X2=2.53
+ $Y2=1.495
r84 44 51 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.53 $Y=1.47
+ $X2=2.53 $Y2=1.495
r85 43 44 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=2.53 $Y=1.19
+ $X2=2.53 $Y2=1.47
r86 42 50 2.87089 $w=2.7e-07 $l=9e-08 $layer=LI1_cond $X=2.53 $Y=0.815 $X2=2.53
+ $Y2=0.905
r87 42 43 11.5244 $w=2.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.53 $Y=0.92
+ $X2=2.53 $Y2=1.19
r88 42 50 0.640246 $w=2.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=0.92
+ $X2=2.53 $Y2=0.905
r89 36 41 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.59
+ $X2=1.695 $Y2=1.59
r90 35 44 4.16041 $w=1.9e-07 $l=1.35e-07 $layer=LI1_cond $X=2.395 $Y=1.59
+ $X2=2.53 $Y2=1.59
r91 35 36 29.7703 $w=1.88e-07 $l=5.1e-07 $layer=LI1_cond $X=2.395 $Y=1.59
+ $X2=1.885 $Y2=1.59
r92 34 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=0.815
+ $X2=1.695 $Y2=0.815
r93 33 42 4.30634 $w=1.8e-07 $l=1.35e-07 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=2.53 $Y2=0.815
r94 33 34 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=2.395 $Y=0.815
+ $X2=1.885 $Y2=0.815
r95 29 41 1.15089 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.695 $Y=1.685
+ $X2=1.695 $Y2=1.59
r96 29 31 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=1.695 $Y=1.685
+ $X2=1.695 $Y2=2.34
r97 25 39 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.695 $Y=0.725
+ $X2=1.695 $Y2=0.815
r98 25 27 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.695 $Y=0.725
+ $X2=1.695 $Y2=0.42
r99 24 38 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.945 $Y=1.58
+ $X2=0.755 $Y2=1.58
r100 23 41 9.12476 $w=1.8e-07 $l=1.94936e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.695 $Y2=1.59
r101 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.945 $Y2=1.58
r102 21 39 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=1.695 $Y2=0.815
r103 21 22 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=0.945 $Y2=0.815
r104 17 38 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=1.665
+ $X2=0.755 $Y2=1.58
r105 17 19 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.755 $Y=1.665
+ $X2=0.755 $Y2=2.34
r106 13 22 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.755 $Y=0.725
+ $X2=0.945 $Y2=0.815
r107 13 15 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=0.755 $Y=0.725
+ $X2=0.755 $Y2=0.42
r108 4 41 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.66
r109 4 31 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2.34
r110 3 38 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.485 $X2=0.78 $Y2=1.66
r111 3 19 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.635
+ $Y=1.485 $X2=0.78 $Y2=2.34
r112 2 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.72 $Y2=0.42
r113 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=0.645
+ $Y=0.235 $X2=0.78 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_4%VGND 1 2 3 10 12 16 20 23 24 26 27 28 38 39
r45 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r46 36 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r47 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r48 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r49 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r50 30 42 4.1239 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r51 30 32 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=1.15
+ $Y2=0
r52 28 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r53 28 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r54 26 35 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.07
+ $Y2=0
r55 26 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.23
+ $Y2=0
r56 25 38 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.53
+ $Y2=0
r57 25 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.23
+ $Y2=0
r58 23 32 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=0 $X2=1.15
+ $Y2=0
r59 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.165 $Y=0 $X2=1.25
+ $Y2=0
r60 22 35 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=2.07
+ $Y2=0
r61 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.25
+ $Y2=0
r62 18 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.085
+ $X2=2.23 $Y2=0
r63 18 20 13.8293 $w=2.48e-07 $l=3e-07 $layer=LI1_cond $X=2.23 $Y=0.085 $X2=2.23
+ $Y2=0.385
r64 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0
r65 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.25 $Y=0.085
+ $X2=1.25 $Y2=0.38
r66 10 42 3.12417 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.197 $Y2=0
r67 10 12 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.262 $Y=0.085
+ $X2=0.262 $Y2=0.38
r68 3 20 182 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.385
r69 2 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.115
+ $Y=0.235 $X2=1.25 $Y2=0.38
r70 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

