* File: sky130_fd_sc_hdll__nor3b_4.pex.spice
* Created: Thu Aug 27 19:16:46 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%C_N 1 3 4 6 7 12 15
c27 4 0 1.57516e-19 $X=0.54 $Y=0.995
r28 12 13 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r29 10 12 31.8678 $w=3.63e-07 $l=2.4e-07 $layer=POLY_cond $X=0.275 $Y=1.202
+ $X2=0.515 $Y2=1.202
r30 7 15 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.18 $X2=0.23
+ $Y2=1.18
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r32 4 13 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r34 1 12 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 43 49 52 56
r71 43 44 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.42 $Y2=1.202
r72 42 52 7.65801 $w=2.08e-07 $l=1.45e-07 $layer=LI1_cond $X=2.22 $Y=1.18
+ $X2=2.075 $Y2=1.18
r73 41 43 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=2.22 $Y=1.202
+ $X2=2.395 $Y2=1.202
r74 41 42 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.22
+ $Y=1.16 $X2=2.22 $Y2=1.16
r75 39 41 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=2.22 $Y2=1.202
r76 38 39 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.9 $Y=1.202
+ $X2=1.925 $Y2=1.202
r77 37 38 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.9 $Y2=1.202
r78 35 37 1.94355 $w=3.72e-07 $l=1.5e-08 $layer=POLY_cond $X=1.44 $Y=1.202
+ $X2=1.455 $Y2=1.202
r79 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.44
+ $Y=1.16 $X2=1.44 $Y2=1.16
r80 33 35 1.2957 $w=3.72e-07 $l=1e-08 $layer=POLY_cond $X=1.43 $Y=1.202 $X2=1.44
+ $Y2=1.202
r81 32 33 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r82 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r83 27 56 0.528139 $w=2.08e-07 $l=1e-08 $layer=LI1_cond $X=2.525 $Y=1.18
+ $X2=2.535 $Y2=1.18
r84 27 42 16.1082 $w=2.08e-07 $l=3.05e-07 $layer=LI1_cond $X=2.525 $Y=1.18
+ $X2=2.22 $Y2=1.18
r85 26 52 0.792208 $w=2.08e-07 $l=1.5e-08 $layer=LI1_cond $X=2.06 $Y=1.18
+ $X2=2.075 $Y2=1.18
r86 26 49 23.5022 $w=2.08e-07 $l=4.45e-07 $layer=LI1_cond $X=2.06 $Y=1.18
+ $X2=1.615 $Y2=1.18
r87 25 49 0.792208 $w=2.08e-07 $l=1.5e-08 $layer=LI1_cond $X=1.6 $Y=1.18
+ $X2=1.615 $Y2=1.18
r88 25 36 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=1.6 $Y=1.18 $X2=1.44
+ $Y2=1.18
r89 22 44 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=0.56
r91 19 43 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r93 16 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r95 13 38 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.9 $Y=0.995
+ $X2=1.9 $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.9 $Y=0.995 $X2=1.9
+ $Y2=0.56
r97 10 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r99 7 33 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r101 4 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r103 1 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 36 39 45
c74 36 0 1.54579e-19 $X=4.23 $Y=1.16
r75 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=4.82 $Y2=1.202
r76 38 39 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=4.325 $Y=1.202
+ $X2=4.795 $Y2=1.202
r77 37 38 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=4.3 $Y=1.202
+ $X2=4.325 $Y2=1.202
r78 36 45 17.1645 $w=2.08e-07 $l=3.25e-07 $layer=LI1_cond $X=4.23 $Y=1.18
+ $X2=3.905 $Y2=1.18
r79 35 37 9.06989 $w=3.72e-07 $l=7e-08 $layer=POLY_cond $X=4.23 $Y=1.202 $X2=4.3
+ $Y2=1.202
r80 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.23
+ $Y=1.16 $X2=4.23 $Y2=1.16
r81 33 35 48.5887 $w=3.72e-07 $l=3.75e-07 $layer=POLY_cond $X=3.855 $Y=1.202
+ $X2=4.23 $Y2=1.202
r82 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.83 $Y=1.202
+ $X2=3.855 $Y2=1.202
r83 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=3.45 $Y=1.202
+ $X2=3.83 $Y2=1.202
r84 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.16 $X2=3.45 $Y2=1.16
r85 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=3.385 $Y=1.202
+ $X2=3.45 $Y2=1.202
r86 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.36 $Y=1.202
+ $X2=3.385 $Y2=1.202
r87 25 45 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=3.9 $Y=1.18 $X2=3.905
+ $Y2=1.18
r88 25 31 23.7662 $w=2.08e-07 $l=4.5e-07 $layer=LI1_cond $X=3.9 $Y=1.18 $X2=3.45
+ $Y2=1.18
r89 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=0.56
r91 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.795 $Y=1.41
+ $X2=4.795 $Y2=1.985
r93 16 38 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.325 $Y=1.41
+ $X2=4.325 $Y2=1.985
r95 13 37 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.3 $Y=0.995
+ $X2=4.3 $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.3 $Y=0.995 $X2=4.3
+ $Y2=0.56
r97 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.855 $Y=1.41
+ $X2=3.855 $Y2=1.985
r99 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r101 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.985
r103 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.36 $Y=0.995
+ $X2=3.36 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%A_27_47# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 35 37 39 41 42 44 45 48 49 54 59 68
c154 68 0 1.54579e-19 $X=6.675 $Y=1.202
r155 68 69 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.675 $Y=1.202
+ $X2=6.7 $Y2=1.202
r156 65 66 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.18 $Y=1.202
+ $X2=6.205 $Y2=1.202
r157 64 65 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=5.735 $Y=1.202
+ $X2=6.18 $Y2=1.202
r158 63 64 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.71 $Y=1.202
+ $X2=5.735 $Y2=1.202
r159 60 61 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.265 $Y2=1.202
r160 55 68 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=6.5 $Y=1.202
+ $X2=6.675 $Y2=1.202
r161 55 66 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=6.5 $Y=1.202
+ $X2=6.205 $Y2=1.202
r162 54 55 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.5
+ $Y=1.16 $X2=6.5 $Y2=1.16
r163 52 63 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=5.33 $Y=1.202
+ $X2=5.71 $Y2=1.202
r164 52 61 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=5.33 $Y=1.202
+ $X2=5.265 $Y2=1.202
r165 51 54 61.7922 $w=2.08e-07 $l=1.17e-06 $layer=LI1_cond $X=5.33 $Y=1.18
+ $X2=6.5 $Y2=1.18
r166 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.33
+ $Y=1.16 $X2=5.33 $Y2=1.16
r167 49 51 9.24242 $w=2.08e-07 $l=1.75e-07 $layer=LI1_cond $X=5.155 $Y=1.18
+ $X2=5.33 $Y2=1.18
r168 47 49 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=5.07 $Y=1.285
+ $X2=5.155 $Y2=1.18
r169 47 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.07 $Y=1.285
+ $X2=5.07 $Y2=1.455
r170 46 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=1.54
+ $X2=0.75 $Y2=1.54
r171 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.985 $Y=1.54
+ $X2=5.07 $Y2=1.455
r172 45 46 270.749 $w=1.68e-07 $l=4.15e-06 $layer=LI1_cond $X=4.985 $Y=1.54
+ $X2=0.835 $Y2=1.54
r173 44 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.455
+ $X2=0.75 $Y2=1.54
r174 43 44 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.75 $Y=0.905
+ $X2=0.75 $Y2=1.455
r175 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.665 $Y=0.82
+ $X2=0.75 $Y2=0.905
r176 41 42 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.665 $Y=0.82
+ $X2=0.445 $Y2=0.82
r177 40 58 4.74967 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.257 $Y2=1.54
r178 39 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=1.54
+ $X2=0.75 $Y2=1.54
r179 39 40 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.665 $Y=1.54
+ $X2=0.405 $Y2=1.54
r180 35 58 2.72785 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=0.257 $Y=1.625
+ $X2=0.257 $Y2=1.54
r181 35 37 26.3695 $w=2.93e-07 $l=6.75e-07 $layer=LI1_cond $X=0.257 $Y=1.625
+ $X2=0.257 $Y2=2.3
r182 31 42 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.277 $Y=0.735
+ $X2=0.445 $Y2=0.82
r183 31 33 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=0.277 $Y=0.735
+ $X2=0.277 $Y2=0.39
r184 28 69 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.7 $Y=0.995
+ $X2=6.7 $Y2=1.202
r185 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.7 $Y=0.995
+ $X2=6.7 $Y2=0.56
r186 25 68 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.202
r187 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.675 $Y=1.41
+ $X2=6.675 $Y2=1.985
r188 22 66 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.202
r189 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.205 $Y=1.41
+ $X2=6.205 $Y2=1.985
r190 19 65 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.18 $Y=0.995
+ $X2=6.18 $Y2=1.202
r191 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.18 $Y=0.995
+ $X2=6.18 $Y2=0.56
r192 16 64 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.202
r193 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.735 $Y=1.41
+ $X2=5.735 $Y2=1.985
r194 13 63 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=1.202
r195 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=0.56
r196 10 61 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.202
r197 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.265 $Y=1.41
+ $X2=5.265 $Y2=1.985
r198 7 60 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r199 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r200 2 58 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r201 2 37 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r202 1 33 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%VPWR 1 2 3 14 16 20 22 26 28 35 36 39 42
+ 45
r93 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r94 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r95 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r96 40 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r97 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r98 35 36 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r99 33 36 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=2.99 $Y=2.72 $X2=7.13
+ $Y2=2.72
r100 33 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r101 32 35 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=7.13 $Y2=2.72
r102 32 33 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r103 30 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.63 $Y2=2.72
r104 30 32 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.755 $Y=2.72
+ $X2=2.99 $Y2=2.72
r105 28 40 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r106 24 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2.72
r107 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.63 $Y=2.635
+ $X2=2.63 $Y2=2.3
r108 23 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=2.72
+ $X2=1.69 $Y2=2.72
r109 22 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=2.63 $Y2=2.72
r110 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.505 $Y=2.72
+ $X2=1.815 $Y2=2.72
r111 18 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r112 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.3
r113 17 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r114 16 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=1.69 $Y2=2.72
r115 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=2.72
+ $X2=0.875 $Y2=2.72
r116 12 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r117 12 14 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r118 3 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=2.3
r119 2 20 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2.3
r120 1 14 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%A_215_297# 1 2 3 4 15 19 21 24 26 27 32
r48 32 35 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.56 $Y=1.88 $X2=4.56
+ $Y2=1.96
r49 27 30 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.62 $Y=1.88 $X2=3.62
+ $Y2=1.96
r50 22 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.745 $Y=1.88
+ $X2=3.62 $Y2=1.88
r51 21 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=1.88
+ $X2=4.56 $Y2=1.88
r52 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.435 $Y=1.88
+ $X2=3.745 $Y2=1.88
r53 20 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=1.88
+ $X2=2.16 $Y2=1.88
r54 19 27 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.495 $Y=1.88
+ $X2=3.62 $Y2=1.88
r55 19 20 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=3.495 $Y=1.88
+ $X2=2.285 $Y2=1.88
r56 16 24 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.88
+ $X2=1.22 $Y2=1.88
r57 15 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=1.88
+ $X2=2.16 $Y2=1.88
r58 15 16 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.88
+ $X2=1.345 $Y2=1.88
r59 4 35 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.415
+ $Y=1.485 $X2=4.56 $Y2=1.96
r60 3 30 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.62 $Y2=1.96
r61 2 26 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.96
r62 1 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%A_605_297# 1 2 3 4 5 16 18 22 24 28 30 34
+ 37 42 46 47
r58 42 44 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.09 $Y=2.3 $X2=4.09
+ $Y2=2.38
r59 37 39 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.15 $Y=2.3 $X2=3.15
+ $Y2=2.38
r60 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.91 $Y=2.295
+ $X2=6.91 $Y2=1.96
r61 31 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.095 $Y=2.38
+ $X2=5.97 $Y2=2.38
r62 30 32 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.785 $Y=2.38
+ $X2=6.91 $Y2=2.295
r63 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.785 $Y=2.38
+ $X2=6.095 $Y2=2.38
r64 26 47 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=2.295
+ $X2=5.97 $Y2=2.38
r65 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.97 $Y=2.295
+ $X2=5.97 $Y2=1.96
r66 25 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.155 $Y=2.38
+ $X2=5.03 $Y2=2.38
r67 24 47 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.845 $Y=2.38
+ $X2=5.97 $Y2=2.38
r68 24 25 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.845 $Y=2.38
+ $X2=5.155 $Y2=2.38
r69 20 46 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=2.295
+ $X2=5.03 $Y2=2.38
r70 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.03 $Y=2.295
+ $X2=5.03 $Y2=1.96
r71 19 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.215 $Y=2.38
+ $X2=4.09 $Y2=2.38
r72 18 46 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.905 $Y=2.38
+ $X2=5.03 $Y2=2.38
r73 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.905 $Y=2.38
+ $X2=4.215 $Y2=2.38
r74 17 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.275 $Y=2.38
+ $X2=3.15 $Y2=2.38
r75 16 44 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.965 $Y=2.38
+ $X2=4.09 $Y2=2.38
r76 16 17 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.965 $Y=2.38
+ $X2=3.275 $Y2=2.38
r77 5 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.765
+ $Y=1.485 $X2=6.91 $Y2=1.96
r78 4 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.825
+ $Y=1.485 $X2=5.97 $Y2=1.96
r79 3 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.885
+ $Y=1.485 $X2=5.03 $Y2=1.96
r80 2 42 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.945
+ $Y=1.485 $X2=4.09 $Y2=2.3
r81 1 37 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.025
+ $Y=1.485 $X2=3.15 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%Y 1 2 3 4 5 6 7 8 27 29 30 33 35 39 41 45
+ 47 51 55 57 61 65 67 69 70 71 72 74 75 77 80 83
c163 30 0 1.57516e-19 $X=1.385 $Y=0.815
r164 80 83 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=7.075 $Y=1.19
+ $X2=7.075 $Y2=1.155
r165 79 80 8.98228 $w=3.38e-07 $l=2.65e-07 $layer=LI1_cond $X=7.075 $Y=1.455
+ $X2=7.075 $Y2=1.19
r166 78 83 8.47385 $w=3.38e-07 $l=2.5e-07 $layer=LI1_cond $X=7.075 $Y=0.905
+ $X2=7.075 $Y2=1.155
r167 68 75 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.605 $Y=0.815
+ $X2=6.415 $Y2=0.815
r168 67 78 7.6914 $w=1.8e-07 $l=2.10238e-07 $layer=LI1_cond $X=6.905 $Y=0.815
+ $X2=7.075 $Y2=0.905
r169 67 68 18.4848 $w=1.78e-07 $l=3e-07 $layer=LI1_cond $X=6.905 $Y=0.815
+ $X2=6.605 $Y2=0.815
r170 66 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.565 $Y=1.54
+ $X2=6.44 $Y2=1.54
r171 65 79 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.905 $Y=1.54
+ $X2=7.075 $Y2=1.455
r172 65 66 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.905 $Y=1.54
+ $X2=6.565 $Y2=1.54
r173 59 75 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.415 $Y=0.725
+ $X2=6.415 $Y2=0.815
r174 59 61 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.415 $Y=0.725
+ $X2=6.415 $Y2=0.39
r175 58 72 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.665 $Y=0.815
+ $X2=5.475 $Y2=0.815
r176 57 75 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.225 $Y=0.815
+ $X2=6.415 $Y2=0.815
r177 57 58 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.225 $Y=0.815
+ $X2=5.665 $Y2=0.815
r178 56 74 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.625 $Y=1.54
+ $X2=5.5 $Y2=1.54
r179 55 77 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.315 $Y=1.54
+ $X2=6.44 $Y2=1.54
r180 55 56 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.315 $Y=1.54
+ $X2=5.625 $Y2=1.54
r181 49 72 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.475 $Y=0.725
+ $X2=5.475 $Y2=0.815
r182 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.475 $Y=0.725
+ $X2=5.475 $Y2=0.39
r183 48 71 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.725 $Y=0.815
+ $X2=4.535 $Y2=0.815
r184 47 72 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=5.475 $Y2=0.815
r185 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.285 $Y=0.815
+ $X2=4.725 $Y2=0.815
r186 43 71 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.535 $Y=0.725
+ $X2=4.535 $Y2=0.815
r187 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.535 $Y=0.725
+ $X2=4.535 $Y2=0.39
r188 42 70 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.785 $Y=0.815
+ $X2=3.595 $Y2=0.815
r189 41 71 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.345 $Y=0.815
+ $X2=4.535 $Y2=0.815
r190 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.345 $Y=0.815
+ $X2=3.785 $Y2=0.815
r191 37 70 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.595 $Y=0.725
+ $X2=3.595 $Y2=0.815
r192 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.595 $Y=0.725
+ $X2=3.595 $Y2=0.39
r193 36 69 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=0.815
+ $X2=2.135 $Y2=0.815
r194 35 70 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.405 $Y=0.815
+ $X2=3.595 $Y2=0.815
r195 35 36 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=3.405 $Y=0.815
+ $X2=2.325 $Y2=0.815
r196 31 69 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.135 $Y=0.725
+ $X2=2.135 $Y2=0.815
r197 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.135 $Y=0.725
+ $X2=2.135 $Y2=0.39
r198 29 69 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=0.815
+ $X2=2.135 $Y2=0.815
r199 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.945 $Y=0.815
+ $X2=1.385 $Y2=0.815
r200 25 30 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=1.195 $Y=0.725
+ $X2=1.385 $Y2=0.815
r201 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.195 $Y=0.725
+ $X2=1.195 $Y2=0.39
r202 8 77 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.295
+ $Y=1.485 $X2=6.44 $Y2=1.62
r203 7 74 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.355
+ $Y=1.485 $X2=5.5 $Y2=1.62
r204 6 61 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.255
+ $Y=0.235 $X2=6.44 $Y2=0.39
r205 5 51 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.39
r206 4 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.375
+ $Y=0.235 $X2=4.56 $Y2=0.39
r207 3 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.435
+ $Y=0.235 $X2=3.62 $Y2=0.39
r208 2 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.975
+ $Y=0.235 $X2=2.16 $Y2=0.39
r209 1 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3B_4%VGND 1 2 3 4 5 6 7 26 28 32 36 40 44 48 51
+ 52 54 55 57 58 60 61 62 83 84 87 90 95 98 100
r118 97 98 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=0.235
+ $X2=3.235 $Y2=0.235
r119 93 97 2.9902 $w=6.38e-07 $l=1.6e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=3.15 $Y2=0.235
r120 93 95 15.6497 $w=6.38e-07 $l=4.45e-07 $layer=LI1_cond $X=2.99 $Y=0.235
+ $X2=2.545 $Y2=0.235
r121 93 94 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r122 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r123 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r124 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r125 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r126 81 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r127 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r128 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r129 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r130 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r131 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r132 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r133 72 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r134 71 98 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=3.91 $Y=0
+ $X2=3.235 $Y2=0
r135 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r136 68 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r137 68 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r138 67 95 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.53 $Y=0 $X2=2.545
+ $Y2=0
r139 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r140 65 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.69
+ $Y2=0
r141 65 67 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=2.53 $Y2=0
r142 62 88 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r143 62 100 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r144 60 80 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.825 $Y=0
+ $X2=6.67 $Y2=0
r145 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.825 $Y=0 $X2=6.91
+ $Y2=0
r146 59 83 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.995 $Y=0
+ $X2=7.13 $Y2=0
r147 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=0 $X2=6.91
+ $Y2=0
r148 57 77 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.885 $Y=0
+ $X2=5.75 $Y2=0
r149 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.885 $Y=0 $X2=5.97
+ $Y2=0
r150 56 80 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.055 $Y=0 $X2=6.67
+ $Y2=0
r151 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=0 $X2=5.97
+ $Y2=0
r152 54 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.945 $Y=0
+ $X2=4.83 $Y2=0
r153 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.945 $Y=0 $X2=5.03
+ $Y2=0
r154 53 77 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.115 $Y=0
+ $X2=5.75 $Y2=0
r155 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.115 $Y=0 $X2=5.03
+ $Y2=0
r156 51 71 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.005 $Y=0 $X2=3.91
+ $Y2=0
r157 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.005 $Y=0 $X2=4.09
+ $Y2=0
r158 50 74 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.175 $Y=0
+ $X2=4.83 $Y2=0
r159 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=0 $X2=4.09
+ $Y2=0
r160 46 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0
r161 46 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.91 $Y=0.085
+ $X2=6.91 $Y2=0.39
r162 42 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0
r163 42 44 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.97 $Y=0.085
+ $X2=5.97 $Y2=0.39
r164 38 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0
r165 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.03 $Y=0.085
+ $X2=5.03 $Y2=0.39
r166 34 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r167 34 36 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.39
r168 30 90 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0
r169 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0.39
r170 29 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.75
+ $Y2=0
r171 28 90 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.69
+ $Y2=0
r172 28 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.835 $Y2=0
r173 24 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r174 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.39
r175 7 48 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=6.775
+ $Y=0.235 $X2=6.91 $Y2=0.39
r176 6 44 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.235 $X2=5.97 $Y2=0.39
r177 5 40 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.895
+ $Y=0.235 $X2=5.03 $Y2=0.39
r178 4 36 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.09 $Y2=0.39
r179 3 97 91 $w=1.7e-07 $l=7.28389e-07 $layer=licon1_NDIFF $count=2 $X=2.495
+ $Y=0.235 $X2=3.15 $Y2=0.39
r180 2 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r181 1 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

