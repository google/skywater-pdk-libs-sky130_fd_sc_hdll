* NGSPICE file created from sky130_fd_sc_hdll__a21o_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 VGND B1 a_84_21# VNB nshort w=650000u l=150000u
+  ad=1.365e+12p pd=1.07e+07u as=4.81e+11p ps=4.08e+06u
M1001 a_523_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.255e+12p pd=1.051e+07u as=1.47e+12p ps=1.294e+07u
M1002 X a_84_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1003 VPWR a_84_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6e+11p ps=5.2e+06u
M1004 VPWR A2 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_84_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_84_21# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_801_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.82e+11p pd=1.86e+06u as=0p ps=0u
M1008 VGND a_84_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_991_47# A1 a_84_21# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1010 VGND A2 a_991_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_523_297# B1 a_84_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1012 VPWR a_84_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_523_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_84_21# B1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VPWR A1 a_523_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND a_84_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_84_21# A1 a_801_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 X a_84_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_84_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

