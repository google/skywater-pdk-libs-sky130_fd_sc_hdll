* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4b_1 A_N B C D VGND VNB VPB VPWR Y
X0 Y a_40_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_40_93# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X3 a_334_47# B a_431_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_40_93# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VGND D a_251_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_251_47# C a_334_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_431_47# a_40_93# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
