* File: sky130_fd_sc_hdll__einvp_1.pex.spice
* Created: Wed Sep  2 08:31:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%TE 3 5 6 7 9 10 12 14 15 16 22
c33 5 0 3.76507e-19 $X=0.495 $Y=1.325
r34 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.16 $X2=0.46 $Y2=1.16
r35 19 21 22.9087 $w=2.63e-07 $l=1.25e-07 $layer=POLY_cond $X=0.46 $Y=1.035
+ $X2=0.46 $Y2=1.16
r36 15 16 7.97386 $w=5.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.34 $Y=1.19
+ $X2=0.34 $Y2=1.53
r37 15 22 0.703576 $w=5.08e-07 $l=3e-08 $layer=LI1_cond $X=0.34 $Y=1.19 $X2=0.34
+ $Y2=1.16
r38 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.945 $Y=0.96
+ $X2=0.945 $Y2=0.56
r39 11 19 15.8942 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.595 $Y=1.035
+ $X2=0.46 $Y2=1.035
r40 10 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.945 $Y2=0.96
r41 10 11 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=0.87 $Y=1.035
+ $X2=0.595 $Y2=1.035
r42 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r43 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r44 5 21 33.1221 $w=2.63e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.46 $Y2=1.16
r45 5 6 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
r46 1 19 22.5691 $w=2.63e-07 $l=7.98436e-08 $layer=POLY_cond $X=0.47 $Y=0.96
+ $X2=0.46 $Y2=1.035
r47 1 3 264.074 $w=1.5e-07 $l=5.15e-07 $layer=POLY_cond $X=0.47 $Y=0.96 $X2=0.47
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%A_27_47# 1 2 7 9 12 16 18 19 20 21 25
c58 21 0 6.83631e-20 $X=0.345 $Y=1.98
c59 20 0 1.52837e-19 $X=0.765 $Y=1.98
c60 19 0 1.55307e-19 $X=0.345 $Y=0.74
c61 7 0 1.1238e-19 $X=1.57 $Y=1.41
r62 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.605
+ $Y=1.16 $X2=1.605 $Y2=1.16
r63 23 25 9.69405 $w=9.23e-07 $l=7.35e-07 $layer=LI1_cond $X=1.227 $Y=1.895
+ $X2=1.227 $Y2=1.16
r64 22 25 4.41838 $w=9.23e-07 $l=3.35e-07 $layer=LI1_cond $X=1.227 $Y=0.825
+ $X2=1.227 $Y2=1.16
r65 20 23 12.3116 $w=1.7e-07 $l=5.02707e-07 $layer=LI1_cond $X=0.765 $Y=1.98
+ $X2=1.227 $Y2=1.895
r66 20 21 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.765 $Y=1.98
+ $X2=0.345 $Y2=1.98
r67 18 22 12.3116 $w=1.7e-07 $l=5.02707e-07 $layer=LI1_cond $X=0.765 $Y=0.74
+ $X2=1.227 $Y2=0.825
r68 18 19 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=0.765 $Y=0.74
+ $X2=0.345 $Y2=0.74
r69 14 21 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=2.065
+ $X2=0.345 $Y2=1.98
r70 14 16 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=2.065
+ $X2=0.215 $Y2=2.275
r71 10 19 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.345 $Y2=0.74
r72 10 12 9.30819 $w=2.58e-07 $l=2.1e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.445
r73 7 26 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.57 $Y=1.41
+ $X2=1.605 $Y2=1.16
r74 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.57 $Y=1.41 $X2=1.57
+ $Y2=1.985
r75 2 16 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.275
r76 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%A 1 3 4 6 7 8 9 14
r29 14 16 35.0907 $w=3.64e-07 $l=2.65e-07 $layer=POLY_cond $X=2.205 $Y=1.202
+ $X2=2.47 $Y2=1.202
r30 13 14 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=2.18 $Y=1.202
+ $X2=2.205 $Y2=1.202
r31 8 9 16.3263 $w=2.38e-07 $l=3.4e-07 $layer=LI1_cond $X=2.505 $Y=1.53
+ $X2=2.505 $Y2=1.87
r32 7 8 17.7668 $w=2.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.505 $Y=1.16
+ $X2=2.505 $Y2=1.53
r33 7 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.16 $X2=2.47 $Y2=1.16
r34 4 14 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.205 $Y=1.41
+ $X2=2.205 $Y2=1.202
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.205 $Y=1.41
+ $X2=2.205 $Y2=1.985
r36 1 13 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.18 $Y=0.995
+ $X2=2.18 $Y2=1.202
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.18 $Y=0.995 $X2=2.18
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%VPWR 1 4 5 8 17 18 23 27
r31 25 27 9.22658 $w=5.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=2.52
+ $X2=1.74 $Y2=2.52
r32 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 22 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r34 21 23 10.1709 $w=5.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.69 $Y=2.52
+ $X2=0.515 $Y2=2.52
r35 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r36 18 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 17 27 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=1.74 $Y2=2.72
r38 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 12 23 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r40 8 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r42 5 21 2.30822 $w=5.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.8 $Y=2.52 $X2=0.69
+ $Y2=2.52
r43 5 7 9.23289 $w=5.68e-07 $l=4.4e-07 $layer=LI1_cond $X=0.8 $Y=2.52 $X2=1.24
+ $Y2=2.52
r44 4 25 3.25249 $w=5.68e-07 $l=1.55e-07 $layer=LI1_cond $X=1.455 $Y=2.52
+ $X2=1.61 $Y2=2.52
r45 4 7 4.51152 $w=5.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.455 $Y=2.52
+ $X2=1.24 $Y2=2.52
r46 1 7 300 $w=1.7e-07 $l=7.8675e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=2.065 $X2=1.24 $Y2=2.355
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%Z 1 2 8 9 10 11 15 24
r34 24 27 3.37077 $w=5.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.285 $Y=0.53
+ $X2=2.44 $Y2=0.53
r35 21 24 4.74082 $w=5.48e-07 $l=2.18e-07 $layer=LI1_cond $X=2.067 $Y=0.53
+ $X2=2.285 $Y2=0.53
r36 15 18 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=2.285 $Y=2.295
+ $X2=2.45 $Y2=2.295
r37 11 18 1.18634 $w=3.38e-07 $l=3.5e-08 $layer=LI1_cond $X=2.485 $Y=2.295
+ $X2=2.45 $Y2=2.295
r38 10 27 0.97861 $w=5.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.485 $Y=0.53
+ $X2=2.44 $Y2=0.53
r39 9 15 4.4064 $w=3.38e-07 $l=1.3e-07 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.285 $Y2=2.295
r40 8 9 7.76859 $w=3.4e-07 $l=2.09428e-07 $layer=LI1_cond $X=2.067 $Y=2.125
+ $X2=2.155 $Y2=2.295
r41 7 21 7.58619 $w=1.75e-07 $l=2.75e-07 $layer=LI1_cond $X=2.067 $Y=0.805
+ $X2=2.067 $Y2=0.53
r42 7 8 83.6571 $w=1.73e-07 $l=1.32e-06 $layer=LI1_cond $X=2.067 $Y=0.805
+ $X2=2.067 $Y2=2.125
r43 2 18 600 $w=1.7e-07 $l=8.89129e-07 $layer=licon1_PDIFF $count=1 $X=2.295
+ $Y=1.485 $X2=2.45 $Y2=2.3
r44 1 27 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.255
+ $Y=0.235 $X2=2.44 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVP_1%VGND 1 4 16 17 21 28
c27 28 0 1.1238e-19 $X=1.5 $Y=0.2
r28 26 28 13.843 $w=5.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.15 $Y=0.2 $X2=1.5
+ $Y2=0.2
r29 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 24 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r31 23 26 9.65256 $w=5.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.2 $X2=1.15
+ $Y2=0.2
r32 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 20 23 0.209838 $w=5.68e-07 $l=1e-08 $layer=LI1_cond $X=0.68 $Y=0.2 $X2=0.69
+ $Y2=0.2
r34 20 21 9.96101 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.68 $Y=0.2
+ $X2=0.515 $Y2=0.2
r35 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r36 14 17 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r37 14 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r38 13 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r39 13 28 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.5
+ $Y2=0
r40 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r41 8 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.515
+ $Y2=0
r42 4 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r44 1 20 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.68 $Y2=0.36
.ends

