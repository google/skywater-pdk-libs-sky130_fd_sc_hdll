* File: sky130_fd_sc_hdll__einvn_1.pex.spice
* Created: Thu Aug 27 19:07:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%TE_B 1 2 3 5 8 10 12 14 15 16 21
r46 20 22 28.2107 $w=2.99e-07 $l=1.75e-07 $layer=POLY_cond $X=0.432 $Y=1.16
+ $X2=0.432 $Y2=1.335
r47 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.405
+ $Y=1.16 $X2=0.405 $Y2=1.16
r48 15 16 9.21954 $w=4.23e-07 $l=3.4e-07 $layer=LI1_cond $X=0.297 $Y=1.19
+ $X2=0.297 $Y2=1.53
r49 15 21 0.813489 $w=4.23e-07 $l=3e-08 $layer=LI1_cond $X=0.297 $Y=1.19
+ $X2=0.297 $Y2=1.16
r50 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r51 11 22 18.89 $w=1.5e-07 $l=1.63e-07 $layer=POLY_cond $X=0.595 $Y=1.335
+ $X2=0.432 $Y2=1.335
r52 10 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.93 $Y=1.335
+ $X2=1.02 $Y2=1.41
r53 10 11 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.93 $Y=1.335
+ $X2=0.595 $Y2=1.335
r54 6 20 38.5562 $w=2.99e-07 $l=2.04316e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.432 $Y2=1.16
r55 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r56 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r57 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r58 1 22 17.3898 $w=2.99e-07 $l=1.01735e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.432 $Y2=1.335
r59 1 2 86.2101 $w=2e-07 $l=2.6e-07 $layer=POLY_cond $X=0.495 $Y=1.41 $X2=0.495
+ $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%A_27_47# 1 2 9 12 14 18 19 20 22 23 24 25
+ 28 29 31 34
c72 28 0 1.38301e-19 $X=1.465 $Y=1.16
r73 29 34 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=1.512 $Y=1.16
+ $X2=1.512 $Y2=0.995
r74 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.16 $X2=1.465 $Y2=1.16
r75 26 28 6.97712 $w=4.78e-07 $l=2.8e-07 $layer=LI1_cond $X=1.36 $Y=1.44
+ $X2=1.36 $Y2=1.16
r76 25 31 36.6314 $w=1.88e-07 $l=6.25e-07 $layer=LI1_cond $X=1.36 $Y=0.71
+ $X2=0.735 $Y2=0.71
r77 25 28 8.846 $w=4.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.36 $Y=0.805
+ $X2=1.36 $Y2=1.16
r78 23 26 8.94461 $w=1.75e-07 $l=2.80143e-07 $layer=LI1_cond $X=1.12 $Y=1.527
+ $X2=1.36 $Y2=1.44
r79 23 24 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.12 $Y=1.527 $X2=0.92
+ $Y2=1.527
r80 21 24 6.82334 $w=1.75e-07 $l=1.29742e-07 $layer=LI1_cond $X=0.827 $Y=1.615
+ $X2=0.92 $Y2=1.527
r81 21 22 16.7862 $w=1.83e-07 $l=2.8e-07 $layer=LI1_cond $X=0.827 $Y=1.615
+ $X2=0.827 $Y2=1.895
r82 19 22 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=0.735 $Y=1.98
+ $X2=0.827 $Y2=1.895
r83 19 20 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.735 $Y=1.98
+ $X2=0.37 $Y2=1.98
r84 18 31 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.37 $Y=0.7
+ $X2=0.735 $Y2=0.7
r85 14 20 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.227 $Y=2.065
+ $X2=0.37 $Y2=1.98
r86 14 16 4.2807 $w=2.85e-07 $l=1e-07 $layer=LI1_cond $X=0.227 $Y=2.065
+ $X2=0.227 $Y2=2.165
r87 10 18 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.227 $Y=0.615
+ $X2=0.37 $Y2=0.7
r88 10 12 6.87422 $w=2.83e-07 $l=1.7e-07 $layer=LI1_cond $X=0.227 $Y=0.615
+ $X2=0.227 $Y2=0.445
r89 9 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.505 $Y=0.56
+ $X2=1.505 $Y2=0.995
r90 2 16 600 $w=1.7e-07 $l=3.77359e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.165
r91 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%A 1 3 4 6 7 8 9 14
c29 4 0 1.38301e-19 $X=2.265 $Y=1.41
r30 14 16 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=2.265 $Y=1.202
+ $X2=2.515 $Y2=1.202
r31 13 14 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.24 $Y=1.202
+ $X2=2.265 $Y2=1.202
r32 8 9 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.552 $Y=1.16
+ $X2=2.552 $Y2=1.53
r33 8 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.515
+ $Y=1.16 $X2=2.515 $Y2=1.16
r34 7 8 14.5819 $w=2.43e-07 $l=3.1e-07 $layer=LI1_cond $X=2.552 $Y=0.85
+ $X2=2.552 $Y2=1.16
r35 4 14 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.265 $Y=1.41
+ $X2=2.265 $Y2=1.202
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.265 $Y=1.41
+ $X2=2.265 $Y2=1.985
r37 1 13 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.24 $Y=0.995
+ $X2=2.24 $Y2=1.202
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.24 $Y=0.995 $X2=2.24
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%VPWR 1 6 8 10 20 21 24
r27 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r28 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r29 18 21 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r30 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r31 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r32 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 15 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.92 $Y=2.72 $X2=0.73
+ $Y2=2.72
r34 15 17 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.92 $Y=2.72
+ $X2=1.15 $Y2=2.72
r35 10 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.54 $Y=2.72 $X2=0.73
+ $Y2=2.72
r36 10 12 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r37 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r38 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r39 4 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r40 4 6 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.36
r41 1 6 600 $w=1.7e-07 $l=5.93949e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.755 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%Z 1 2 7 9 11 13 14 26 32 39
r37 42 44 7.21165 $w=6.78e-07 $l=4.1e-07 $layer=LI1_cond $X=2.09 $Y=2.125
+ $X2=2.5 $Y2=2.125
r38 14 44 0.439735 $w=6.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.525 $Y=2.125
+ $X2=2.5 $Y2=2.125
r39 13 26 0.847385 $w=3.38e-07 $l=2.5e-08 $layer=LI1_cond $X=2.525 $Y=0.425
+ $X2=2.5 $Y2=0.425
r40 11 42 0.439735 $w=6.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.065 $Y=2.125
+ $X2=2.09 $Y2=2.125
r41 11 42 6.92279 $w=2.4e-07 $l=3.4e-07 $layer=LI1_cond $X=2.09 $Y=1.785
+ $X2=2.09 $Y2=2.125
r42 11 39 0.0879469 $w=6.78e-07 $l=5e-09 $layer=LI1_cond $X=2.065 $Y=2.125
+ $X2=2.06 $Y2=2.125
r43 9 39 8.00317 $w=6.78e-07 $l=4.55e-07 $layer=LI1_cond $X=1.605 $Y=2.125
+ $X2=2.06 $Y2=2.125
r44 9 32 1.75894 $w=6.78e-07 $l=1e-07 $layer=LI1_cond $X=1.605 $Y=2.125
+ $X2=1.505 $Y2=2.125
r45 8 11 34.6007 $w=4.08e-07 $l=1.19e-06 $layer=LI1_cond $X=2.09 $Y=0.595
+ $X2=2.09 $Y2=1.785
r46 7 26 9.82966 $w=3.38e-07 $l=2.9e-07 $layer=LI1_cond $X=2.21 $Y=0.425 $X2=2.5
+ $Y2=0.425
r47 7 8 7.08339 $w=3.4e-07 $l=2.22036e-07 $layer=LI1_cond $X=2.21 $Y=0.425
+ $X2=2.09 $Y2=0.595
r48 2 44 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.355
+ $Y=1.485 $X2=2.5 $Y2=1.96
r49 1 26 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=2.315
+ $Y=0.235 $X2=2.5 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_1%VGND 1 4 16 17 22 28
r28 26 28 15.9104 $w=5.28e-07 $l=4.4e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.59 $Y2=0.18
r29 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 24 26 0.45135 $w=5.28e-07 $l=2e-08 $layer=LI1_cond $X=1.13 $Y=0.18 $X2=1.15
+ $Y2=0.18
r31 21 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r32 20 24 9.92971 $w=5.28e-07 $l=4.4e-07 $layer=LI1_cond $X=0.69 $Y=0.18
+ $X2=1.13 $Y2=0.18
r33 20 22 9.36586 $w=5.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.69 $Y=0.18
+ $X2=0.54 $Y2=0.18
r34 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r35 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r36 14 17 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r37 14 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r38 13 16 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r39 13 28 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.59
+ $Y2=0
r40 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r41 8 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.54
+ $Y2=0
r42 4 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 4 8 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r44 1 24 91 $w=1.7e-07 $l=5.94222e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=1.13 $Y2=0.36
.ends

