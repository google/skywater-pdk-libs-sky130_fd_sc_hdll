* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4_1 A B C D VGND VNB VPB VPWR Y
M1000 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=8.7e+11p pd=7.74e+06u as=6.4e+11p ps=5.28e+06u
M1001 a_213_47# C a_119_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=2.08e+11p ps=1.94e+06u
M1002 Y A a_297_47# VNB nshort w=650000u l=150000u
+  ad=2.275e+11p pd=2e+06u as=2.47e+11p ps=2.06e+06u
M1003 a_297_47# B a_213_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_119_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1007 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
