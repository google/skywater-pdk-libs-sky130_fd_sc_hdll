* File: sky130_fd_sc_hdll__a31o_2.pxi.spice
* Created: Wed Sep  2 08:19:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31O_2%A_79_21# N_A_79_21#_M1002_d N_A_79_21#_M1007_d
+ N_A_79_21#_c_55_n N_A_79_21#_M1001_g N_A_79_21#_c_59_n N_A_79_21#_M1000_g
+ N_A_79_21#_c_60_n N_A_79_21#_M1005_g N_A_79_21#_c_56_n N_A_79_21#_M1009_g
+ N_A_79_21#_c_61_n N_A_79_21#_c_65_p N_A_79_21#_c_106_p N_A_79_21#_c_57_n
+ N_A_79_21#_c_84_p N_A_79_21#_c_85_p N_A_79_21#_c_72_p N_A_79_21#_c_86_p
+ N_A_79_21#_c_58_n PM_SKY130_FD_SC_HDLL__A31O_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__A31O_2%A3 N_A3_c_145_n N_A3_M1008_g N_A3_c_146_n
+ N_A3_M1011_g A3 A3 PM_SKY130_FD_SC_HDLL__A31O_2%A3
x_PM_SKY130_FD_SC_HDLL__A31O_2%A2 N_A2_c_179_n N_A2_M1010_g N_A2_c_180_n
+ N_A2_M1006_g A2 PM_SKY130_FD_SC_HDLL__A31O_2%A2
x_PM_SKY130_FD_SC_HDLL__A31O_2%A1 N_A1_c_209_n N_A1_M1002_g N_A1_c_210_n
+ N_A1_M1004_g A1 PM_SKY130_FD_SC_HDLL__A31O_2%A1
x_PM_SKY130_FD_SC_HDLL__A31O_2%B1 N_B1_c_242_n N_B1_M1007_g N_B1_c_239_n
+ N_B1_M1003_g B1 B1 N_B1_c_241_n PM_SKY130_FD_SC_HDLL__A31O_2%B1
x_PM_SKY130_FD_SC_HDLL__A31O_2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d N_VPWR_M1006_d
+ N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n N_VPWR_c_275_n
+ VPWR N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_270_n N_VPWR_c_279_n
+ N_VPWR_c_280_n PM_SKY130_FD_SC_HDLL__A31O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A31O_2%X N_X_M1001_s N_X_M1000_s N_X_c_331_n N_X_c_342_n
+ N_X_c_347_n N_X_c_349_n X X X X N_X_c_333_n N_X_c_335_n
+ PM_SKY130_FD_SC_HDLL__A31O_2%X
x_PM_SKY130_FD_SC_HDLL__A31O_2%A_305_297# N_A_305_297#_M1008_d
+ N_A_305_297#_M1004_d N_A_305_297#_c_383_n N_A_305_297#_c_390_n
+ N_A_305_297#_c_384_n N_A_305_297#_c_385_n N_A_305_297#_c_388_n
+ PM_SKY130_FD_SC_HDLL__A31O_2%A_305_297#
x_PM_SKY130_FD_SC_HDLL__A31O_2%VGND N_VGND_M1001_d N_VGND_M1009_d N_VGND_M1003_d
+ N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n N_VGND_c_413_n VGND
+ N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n N_VGND_c_417_n
+ PM_SKY130_FD_SC_HDLL__A31O_2%VGND
cc_1 VNB N_A_79_21#_c_55_n 0.0191307f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_56_n 0.0165471f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A_79_21#_c_57_n 0.00324285f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.42
cc_4 VNB N_A_79_21#_c_58_n 0.0375994f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_A3_c_145_n 0.0247825f $X=-0.19 $Y=-0.24 $X2=2.485 $Y2=0.235
cc_6 VNB N_A3_c_146_n 0.0168741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB A3 0.00154476f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_8 VNB N_A2_c_179_n 0.016791f $X=-0.19 $Y=-0.24 $X2=2.485 $Y2=0.235
cc_9 VNB N_A2_c_180_n 0.0236908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A2 0.00280954f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_11 VNB N_A1_c_209_n 0.0186185f $X=-0.19 $Y=-0.24 $X2=2.485 $Y2=0.235
cc_12 VNB N_A1_c_210_n 0.0265701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A1 7.47956e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB N_B1_c_239_n 0.0212215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB B1 0.0230379f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_B1_c_241_n 0.0433701f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_17 VNB N_VPWR_c_270_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_331_n 0.00103514f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_19 VNB X 0.0212588f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.245
cc_20 VNB N_X_c_333_n 0.00764178f $X=-0.19 $Y=-0.24 $X2=3.26 $Y2=1.665
cc_21 VNB N_VGND_c_410_n 0.0102396f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_22 VNB N_VGND_c_411_n 0.0120786f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_23 VNB N_VGND_c_412_n 0.0143677f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_24 VNB N_VGND_c_413_n 0.0184663f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_25 VNB N_VGND_c_414_n 0.0139026f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.495
cc_26 VNB N_VGND_c_415_n 0.052025f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.42
cc_27 VNB N_VGND_c_416_n 0.00872199f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=1.58
cc_28 VNB N_VGND_c_417_n 0.20222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A_79_21#_c_59_n 0.0188133f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_A_79_21#_c_60_n 0.0159335f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_31 VPB N_A_79_21#_c_61_n 0.00155146f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.495
cc_32 VPB N_A_79_21#_c_57_n 0.00175777f $X=-0.19 $Y=1.305 $X2=2.87 $Y2=0.42
cc_33 VPB N_A_79_21#_c_58_n 0.0197989f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_34 VPB N_A3_c_145_n 0.0265631f $X=-0.19 $Y=1.305 $X2=2.485 $Y2=0.235
cc_35 VPB A3 0.00262016f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_36 VPB N_A2_c_180_n 0.0274282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A2 0.00153297f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_38 VPB N_A1_c_210_n 0.0279536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB A1 7.41849e-19 $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_40 VPB N_B1_c_242_n 0.0212613f $X=-0.19 $Y=1.305 $X2=2.485 $Y2=0.235
cc_41 VPB B1 0.00967422f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_42 VPB N_B1_c_241_n 0.0193105f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_43 VPB N_VPWR_c_271_n 0.011108f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_44 VPB N_VPWR_c_272_n 0.00457488f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_45 VPB N_VPWR_c_273_n 0.0023174f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_46 VPB N_VPWR_c_274_n 0.0195799f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_47 VPB N_VPWR_c_275_n 0.00561441f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.58
cc_48 VPB N_VPWR_c_276_n 0.0154084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_277_n 0.0394474f $X=-0.19 $Y=1.305 $X2=0.68 $Y2=1.16
cc_50 VPB N_VPWR_c_270_n 0.0519839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_279_n 0.00426507f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_52 VPB N_VPWR_c_280_n 0.006319f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB X 0.0223432f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.245
cc_54 VPB N_X_c_335_n 0.00784838f $X=-0.19 $Y=1.305 $X2=3.26 $Y2=1.96
cc_55 N_A_79_21#_c_60_n N_A3_c_145_n 0.0243735f $X=0.965 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_56 N_A_79_21#_c_65_p N_A3_c_145_n 0.0167303f $X=2.785 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_57 N_A_79_21#_c_58_n N_A3_c_145_n 0.0258832f $X=0.965 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_58 N_A_79_21#_c_56_n N_A3_c_146_n 0.0206191f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_55_n A3 6.16843e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_56_n A3 0.00708435f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_61_n A3 0.00336796f $X=0.6 $Y=1.495 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_65_p A3 0.0348559f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_72_p A3 0.0123121f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_58_n A3 0.0126526f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_65_p N_A2_c_180_n 0.0156645f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_65_p A2 0.0173292f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_57_n A2 4.17699e-19 $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_57_n N_A1_c_209_n 0.0045847f $X=2.87 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_69 N_A_79_21#_c_65_p N_A1_c_210_n 0.0157082f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_57_n N_A1_c_210_n 0.0051544f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_71 N_A_79_21#_M1002_d A1 0.00528447f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_65_p A1 0.0155046f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_57_n A1 0.0675388f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_57_n N_B1_c_242_n 0.00436023f $X=2.87 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_79_21#_c_84_p N_B1_c_242_n 0.0135581f $X=3.175 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_79_21#_c_85_p N_B1_c_242_n 0.0209477f $X=3.26 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_79_21#_c_86_p N_B1_c_242_n 0.00700657f $X=2.87 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_79_21#_c_57_n N_B1_c_239_n 0.00312459f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_57_n B1 0.0247335f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_84_p B1 0.0128562f $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_57_n N_B1_c_241_n 0.0163471f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_84_p N_B1_c_241_n 0.00576715f $X=3.175 $Y=1.58 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_65_p N_VPWR_M1005_d 0.00366967f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_65_p N_VPWR_M1006_d 0.00854556f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_59_n N_VPWR_c_272_n 0.00337796f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_59_n N_VPWR_c_273_n 7.4903e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_60_n N_VPWR_c_273_n 0.0150044f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_65_p N_VPWR_c_273_n 0.0192076f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_59_n N_VPWR_c_276_n 0.00523784f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_60_n N_VPWR_c_276_n 0.00427505f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_85_p N_VPWR_c_277_n 0.0118139f $X=3.26 $Y=1.96 $X2=0 $Y2=0
cc_92 N_A_79_21#_M1007_d N_VPWR_c_270_n 0.00829902f $X=3.055 $Y=1.485 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_59_n N_VPWR_c_270_n 0.00769802f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_60_n N_VPWR_c_270_n 0.00732977f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_85_p N_VPWR_c_270_n 0.00646998f $X=3.26 $Y=1.96 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_65_p N_X_M1000_s 0.00242592f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_106_p N_X_M1000_s 4.25287e-19 $X=0.685 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_55_n N_X_c_331_n 0.0169534f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_56_n N_X_c_331_n 0.00255012f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_72_p N_X_c_331_n 0.0186002f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_58_n N_X_c_331_n 0.00454345f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_59_n N_X_c_342_n 0.0181701f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_60_n N_X_c_342_n 0.00141217f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_65_p N_X_c_342_n 0.0104749f $X=2.785 $Y=1.58 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_106_p N_X_c_342_n 0.00863034f $X=0.685 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_58_n N_X_c_342_n 3.69869e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_55_n N_X_c_347_n 0.00581948f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_56_n N_X_c_347_n 0.00573592f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_59_n N_X_c_349_n 0.00492036f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_60_n N_X_c_349_n 0.00170979f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_55_n X 0.0179588f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_59_n X 0.0128144f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_61_n X 0.0183937f $X=0.6 $Y=1.495 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_106_p X 0.0137498f $X=0.685 $Y=1.58 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_72_p X 0.0130898f $X=0.68 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_65_p N_A_305_297#_M1008_d 0.00820916f $X=2.785 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_117 N_A_79_21#_c_65_p N_A_305_297#_M1004_d 0.00778023f $X=2.785 $Y=1.58 $X2=0
+ $Y2=0
cc_118 N_A_79_21#_c_86_p N_A_305_297#_M1004_d 3.5412e-19 $X=2.87 $Y=1.58 $X2=0
+ $Y2=0
cc_119 N_A_79_21#_c_65_p N_A_305_297#_c_383_n 0.0191431f $X=2.785 $Y=1.58 $X2=0
+ $Y2=0
cc_120 N_A_79_21#_c_65_p N_A_305_297#_c_384_n 0.0417264f $X=2.785 $Y=1.58 $X2=0
+ $Y2=0
cc_121 N_A_79_21#_c_65_p N_A_305_297#_c_385_n 0.0160491f $X=2.785 $Y=1.58 $X2=0
+ $Y2=0
cc_122 N_A_79_21#_c_85_p N_A_305_297#_c_385_n 0.00908335f $X=3.26 $Y=1.96 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_c_86_p N_A_305_297#_c_385_n 0.00453367f $X=2.87 $Y=1.58 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_c_85_p N_A_305_297#_c_388_n 0.0210128f $X=3.26 $Y=1.96 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_55_n N_VGND_c_411_n 0.00830113f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_56_n N_VGND_c_411_n 4.82686e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_55_n N_VGND_c_414_n 0.00348405f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_56_n N_VGND_c_414_n 0.00351231f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_57_n N_VGND_c_415_n 0.0116048f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_55_n N_VGND_c_416_n 5.13253e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_56_n N_VGND_c_416_n 0.00971119f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_79_21#_M1002_d N_VGND_c_417_n 0.012015f $X=2.485 $Y=0.235 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_55_n N_VGND_c_417_n 0.0043436f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_56_n N_VGND_c_417_n 0.00631413f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_57_n N_VGND_c_417_n 0.00646998f $X=2.87 $Y=0.42 $X2=0 $Y2=0
cc_136 N_A3_c_146_n N_A2_c_179_n 0.0412289f $X=1.46 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_137 N_A3_c_145_n N_A2_c_180_n 0.0474726f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_138 A3 N_A2_c_180_n 0.00113056f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A3_c_145_n A2 0.00101541f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A3_c_146_n A2 0.00244571f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_141 A3 A2 0.0191206f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_142 N_A3_c_145_n N_VPWR_c_273_n 0.00596005f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A3_c_145_n N_VPWR_c_274_n 0.00601503f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A3_c_145_n N_VPWR_c_270_n 0.0100936f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_145 A3 N_X_c_331_n 0.00866452f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_146 N_A3_c_145_n N_A_305_297#_c_383_n 0.00336202f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A3_c_145_n N_A_305_297#_c_390_n 0.00655764f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_148 A3 N_VGND_M1009_d 0.00309516f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A3_c_146_n N_VGND_c_415_n 0.00585385f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A3_c_145_n N_VGND_c_416_n 3.35359e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A3_c_146_n N_VGND_c_416_n 0.00325898f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_152 A3 N_VGND_c_416_n 0.0123749f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A3_c_146_n N_VGND_c_417_n 0.0106542f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_154 A3 N_VGND_c_417_n 0.00179833f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A2_c_179_n N_A1_c_209_n 0.0267356f $X=1.88 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_156 A2 N_A1_c_209_n 0.0064626f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_157 N_A2_c_180_n N_A1_c_210_n 0.0547948f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_179_n A1 5.28842e-19 $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_180_n A1 3.6629e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_160 A2 A1 0.0540197f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_161 N_A2_c_180_n N_VPWR_c_274_n 0.00523784f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_180_n N_VPWR_c_275_n 0.00335717f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_180_n N_VPWR_c_270_n 0.00707245f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_180_n N_A_305_297#_c_384_n 0.0121189f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A2_c_179_n N_VGND_c_415_n 0.00520302f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_166 A2 N_VGND_c_415_n 0.00790477f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_167 A2 N_VGND_c_416_n 0.00219626f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_168 N_A2_c_179_n N_VGND_c_417_n 0.00935289f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_169 A2 N_VGND_c_417_n 0.00855668f $X=1.985 $Y=0.425 $X2=0 $Y2=0
cc_170 A2 A_391_47# 0.00700281f $X=1.985 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_171 N_A1_c_210_n N_B1_c_242_n 0.0275932f $X=2.435 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_172 N_A1_c_209_n N_B1_c_239_n 0.0122621f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A1_c_210_n N_B1_c_241_n 0.0233951f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_174 A1 N_B1_c_241_n 3.28305e-19 $X=2.41 $Y=0.425 $X2=0 $Y2=0
cc_175 N_A1_c_210_n N_VPWR_c_275_n 0.00349223f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A1_c_210_n N_VPWR_c_277_n 0.00522999f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A1_c_210_n N_VPWR_c_270_n 0.0071634f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A1_c_210_n N_A_305_297#_c_384_n 0.0145195f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A1_c_210_n N_A_305_297#_c_388_n 0.00708501f $X=2.435 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A1_c_209_n N_VGND_c_415_n 0.00455696f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_181 A1 N_VGND_c_415_n 0.0067485f $X=2.41 $Y=0.425 $X2=0 $Y2=0
cc_182 N_A1_c_209_n N_VGND_c_417_n 0.00807669f $X=2.41 $Y=0.995 $X2=0 $Y2=0
cc_183 A1 N_VGND_c_417_n 0.00752092f $X=2.41 $Y=0.425 $X2=0 $Y2=0
cc_184 N_B1_c_242_n N_VPWR_c_277_n 0.00674661f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B1_c_242_n N_VPWR_c_270_n 0.0133315f $X=2.965 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B1_c_242_n N_A_305_297#_c_385_n 0.00262889f $X=2.965 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_B1_c_242_n N_A_305_297#_c_388_n 0.00600985f $X=2.965 $Y=1.41 $X2=0
+ $Y2=0
cc_188 B1 N_VGND_M1003_d 0.0029656f $X=3.21 $Y=0.765 $X2=0 $Y2=0
cc_189 B1 N_VGND_c_412_n 0.00109862f $X=3.21 $Y=0.765 $X2=0 $Y2=0
cc_190 N_B1_c_239_n N_VGND_c_413_n 0.00478506f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_191 B1 N_VGND_c_413_n 0.0198424f $X=3.21 $Y=0.765 $X2=0 $Y2=0
cc_192 N_B1_c_241_n N_VGND_c_413_n 9.77692e-19 $X=3.08 $Y=1.202 $X2=0 $Y2=0
cc_193 N_B1_c_239_n N_VGND_c_415_n 0.00585385f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_194 N_B1_c_239_n N_VGND_c_417_n 0.0120436f $X=3.08 $Y=0.995 $X2=0 $Y2=0
cc_195 B1 N_VGND_c_417_n 0.00306869f $X=3.21 $Y=0.765 $X2=0 $Y2=0
cc_196 N_VPWR_c_270_n N_X_M1000_s 0.00467205f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_197 N_VPWR_c_273_n N_X_c_342_n 0.0139456f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_198 N_VPWR_c_276_n N_X_c_342_n 0.00309089f $X=0.985 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_c_270_n N_X_c_342_n 0.0060752f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_273_n N_X_c_349_n 0.0336782f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_201 N_VPWR_c_276_n N_X_c_349_n 0.0117479f $X=0.985 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_270_n N_X_c_349_n 0.00645703f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_M1000_d X 0.00619658f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_204 N_VPWR_M1000_d N_X_c_335_n 0.00308968f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_205 N_VPWR_c_271_n N_X_c_335_n 7.73122e-19 $X=0.26 $Y=2.635 $X2=0 $Y2=0
cc_206 N_VPWR_c_272_n N_X_c_335_n 0.0179856f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_207 N_VPWR_c_270_n N_X_c_335_n 0.00220706f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_208 N_VPWR_c_270_n N_A_305_297#_M1008_d 0.00262984f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_209 N_VPWR_c_270_n N_A_305_297#_M1004_d 0.00311683f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_273_n N_A_305_297#_c_383_n 0.0139118f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_211 N_VPWR_c_273_n N_A_305_297#_c_390_n 0.032099f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_212 N_VPWR_c_274_n N_A_305_297#_c_390_n 0.0148159f $X=2.015 $Y=2.72 $X2=0
+ $Y2=0
cc_213 N_VPWR_c_270_n N_A_305_297#_c_390_n 0.0108685f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_M1006_d N_A_305_297#_c_384_n 0.00487505f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_274_n N_A_305_297#_c_384_n 0.00308517f $X=2.015 $Y=2.72 $X2=0
+ $Y2=0
cc_216 N_VPWR_c_275_n N_A_305_297#_c_384_n 0.0184247f $X=2.18 $Y=2.26 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_277_n N_A_305_297#_c_384_n 0.00293179f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_218 N_VPWR_c_270_n N_A_305_297#_c_384_n 0.0127596f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_219 N_VPWR_c_275_n N_A_305_297#_c_388_n 0.0158699f $X=2.18 $Y=2.26 $X2=0
+ $Y2=0
cc_220 N_VPWR_c_277_n N_A_305_297#_c_388_n 0.0154672f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_221 N_VPWR_c_270_n N_A_305_297#_c_388_n 0.0114786f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_222 N_X_c_333_n N_VGND_M1001_d 0.00334111f $X=0.217 $Y=0.885 $X2=-0.19
+ $Y2=-0.24
cc_223 N_X_c_331_n N_VGND_c_411_n 0.00143691f $X=0.645 $Y=0.8 $X2=0 $Y2=0
cc_224 N_X_c_347_n N_VGND_c_411_n 0.0127288f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_225 N_X_c_333_n N_VGND_c_411_n 0.0151594f $X=0.217 $Y=0.885 $X2=0 $Y2=0
cc_226 N_X_c_331_n N_VGND_c_414_n 0.00271566f $X=0.645 $Y=0.8 $X2=0 $Y2=0
cc_227 N_X_c_347_n N_VGND_c_414_n 0.0117479f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_228 N_X_c_347_n N_VGND_c_416_n 0.0143868f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_229 N_X_M1001_s N_VGND_c_417_n 0.0069264f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_230 N_X_c_331_n N_VGND_c_417_n 0.00559444f $X=0.645 $Y=0.8 $X2=0 $Y2=0
cc_231 N_X_c_347_n N_VGND_c_417_n 0.00645703f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_232 N_X_c_333_n N_VGND_c_417_n 0.0013612f $X=0.217 $Y=0.885 $X2=0 $Y2=0
cc_233 N_VGND_c_417_n A_307_47# 0.0115413f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_234 N_VGND_c_417_n A_391_47# 0.00948296f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
