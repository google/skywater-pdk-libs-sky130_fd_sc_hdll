* File: sky130_fd_sc_hdll__inputiso0p_1.pex.spice
* Created: Thu Aug 27 19:08:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%SLEEP 2 3 5 8 10 11 12 17
c33 17 0 1.89169e-19 $X=0.36 $Y=1.16
c34 10 0 1.01663e-19 $X=0.23 $Y=0.85
r35 17 20 36.8359 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=1.325
r36 17 19 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=0.995
r37 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r38 11 12 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.53
r39 11 18 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.16
r40 10 18 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.295 $Y=0.85
+ $X2=0.295 $Y2=1.16
r41 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.445
+ $X2=0.52 $Y2=0.995
r42 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r43 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r44 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_27_413# 1 2 8 9 11 12 16 20 22 23
+ 26 29 34 37
c71 37 0 1.01663e-19 $X=1 $Y=0.88
c72 22 0 1.89169e-19 $X=0.645 $Y=1.9
c73 12 0 1.77329e-20 $X=1.385 $Y=0.88
r74 35 40 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1 $Y=0.97 $X2=1
+ $Y2=1.135
r75 35 37 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1 $Y=0.97 $X2=1
+ $Y2=0.88
r76 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=0.97
+ $X2=1 $Y2=0.97
r77 32 34 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=0.77 $Y=0.97 $X2=1
+ $Y2=0.97
r78 30 32 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.765 $Y=0.97
+ $X2=0.77 $Y2=0.97
r79 28 32 2.36532 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=0.77 $Y=1.135
+ $X2=0.77 $Y2=0.97
r80 28 29 29.9635 $w=2.48e-07 $l=6.5e-07 $layer=LI1_cond $X=0.77 $Y=1.135
+ $X2=0.77 $Y2=1.785
r81 24 30 2.60351 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=0.805
+ $X2=0.765 $Y2=0.97
r82 24 26 17.2866 $w=2.38e-07 $l=3.6e-07 $layer=LI1_cond $X=0.765 $Y=0.805
+ $X2=0.765 $Y2=0.445
r83 22 29 6.8319 $w=2.3e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.645 $Y=1.9
+ $X2=0.77 $Y2=1.785
r84 22 23 15.0319 $w=2.28e-07 $l=3e-07 $layer=LI1_cond $X=0.645 $Y=1.9 $X2=0.345
+ $Y2=1.9
r85 18 23 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.345 $Y2=1.9
r86 18 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=2.225
r87 14 16 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.46 $Y=0.805
+ $X2=1.46 $Y2=0.445
r88 13 37 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.135 $Y=0.88 $X2=1
+ $Y2=0.88
r89 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.385 $Y=0.88
+ $X2=1.46 $Y2=0.805
r90 12 13 128.191 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=1.385 $Y=0.88
+ $X2=1.135 $Y2=0.88
r91 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.965 $Y=1.99
+ $X2=0.965 $Y2=2.275
r92 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.89 $X2=0.965
+ $Y2=1.99
r93 8 40 250.341 $w=2e-07 $l=7.55e-07 $layer=POLY_cond $X=0.965 $Y=1.89
+ $X2=0.965 $Y2=1.135
r94 2 20 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.225
r95 1 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A 1 3 6 8 12 16
c38 8 0 1.77329e-20 $X=1.605 $Y=1.785
r39 13 16 4.83283 $w=3.08e-07 $l=1.3e-07 $layer=LI1_cond $X=1.67 $Y=1.8 $X2=1.54
+ $Y2=1.8
r40 12 14 19.8082 $w=3.65e-07 $l=1.5e-07 $layer=POLY_cond $X=1.67 $Y=1.777
+ $X2=1.82 $Y2=1.777
r41 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.73 $X2=1.67 $Y2=1.73
r42 10 12 28.3918 $w=3.65e-07 $l=2.15e-07 $layer=POLY_cond $X=1.455 $Y=1.777
+ $X2=1.67 $Y2=1.777
r43 8 13 0.743512 $w=3.08e-07 $l=2e-08 $layer=LI1_cond $X=1.69 $Y=1.8 $X2=1.67
+ $Y2=1.8
r44 4 14 23.6381 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=1.82 $Y=1.565
+ $X2=1.82 $Y2=1.777
r45 4 6 574.298 $w=1.5e-07 $l=1.12e-06 $layer=POLY_cond $X=1.82 $Y=1.565
+ $X2=1.82 $Y2=0.445
r46 1 10 19.2931 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=1.455 $Y=1.99
+ $X2=1.455 $Y2=1.777
r47 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.455 $Y=1.99
+ $X2=1.455 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%A_211_413# 1 2 7 9 10 12 15 18 19 21
+ 27
r56 27 28 10.6087 $w=2.53e-07 $l=2.2e-07 $layer=LI1_cond $X=1.25 $Y=0.44
+ $X2=1.47 $Y2=0.44
r57 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.39
+ $Y=1.16 $X2=2.39 $Y2=1.16
r58 19 25 12.5903 $w=4.04e-07 $l=4.50943e-07 $layer=LI1_cond $X=1.885 $Y=1.135
+ $X2=1.47 $Y2=1.21
r59 19 21 15.3154 $w=3.78e-07 $l=5.05e-07 $layer=LI1_cond $X=1.885 $Y=1.135
+ $X2=2.39 $Y2=1.135
r60 18 25 3.784 $w=2.4e-07 $l=2.65e-07 $layer=LI1_cond $X=1.47 $Y=0.945 $X2=1.47
+ $Y2=1.21
r61 17 28 1.0361 $w=2.4e-07 $l=1.7e-07 $layer=LI1_cond $X=1.47 $Y=0.61 $X2=1.47
+ $Y2=0.44
r62 17 18 16.0862 $w=2.38e-07 $l=3.35e-07 $layer=LI1_cond $X=1.47 $Y=0.61
+ $X2=1.47 $Y2=0.945
r63 13 25 8.15347 $w=4.04e-07 $l=3.80066e-07 $layer=LI1_cond $X=1.2 $Y=1.475
+ $X2=1.47 $Y2=1.21
r64 13 15 32.0123 $w=2.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.2 $Y=1.475 $X2=1.2
+ $Y2=2.225
r65 10 22 40.2498 $w=2.92e-07 $l=2.12485e-07 $layer=POLY_cond $X=2.495 $Y=0.985
+ $X2=2.412 $Y2=1.16
r66 10 12 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.495 $Y=0.985
+ $X2=2.495 $Y2=0.56
r67 7 22 48.3126 $w=2.92e-07 $l=2.77489e-07 $layer=POLY_cond $X=2.47 $Y=1.41
+ $X2=2.412 $Y2=1.16
r68 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.47 $Y=1.41 $X2=2.47
+ $Y2=1.985
r69 2 15 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=2.065 $X2=1.21 $Y2=2.225
r70 1 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VPWR 1 2 9 13 15 22 23 26 31 37
r39 35 37 12.0988 $w=6.38e-07 $l=2.55e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=2.325 $Y2=2.485
r40 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 33 35 6.16728 $w=6.38e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.485
+ $X2=2.07 $Y2=2.485
r42 30 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 29 33 2.42953 $w=6.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=2.485
+ $X2=1.74 $Y2=2.485
r44 29 31 8.17421 $w=6.38e-07 $l=4.5e-08 $layer=LI1_cond $X=1.61 $Y=2.485
+ $X2=1.565 $Y2=2.485
r45 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r46 27 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r47 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 23 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r49 22 37 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.325 $Y2=2.72
r50 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r51 15 26 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r52 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 13 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 12 26 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r56 12 31 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.565 $Y2=2.72
r57 7 26 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r58 7 9 11.0695 $w=3.78e-07 $l=3.65e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.27
r59 2 33 600 $w=1.7e-07 $l=3.49142e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=2.065 $X2=1.74 $Y2=2.33
r60 1 9 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%X 1 2 9 10 11 22
r16 19 22 51.0182 $w=1.73e-07 $l=8.05e-07 $layer=LI1_cond $X=2.992 $Y=0.775
+ $X2=2.992 $Y2=1.58
r17 10 11 7.80051 $w=5.73e-07 $l=3.75e-07 $layer=LI1_cond $X=2.792 $Y=1.835
+ $X2=2.792 $Y2=2.21
r18 10 22 11.6583 $w=5.73e-07 $l=2.55e-07 $layer=LI1_cond $X=2.792 $Y=1.835
+ $X2=2.792 $Y2=1.58
r19 9 19 11.6809 $w=4.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.85 $Y=0.51
+ $X2=2.85 $Y2=0.775
r20 2 10 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=2.56
+ $Y=1.485 $X2=2.705 $Y2=1.835
r21 1 9 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.57
+ $Y=0.235 $X2=2.705 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__INPUTISO0P_1%VGND 1 2 7 9 13 15 17 24 25 31
r35 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r36 25 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r37 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r38 22 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.235
+ $Y2=0
r39 22 24 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=2.4 $Y=0 $X2=2.99
+ $Y2=0
r40 21 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r41 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r42 18 28 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r43 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r44 17 31 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.235
+ $Y2=0
r45 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=0.69
+ $Y2=0
r46 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r47 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r48 11 31 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0
r49 11 13 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.235 $Y=0.085
+ $X2=2.235 $Y2=0.47
r50 7 28 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r51 7 9 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.445
r52 2 13 182 $w=1.7e-07 $l=4.42154e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.235 $Y2=0.47
r53 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

