# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__ebufn_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__ebufn_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.430000 1.615000 ;
    END
  END A
  PIN TE_B
    ANTENNAGATEAREA  1.631100 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.020000 0.620000 1.405000 0.995000 ;
        RECT 1.020000 0.995000 1.530000 1.325000 ;
        RECT 1.020000 1.325000 1.405000 1.695000 ;
    END
  END TE_B
  PIN VGND
    ANTENNADIFFAREA  1.417000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 11.040000 0.085000 ;
        RECT 0.085000  0.085000  0.445000 0.825000 ;
        RECT 1.020000  0.085000  1.405000 0.445000 ;
        RECT 2.855000  0.085000  3.285000 0.485000 ;
        RECT 3.895000  0.085000  4.325000 0.485000 ;
        RECT 4.935000  0.085000  5.365000 0.485000 ;
        RECT 5.975000  0.085000  6.405000 0.485000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.958400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 11.040000 2.805000 ;
        RECT 0.085000 1.785000  0.445000 2.635000 ;
        RECT 1.020000 1.865000  1.405000 2.635000 ;
        RECT 2.565000 2.235000  2.995000 2.635000 ;
        RECT 3.605000 2.235000  4.035000 2.635000 ;
        RECT 4.645000 2.235000  5.075000 2.635000 ;
        RECT 5.685000 2.235000  6.115000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  2.145000 1.445000 10.925000 1.725000 ;
        RECT  7.225000 0.615000 10.925000 0.855000 ;
        RECT 10.675000 0.855000 10.925000 1.445000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT 0.650000 0.280000  0.850000 1.615000 ;
      RECT 0.665000 1.615000  0.850000 2.465000 ;
      RECT 1.575000 0.255000  2.135000 0.825000 ;
      RECT 1.575000 1.495000  1.975000 2.465000 ;
      RECT 1.750000 0.825000  2.135000 1.025000 ;
      RECT 1.750000 1.025000  6.875000 1.275000 ;
      RECT 1.750000 1.275000  1.975000 1.495000 ;
      RECT 2.145000 1.895000 10.925000 2.065000 ;
      RECT 2.145000 2.065000  2.395000 2.465000 ;
      RECT 2.305000 0.255000  2.685000 0.655000 ;
      RECT 2.305000 0.655000  7.055000 0.855000 ;
      RECT 3.215000 2.065000  3.385000 2.465000 ;
      RECT 3.505000 0.275000  3.725000 0.655000 ;
      RECT 4.255000 2.065000  4.425000 2.465000 ;
      RECT 4.545000 0.255000  4.765000 0.655000 ;
      RECT 5.295000 2.065000  5.465000 2.465000 ;
      RECT 5.585000 0.275000  5.805000 0.655000 ;
      RECT 6.335000 2.065000 10.925000 2.465000 ;
      RECT 6.625000 0.255000 10.925000 0.445000 ;
      RECT 6.625000 0.445000  7.055000 0.655000 ;
      RECT 7.125000 1.025000 10.455000 1.275000 ;
    LAYER mcon ;
      RECT 0.655000 1.060000 0.825000 1.230000 ;
      RECT 7.630000 1.060000 7.800000 1.230000 ;
    LAYER met1 ;
      RECT 0.545000 1.030000 0.885000 1.120000 ;
      RECT 0.545000 1.120000 7.860000 1.260000 ;
      RECT 7.520000 1.030000 7.860000 1.120000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__ebufn_8
