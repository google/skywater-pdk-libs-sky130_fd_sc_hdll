* File: sky130_fd_sc_hdll__and3b_1.spice
* Created: Wed Sep  2 08:22:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and3b_1.pex.spice"
.subckt sky130_fd_sc_hdll__and3b_1  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_117_413#_M1006_d N_A_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 A_317_53# N_A_117_413#_M1000_g N_A_225_311#_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1197 PD=0.74 PS=1.41 NRD=30 NRS=5.712 M=1 R=2.8
+ SA=75000.2 SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 A_411_53# N_B_M1007_g A_317_53# VNB NSHORT L=0.15 W=0.42 AD=0.05355
+ AS=0.0672 PD=0.675 PS=0.74 NRD=20.712 NRS=30 M=1 R=2.8 SA=75000.7 SB=75001.4
+ A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_C_M1009_g A_411_53# VNB NSHORT L=0.15 W=0.42 AD=0.133556
+ AS=0.05355 PD=1.00093 PS=0.675 NRD=97.14 NRS=20.712 M=1 R=2.8 SA=75001.1
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_225_311#_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.206694 PD=1.82 PS=1.54907 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75001.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_117_413#_M1002_d N_A_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_117_413#_M1005_g N_A_225_311#_M1005_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1003 N_A_225_311#_M1003_d N_B_M1003_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.078575 AS=0.0609 PD=0.835 PS=0.71 NRD=25.7873 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_C_M1004_g N_A_225_311#_M1003_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.105325 AS=0.078575 PD=0.872535 PS=0.835 NRD=91.8217 NRS=4.6886 M=1
+ R=2.33333 SA=90001 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1008 N_X_M1008_d N_A_225_311#_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.250775 PD=2.54 PS=2.07746 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_13 B B PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and3b_1.pxi.spice"
*
.ends
*
*
