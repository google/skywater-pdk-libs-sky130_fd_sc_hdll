* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb16to1_4 D[15] D[14] D[13] D[12] D[11] D[10] D[9] D[8]
+ D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[15] S[14] S[13] S[12] S[11] S[10] S[9]
+ S[8] S[7] S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
X0 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Z S[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 VGND D[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_9250_599# S[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X4 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR D[7] a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_6937_918# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X8 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND D[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Z a_4006_599# a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 VPWR D[13] a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_6937_66# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z S[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X15 Z S[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X16 VGND S[8] a_559_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X18 Z a_9250_599# a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 a_7939_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 VPWR S[8] a_559_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X21 VGND D[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND D[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR D[12] a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Z a_8379_265# a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X25 VGND D[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_4269_918# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Z S[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X28 Z a_3135_793# a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X29 Z a_5803_793# a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X30 a_559_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_7939_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_117_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VPWR D[11] a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_1430_599# S[9] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X36 a_3135_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 a_7937_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 a_9463_613# a_9250_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X40 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 a_9463_311# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X44 Z a_559_793# a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X45 a_5361_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 VPWR S[14] a_8379_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X47 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X48 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_559_793# S[8] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X51 a_2693_591# a_3135_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X52 VGND S[3] a_4006_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X53 VPWR D[8] a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 Z S[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 a_4219_613# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X56 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 a_3135_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X58 Z S[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X59 VGND S[14] a_8379_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X60 a_2695_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X61 a_9463_613# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 VPWR D[6] a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X63 Z S[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 VGND S[13] a_6674_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X65 a_4269_918# D[11] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X66 Z S[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X67 Z S[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X68 a_117_591# a_559_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_1430_325# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X70 a_6887_311# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X71 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X72 a_2693_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X73 VPWR S[2] a_3135_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X74 VGND S[0] a_559_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X75 Z a_6674_599# a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X77 VGND S[12] a_5803_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X78 a_4006_599# S[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X79 VGND S[4] a_5803_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X80 a_6674_325# S[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X81 a_5803_793# S[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X82 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X83 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X84 Z S[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X85 VPWR D[5] a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X86 a_4006_325# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X87 VPWR D[9] a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X88 VGND D[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X89 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X90 a_5361_297# a_5803_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X91 a_4006_599# S[11] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X92 VPWR D[10] a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X93 a_8379_793# S[14] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X94 a_6937_66# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X95 a_9250_325# S[7] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X96 Z S[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X97 a_1643_613# a_1430_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X98 a_9513_66# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X99 VGND D[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X100 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X101 a_6937_66# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X102 VPWR S[5] a_6674_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X103 VPWR S[12] a_5803_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X104 VPWR D[14] a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X105 VPWR D[4] a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X106 Z a_8379_793# a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X107 VGND D[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X108 a_5363_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X109 Z S[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X110 a_9513_918# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X111 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X112 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X113 VPWR S[15] a_9250_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X114 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X115 a_559_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X116 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X117 VGND D[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X118 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X119 a_5361_297# a_5803_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X120 Z S[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X121 VGND S[15] a_9250_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X122 VGND D[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X123 a_4219_613# a_4006_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X124 a_7939_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 a_6887_613# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X126 Z a_3135_793# a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X127 VPWR S[3] a_4006_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X128 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X129 a_5361_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X130 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X131 VGND D[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X132 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X133 a_8379_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X134 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X135 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X136 VGND S[7] a_9250_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X137 Z S[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X138 Z a_5803_265# a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X139 a_9513_918# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 a_9463_311# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X141 a_7937_297# a_8379_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X142 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X143 VGND S[1] a_1430_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X144 a_9463_311# a_9250_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X145 a_6937_918# S[13] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X146 a_7937_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X147 a_9513_918# D[15] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X148 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X149 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 VGND S[9] a_1430_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X151 a_9250_599# S[15] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X152 VGND S[2] a_3135_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X153 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X154 a_2695_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X155 VPWR D[12] a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X156 VGND D[10] a_2695_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X157 a_6887_311# a_6674_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X158 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X159 a_117_591# D[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X160 a_2693_591# D[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X161 VPWR D[11] a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X162 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X163 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X164 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X165 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X166 a_1693_918# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X167 a_6937_918# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X168 a_5361_591# a_5803_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X169 Z S[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X170 VPWR D[15] a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X171 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X172 a_3135_793# S[10] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X173 Z a_559_793# a_117_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X174 VPWR S[1] a_1430_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X175 a_6674_325# S[5] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X176 VPWR D[6] a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X177 a_7939_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X178 a_5803_265# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X179 Z a_6674_325# a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X180 a_3135_793# S[10] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X181 VGND D[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X182 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X183 a_8379_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X184 Z S[8] a_119_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X185 a_1430_599# S[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X186 a_4219_613# D[11] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X187 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X188 Z a_9250_325# a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X189 a_7939_911# S[14] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X190 a_2695_911# D[10] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X191 VPWR S[10] a_3135_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X192 Z a_4006_599# a_4219_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X193 a_5361_591# a_5803_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X194 a_9250_325# S[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X195 a_6887_311# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X196 a_1643_613# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X197 a_6674_599# S[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X198 Z S[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X199 a_5363_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X200 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X201 a_6887_311# a_6674_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X202 a_9513_918# S[15] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X203 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X204 a_9513_66# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X205 Z a_1430_599# a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X206 VGND D[11] a_4269_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X207 a_7939_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X208 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X209 a_6937_918# D[13] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X210 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X211 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X212 Z S[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X213 Z a_8379_265# a_7937_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X214 VGND D[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X215 a_4269_918# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X216 Z S[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X217 Z a_5803_793# a_5361_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X218 VPWR D[9] a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X219 VPWR S[13] a_6674_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X220 a_7937_591# a_8379_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X221 a_119_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X222 VPWR S[0] a_559_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X223 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X224 Z S[6] a_7939_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X225 a_7937_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X226 VGND D[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X227 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X228 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X229 a_7939_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X230 a_1643_613# a_1430_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X231 VGND D[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X232 a_9463_613# a_9250_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X233 VGND S[6] a_8379_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X234 a_559_793# S[8] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X235 a_5361_591# D[12] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X236 VPWR D[13] a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X237 a_7937_297# a_8379_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X238 VPWR D[4] a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X239 a_2693_591# a_3135_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X240 a_1693_918# S[9] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X241 a_5363_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X242 a_6887_613# a_6674_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X243 Z S[15] a_9513_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X244 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X245 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X246 VPWR S[11] a_4006_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X247 a_7939_911# D[14] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X248 VPWR D[15] a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X249 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X250 VPWR S[6] a_8379_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X251 a_5363_47# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X252 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X253 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X254 a_9513_66# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X255 VGND D[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X256 a_1430_325# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X257 VPWR D[7] a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X258 a_1693_918# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X259 a_8379_793# S[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X260 VGND D[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X261 a_9513_66# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X262 Z a_9250_325# a_9463_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X263 Z a_6674_599# a_6887_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X264 a_5363_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X265 a_5363_47# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X266 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X267 VGND D[12] a_5363_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X268 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X269 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X270 Z a_5803_265# a_5361_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X271 a_119_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X272 VGND S[11] a_4006_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X273 a_6674_599# S[13] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X274 Z a_9250_599# a_9463_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X275 Z S[9] a_1693_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X276 VPWR D[10] a_2693_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X277 VGND D[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X278 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X279 a_4006_325# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X280 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X281 a_9463_311# a_9250_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X282 a_5803_265# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X283 a_5803_793# S[12] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X284 a_7937_591# D[14] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X285 a_2695_911# S[10] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X286 a_6887_613# a_6674_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X287 a_9463_613# D[15] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X288 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X289 VGND D[4] a_5363_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X290 Z S[13] a_6937_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X291 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X292 VGND D[7] a_9513_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X293 a_1693_918# D[9] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X294 VGND S[10] a_3135_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X295 a_117_591# a_559_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X296 a_6937_66# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X297 Z a_8379_793# a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X298 Z S[5] a_6937_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X299 a_119_911# S[8] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X300 a_1643_613# D[9] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X301 VGND S[5] a_6674_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X302 a_4269_918# S[11] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X303 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X304 VPWR S[9] a_1430_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X305 VPWR S[4] a_5803_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X306 Z a_1430_599# a_1643_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X307 VPWR D[14] a_7937_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X308 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X309 a_5363_911# D[12] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X310 a_4219_613# a_4006_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X311 a_6887_613# D[13] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X312 a_119_911# D[8] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X313 VPWR S[7] a_9250_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X314 VPWR D[5] a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X315 a_5361_297# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X316 a_5363_911# S[12] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X317 a_7937_591# a_8379_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X318 VGND D[14] a_7939_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X319 Z a_6674_325# a_6887_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
