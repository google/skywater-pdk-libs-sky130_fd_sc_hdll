* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=3.9325e+11p ps=3.81e+06u
M1001 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A2 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.2e+11p pd=5.84e+06u as=2.3e+11p ps=2.46e+06u
M1003 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=6.2e+11p pd=5.24e+06u as=0p ps=0u
M1004 Y C1 a_304_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=2.46e+06u as=2.4375e+11p ps=2.05e+06u
M1005 a_118_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_304_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
