* File: sky130_fd_sc_hdll__diode_4.spice
* Created: Thu Aug 27 19:05:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__diode_4.pex.spice"
.subckt sky130_fd_sc_hdll__diode_4  VNB VPB DIODE VGND VPWR
* 
* DIODE	DIODE
* VPB	VPB
* VNB	VNB
D0_noxref VNB N_DIODE_D0_noxref_neg NDIODE  AREA=1.0557 PJ=4.44 M=1
+ AHFTEMPPERIM=4.44
DX1_noxref VNB VPB NWDIODE A=3.5631 P=7.65
*
.include "sky130_fd_sc_hdll__diode_4.pxi.spice"
*
.ends
*
*
