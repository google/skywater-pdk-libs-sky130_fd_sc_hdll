* File: sky130_fd_sc_hdll__inv_16.pxi.spice
* Created: Wed Sep  2 08:32:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_16%A N_A_c_128_n N_A_M1000_g N_A_c_110_n N_A_M1004_g
+ N_A_c_129_n N_A_M1001_g N_A_c_111_n N_A_M1006_g N_A_c_130_n N_A_M1002_g
+ N_A_c_112_n N_A_M1007_g N_A_c_131_n N_A_M1003_g N_A_c_113_n N_A_M1008_g
+ N_A_c_132_n N_A_M1005_g N_A_c_114_n N_A_M1009_g N_A_c_133_n N_A_M1010_g
+ N_A_c_115_n N_A_M1014_g N_A_c_134_n N_A_M1011_g N_A_c_116_n N_A_M1016_g
+ N_A_c_135_n N_A_M1012_g N_A_c_117_n N_A_M1017_g N_A_c_136_n N_A_M1013_g
+ N_A_c_118_n N_A_M1019_g N_A_c_137_n N_A_M1015_g N_A_c_119_n N_A_M1021_g
+ N_A_c_138_n N_A_M1018_g N_A_c_120_n N_A_M1023_g N_A_c_139_n N_A_M1020_g
+ N_A_c_121_n N_A_M1025_g N_A_c_140_n N_A_M1022_g N_A_c_122_n N_A_M1026_g
+ N_A_c_141_n N_A_M1024_g N_A_c_123_n N_A_M1027_g N_A_c_142_n N_A_M1028_g
+ N_A_c_124_n N_A_M1029_g N_A_c_143_n N_A_M1031_g N_A_c_125_n N_A_M1030_g A A A
+ A A A N_A_c_126_n N_A_c_127_n A A A A A PM_SKY130_FD_SC_HDLL__INV_16%A
x_PM_SKY130_FD_SC_HDLL__INV_16%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_M1010_d N_VPWR_M1012_d N_VPWR_M1015_d N_VPWR_M1020_d N_VPWR_M1024_d
+ N_VPWR_M1031_d N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n
+ N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n N_VPWR_c_407_n N_VPWR_c_408_n
+ N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n N_VPWR_c_412_n N_VPWR_c_413_n
+ N_VPWR_c_414_n N_VPWR_c_415_n N_VPWR_c_416_n N_VPWR_c_417_n N_VPWR_c_418_n
+ N_VPWR_c_419_n N_VPWR_c_420_n N_VPWR_c_421_n N_VPWR_c_422_n N_VPWR_c_423_n
+ N_VPWR_c_424_n N_VPWR_c_425_n VPWR N_VPWR_c_426_n N_VPWR_c_399_n
+ PM_SKY130_FD_SC_HDLL__INV_16%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_16%Y N_Y_M1004_d N_Y_M1007_d N_Y_M1009_d N_Y_M1016_d
+ N_Y_M1019_d N_Y_M1023_d N_Y_M1026_d N_Y_M1029_d N_Y_M1000_s N_Y_M1002_s
+ N_Y_M1005_s N_Y_M1011_s N_Y_M1013_s N_Y_M1018_s N_Y_M1022_s N_Y_M1028_s
+ N_Y_c_549_n N_Y_c_550_n N_Y_c_554_n N_Y_c_533_n N_Y_c_534_n N_Y_c_564_n
+ N_Y_c_568_n N_Y_c_570_n N_Y_c_535_n N_Y_c_578_n N_Y_c_582_n N_Y_c_584_n
+ N_Y_c_536_n N_Y_c_592_n N_Y_c_596_n N_Y_c_598_n N_Y_c_537_n N_Y_c_606_n
+ N_Y_c_610_n N_Y_c_612_n N_Y_c_538_n N_Y_c_620_n N_Y_c_624_n N_Y_c_626_n
+ N_Y_c_539_n N_Y_c_634_n N_Y_c_638_n N_Y_c_640_n N_Y_c_540_n N_Y_c_646_n
+ N_Y_c_648_n N_Y_c_650_n N_Y_c_541_n N_Y_c_656_n N_Y_c_542_n N_Y_c_663_n
+ N_Y_c_543_n N_Y_c_670_n N_Y_c_544_n N_Y_c_677_n N_Y_c_545_n N_Y_c_684_n
+ N_Y_c_546_n N_Y_c_690_n N_Y_c_693_n Y Y PM_SKY130_FD_SC_HDLL__INV_16%Y
x_PM_SKY130_FD_SC_HDLL__INV_16%VGND N_VGND_M1004_s N_VGND_M1006_s N_VGND_M1008_s
+ N_VGND_M1014_s N_VGND_M1017_s N_VGND_M1021_s N_VGND_M1025_s N_VGND_M1027_s
+ N_VGND_M1030_s N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n N_VGND_c_831_n
+ N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n N_VGND_c_836_n
+ N_VGND_c_837_n N_VGND_c_838_n N_VGND_c_839_n N_VGND_c_840_n N_VGND_c_841_n
+ N_VGND_c_842_n N_VGND_c_843_n N_VGND_c_844_n N_VGND_c_845_n N_VGND_c_846_n
+ N_VGND_c_847_n N_VGND_c_848_n N_VGND_c_849_n N_VGND_c_850_n N_VGND_c_851_n
+ N_VGND_c_852_n N_VGND_c_853_n VGND N_VGND_c_854_n N_VGND_c_855_n
+ PM_SKY130_FD_SC_HDLL__INV_16%VGND
cc_1 VNB N_A_c_110_n 0.0223575f $X=-0.19 $Y=-0.24 $X2=0.585 $Y2=0.995
cc_2 VNB N_A_c_111_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_3 VNB N_A_c_112_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.995
cc_4 VNB N_A_c_113_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=0.995
cc_5 VNB N_A_c_114_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=0.995
cc_6 VNB N_A_c_115_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=0.995
cc_7 VNB N_A_c_116_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=0.995
cc_8 VNB N_A_c_117_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=3.875 $Y2=0.995
cc_9 VNB N_A_c_118_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=4.345 $Y2=0.995
cc_10 VNB N_A_c_119_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=4.815 $Y2=0.995
cc_11 VNB N_A_c_120_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=5.285 $Y2=0.995
cc_12 VNB N_A_c_121_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=5.755 $Y2=0.995
cc_13 VNB N_A_c_122_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=6.225 $Y2=0.995
cc_14 VNB N_A_c_123_n 0.0167268f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.995
cc_15 VNB N_A_c_124_n 0.015981f $X=-0.19 $Y=-0.24 $X2=7.165 $Y2=0.995
cc_16 VNB N_A_c_125_n 0.0224185f $X=-0.19 $Y=-0.24 $X2=7.635 $Y2=0.995
cc_17 VNB N_A_c_126_n 0.0109395f $X=-0.19 $Y=-0.24 $X2=5.96 $Y2=1.16
cc_18 VNB N_A_c_127_n 0.340452f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.202
cc_19 VNB N_VPWR_c_399_n 0.345644f $X=-0.19 $Y=-0.24 $X2=1.995 $Y2=1.202
cc_20 VNB N_Y_c_533_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=4.79 $Y2=1.985
cc_21 VNB N_Y_c_534_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=4.815 $Y2=0.995
cc_22 VNB N_Y_c_535_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=5.73 $Y2=1.985
cc_23 VNB N_Y_c_536_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=6.67 $Y2=1.985
cc_24 VNB N_Y_c_537_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.985
cc_25 VNB N_Y_c_538_n 0.00264996f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_539_n 0.00277027f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.202
cc_27 VNB N_Y_c_540_n 0.00286256f $X=-0.19 $Y=-0.24 $X2=4.345 $Y2=1.202
cc_28 VNB N_Y_c_541_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.202
cc_29 VNB N_Y_c_542_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=7.635 $Y2=1.202
cc_30 VNB N_Y_c_543_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_544_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=1.255 $Y2=1.19
cc_32 VNB N_Y_c_545_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=2.29 $Y2=1.19
cc_33 VNB N_Y_c_546_n 0.00335997f $X=-0.19 $Y=-0.24 $X2=3.295 $Y2=1.19
cc_34 VNB Y 0.00216435f $X=-0.19 $Y=-0.24 $X2=4.845 $Y2=1.19
cc_35 VNB N_VGND_c_828_n 0.0123634f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=0.995
cc_36 VNB N_VGND_c_829_n 0.0299645f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=0.56
cc_37 VNB N_VGND_c_830_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=2.935 $Y2=0.995
cc_38 VNB N_VGND_c_831_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=3.38 $Y2=1.985
cc_39 VNB N_VGND_c_832_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=3.405 $Y2=0.56
cc_40 VNB N_VGND_c_833_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=3.875 $Y2=0.995
cc_41 VNB N_VGND_c_834_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=4.32 $Y2=1.985
cc_42 VNB N_VGND_c_835_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=4.345 $Y2=0.56
cc_43 VNB N_VGND_c_836_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=4.815 $Y2=0.995
cc_44 VNB N_VGND_c_837_n 0.0131823f $X=-0.19 $Y=-0.24 $X2=5.26 $Y2=1.985
cc_45 VNB N_VGND_c_838_n 0.0198983f $X=-0.19 $Y=-0.24 $X2=5.285 $Y2=0.56
cc_46 VNB N_VGND_c_839_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=5.285 $Y2=0.56
cc_47 VNB N_VGND_c_840_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=5.73 $Y2=1.985
cc_48 VNB N_VGND_c_841_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=5.73 $Y2=1.985
cc_49 VNB N_VGND_c_842_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=5.755 $Y2=0.56
cc_50 VNB N_VGND_c_843_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=5.755 $Y2=0.56
cc_51 VNB N_VGND_c_844_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=6.2 $Y2=1.985
cc_52 VNB N_VGND_c_845_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=6.2 $Y2=1.985
cc_53 VNB N_VGND_c_846_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=6.225 $Y2=0.56
cc_54 VNB N_VGND_c_847_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=6.225 $Y2=0.56
cc_55 VNB N_VGND_c_848_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=6.67 $Y2=1.985
cc_56 VNB N_VGND_c_849_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=6.67 $Y2=1.985
cc_57 VNB N_VGND_c_850_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.56
cc_58 VNB N_VGND_c_851_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=6.695 $Y2=0.56
cc_59 VNB N_VGND_c_852_n 0.0200866f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.985
cc_60 VNB N_VGND_c_853_n 0.0040393f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.985
cc_61 VNB N_VGND_c_854_n 0.0120081f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.202
cc_62 VNB N_VGND_c_855_n 0.401764f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.202
cc_63 VPB N_A_c_128_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.41
cc_64 VPB N_A_c_129_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_65 VPB N_A_c_130_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.41
cc_66 VPB N_A_c_131_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.41
cc_67 VPB N_A_c_132_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.44 $Y2=1.41
cc_68 VPB N_A_c_133_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.91 $Y2=1.41
cc_69 VPB N_A_c_134_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.38 $Y2=1.41
cc_70 VPB N_A_c_135_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.85 $Y2=1.41
cc_71 VPB N_A_c_136_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.32 $Y2=1.41
cc_72 VPB N_A_c_137_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.79 $Y2=1.41
cc_73 VPB N_A_c_138_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.26 $Y2=1.41
cc_74 VPB N_A_c_139_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.73 $Y2=1.41
cc_75 VPB N_A_c_140_n 0.0162635f $X=-0.19 $Y=1.305 $X2=6.2 $Y2=1.41
cc_76 VPB N_A_c_141_n 0.0162499f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_77 VPB N_A_c_142_n 0.0155986f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.41
cc_78 VPB N_A_c_143_n 0.0207627f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.41
cc_79 VPB N_A_c_126_n 0.00197941f $X=-0.19 $Y=1.305 $X2=5.96 $Y2=1.16
cc_80 VPB N_A_c_127_n 0.220237f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.202
cc_81 VPB N_VPWR_c_400_n 0.0125908f $X=-0.19 $Y=1.305 $X2=2.465 $Y2=0.995
cc_82 VPB N_VPWR_c_401_n 0.0061958f $X=-0.19 $Y=1.305 $X2=2.465 $Y2=0.56
cc_83 VPB N_VPWR_c_402_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.935 $Y2=0.56
cc_84 VPB N_VPWR_c_403_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.405 $Y2=0.995
cc_85 VPB N_VPWR_c_404_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.85 $Y2=1.985
cc_86 VPB N_VPWR_c_405_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.875 $Y2=0.56
cc_87 VPB N_VPWR_c_406_n 0.00469739f $X=-0.19 $Y=1.305 $X2=4.345 $Y2=0.995
cc_88 VPB N_VPWR_c_407_n 0.00469739f $X=-0.19 $Y=1.305 $X2=4.79 $Y2=1.985
cc_89 VPB N_VPWR_c_408_n 0.00469739f $X=-0.19 $Y=1.305 $X2=4.815 $Y2=0.56
cc_90 VPB N_VPWR_c_409_n 0.00496839f $X=-0.19 $Y=1.305 $X2=5.285 $Y2=0.995
cc_91 VPB N_VPWR_c_410_n 0.0206409f $X=-0.19 $Y=1.305 $X2=5.73 $Y2=1.41
cc_92 VPB N_VPWR_c_411_n 0.00324069f $X=-0.19 $Y=1.305 $X2=5.73 $Y2=1.985
cc_93 VPB N_VPWR_c_412_n 0.0206409f $X=-0.19 $Y=1.305 $X2=5.755 $Y2=0.995
cc_94 VPB N_VPWR_c_413_n 0.00324069f $X=-0.19 $Y=1.305 $X2=5.755 $Y2=0.56
cc_95 VPB N_VPWR_c_414_n 0.0206409f $X=-0.19 $Y=1.305 $X2=6.2 $Y2=1.41
cc_96 VPB N_VPWR_c_415_n 0.00324069f $X=-0.19 $Y=1.305 $X2=6.2 $Y2=1.985
cc_97 VPB N_VPWR_c_416_n 0.0206409f $X=-0.19 $Y=1.305 $X2=6.225 $Y2=0.995
cc_98 VPB N_VPWR_c_417_n 0.00324069f $X=-0.19 $Y=1.305 $X2=6.225 $Y2=0.56
cc_99 VPB N_VPWR_c_418_n 0.0206409f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_100 VPB N_VPWR_c_419_n 0.00324069f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.985
cc_101 VPB N_VPWR_c_420_n 0.0206409f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=0.995
cc_102 VPB N_VPWR_c_421_n 0.00324069f $X=-0.19 $Y=1.305 $X2=6.695 $Y2=0.56
cc_103 VPB N_VPWR_c_422_n 0.0206409f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.41
cc_104 VPB N_VPWR_c_423_n 0.00324069f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.985
cc_105 VPB N_VPWR_c_424_n 0.0206409f $X=-0.19 $Y=1.305 $X2=7.165 $Y2=0.995
cc_106 VPB N_VPWR_c_425_n 0.00401341f $X=-0.19 $Y=1.305 $X2=7.165 $Y2=0.56
cc_107 VPB N_VPWR_c_426_n 0.0120081f $X=-0.19 $Y=1.305 $X2=1.97 $Y2=1.202
cc_108 VPB N_VPWR_c_399_n 0.056908f $X=-0.19 $Y=1.305 $X2=1.995 $Y2=1.202
cc_109 VPB Y 0.00186291f $X=-0.19 $Y=1.305 $X2=4.845 $Y2=1.19
cc_110 N_A_c_128_n N_VPWR_c_401_n 0.00777746f $X=0.56 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_126_n N_VPWR_c_401_n 0.0168032f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_c_127_n N_VPWR_c_401_n 0.0049041f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_113 N_A_c_129_n N_VPWR_c_402_n 0.0052072f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_130_n N_VPWR_c_402_n 0.004751f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_131_n N_VPWR_c_403_n 0.0052072f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_132_n N_VPWR_c_403_n 0.004751f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_133_n N_VPWR_c_404_n 0.0052072f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_134_n N_VPWR_c_404_n 0.004751f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_135_n N_VPWR_c_405_n 0.0052072f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_136_n N_VPWR_c_405_n 0.004751f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_137_n N_VPWR_c_406_n 0.0052072f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_c_138_n N_VPWR_c_406_n 0.004751f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_139_n N_VPWR_c_407_n 0.0052072f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_140_n N_VPWR_c_407_n 0.004751f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_141_n N_VPWR_c_408_n 0.0052072f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_142_n N_VPWR_c_408_n 0.004751f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_143_n N_VPWR_c_409_n 0.00707238f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_128_n N_VPWR_c_410_n 0.00597712f $X=0.56 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_129_n N_VPWR_c_410_n 0.00673617f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_130_n N_VPWR_c_412_n 0.00597712f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_131_n N_VPWR_c_412_n 0.00673617f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_132_n N_VPWR_c_414_n 0.00597712f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_133_n N_VPWR_c_414_n 0.00673617f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_134_n N_VPWR_c_416_n 0.00597712f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_135_n N_VPWR_c_416_n 0.00673617f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_136_n N_VPWR_c_418_n 0.00597712f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_c_137_n N_VPWR_c_418_n 0.00673617f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_138_n N_VPWR_c_420_n 0.00597712f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_139_n N_VPWR_c_420_n 0.00673617f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_140_n N_VPWR_c_422_n 0.00597712f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_141_n N_VPWR_c_422_n 0.00673617f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_142_n N_VPWR_c_424_n 0.00597712f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_143_n N_VPWR_c_424_n 0.00673617f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_128_n N_VPWR_c_399_n 0.0109611f $X=0.56 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_129_n N_VPWR_c_399_n 0.0118438f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_130_n N_VPWR_c_399_n 0.00999457f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_131_n N_VPWR_c_399_n 0.0118438f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_132_n N_VPWR_c_399_n 0.00999457f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_133_n N_VPWR_c_399_n 0.0118438f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_134_n N_VPWR_c_399_n 0.00999457f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_135_n N_VPWR_c_399_n 0.0118438f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_136_n N_VPWR_c_399_n 0.00999457f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_137_n N_VPWR_c_399_n 0.0118438f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_138_n N_VPWR_c_399_n 0.00999457f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_139_n N_VPWR_c_399_n 0.0118438f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_140_n N_VPWR_c_399_n 0.00999457f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_141_n N_VPWR_c_399_n 0.0118438f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_142_n N_VPWR_c_399_n 0.00999457f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_143_n N_VPWR_c_399_n 0.012882f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_110_n N_Y_c_549_n 0.00724548f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_128_n N_Y_c_550_n 0.00350242f $X=0.56 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_c_129_n N_Y_c_550_n 5.87864e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_c_126_n N_Y_c_550_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_c_127_n N_Y_c_550_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_165 N_A_c_128_n N_Y_c_554_n 0.0121679f $X=0.56 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_129_n N_Y_c_554_n 0.0106251f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_130_n N_Y_c_554_n 6.24674e-19 $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_111_n N_Y_c_533_n 0.0111881f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_112_n N_Y_c_533_n 0.00640878f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_126_n N_Y_c_533_n 0.0405394f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_127_n N_Y_c_533_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_c_110_n N_Y_c_534_n 0.00487025f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_126_n N_Y_c_534_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A_c_127_n N_Y_c_534_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_c_129_n N_Y_c_564_n 0.0138566f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_130_n N_Y_c_564_n 0.0101493f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_126_n N_Y_c_564_n 0.0339162f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_c_127_n N_Y_c_564_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_179 N_A_c_111_n N_Y_c_568_n 5.79378e-19 $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_112_n N_Y_c_568_n 0.00837042f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_129_n N_Y_c_570_n 6.48386e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_130_n N_Y_c_570_n 0.0130707f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_131_n N_Y_c_570_n 0.0106251f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_132_n N_Y_c_570_n 6.24674e-19 $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_113_n N_Y_c_535_n 0.0111881f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_114_n N_Y_c_535_n 0.00640878f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_126_n N_Y_c_535_n 0.0405394f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_c_127_n N_Y_c_535_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_189 N_A_c_131_n N_Y_c_578_n 0.0138566f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_132_n N_Y_c_578_n 0.0101493f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_126_n N_Y_c_578_n 0.0339162f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_c_127_n N_Y_c_578_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_193 N_A_c_113_n N_Y_c_582_n 5.79378e-19 $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_114_n N_Y_c_582_n 0.00837042f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_131_n N_Y_c_584_n 6.48386e-19 $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_132_n N_Y_c_584_n 0.0130707f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_133_n N_Y_c_584_n 0.0106251f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_134_n N_Y_c_584_n 6.24674e-19 $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_115_n N_Y_c_536_n 0.0111881f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_116_n N_Y_c_536_n 0.00640878f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_126_n N_Y_c_536_n 0.0405394f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_202 N_A_c_127_n N_Y_c_536_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_203 N_A_c_133_n N_Y_c_592_n 0.0138566f $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_c_134_n N_Y_c_592_n 0.0101493f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_126_n N_Y_c_592_n 0.0339162f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_c_127_n N_Y_c_592_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_207 N_A_c_115_n N_Y_c_596_n 5.79378e-19 $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_c_116_n N_Y_c_596_n 0.00837042f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_133_n N_Y_c_598_n 6.48386e-19 $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_134_n N_Y_c_598_n 0.0130707f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_135_n N_Y_c_598_n 0.0106251f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_136_n N_Y_c_598_n 6.24674e-19 $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_c_117_n N_Y_c_537_n 0.0111881f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_118_n N_Y_c_537_n 0.00640878f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_c_126_n N_Y_c_537_n 0.0405394f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_c_127_n N_Y_c_537_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A_c_135_n N_Y_c_606_n 0.0138566f $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_136_n N_Y_c_606_n 0.0101493f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_c_126_n N_Y_c_606_n 0.0339162f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_c_127_n N_Y_c_606_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_221 N_A_c_117_n N_Y_c_610_n 5.79378e-19 $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_118_n N_Y_c_610_n 0.00837042f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_135_n N_Y_c_612_n 6.48386e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_136_n N_Y_c_612_n 0.0130707f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_137_n N_Y_c_612_n 0.0106251f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_138_n N_Y_c_612_n 6.24674e-19 $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_c_119_n N_Y_c_538_n 0.0111881f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_c_120_n N_Y_c_538_n 0.00640878f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A_c_126_n N_Y_c_538_n 0.0405394f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_c_127_n N_Y_c_538_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_231 N_A_c_137_n N_Y_c_620_n 0.0138566f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_c_138_n N_Y_c_620_n 0.0101493f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_c_126_n N_Y_c_620_n 0.0339162f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_c_127_n N_Y_c_620_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_235 N_A_c_119_n N_Y_c_624_n 5.79378e-19 $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_120_n N_Y_c_624_n 0.00837042f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_c_137_n N_Y_c_626_n 6.48386e-19 $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A_c_138_n N_Y_c_626_n 0.0130707f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_139_n N_Y_c_626_n 0.0106251f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_c_140_n N_Y_c_626_n 6.24674e-19 $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_c_121_n N_Y_c_539_n 0.0111881f $X=5.755 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_122_n N_Y_c_539_n 0.00728451f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_126_n N_Y_c_539_n 0.0338085f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_c_127_n N_Y_c_539_n 0.00346f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_245 N_A_c_139_n N_Y_c_634_n 0.0138566f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_140_n N_Y_c_634_n 0.0113102f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_126_n N_Y_c_634_n 0.0276305f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_127_n N_Y_c_634_n 0.0063804f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_249 N_A_c_121_n N_Y_c_638_n 5.79378e-19 $X=5.755 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_122_n N_Y_c_638_n 0.00837042f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_139_n N_Y_c_640_n 6.48386e-19 $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_140_n N_Y_c_640_n 0.0130707f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_141_n N_Y_c_640_n 0.0106251f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_142_n N_Y_c_640_n 6.24674e-19 $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_123_n N_Y_c_540_n 0.0130722f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_c_127_n N_Y_c_540_n 0.00416659f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_257 N_A_c_141_n N_Y_c_646_n 0.0158202f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_127_n N_Y_c_646_n 0.00650521f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_259 N_A_c_123_n N_Y_c_648_n 5.79378e-19 $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_124_n N_Y_c_648_n 0.00837042f $X=7.165 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_c_141_n N_Y_c_650_n 6.48386e-19 $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_142_n N_Y_c_650_n 0.0130707f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_143_n N_Y_c_650_n 0.0153658f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_112_n N_Y_c_541_n 0.00281161f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_c_126_n N_Y_c_541_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_c_127_n N_Y_c_541_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_267 N_A_c_130_n N_Y_c_656_n 0.00213487f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_131_n N_Y_c_656_n 5.87864e-19 $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_126_n N_Y_c_656_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_c_127_n N_Y_c_656_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_271 N_A_c_114_n N_Y_c_542_n 0.00281161f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_c_126_n N_Y_c_542_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_c_127_n N_Y_c_542_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_274 N_A_c_132_n N_Y_c_663_n 0.00213487f $X=2.44 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_133_n N_Y_c_663_n 5.87864e-19 $X=2.91 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_126_n N_Y_c_663_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_277 N_A_c_127_n N_Y_c_663_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_278 N_A_c_116_n N_Y_c_543_n 0.00281161f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_126_n N_Y_c_543_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_280 N_A_c_127_n N_Y_c_543_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_281 N_A_c_134_n N_Y_c_670_n 0.00213487f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_282 N_A_c_135_n N_Y_c_670_n 5.87864e-19 $X=3.85 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A_c_126_n N_Y_c_670_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_284 N_A_c_127_n N_Y_c_670_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_285 N_A_c_118_n N_Y_c_544_n 0.00281161f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_c_126_n N_Y_c_544_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_c_127_n N_Y_c_544_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_288 N_A_c_136_n N_Y_c_677_n 0.00213487f $X=4.32 $Y=1.41 $X2=0 $Y2=0
cc_289 N_A_c_137_n N_Y_c_677_n 5.87864e-19 $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A_c_126_n N_Y_c_677_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_c_127_n N_Y_c_677_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_292 N_A_c_120_n N_Y_c_545_n 0.00281161f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_c_126_n N_Y_c_545_n 0.0308883f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_c_127_n N_Y_c_545_n 0.00358305f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_295 N_A_c_138_n N_Y_c_684_n 0.00213487f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_c_139_n N_Y_c_684_n 5.87864e-19 $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A_c_126_n N_Y_c_684_n 0.024137f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_c_127_n N_Y_c_684_n 0.00654533f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_299 N_A_c_122_n N_Y_c_546_n 0.00373419f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_c_127_n N_Y_c_546_n 0.0045214f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_301 N_A_c_140_n N_Y_c_690_n 0.00292575f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_c_141_n N_Y_c_690_n 8.05641e-19 $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_c_127_n N_Y_c_690_n 0.00756182f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_304 N_A_c_142_n N_Y_c_693_n 0.0106681f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_c_143_n N_Y_c_693_n 0.00800284f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A_c_141_n Y 0.00177416f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_c_123_n Y 0.00213489f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_142_n Y 0.00265828f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_c_124_n Y 0.00995572f $X=7.165 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_c_143_n Y 0.00467389f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_c_125_n Y 0.00345209f $X=7.635 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_c_127_n Y 0.0686064f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_313 N_A_c_110_n N_VGND_c_829_n 0.00614891f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_c_126_n N_VGND_c_829_n 0.0169352f $X=5.96 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A_c_127_n N_VGND_c_829_n 0.0057967f $X=7.61 $Y=1.202 $X2=0 $Y2=0
cc_316 N_A_c_111_n N_VGND_c_830_n 0.00276126f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_c_112_n N_VGND_c_830_n 0.0035663f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A_c_113_n N_VGND_c_831_n 0.00276126f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_114_n N_VGND_c_831_n 0.0035663f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_115_n N_VGND_c_832_n 0.00276126f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_c_116_n N_VGND_c_832_n 0.0035663f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_c_117_n N_VGND_c_833_n 0.00276126f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_c_118_n N_VGND_c_833_n 0.0035663f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_c_119_n N_VGND_c_834_n 0.00276126f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_c_120_n N_VGND_c_834_n 0.0035663f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_c_121_n N_VGND_c_835_n 0.00276126f $X=5.755 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_c_122_n N_VGND_c_835_n 0.0035663f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_c_123_n N_VGND_c_836_n 0.00276126f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_c_124_n N_VGND_c_836_n 0.0035663f $X=7.165 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_c_125_n N_VGND_c_837_n 0.00444548f $X=7.635 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_c_110_n N_VGND_c_838_n 0.00465454f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_c_111_n N_VGND_c_838_n 0.00436487f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_c_112_n N_VGND_c_840_n 0.00395968f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_c_113_n N_VGND_c_840_n 0.00436487f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_c_114_n N_VGND_c_842_n 0.00395968f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A_c_115_n N_VGND_c_842_n 0.00436487f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A_c_116_n N_VGND_c_844_n 0.00395968f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_c_117_n N_VGND_c_844_n 0.00436487f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A_c_118_n N_VGND_c_846_n 0.00395968f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_340 N_A_c_119_n N_VGND_c_846_n 0.00436487f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_341 N_A_c_120_n N_VGND_c_848_n 0.00395968f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A_c_121_n N_VGND_c_848_n 0.00436487f $X=5.755 $Y=0.995 $X2=0 $Y2=0
cc_343 N_A_c_122_n N_VGND_c_850_n 0.00395968f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_344 N_A_c_123_n N_VGND_c_850_n 0.00436487f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_345 N_A_c_124_n N_VGND_c_852_n 0.00395904f $X=7.165 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A_c_125_n N_VGND_c_852_n 0.00585385f $X=7.635 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A_c_110_n N_VGND_c_855_n 0.0089497f $X=0.585 $Y=0.995 $X2=0 $Y2=0
cc_348 N_A_c_111_n N_VGND_c_855_n 0.0061161f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A_c_112_n N_VGND_c_855_n 0.0058034f $X=1.525 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A_c_113_n N_VGND_c_855_n 0.0061161f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A_c_114_n N_VGND_c_855_n 0.0058034f $X=2.465 $Y=0.995 $X2=0 $Y2=0
cc_352 N_A_c_115_n N_VGND_c_855_n 0.0061161f $X=2.935 $Y=0.995 $X2=0 $Y2=0
cc_353 N_A_c_116_n N_VGND_c_855_n 0.0058034f $X=3.405 $Y=0.995 $X2=0 $Y2=0
cc_354 N_A_c_117_n N_VGND_c_855_n 0.0061161f $X=3.875 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A_c_118_n N_VGND_c_855_n 0.0058034f $X=4.345 $Y=0.995 $X2=0 $Y2=0
cc_356 N_A_c_119_n N_VGND_c_855_n 0.0061161f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A_c_120_n N_VGND_c_855_n 0.0058034f $X=5.285 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A_c_121_n N_VGND_c_855_n 0.0061161f $X=5.755 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A_c_122_n N_VGND_c_855_n 0.0058034f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A_c_123_n N_VGND_c_855_n 0.0061161f $X=6.695 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A_c_124_n N_VGND_c_855_n 0.00580225f $X=7.165 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A_c_125_n N_VGND_c_855_n 0.011749f $X=7.635 $Y=0.995 $X2=0 $Y2=0
cc_363 N_VPWR_c_399_n N_Y_M1000_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_399_n N_Y_M1002_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_365 N_VPWR_c_399_n N_Y_M1005_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_366 N_VPWR_c_399_n N_Y_M1011_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_367 N_VPWR_c_399_n N_Y_M1013_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_399_n N_Y_M1018_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_c_399_n N_Y_M1022_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_399_n N_Y_M1028_s 0.00231261f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_401_n N_Y_c_550_n 0.0135612f $X=0.325 $Y=1.65 $X2=0 $Y2=0
cc_372 N_VPWR_c_401_n N_Y_c_554_n 0.0606207f $X=0.325 $Y=1.65 $X2=0 $Y2=0
cc_373 N_VPWR_c_402_n N_Y_c_554_n 0.0385613f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_374 N_VPWR_c_410_n N_Y_c_554_n 0.0223557f $X=1.18 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_c_399_n N_Y_c_554_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_M1001_d N_Y_c_564_n 0.00329096f $X=1.12 $Y=1.485 $X2=0 $Y2=0
cc_377 N_VPWR_c_402_n N_Y_c_564_n 0.0136682f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_378 N_VPWR_c_402_n N_Y_c_570_n 0.0470327f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_379 N_VPWR_c_403_n N_Y_c_570_n 0.0385613f $X=2.205 $Y=2 $X2=0 $Y2=0
cc_380 N_VPWR_c_412_n N_Y_c_570_n 0.0223557f $X=2.12 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_399_n N_Y_c_570_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_M1003_d N_Y_c_578_n 0.00329096f $X=2.06 $Y=1.485 $X2=0 $Y2=0
cc_383 N_VPWR_c_403_n N_Y_c_578_n 0.0136682f $X=2.205 $Y=2 $X2=0 $Y2=0
cc_384 N_VPWR_c_403_n N_Y_c_584_n 0.0470327f $X=2.205 $Y=2 $X2=0 $Y2=0
cc_385 N_VPWR_c_404_n N_Y_c_584_n 0.0385613f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_386 N_VPWR_c_414_n N_Y_c_584_n 0.0223557f $X=3.06 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_399_n N_Y_c_584_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1010_d N_Y_c_592_n 0.00329096f $X=3 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_404_n N_Y_c_592_n 0.0136682f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_390 N_VPWR_c_404_n N_Y_c_598_n 0.0470327f $X=3.145 $Y=2 $X2=0 $Y2=0
cc_391 N_VPWR_c_405_n N_Y_c_598_n 0.0385613f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_392 N_VPWR_c_416_n N_Y_c_598_n 0.0223557f $X=4 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_399_n N_Y_c_598_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1012_d N_Y_c_606_n 0.00329096f $X=3.94 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_405_n N_Y_c_606_n 0.0136682f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_405_n N_Y_c_612_n 0.0470327f $X=4.085 $Y=2 $X2=0 $Y2=0
cc_397 N_VPWR_c_406_n N_Y_c_612_n 0.0385613f $X=5.025 $Y=2 $X2=0 $Y2=0
cc_398 N_VPWR_c_418_n N_Y_c_612_n 0.0223557f $X=4.94 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_399_n N_Y_c_612_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_M1015_d N_Y_c_620_n 0.00329096f $X=4.88 $Y=1.485 $X2=0 $Y2=0
cc_401 N_VPWR_c_406_n N_Y_c_620_n 0.0136682f $X=5.025 $Y=2 $X2=0 $Y2=0
cc_402 N_VPWR_c_406_n N_Y_c_626_n 0.0470327f $X=5.025 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_407_n N_Y_c_626_n 0.0385613f $X=5.965 $Y=2 $X2=0 $Y2=0
cc_404 N_VPWR_c_420_n N_Y_c_626_n 0.0223557f $X=5.88 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_c_399_n N_Y_c_626_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_M1020_d N_Y_c_634_n 0.00329096f $X=5.82 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_c_407_n N_Y_c_634_n 0.0136682f $X=5.965 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_407_n N_Y_c_640_n 0.0470327f $X=5.965 $Y=2 $X2=0 $Y2=0
cc_409 N_VPWR_c_408_n N_Y_c_640_n 0.0385613f $X=6.905 $Y=2 $X2=0 $Y2=0
cc_410 N_VPWR_c_422_n N_Y_c_640_n 0.0223557f $X=6.82 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_c_399_n N_Y_c_640_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_M1024_d N_Y_c_646_n 0.00410773f $X=6.76 $Y=1.485 $X2=0 $Y2=0
cc_413 N_VPWR_c_408_n N_Y_c_646_n 0.0136682f $X=6.905 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_408_n N_Y_c_650_n 0.0470327f $X=6.905 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_409_n N_Y_c_650_n 0.0391697f $X=7.845 $Y=2 $X2=0 $Y2=0
cc_416 N_VPWR_c_424_n N_Y_c_650_n 0.0223557f $X=7.76 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_c_399_n N_Y_c_650_n 0.0140101f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_418 N_Y_c_533_n N_VGND_M1006_s 0.0025045f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_419 N_Y_c_535_n N_VGND_M1008_s 0.0025045f $X=2.46 $Y=0.81 $X2=0 $Y2=0
cc_420 N_Y_c_536_n N_VGND_M1014_s 0.0025045f $X=3.4 $Y=0.81 $X2=0 $Y2=0
cc_421 N_Y_c_537_n N_VGND_M1017_s 0.0025045f $X=4.34 $Y=0.81 $X2=0 $Y2=0
cc_422 N_Y_c_538_n N_VGND_M1021_s 0.0025045f $X=5.28 $Y=0.81 $X2=0 $Y2=0
cc_423 N_Y_c_539_n N_VGND_M1025_s 0.0025045f $X=6.22 $Y=0.81 $X2=0 $Y2=0
cc_424 N_Y_c_540_n N_VGND_M1027_s 0.00214188f $X=7.015 $Y=0.81 $X2=0 $Y2=0
cc_425 Y N_VGND_M1027_s 3.59126e-19 $X=7.335 $Y=0.765 $X2=0 $Y2=0
cc_426 N_Y_c_549_n N_VGND_c_829_n 0.0350772f $X=0.795 $Y=0.38 $X2=0 $Y2=0
cc_427 N_Y_c_534_n N_VGND_c_829_n 0.013649f $X=0.96 $Y=0.81 $X2=0 $Y2=0
cc_428 N_Y_c_533_n N_VGND_c_830_n 0.0127393f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_429 N_Y_c_568_n N_VGND_c_830_n 0.0216501f $X=1.735 $Y=0.38 $X2=0 $Y2=0
cc_430 N_Y_c_535_n N_VGND_c_831_n 0.0127393f $X=2.46 $Y=0.81 $X2=0 $Y2=0
cc_431 N_Y_c_582_n N_VGND_c_831_n 0.0216501f $X=2.675 $Y=0.38 $X2=0 $Y2=0
cc_432 N_Y_c_536_n N_VGND_c_832_n 0.0127393f $X=3.4 $Y=0.81 $X2=0 $Y2=0
cc_433 N_Y_c_596_n N_VGND_c_832_n 0.0216501f $X=3.615 $Y=0.38 $X2=0 $Y2=0
cc_434 N_Y_c_537_n N_VGND_c_833_n 0.0127393f $X=4.34 $Y=0.81 $X2=0 $Y2=0
cc_435 N_Y_c_610_n N_VGND_c_833_n 0.0216501f $X=4.555 $Y=0.38 $X2=0 $Y2=0
cc_436 N_Y_c_538_n N_VGND_c_834_n 0.0127393f $X=5.28 $Y=0.81 $X2=0 $Y2=0
cc_437 N_Y_c_624_n N_VGND_c_834_n 0.0216501f $X=5.495 $Y=0.38 $X2=0 $Y2=0
cc_438 N_Y_c_539_n N_VGND_c_835_n 0.0127393f $X=6.22 $Y=0.81 $X2=0 $Y2=0
cc_439 N_Y_c_638_n N_VGND_c_835_n 0.0216501f $X=6.435 $Y=0.38 $X2=0 $Y2=0
cc_440 N_Y_c_540_n N_VGND_c_836_n 0.0127393f $X=7.015 $Y=0.81 $X2=0 $Y2=0
cc_441 N_Y_c_648_n N_VGND_c_836_n 0.0216501f $X=7.375 $Y=0.38 $X2=0 $Y2=0
cc_442 N_Y_c_549_n N_VGND_c_838_n 0.023074f $X=0.795 $Y=0.38 $X2=0 $Y2=0
cc_443 N_Y_c_533_n N_VGND_c_838_n 0.00260993f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_444 N_Y_c_533_n N_VGND_c_840_n 0.0020445f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_445 N_Y_c_568_n N_VGND_c_840_n 0.023074f $X=1.735 $Y=0.38 $X2=0 $Y2=0
cc_446 N_Y_c_535_n N_VGND_c_840_n 0.00260993f $X=2.46 $Y=0.81 $X2=0 $Y2=0
cc_447 N_Y_c_535_n N_VGND_c_842_n 0.0020445f $X=2.46 $Y=0.81 $X2=0 $Y2=0
cc_448 N_Y_c_582_n N_VGND_c_842_n 0.023074f $X=2.675 $Y=0.38 $X2=0 $Y2=0
cc_449 N_Y_c_536_n N_VGND_c_842_n 0.00260993f $X=3.4 $Y=0.81 $X2=0 $Y2=0
cc_450 N_Y_c_536_n N_VGND_c_844_n 0.0020445f $X=3.4 $Y=0.81 $X2=0 $Y2=0
cc_451 N_Y_c_596_n N_VGND_c_844_n 0.023074f $X=3.615 $Y=0.38 $X2=0 $Y2=0
cc_452 N_Y_c_537_n N_VGND_c_844_n 0.00260993f $X=4.34 $Y=0.81 $X2=0 $Y2=0
cc_453 N_Y_c_537_n N_VGND_c_846_n 0.0020445f $X=4.34 $Y=0.81 $X2=0 $Y2=0
cc_454 N_Y_c_610_n N_VGND_c_846_n 0.023074f $X=4.555 $Y=0.38 $X2=0 $Y2=0
cc_455 N_Y_c_538_n N_VGND_c_846_n 0.00260993f $X=5.28 $Y=0.81 $X2=0 $Y2=0
cc_456 N_Y_c_538_n N_VGND_c_848_n 0.0020445f $X=5.28 $Y=0.81 $X2=0 $Y2=0
cc_457 N_Y_c_624_n N_VGND_c_848_n 0.023074f $X=5.495 $Y=0.38 $X2=0 $Y2=0
cc_458 N_Y_c_539_n N_VGND_c_848_n 0.00260993f $X=6.22 $Y=0.81 $X2=0 $Y2=0
cc_459 N_Y_c_539_n N_VGND_c_850_n 0.0020445f $X=6.22 $Y=0.81 $X2=0 $Y2=0
cc_460 N_Y_c_638_n N_VGND_c_850_n 0.023074f $X=6.435 $Y=0.38 $X2=0 $Y2=0
cc_461 N_Y_c_540_n N_VGND_c_850_n 0.00260993f $X=7.015 $Y=0.81 $X2=0 $Y2=0
cc_462 N_Y_c_540_n N_VGND_c_852_n 3.57378e-19 $X=7.015 $Y=0.81 $X2=0 $Y2=0
cc_463 N_Y_c_648_n N_VGND_c_852_n 0.0231393f $X=7.375 $Y=0.38 $X2=0 $Y2=0
cc_464 Y N_VGND_c_852_n 0.0018043f $X=7.335 $Y=0.765 $X2=0 $Y2=0
cc_465 N_Y_M1004_d N_VGND_c_855_n 0.0026371f $X=0.66 $Y=0.235 $X2=0 $Y2=0
cc_466 N_Y_M1007_d N_VGND_c_855_n 0.0026371f $X=1.6 $Y=0.235 $X2=0 $Y2=0
cc_467 N_Y_M1009_d N_VGND_c_855_n 0.0026371f $X=2.54 $Y=0.235 $X2=0 $Y2=0
cc_468 N_Y_M1016_d N_VGND_c_855_n 0.0026371f $X=3.48 $Y=0.235 $X2=0 $Y2=0
cc_469 N_Y_M1019_d N_VGND_c_855_n 0.0026371f $X=4.42 $Y=0.235 $X2=0 $Y2=0
cc_470 N_Y_M1023_d N_VGND_c_855_n 0.0026371f $X=5.36 $Y=0.235 $X2=0 $Y2=0
cc_471 N_Y_M1026_d N_VGND_c_855_n 0.0026371f $X=6.3 $Y=0.235 $X2=0 $Y2=0
cc_472 N_Y_M1029_d N_VGND_c_855_n 0.00324782f $X=7.24 $Y=0.235 $X2=0 $Y2=0
cc_473 N_Y_c_549_n N_VGND_c_855_n 0.0141066f $X=0.795 $Y=0.38 $X2=0 $Y2=0
cc_474 N_Y_c_533_n N_VGND_c_855_n 0.00988931f $X=1.52 $Y=0.81 $X2=0 $Y2=0
cc_475 N_Y_c_568_n N_VGND_c_855_n 0.0141066f $X=1.735 $Y=0.38 $X2=0 $Y2=0
cc_476 N_Y_c_535_n N_VGND_c_855_n 0.00988931f $X=2.46 $Y=0.81 $X2=0 $Y2=0
cc_477 N_Y_c_582_n N_VGND_c_855_n 0.0141066f $X=2.675 $Y=0.38 $X2=0 $Y2=0
cc_478 N_Y_c_536_n N_VGND_c_855_n 0.00988931f $X=3.4 $Y=0.81 $X2=0 $Y2=0
cc_479 N_Y_c_596_n N_VGND_c_855_n 0.0141066f $X=3.615 $Y=0.38 $X2=0 $Y2=0
cc_480 N_Y_c_537_n N_VGND_c_855_n 0.00988931f $X=4.34 $Y=0.81 $X2=0 $Y2=0
cc_481 N_Y_c_610_n N_VGND_c_855_n 0.0141066f $X=4.555 $Y=0.38 $X2=0 $Y2=0
cc_482 N_Y_c_538_n N_VGND_c_855_n 0.00988931f $X=5.28 $Y=0.81 $X2=0 $Y2=0
cc_483 N_Y_c_624_n N_VGND_c_855_n 0.0141066f $X=5.495 $Y=0.38 $X2=0 $Y2=0
cc_484 N_Y_c_539_n N_VGND_c_855_n 0.00988931f $X=6.22 $Y=0.81 $X2=0 $Y2=0
cc_485 N_Y_c_638_n N_VGND_c_855_n 0.0141066f $X=6.435 $Y=0.38 $X2=0 $Y2=0
cc_486 N_Y_c_540_n N_VGND_c_855_n 0.0063975f $X=7.015 $Y=0.81 $X2=0 $Y2=0
cc_487 N_Y_c_648_n N_VGND_c_855_n 0.0141237f $X=7.375 $Y=0.38 $X2=0 $Y2=0
cc_488 Y N_VGND_c_855_n 0.00371433f $X=7.335 $Y=0.765 $X2=0 $Y2=0
