* File: sky130_fd_sc_hdll__einvn_1.pxi.spice
* Created: Wed Sep  2 08:31:04 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVN_1%TE_B N_TE_B_c_43_n N_TE_B_c_48_n N_TE_B_c_49_n
+ N_TE_B_M1001_g N_TE_B_M1002_g N_TE_B_c_45_n N_TE_B_c_51_n N_TE_B_M1004_g TE_B
+ TE_B N_TE_B_c_46_n PM_SKY130_FD_SC_HDLL__EINVN_1%TE_B
x_PM_SKY130_FD_SC_HDLL__EINVN_1%A_27_47# N_A_27_47#_M1002_s N_A_27_47#_M1001_s
+ N_A_27_47#_M1000_g N_A_27_47#_c_89_n N_A_27_47#_c_95_n N_A_27_47#_c_90_n
+ N_A_27_47#_c_103_n N_A_27_47#_c_96_n N_A_27_47#_c_108_n N_A_27_47#_c_97_n
+ N_A_27_47#_c_98_n N_A_27_47#_c_116_n N_A_27_47#_c_91_n N_A_27_47#_c_92_n
+ N_A_27_47#_c_93_n N_A_27_47#_c_94_n PM_SKY130_FD_SC_HDLL__EINVN_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVN_1%A N_A_c_161_n N_A_M1005_g N_A_c_164_n
+ N_A_M1003_g A A A N_A_c_163_n PM_SKY130_FD_SC_HDLL__EINVN_1%A
x_PM_SKY130_FD_SC_HDLL__EINVN_1%VPWR N_VPWR_M1001_d N_VPWR_c_191_n VPWR
+ N_VPWR_c_192_n N_VPWR_c_193_n N_VPWR_c_190_n N_VPWR_c_195_n
+ PM_SKY130_FD_SC_HDLL__EINVN_1%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVN_1%Z N_Z_M1005_d N_Z_M1003_d N_Z_c_226_n Z Z Z Z Z
+ Z Z PM_SKY130_FD_SC_HDLL__EINVN_1%Z
x_PM_SKY130_FD_SC_HDLL__EINVN_1%VGND N_VGND_M1002_d VGND N_VGND_c_258_n
+ N_VGND_c_259_n N_VGND_c_260_n N_VGND_c_261_n
+ PM_SKY130_FD_SC_HDLL__EINVN_1%VGND
cc_1 VNB N_TE_B_c_43_n 0.0327928f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_TE_B_M1002_g 0.0426796f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_3 VNB N_TE_B_c_45_n 0.0193191f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.335
cc_4 VNB N_TE_B_c_46_n 0.0168719f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_5 VNB N_A_27_47#_c_89_n 0.0141471f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.41
cc_6 VNB N_A_27_47#_c_90_n 0.0101961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_91_n 0.00663899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_92_n 0.036323f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_93_n 0.00139297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_94_n 0.0200495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_161_n 0.021023f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB A 0.0206302f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_13 VNB N_A_c_163_n 0.0405042f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.985
cc_14 VNB N_VPWR_c_190_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_15 VNB Z 0.00380052f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.335
cc_16 VNB Z 0.0152064f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.985
cc_17 VNB N_VGND_c_258_n 0.0315501f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_18 VNB N_VGND_c_259_n 0.162102f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_260_n 0.014818f $X=-0.19 $Y=-0.24 $X2=0.432 $Y2=1.335
cc_20 VNB N_VGND_c_261_n 0.021551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_TE_B_c_43_n 0.00906422f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_22 VPB N_TE_B_c_48_n 0.017843f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_23 VPB N_TE_B_c_49_n 0.0294942f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_24 VPB N_TE_B_c_45_n 0.0121082f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.335
cc_25 VPB N_TE_B_c_51_n 0.0195778f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.41
cc_26 VPB N_TE_B_c_46_n 0.0201207f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_27 VPB N_A_27_47#_c_95_n 0.0156843f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.985
cc_28 VPB N_A_27_47#_c_96_n 0.0076959f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_29 VPB N_A_27_47#_c_97_n 6.61338e-19 $X=-0.19 $Y=1.305 $X2=0.297 $Y2=1.16
cc_30 VPB N_A_27_47#_c_98_n 0.00237273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_27_47#_c_91_n 0.00239242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_47#_c_92_n 0.0120311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_c_164_n 0.0225104f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_34 VPB A 0.0128119f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_35 VPB N_A_c_163_n 0.0168885f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.985
cc_36 VPB N_VPWR_c_191_n 0.00299909f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_37 VPB N_VPWR_c_192_n 0.0148836f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.335
cc_38 VPB N_VPWR_c_193_n 0.0485615f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_39 VPB N_VPWR_c_190_n 0.0443787f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_40 VPB N_VPWR_c_195_n 0.00594495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB Z 0.00228085f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.335
cc_42 VPB Z 0.0296293f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.985
cc_43 N_TE_B_c_43_n N_A_27_47#_c_90_n 6.91349e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_TE_B_c_46_n N_A_27_47#_c_90_n 0.0261211f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_45 N_TE_B_c_49_n N_A_27_47#_c_103_n 0.0149473f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_46 N_TE_B_c_45_n N_A_27_47#_c_103_n 0.00121726f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_47 N_TE_B_c_46_n N_A_27_47#_c_103_n 0.00950979f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_48 N_TE_B_c_43_n N_A_27_47#_c_96_n 3.10924e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_49 N_TE_B_c_46_n N_A_27_47#_c_96_n 0.0248947f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_50 N_TE_B_c_48_n N_A_27_47#_c_108_n 0.00183873f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_51 N_TE_B_c_49_n N_A_27_47#_c_108_n 0.00278004f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_52 N_TE_B_c_46_n N_A_27_47#_c_108_n 0.00665669f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_53 N_TE_B_c_45_n N_A_27_47#_c_97_n 2.77516e-19 $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_54 N_TE_B_c_51_n N_A_27_47#_c_97_n 0.020203f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_55 N_TE_B_c_48_n N_A_27_47#_c_98_n 0.00150938f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_56 N_TE_B_c_45_n N_A_27_47#_c_98_n 0.00333143f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_57 N_TE_B_c_46_n N_A_27_47#_c_98_n 0.0119344f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_58 N_TE_B_M1002_g N_A_27_47#_c_116_n 8.06856e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_59 N_TE_B_c_45_n N_A_27_47#_c_116_n 0.00789825f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_60 N_TE_B_M1002_g N_A_27_47#_c_91_n 0.00955669f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_61 N_TE_B_c_45_n N_A_27_47#_c_91_n 0.00455883f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_62 N_TE_B_c_51_n N_A_27_47#_c_91_n 9.39224e-19 $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_63 N_TE_B_c_46_n N_A_27_47#_c_91_n 0.0152387f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_64 N_TE_B_c_45_n N_A_27_47#_c_92_n 0.00424579f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_65 N_TE_B_c_43_n N_A_27_47#_c_93_n 4.66638e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_TE_B_M1002_g N_A_27_47#_c_93_n 0.0169554f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_67 N_TE_B_c_45_n N_A_27_47#_c_93_n 0.00392316f $X=0.93 $Y=1.335 $X2=0 $Y2=0
cc_68 N_TE_B_c_46_n N_A_27_47#_c_93_n 0.011171f $X=0.405 $Y=1.16 $X2=0 $Y2=0
cc_69 N_TE_B_c_49_n N_VPWR_c_191_n 0.00983058f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_70 N_TE_B_c_51_n N_VPWR_c_191_n 0.00329012f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_71 N_TE_B_c_49_n N_VPWR_c_192_n 0.00384491f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_72 N_TE_B_c_51_n N_VPWR_c_193_n 0.00702461f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_73 N_TE_B_c_49_n N_VPWR_c_190_n 0.00545975f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_74 N_TE_B_c_51_n N_VPWR_c_190_n 0.0139274f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_75 N_TE_B_c_51_n Z 0.0172382f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_76 N_TE_B_M1002_g N_VGND_c_259_n 0.0042776f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_77 N_TE_B_M1002_g N_VGND_c_260_n 0.00266649f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_78 N_TE_B_M1002_g N_VGND_c_261_n 0.0112582f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_91_n N_A_c_161_n 4.13669e-19 $X=1.465 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_47#_c_94_n N_A_c_161_n 0.0130391f $X=1.512 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_27_47#_c_97_n N_A_c_164_n 8.81552e-19 $X=1.12 $Y=1.527 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_91_n N_A_c_163_n 6.94707e-19 $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_92_n N_A_c_163_n 0.0069166f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_103_n N_VPWR_M1001_d 0.0058167f $X=0.735 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_27_47#_c_108_n N_VPWR_M1001_d 0.00363839f $X=0.827 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_27_47#_c_98_n N_VPWR_M1001_d 0.00136109f $X=0.92 $Y=1.527 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_27_47#_c_103_n N_VPWR_c_191_n 0.0218593f $X=0.735 $Y=1.98 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_95_n N_VPWR_c_192_n 0.0189983f $X=0.227 $Y=2.065 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_103_n N_VPWR_c_192_n 0.00241908f $X=0.735 $Y=1.98 $X2=0 $Y2=0
cc_90 N_A_27_47#_M1001_s N_VPWR_c_190_n 0.002313f $X=0.135 $Y=1.845 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_95_n N_VPWR_c_190_n 0.0108489f $X=0.227 $Y=2.065 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_103_n N_VPWR_c_190_n 0.00578679f $X=0.735 $Y=1.98 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_97_n A_222_297# 0.0164657f $X=1.12 $Y=1.527 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_27_47#_c_94_n N_Z_c_226_n 0.00447459f $X=1.512 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_97_n Z 0.00836614f $X=1.12 $Y=1.527 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_91_n Z 0.0273348f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_92_n Z 0.00302888f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_94_n Z 0.00192642f $X=1.512 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_97_n Z 0.0179488f $X=1.12 $Y=1.527 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_92_n Z 0.00392927f $X=1.465 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_116_n N_VGND_M1002_d 0.0184931f $X=1.36 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_27_47#_c_91_n N_VGND_M1002_d 0.00235026f $X=1.465 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_27_47#_c_93_n N_VGND_M1002_d 0.00180161f $X=0.735 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_27_47#_M1002_s N_VGND_c_259_n 0.00278465f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_c_89_n N_VGND_c_259_n 0.0108288f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_116_n N_VGND_c_259_n 2.65731e-19 $X=1.36 $Y=0.805 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_93_n N_VGND_c_259_n 0.00920837f $X=0.735 $Y=0.71 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_89_n N_VGND_c_260_n 0.019607f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_93_n N_VGND_c_260_n 0.00252163f $X=0.735 $Y=0.71 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_89_n N_VGND_c_261_n 0.0154094f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_93_n N_VGND_c_261_n 0.0691774f $X=0.735 $Y=0.71 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_94_n N_VGND_c_261_n 0.0207421f $X=1.512 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_c_164_n N_VPWR_c_193_n 0.00429453f $X=2.265 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_164_n N_VPWR_c_190_n 0.00830809f $X=2.265 $Y=1.41 $X2=0 $Y2=0
cc_115 A N_Z_M1005_d 0.00371964f $X=2.44 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_116 A N_Z_M1003_d 0.00446811f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_117 N_A_c_161_n N_Z_c_226_n 0.00649803f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_161_n Z 0.0158782f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_c_164_n Z 0.017094f $X=2.265 $Y=1.41 $X2=0 $Y2=0
cc_120 A Z 0.0511712f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_121 N_A_c_163_n Z 0.013627f $X=2.265 $Y=1.202 $X2=0 $Y2=0
cc_122 N_A_c_161_n Z 0.00910094f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_123 A Z 0.0201989f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_124 N_A_c_163_n Z 0.00387543f $X=2.265 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_c_164_n Z 0.0370161f $X=2.265 $Y=1.41 $X2=0 $Y2=0
cc_126 A Z 0.0219813f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_127 N_A_c_163_n Z 0.00223631f $X=2.265 $Y=1.202 $X2=0 $Y2=0
cc_128 N_A_c_161_n N_VGND_c_258_n 0.00357815f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_161_n N_VGND_c_259_n 0.00686814f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_161_n N_VGND_c_261_n 0.00135425f $X=2.24 $Y=0.995 $X2=0 $Y2=0
cc_131 N_VPWR_c_190_n A_222_297# 0.0187386f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_132 N_VPWR_c_190_n N_Z_M1003_d 0.00217543f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_193_n Z 0.0847414f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_190_n Z 0.0481744f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 A_222_297# Z 0.00956008f $X=1.11 $Y=1.485 $X2=0.227 $Y2=0.445
cc_136 A_222_297# Z 0.0556527f $X=1.11 $Y=1.485 $X2=0.227 $Y2=2.065
cc_137 N_Z_c_226_n N_VGND_c_258_n 0.0147948f $X=2.21 $Y=0.425 $X2=0 $Y2=0
cc_138 Z N_VGND_c_258_n 0.0289189f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_139 N_Z_M1005_d N_VGND_c_259_n 0.00250339f $X=2.315 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Z_c_226_n N_VGND_c_259_n 0.00903703f $X=2.21 $Y=0.425 $X2=0 $Y2=0
cc_141 Z N_VGND_c_259_n 0.0170352f $X=2.44 $Y=0.425 $X2=0 $Y2=0
cc_142 N_Z_c_226_n A_316_47# 0.00663916f $X=2.21 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_143 Z A_316_47# 0.00395336f $X=1.98 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_144 N_VGND_c_259_n A_316_47# 0.0175224f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
