* File: sky130_fd_sc_hdll__xnor3_1.pxi.spice
* Created: Wed Sep  2 08:53:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_83_21# N_A_83_21#_M1002_d N_A_83_21#_M1015_d
+ N_A_83_21#_c_152_n N_A_83_21#_M1012_g N_A_83_21#_c_153_n N_A_83_21#_M1000_g
+ N_A_83_21#_c_154_n N_A_83_21#_c_159_n N_A_83_21#_c_165_p N_A_83_21#_c_201_p
+ N_A_83_21#_c_170_p N_A_83_21#_c_205_p N_A_83_21#_c_155_n N_A_83_21#_c_160_n
+ N_A_83_21#_c_156_n N_A_83_21#_c_161_n N_A_83_21#_c_162_n N_A_83_21#_c_174_p
+ N_A_83_21#_c_230_p N_A_83_21#_c_177_p N_A_83_21#_c_157_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%A_83_21#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%C N_C_c_251_n N_C_M1020_g N_C_M1017_g
+ N_C_c_252_n N_C_M1015_g N_C_c_253_n N_C_M1002_g N_C_c_254_n N_C_c_255_n C
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%C
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_226_93# N_A_226_93#_M1020_d
+ N_A_226_93#_M1017_d N_A_226_93#_c_311_n N_A_226_93#_M1021_g
+ N_A_226_93#_c_312_n N_A_226_93#_M1013_g N_A_226_93#_c_326_n
+ N_A_226_93#_c_313_n N_A_226_93#_c_317_n N_A_226_93#_c_318_n
+ N_A_226_93#_c_319_n N_A_226_93#_c_314_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%A_226_93#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_783_297# N_A_783_297#_M1008_d
+ N_A_783_297#_M1004_d N_A_783_297#_c_395_n N_A_783_297#_M1018_g
+ N_A_783_297#_M1016_g N_A_783_297#_c_382_n N_A_783_297#_c_397_n
+ N_A_783_297#_M1005_g N_A_783_297#_M1001_g N_A_783_297#_c_383_n
+ N_A_783_297#_c_384_n N_A_783_297#_c_400_n N_A_783_297#_c_385_n
+ N_A_783_297#_c_386_n N_A_783_297#_c_404_p N_A_783_297#_c_387_n
+ N_A_783_297#_c_388_n N_A_783_297#_c_389_n N_A_783_297#_c_390_n
+ N_A_783_297#_c_391_n N_A_783_297#_c_392_n N_A_783_297#_c_393_n
+ N_A_783_297#_c_394_n PM_SKY130_FD_SC_HDLL__XNOR3_1%A_783_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%B N_B_c_570_n N_B_M1004_g N_B_M1008_g
+ N_B_c_563_n N_B_c_564_n N_B_M1010_g N_B_M1006_g N_B_c_573_n N_B_c_574_n
+ N_B_M1019_g N_B_c_575_n N_B_c_576_n N_B_M1011_g N_B_c_566_n N_B_c_579_n
+ N_B_c_567_n N_B_c_568_n B B N_B_c_569_n PM_SKY130_FD_SC_HDLL__XNOR3_1%B
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A N_A_c_698_n N_A_M1014_g N_A_c_699_n
+ N_A_M1009_g A A PM_SKY130_FD_SC_HDLL__XNOR3_1%A
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_901_297# N_A_901_297#_M1006_s
+ N_A_901_297#_M1001_d N_A_901_297#_M1010_s N_A_901_297#_M1005_d
+ N_A_901_297#_c_736_n N_A_901_297#_M1007_g N_A_901_297#_c_737_n
+ N_A_901_297#_M1003_g N_A_901_297#_c_738_n N_A_901_297#_c_746_n
+ N_A_901_297#_c_739_n N_A_901_297#_c_740_n N_A_901_297#_c_741_n
+ N_A_901_297#_c_748_n N_A_901_297#_c_758_n N_A_901_297#_c_742_n
+ N_A_901_297#_c_743_n N_A_901_297#_c_771_n N_A_901_297#_c_772_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%A_901_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%X N_X_M1012_s N_X_M1000_s N_X_c_866_n
+ N_X_c_868_n X N_X_c_869_n PM_SKY130_FD_SC_HDLL__XNOR3_1%X
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%VPWR N_VPWR_M1000_d N_VPWR_M1004_s
+ N_VPWR_M1014_d N_VPWR_c_888_n N_VPWR_c_889_n VPWR N_VPWR_c_890_n
+ N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_887_n N_VPWR_c_894_n N_VPWR_c_895_n
+ N_VPWR_c_896_n N_VPWR_c_897_n PM_SKY130_FD_SC_HDLL__XNOR3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_351_325# N_A_351_325#_M1013_d
+ N_A_351_325#_M1006_d N_A_351_325#_M1015_s N_A_351_325#_M1011_d
+ N_A_351_325#_c_985_n N_A_351_325#_c_979_n N_A_351_325#_c_980_n
+ N_A_351_325#_c_981_n N_A_351_325#_c_987_n N_A_351_325#_c_988_n
+ N_A_351_325#_c_989_n N_A_351_325#_c_990_n N_A_351_325#_c_982_n
+ N_A_351_325#_c_992_n N_A_351_325#_c_1028_n N_A_351_325#_c_983_n
+ N_A_351_325#_c_993_n N_A_351_325#_c_984_n N_A_351_325#_c_994_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%A_351_325#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_375_49# N_A_375_49#_M1002_s
+ N_A_375_49#_M1019_d N_A_375_49#_M1021_d N_A_375_49#_M1010_d
+ N_A_375_49#_c_1144_n N_A_375_49#_c_1132_n N_A_375_49#_c_1136_n
+ N_A_375_49#_c_1173_n N_A_375_49#_c_1137_n N_A_375_49#_c_1133_n
+ N_A_375_49#_c_1252_p N_A_375_49#_c_1186_n N_A_375_49#_c_1187_n
+ N_A_375_49#_c_1134_n N_A_375_49#_c_1208_n N_A_375_49#_c_1139_n
+ N_A_375_49#_c_1140_n N_A_375_49#_c_1141_n N_A_375_49#_c_1142_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%A_375_49#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%A_1184_297# N_A_1184_297#_M1016_d
+ N_A_1184_297#_M1003_d N_A_1184_297#_M1018_d N_A_1184_297#_M1007_d
+ N_A_1184_297#_c_1268_n N_A_1184_297#_c_1280_n N_A_1184_297#_c_1272_n
+ N_A_1184_297#_c_1269_n N_A_1184_297#_c_1281_n N_A_1184_297#_c_1274_n
+ N_A_1184_297#_c_1270_n PM_SKY130_FD_SC_HDLL__XNOR3_1%A_1184_297#
x_PM_SKY130_FD_SC_HDLL__XNOR3_1%VGND N_VGND_M1012_d N_VGND_M1008_s
+ N_VGND_M1009_d N_VGND_c_1334_n N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n
+ N_VGND_c_1338_n VGND N_VGND_c_1339_n N_VGND_c_1340_n N_VGND_c_1341_n
+ N_VGND_c_1342_n N_VGND_c_1343_n N_VGND_c_1344_n
+ PM_SKY130_FD_SC_HDLL__XNOR3_1%VGND
cc_1 VNB N_A_83_21#_c_152_n 0.020956f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_83_21#_c_153_n 0.0298591f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_3 VNB N_A_83_21#_c_154_n 0.00109789f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_4 VNB N_A_83_21#_c_155_n 0.00138296f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.695
cc_5 VNB N_A_83_21#_c_156_n 0.00216101f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.34
cc_6 VNB N_A_83_21#_c_157_n 0.0163051f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.355
cc_7 VNB N_C_c_251_n 0.0198604f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=0.245
cc_8 VNB N_C_c_252_n 0.0145755f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_9 VNB N_C_c_253_n 0.0217833f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_10 VNB N_C_c_254_n 0.0118432f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_11 VNB N_C_c_255_n 0.0544628f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.33
cc_12 VNB N_A_226_93#_c_311_n 0.0252181f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_13 VNB N_A_226_93#_c_312_n 0.0208877f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_14 VNB N_A_226_93#_c_313_n 0.0026062f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.33
cc_15 VNB N_A_226_93#_c_314_n 0.00274123f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.34
cc_16 VNB N_A_783_297#_M1016_g 0.0360077f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_17 VNB N_A_783_297#_c_382_n 0.00169947f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_18 VNB N_A_783_297#_c_383_n 0.0288368f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.96
cc_19 VNB N_A_783_297#_c_384_n 0.0176837f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.96
cc_20 VNB N_A_783_297#_c_385_n 0.00239744f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.355
cc_21 VNB N_A_783_297#_c_386_n 0.00792514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_783_297#_c_387_n 0.0128101f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.355
cc_23 VNB N_A_783_297#_c_388_n 0.00136794f $X=-0.19 $Y=-0.24 $X2=0.592 $Y2=1.16
cc_24 VNB N_A_783_297#_c_389_n 0.00305152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_783_297#_c_390_n 0.00216737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_783_297#_c_391_n 0.00613074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_783_297#_c_392_n 0.0286332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_783_297#_c_393_n 0.0195573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_783_297#_c_394_n 0.00256224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_B_M1008_g 0.0302339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_B_c_563_n 0.0558482f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_32 VNB N_B_c_564_n 0.0317672f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_33 VNB N_B_M1006_g 0.0287454f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_34 VNB N_B_c_566_n 0.010365f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=2.32
cc_35 VNB N_B_c_567_n 0.00131136f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.355
cc_36 VNB N_B_c_568_n 0.0298426f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.37
cc_37 VNB N_B_c_569_n 0.0212173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_c_698_n 0.0264354f $X=-0.19 $Y=-0.24 $X2=2.345 $Y2=0.245
cc_39 VNB N_A_c_699_n 0.0204396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB A 0.00736307f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_41 VNB N_A_901_297#_c_736_n 0.0299974f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.865
cc_42 VNB N_A_901_297#_c_737_n 0.0219434f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_43 VNB N_A_901_297#_c_738_n 0.00634916f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=0.78
cc_44 VNB N_A_901_297#_c_739_n 0.00633318f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=2.235
cc_45 VNB N_A_901_297#_c_740_n 0.00201667f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.34
cc_46 VNB N_A_901_297#_c_741_n 0.00462287f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.34
cc_47 VNB N_A_901_297#_c_742_n 0.00212326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_901_297#_c_743_n 0.00497895f $X=-0.19 $Y=-0.24 $X2=0.592 $Y2=1.16
cc_49 VNB N_X_c_866_n 0.042291f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_50 VNB N_VPWR_c_887_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_351_325#_c_979_n 0.0107596f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_52 VNB N_A_351_325#_c_980_n 0.0137602f $X=-0.19 $Y=-0.24 $X2=1.1 $Y2=1.96
cc_53 VNB N_A_351_325#_c_981_n 0.00281469f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.425
cc_54 VNB N_A_351_325#_c_982_n 0.00223628f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=2.32
cc_55 VNB N_A_351_325#_c_983_n 0.0104576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_351_325#_c_984_n 2.7378e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_375_49#_c_1132_n 0.00887988f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_58 VNB N_A_375_49#_c_1133_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.425
cc_59 VNB N_A_375_49#_c_1134_n 0.00622338f $X=-0.19 $Y=-0.24 $X2=2.37 $Y2=0.355
cc_60 VNB N_A_1184_297#_c_1268_n 0.00788636f $X=-0.19 $Y=-0.24 $X2=0.635
+ $Y2=1.16
cc_61 VNB N_A_1184_297#_c_1269_n 0.0307904f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=2.045
cc_62 VNB N_A_1184_297#_c_1270_n 0.0135316f $X=-0.19 $Y=-0.24 $X2=2.49 $Y2=0.37
cc_63 VNB N_VGND_c_1334_n 0.00251453f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_64 VNB N_VGND_c_1335_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_65 VNB N_VGND_c_1336_n 0.00637017f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=0.78
cc_66 VNB N_VGND_c_1337_n 0.0678678f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.96
cc_67 VNB N_VGND_c_1338_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.425
cc_68 VNB N_VGND_c_1339_n 0.0154693f $X=-0.19 $Y=-0.24 $X2=1.21 $Y2=2.235
cc_69 VNB N_VGND_c_1340_n 0.109622f $X=-0.19 $Y=-0.24 $X2=2.17 $Y2=0.355
cc_70 VNB N_VGND_c_1341_n 0.0207369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1342_n 0.46301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1343_n 0.0043801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1344_n 0.00881997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_A_83_21#_c_153_n 0.0324414f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_75 VPB N_A_83_21#_c_159_n 0.00153829f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.875
cc_76 VPB N_A_83_21#_c_160_n 0.0038652f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=2.235
cc_77 VPB N_A_83_21#_c_161_n 0.00112766f $X=-0.19 $Y=1.305 $X2=1.32 $Y2=2.32
cc_78 VPB N_A_83_21#_c_162_n 0.0124849f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=2.32
cc_79 VPB N_C_M1017_g 0.0314008f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.995
cc_80 VPB N_C_c_252_n 0.0408591f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_81 VPB N_C_c_254_n 0.00696929f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_82 VPB N_C_c_255_n 0.0248178f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.33
cc_83 VPB N_A_226_93#_c_311_n 0.0344462f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.995
cc_84 VPB N_A_226_93#_c_313_n 0.00441836f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.33
cc_85 VPB N_A_226_93#_c_317_n 0.00959494f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=0.78
cc_86 VPB N_A_226_93#_c_318_n 0.00173389f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.96
cc_87 VPB N_A_226_93#_c_319_n 0.00184072f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.425
cc_88 VPB N_A_226_93#_c_314_n 2.68423e-19 $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.34
cc_89 VPB N_A_783_297#_c_395_n 0.0204513f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.995
cc_90 VPB N_A_783_297#_c_382_n 0.0104623f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=1.16
cc_91 VPB N_A_783_297#_c_397_n 0.0241571f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_92 VPB N_A_783_297#_c_383_n 0.0104543f $X=-0.19 $Y=1.305 $X2=1.1 $Y2=1.96
cc_93 VPB N_A_783_297#_c_384_n 0.00765838f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.96
cc_94 VPB N_A_783_297#_c_400_n 0.00601461f $X=-0.19 $Y=1.305 $X2=1.21 $Y2=2.235
cc_95 VPB N_A_783_297#_c_394_n 0.00321756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_B_c_570_n 0.0216593f $X=-0.19 $Y=1.305 $X2=2.345 $Y2=0.245
cc_97 VPB N_B_c_564_n 0.00748587f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_98 VPB N_B_M1010_g 0.0155244f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=0.865
cc_99 VPB N_B_c_573_n 0.124505f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.33
cc_100 VPB N_B_c_574_n 0.0170126f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.875
cc_101 VPB N_B_c_575_n 0.0101708f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.425
cc_102 VPB N_B_c_576_n 0.00717497f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.695
cc_103 VPB N_B_M1011_g 0.0130994f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.34
cc_104 VPB N_B_c_566_n 0.00875008f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=2.32
cc_105 VPB N_B_c_579_n 0.00204456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_B_c_567_n 9.77983e-19 $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.355
cc_107 VPB N_B_c_568_n 0.00525711f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.37
cc_108 VPB B 0.00802749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_c_698_n 0.0299898f $X=-0.19 $Y=1.305 $X2=2.345 $Y2=0.245
cc_110 VPB A 0.00388732f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.995
cc_111 VPB N_A_901_297#_c_736_n 0.0318269f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=0.865
cc_112 VPB N_A_901_297#_c_738_n 0.00274744f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=0.78
cc_113 VPB N_A_901_297#_c_746_n 0.00189028f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.96
cc_114 VPB N_A_901_297#_c_741_n 3.16686e-19 $X=-0.19 $Y=1.305 $X2=1.205 $Y2=0.34
cc_115 VPB N_A_901_297#_c_748_n 0.00207619f $X=-0.19 $Y=1.305 $X2=1.32 $Y2=2.32
cc_116 VPB N_X_c_866_n 0.00689512f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_117 VPB N_X_c_868_n 0.00673866f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_118 VPB N_X_c_869_n 0.0342476f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_119 VPB N_VPWR_c_888_n 0.00693804f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_120 VPB N_VPWR_c_889_n 0.00743637f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_121 VPB N_VPWR_c_890_n 0.0155059f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=0.78
cc_122 VPB N_VPWR_c_891_n 0.0625838f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.695
cc_123 VPB N_VPWR_c_892_n 0.0165566f $X=-0.19 $Y=1.305 $X2=0.592 $Y2=1.16
cc_124 VPB N_VPWR_c_887_n 0.0709586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_VPWR_c_894_n 0.00589444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_895_n 0.00513206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_896_n 0.0965956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_897_n 0.0123397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_351_325#_c_985_n 0.0110171f $X=-0.19 $Y=1.305 $X2=0.635 $Y2=0.865
cc_130 VPB N_A_351_325#_c_981_n 0.00805098f $X=-0.19 $Y=1.305 $X2=1.095
+ $Y2=0.425
cc_131 VPB N_A_351_325#_c_987_n 0.00296592f $X=-0.19 $Y=1.305 $X2=1.095
+ $Y2=0.695
cc_132 VPB N_A_351_325#_c_988_n 0.00293344f $X=-0.19 $Y=1.305 $X2=2.17 $Y2=0.34
cc_133 VPB N_A_351_325#_c_989_n 0.0106403f $X=-0.19 $Y=1.305 $X2=1.205 $Y2=0.34
cc_134 VPB N_A_351_325#_c_990_n 0.00172555f $X=-0.19 $Y=1.305 $X2=1.32 $Y2=2.32
cc_135 VPB N_A_351_325#_c_982_n 0.00149669f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=2.32
cc_136 VPB N_A_351_325#_c_992_n 0.024643f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.355
cc_137 VPB N_A_351_325#_c_993_n 3.60787e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_351_325#_c_994_n 3.41339e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_375_49#_c_1132_n 0.00148953f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_140 VPB N_A_375_49#_c_1136_n 0.00271724f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_141 VPB N_A_375_49#_c_1137_n 8.62277e-19 $X=-0.19 $Y=1.305 $X2=0.755 $Y2=0.78
cc_142 VPB N_A_375_49#_c_1133_n 0.0021572f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.425
cc_143 VPB N_A_375_49#_c_1139_n 0.0147524f $X=-0.19 $Y=1.305 $X2=2.49 $Y2=0.37
cc_144 VPB N_A_375_49#_c_1140_n 0.00333347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_375_49#_c_1141_n 0.008761f $X=-0.19 $Y=1.305 $X2=0.592 $Y2=1.16
cc_146 VPB N_A_375_49#_c_1142_n 0.00154407f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_1184_297#_c_1268_n 0.00468751f $X=-0.19 $Y=1.305 $X2=0.635
+ $Y2=1.16
cc_148 VPB N_A_1184_297#_c_1272_n 0.0147295f $X=-0.19 $Y=1.305 $X2=0.755
+ $Y2=1.96
cc_149 VPB N_A_1184_297#_c_1269_n 0.0229985f $X=-0.19 $Y=1.305 $X2=1.21
+ $Y2=2.045
cc_150 VPB N_A_1184_297#_c_1274_n 0.0101148f $X=-0.19 $Y=1.305 $X2=2.415
+ $Y2=2.32
cc_151 N_A_83_21#_c_152_n N_C_c_251_n 0.0133179f $X=0.49 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_83_21#_c_154_n N_C_c_251_n 0.00139501f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_83_21#_c_165_p N_C_c_251_n 0.0120994f $X=0.985 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_83_21#_c_155_n N_C_c_251_n 0.0106802f $X=1.095 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_83_21#_c_156_n N_C_c_251_n 0.00609535f $X=1.205 $Y=0.34 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_83_21#_c_153_n N_C_M1017_g 0.0216907f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_83_21#_c_159_n N_C_M1017_g 0.00555142f $X=0.645 $Y=1.875 $X2=0 $Y2=0
cc_158 N_A_83_21#_c_170_p N_C_M1017_g 0.0132115f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_159 N_A_83_21#_c_160_n N_C_M1017_g 0.00742917f $X=1.21 $Y=2.235 $X2=0 $Y2=0
cc_160 N_A_83_21#_c_161_n N_C_M1017_g 0.00743853f $X=1.32 $Y=2.32 $X2=0 $Y2=0
cc_161 N_A_83_21#_c_162_n N_C_c_252_n 0.0112964f $X=2.415 $Y=2.32 $X2=0 $Y2=0
cc_162 N_A_83_21#_c_174_p N_C_c_253_n 0.0106037f $X=2.37 $Y=0.355 $X2=0 $Y2=0
cc_163 N_A_83_21#_c_153_n N_C_c_254_n 0.0253799f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_83_21#_c_154_n N_C_c_254_n 0.00159638f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_83_21#_c_177_p N_C_c_254_n 8.8646e-19 $X=0.635 $Y=1.33 $X2=0 $Y2=0
cc_166 N_A_83_21#_c_157_n N_C_c_255_n 0.0111296f $X=2.17 $Y=0.355 $X2=0 $Y2=0
cc_167 N_A_83_21#_c_157_n C 0.00344638f $X=2.17 $Y=0.355 $X2=0 $Y2=0
cc_168 N_A_83_21#_c_165_p N_A_226_93#_M1020_d 0.00226213f $X=0.985 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_169 N_A_83_21#_c_155_n N_A_226_93#_M1020_d 0.00618081f $X=1.095 $Y=0.695
+ $X2=-0.19 $Y2=-0.24
cc_170 N_A_83_21#_c_170_p N_A_226_93#_M1017_d 0.00416203f $X=1.1 $Y=1.96 $X2=0
+ $Y2=0
cc_171 N_A_83_21#_c_160_n N_A_226_93#_M1017_d 0.00266846f $X=1.21 $Y=2.235 $X2=0
+ $Y2=0
cc_172 N_A_83_21#_c_162_n N_A_226_93#_c_311_n 0.0116412f $X=2.415 $Y=2.32 $X2=0
+ $Y2=0
cc_173 N_A_83_21#_c_165_p N_A_226_93#_c_326_n 0.00409956f $X=0.985 $Y=0.78 $X2=0
+ $Y2=0
cc_174 N_A_83_21#_c_170_p N_A_226_93#_c_326_n 0.0200253f $X=1.1 $Y=1.96 $X2=0
+ $Y2=0
cc_175 N_A_83_21#_c_162_n N_A_226_93#_c_326_n 0.00176797f $X=2.415 $Y=2.32 $X2=0
+ $Y2=0
cc_176 N_A_83_21#_c_153_n N_A_226_93#_c_313_n 6.59446e-19 $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_83_21#_c_154_n N_A_226_93#_c_313_n 0.0181f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_83_21#_c_165_p N_A_226_93#_c_313_n 0.0138474f $X=0.985 $Y=0.78 $X2=0
+ $Y2=0
cc_179 N_A_83_21#_c_155_n N_A_226_93#_c_313_n 0.00736858f $X=1.095 $Y=0.695
+ $X2=0 $Y2=0
cc_180 N_A_83_21#_c_157_n N_A_226_93#_c_313_n 0.0130244f $X=2.17 $Y=0.355 $X2=0
+ $Y2=0
cc_181 N_A_83_21#_M1015_d N_A_226_93#_c_317_n 0.00779963f $X=2.27 $Y=1.625 $X2=0
+ $Y2=0
cc_182 N_A_83_21#_c_162_n N_A_226_93#_c_317_n 0.0039224f $X=2.415 $Y=2.32 $X2=0
+ $Y2=0
cc_183 N_A_83_21#_M1015_d N_A_226_93#_c_318_n 5.89264e-19 $X=2.27 $Y=1.625 $X2=0
+ $Y2=0
cc_184 N_A_83_21#_c_162_n N_A_226_93#_c_319_n 0.00633062f $X=2.415 $Y=2.32 $X2=0
+ $Y2=0
cc_185 N_A_83_21#_c_152_n N_X_c_866_n 0.0182824f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_83_21#_c_153_n N_X_c_866_n 6.56726e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_83_21#_c_154_n N_X_c_866_n 0.0351422f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_188 N_A_83_21#_c_159_n N_X_c_866_n 0.00752799f $X=0.645 $Y=1.875 $X2=0 $Y2=0
cc_189 N_A_83_21#_c_201_p N_X_c_866_n 0.0137849f $X=0.755 $Y=0.78 $X2=0 $Y2=0
cc_190 N_A_83_21#_c_155_n N_X_c_866_n 0.00438168f $X=1.095 $Y=0.695 $X2=0 $Y2=0
cc_191 N_A_83_21#_c_153_n N_X_c_868_n 0.00725258f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_83_21#_c_159_n N_X_c_868_n 0.0323512f $X=0.645 $Y=1.875 $X2=0 $Y2=0
cc_193 N_A_83_21#_c_205_p N_X_c_869_n 0.0138426f $X=0.755 $Y=1.96 $X2=0 $Y2=0
cc_194 N_A_83_21#_c_159_n N_VPWR_M1000_d 0.00451219f $X=0.645 $Y=1.875 $X2=-0.19
+ $Y2=-0.24
cc_195 N_A_83_21#_c_170_p N_VPWR_M1000_d 0.00859265f $X=1.1 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A_83_21#_c_205_p N_VPWR_M1000_d 9.86211e-19 $X=0.755 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_197 N_A_83_21#_c_153_n N_VPWR_c_888_n 0.0126469f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_83_21#_c_170_p N_VPWR_c_888_n 0.0126548f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_199 N_A_83_21#_c_205_p N_VPWR_c_888_n 0.0133756f $X=0.755 $Y=1.96 $X2=0 $Y2=0
cc_200 N_A_83_21#_c_160_n N_VPWR_c_888_n 0.00145799f $X=1.21 $Y=2.235 $X2=0
+ $Y2=0
cc_201 N_A_83_21#_c_161_n N_VPWR_c_888_n 0.0137789f $X=1.32 $Y=2.32 $X2=0 $Y2=0
cc_202 N_A_83_21#_c_153_n N_VPWR_c_890_n 0.00427505f $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_83_21#_c_170_p N_VPWR_c_891_n 0.00233941f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_204 N_A_83_21#_c_161_n N_VPWR_c_891_n 0.0109705f $X=1.32 $Y=2.32 $X2=0 $Y2=0
cc_205 N_A_83_21#_c_162_n N_VPWR_c_891_n 0.0597844f $X=2.415 $Y=2.32 $X2=0 $Y2=0
cc_206 N_A_83_21#_c_153_n N_VPWR_c_887_n 0.00825932f $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_83_21#_c_170_p N_VPWR_c_887_n 0.00553584f $X=1.1 $Y=1.96 $X2=0 $Y2=0
cc_208 N_A_83_21#_c_205_p N_VPWR_c_887_n 9.98534e-19 $X=0.755 $Y=1.96 $X2=0
+ $Y2=0
cc_209 N_A_83_21#_c_161_n N_VPWR_c_887_n 0.00809357f $X=1.32 $Y=2.32 $X2=0 $Y2=0
cc_210 N_A_83_21#_c_162_n N_VPWR_c_887_n 0.0473531f $X=2.415 $Y=2.32 $X2=0 $Y2=0
cc_211 N_A_83_21#_c_162_n N_A_351_325#_M1015_s 0.00736441f $X=2.415 $Y=2.32
+ $X2=0 $Y2=0
cc_212 N_A_83_21#_M1015_d N_A_351_325#_c_985_n 0.00509381f $X=2.27 $Y=1.625
+ $X2=0 $Y2=0
cc_213 N_A_83_21#_c_170_p N_A_351_325#_c_985_n 0.00831987f $X=1.1 $Y=1.96 $X2=0
+ $Y2=0
cc_214 N_A_83_21#_c_160_n N_A_351_325#_c_985_n 9.56599e-19 $X=1.21 $Y=2.235
+ $X2=0 $Y2=0
cc_215 N_A_83_21#_c_162_n N_A_351_325#_c_985_n 0.0571361f $X=2.415 $Y=2.32 $X2=0
+ $Y2=0
cc_216 N_A_83_21#_c_157_n N_A_375_49#_M1002_s 0.00652268f $X=2.17 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_217 N_A_83_21#_M1002_d N_A_375_49#_c_1144_n 0.00732564f $X=2.345 $Y=0.245
+ $X2=0 $Y2=0
cc_218 N_A_83_21#_c_230_p N_A_375_49#_c_1144_n 0.0127434f $X=2.49 $Y=0.37 $X2=0
+ $Y2=0
cc_219 N_A_83_21#_c_174_p N_A_375_49#_c_1134_n 0.0127434f $X=2.37 $Y=0.355 $X2=0
+ $Y2=0
cc_220 N_A_83_21#_c_157_n N_A_375_49#_c_1134_n 0.0181831f $X=2.17 $Y=0.355 $X2=0
+ $Y2=0
cc_221 N_A_83_21#_c_154_n N_VGND_M1012_d 2.82564e-19 $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_222 N_A_83_21#_c_165_p N_VGND_M1012_d 0.00889686f $X=0.985 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_223 N_A_83_21#_c_201_p N_VGND_M1012_d 0.00149651f $X=0.755 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_224 N_A_83_21#_c_152_n N_VGND_c_1334_n 0.0143349f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_83_21#_c_153_n N_VGND_c_1334_n 7.15202e-19 $X=0.515 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_83_21#_c_165_p N_VGND_c_1334_n 0.0045481f $X=0.985 $Y=0.78 $X2=0
+ $Y2=0
cc_227 N_A_83_21#_c_201_p N_VGND_c_1334_n 0.0153068f $X=0.755 $Y=0.78 $X2=0
+ $Y2=0
cc_228 N_A_83_21#_c_155_n N_VGND_c_1334_n 0.00744451f $X=1.095 $Y=0.695 $X2=0
+ $Y2=0
cc_229 N_A_83_21#_c_156_n N_VGND_c_1334_n 0.0142743f $X=1.205 $Y=0.34 $X2=0
+ $Y2=0
cc_230 N_A_83_21#_c_165_p N_VGND_c_1337_n 0.00219715f $X=0.985 $Y=0.78 $X2=0
+ $Y2=0
cc_231 N_A_83_21#_c_156_n N_VGND_c_1337_n 0.0156439f $X=1.205 $Y=0.34 $X2=0
+ $Y2=0
cc_232 N_A_83_21#_c_157_n N_VGND_c_1337_n 0.0885651f $X=2.17 $Y=0.355 $X2=0
+ $Y2=0
cc_233 N_A_83_21#_c_152_n N_VGND_c_1339_n 0.00388479f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_234 N_A_83_21#_c_152_n N_VGND_c_1342_n 0.00774695f $X=0.49 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_83_21#_c_165_p N_VGND_c_1342_n 0.00486078f $X=0.985 $Y=0.78 $X2=0
+ $Y2=0
cc_236 N_A_83_21#_c_201_p N_VGND_c_1342_n 0.00106517f $X=0.755 $Y=0.78 $X2=0
+ $Y2=0
cc_237 N_A_83_21#_c_156_n N_VGND_c_1342_n 0.00844855f $X=1.205 $Y=0.34 $X2=0
+ $Y2=0
cc_238 N_A_83_21#_c_157_n N_VGND_c_1342_n 0.0533662f $X=2.17 $Y=0.355 $X2=0
+ $Y2=0
cc_239 N_C_c_252_n N_A_226_93#_c_311_n 0.0592216f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_240 C N_A_226_93#_c_311_n 2.68329e-19 $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_241 N_C_c_253_n N_A_226_93#_c_312_n 0.0213405f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_242 N_C_M1017_g N_A_226_93#_c_326_n 0.011319f $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_243 N_C_c_255_n N_A_226_93#_c_326_n 0.00634718f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_244 N_C_c_251_n N_A_226_93#_c_313_n 0.0043646f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_245 N_C_M1017_g N_A_226_93#_c_313_n 0.00203559f $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_246 N_C_c_252_n N_A_226_93#_c_313_n 0.00508695f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_247 N_C_c_253_n N_A_226_93#_c_313_n 0.00235914f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_248 N_C_c_254_n N_A_226_93#_c_313_n 0.0020376f $X=1.08 $Y=1.202 $X2=0 $Y2=0
cc_249 N_C_c_255_n N_A_226_93#_c_313_n 0.026637f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_250 C N_A_226_93#_c_313_n 0.018733f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_251 N_C_c_252_n N_A_226_93#_c_317_n 0.017213f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_252 N_C_c_255_n N_A_226_93#_c_317_n 0.0140512f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_253 C N_A_226_93#_c_317_n 0.0378363f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_254 N_C_c_252_n N_A_226_93#_c_318_n 0.00427971f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_255 N_C_c_252_n N_A_226_93#_c_314_n 0.00353238f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_256 C N_A_226_93#_c_314_n 0.0207305f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_257 N_C_M1017_g N_VPWR_c_888_n 0.00202848f $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_258 N_C_M1017_g N_VPWR_c_891_n 0.00514356f $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_259 N_C_c_252_n N_VPWR_c_891_n 0.00427564f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_260 N_C_M1017_g N_VPWR_c_887_n 0.00682402f $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_261 N_C_c_252_n N_VPWR_c_887_n 0.00784458f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_262 N_C_M1017_g N_A_351_325#_c_985_n 9.4239e-19 $X=1.08 $Y=1.805 $X2=0 $Y2=0
cc_263 N_C_c_252_n N_A_351_325#_c_985_n 0.0102234f $X=2.18 $Y=1.55 $X2=0 $Y2=0
cc_264 N_C_c_253_n N_A_375_49#_c_1144_n 0.0082764f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_265 C N_A_375_49#_c_1144_n 0.00489958f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_266 N_C_c_253_n N_A_375_49#_c_1134_n 0.00382666f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_267 N_C_c_255_n N_A_375_49#_c_1134_n 0.00656019f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_268 C N_A_375_49#_c_1134_n 0.028934f $X=1.985 $Y=1.105 $X2=0 $Y2=0
cc_269 N_C_c_251_n N_VGND_c_1334_n 0.00138119f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_270 N_C_c_251_n N_VGND_c_1337_n 8.79444e-19 $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_271 N_C_c_253_n N_VGND_c_1337_n 0.00357877f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_272 N_C_c_253_n N_VGND_c_1342_n 0.0068382f $X=2.27 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_226_93#_c_311_n N_VPWR_c_889_n 0.00632978f $X=2.715 $Y=1.41 $X2=0
+ $Y2=0
cc_274 N_A_226_93#_c_311_n N_VPWR_c_891_n 0.00412251f $X=2.715 $Y=1.41 $X2=0
+ $Y2=0
cc_275 N_A_226_93#_c_311_n N_VPWR_c_887_n 0.00595559f $X=2.715 $Y=1.41 $X2=0
+ $Y2=0
cc_276 N_A_226_93#_c_317_n N_A_351_325#_M1015_s 0.00373918f $X=2.5 $Y=1.62 $X2=0
+ $Y2=0
cc_277 N_A_226_93#_c_311_n N_A_351_325#_c_985_n 0.0182967f $X=2.715 $Y=1.41
+ $X2=0 $Y2=0
cc_278 N_A_226_93#_c_317_n N_A_351_325#_c_985_n 0.0556467f $X=2.5 $Y=1.62 $X2=0
+ $Y2=0
cc_279 N_A_226_93#_c_314_n N_A_351_325#_c_985_n 0.00386917f $X=2.69 $Y=1.16
+ $X2=0 $Y2=0
cc_280 N_A_226_93#_c_312_n N_A_351_325#_c_980_n 0.00496015f $X=2.76 $Y=0.995
+ $X2=0 $Y2=0
cc_281 N_A_226_93#_c_311_n N_A_351_325#_c_981_n 0.00449957f $X=2.715 $Y=1.41
+ $X2=0 $Y2=0
cc_282 N_A_226_93#_c_311_n N_A_375_49#_c_1144_n 0.00296047f $X=2.715 $Y=1.41
+ $X2=0 $Y2=0
cc_283 N_A_226_93#_c_312_n N_A_375_49#_c_1144_n 0.0140125f $X=2.76 $Y=0.995
+ $X2=0 $Y2=0
cc_284 N_A_226_93#_c_314_n N_A_375_49#_c_1144_n 0.0192251f $X=2.69 $Y=1.16 $X2=0
+ $Y2=0
cc_285 N_A_226_93#_c_311_n N_A_375_49#_c_1132_n 0.0089074f $X=2.715 $Y=1.41
+ $X2=0 $Y2=0
cc_286 N_A_226_93#_c_312_n N_A_375_49#_c_1132_n 0.00688718f $X=2.76 $Y=0.995
+ $X2=0 $Y2=0
cc_287 N_A_226_93#_c_318_n N_A_375_49#_c_1132_n 0.00218396f $X=2.585 $Y=1.535
+ $X2=0 $Y2=0
cc_288 N_A_226_93#_c_314_n N_A_375_49#_c_1132_n 0.0247426f $X=2.69 $Y=1.16 $X2=0
+ $Y2=0
cc_289 N_A_226_93#_c_312_n N_A_375_49#_c_1134_n 5.22054e-19 $X=2.76 $Y=0.995
+ $X2=0 $Y2=0
cc_290 N_A_226_93#_c_313_n N_A_375_49#_c_1134_n 0.0151384f $X=1.46 $Y=0.76 $X2=0
+ $Y2=0
cc_291 N_A_226_93#_c_317_n N_A_375_49#_c_1140_n 5.94479e-19 $X=2.5 $Y=1.62 $X2=0
+ $Y2=0
cc_292 N_A_226_93#_c_318_n N_A_375_49#_c_1140_n 6.54862e-19 $X=2.585 $Y=1.535
+ $X2=0 $Y2=0
cc_293 N_A_226_93#_c_311_n N_A_375_49#_c_1141_n 0.00719438f $X=2.715 $Y=1.41
+ $X2=0 $Y2=0
cc_294 N_A_226_93#_c_317_n N_A_375_49#_c_1141_n 0.0102953f $X=2.5 $Y=1.62 $X2=0
+ $Y2=0
cc_295 N_A_226_93#_c_318_n N_A_375_49#_c_1141_n 0.00669828f $X=2.585 $Y=1.535
+ $X2=0 $Y2=0
cc_296 N_A_226_93#_c_312_n N_VGND_c_1337_n 0.0042361f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_297 N_A_226_93#_c_312_n N_VGND_c_1342_n 0.00742704f $X=2.76 $Y=0.995 $X2=0
+ $Y2=0
cc_298 N_A_783_297#_c_400_n N_B_c_570_n 0.00852064f $X=4.22 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_783_297#_c_394_n N_B_c_570_n 8.18494e-19 $X=4.28 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_783_297#_c_404_p N_B_M1008_g 0.00381578f $X=4.305 $Y=0.85 $X2=0 $Y2=0
cc_301 N_A_783_297#_c_394_n N_B_M1008_g 0.0178285f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_302 N_A_783_297#_c_386_n N_B_c_563_n 0.0050801f $X=5.495 $Y=0.85 $X2=0 $Y2=0
cc_303 N_A_783_297#_c_394_n N_B_c_563_n 0.0122706f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_304 N_A_783_297#_c_400_n N_B_c_564_n 0.00748737f $X=4.22 $Y=1.58 $X2=0 $Y2=0
cc_305 N_A_783_297#_c_394_n N_B_c_564_n 0.00955042f $X=4.28 $Y=0.74 $X2=0 $Y2=0
cc_306 N_A_783_297#_c_395_n N_B_M1010_g 0.0119272f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_783_297#_M1016_g N_B_M1006_g 0.0102876f $X=5.855 $Y=0.455 $X2=0 $Y2=0
cc_308 N_A_783_297#_c_383_n N_B_M1006_g 0.021209f $X=5.73 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A_783_297#_c_385_n N_B_M1006_g 0.00188578f $X=5.62 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A_783_297#_c_386_n N_B_M1006_g 0.00148554f $X=5.495 $Y=0.85 $X2=0 $Y2=0
cc_311 N_A_783_297#_c_388_n N_B_M1006_g 6.75018e-19 $X=5.785 $Y=0.85 $X2=0 $Y2=0
cc_312 N_A_783_297#_c_389_n N_B_M1006_g 0.00122796f $X=5.64 $Y=0.85 $X2=0 $Y2=0
cc_313 N_A_783_297#_c_395_n N_B_c_573_n 0.0105804f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_783_297#_c_397_n N_B_c_573_n 0.00616735f $X=7.32 $Y=1.57 $X2=0 $Y2=0
cc_315 N_A_783_297#_c_382_n N_B_c_575_n 0.00407979f $X=7.32 $Y=1.47 $X2=0 $Y2=0
cc_316 N_A_783_297#_c_397_n N_B_c_576_n 0.00407979f $X=7.32 $Y=1.57 $X2=0 $Y2=0
cc_317 N_A_783_297#_c_397_n N_B_M1011_g 0.0249809f $X=7.32 $Y=1.57 $X2=0 $Y2=0
cc_318 N_A_783_297#_c_384_n N_B_c_566_n 0.00181049f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_319 N_A_783_297#_c_382_n N_B_c_567_n 9.03117e-19 $X=7.32 $Y=1.47 $X2=0 $Y2=0
cc_320 N_A_783_297#_c_387_n N_B_c_567_n 0.00731236f $X=6.975 $Y=0.85 $X2=0 $Y2=0
cc_321 N_A_783_297#_c_391_n N_B_c_567_n 0.021521f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_322 N_A_783_297#_c_392_n N_B_c_567_n 2.70696e-19 $X=7.24 $Y=1.11 $X2=0 $Y2=0
cc_323 N_A_783_297#_c_382_n N_B_c_568_n 0.00185712f $X=7.32 $Y=1.47 $X2=0 $Y2=0
cc_324 N_A_783_297#_c_384_n N_B_c_568_n 0.00774709f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_325 N_A_783_297#_c_387_n N_B_c_568_n 0.00133312f $X=6.975 $Y=0.85 $X2=0 $Y2=0
cc_326 N_A_783_297#_c_391_n N_B_c_568_n 0.00172718f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_327 N_A_783_297#_c_392_n N_B_c_568_n 0.0173414f $X=7.24 $Y=1.11 $X2=0 $Y2=0
cc_328 N_A_783_297#_c_382_n B 0.00133275f $X=7.32 $Y=1.47 $X2=0 $Y2=0
cc_329 N_A_783_297#_c_397_n B 0.00483815f $X=7.32 $Y=1.57 $X2=0 $Y2=0
cc_330 N_A_783_297#_c_387_n B 0.00414594f $X=6.975 $Y=0.85 $X2=0 $Y2=0
cc_331 N_A_783_297#_c_390_n B 0.00235209f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_332 N_A_783_297#_c_391_n B 0.0183366f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_333 N_A_783_297#_c_392_n B 8.1069e-19 $X=7.24 $Y=1.11 $X2=0 $Y2=0
cc_334 N_A_783_297#_M1016_g N_B_c_569_n 0.00774709f $X=5.855 $Y=0.455 $X2=0
+ $Y2=0
cc_335 N_A_783_297#_c_387_n N_B_c_569_n 0.0073961f $X=6.975 $Y=0.85 $X2=0 $Y2=0
cc_336 N_A_783_297#_c_390_n N_B_c_569_n 0.00141075f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_337 N_A_783_297#_c_391_n N_B_c_569_n 0.00206736f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_338 N_A_783_297#_c_392_n N_B_c_569_n 0.00135765f $X=7.24 $Y=1.11 $X2=0 $Y2=0
cc_339 N_A_783_297#_c_393_n N_B_c_569_n 0.0136423f $X=7.262 $Y=0.945 $X2=0 $Y2=0
cc_340 N_A_783_297#_c_382_n N_A_c_698_n 0.00765017f $X=7.32 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_341 N_A_783_297#_c_397_n N_A_c_698_n 0.0315589f $X=7.32 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_342 N_A_783_297#_c_391_n N_A_c_698_n 6.31262e-19 $X=7.12 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_343 N_A_783_297#_c_392_n N_A_c_698_n 0.020199f $X=7.24 $Y=1.11 $X2=-0.19
+ $Y2=-0.24
cc_344 N_A_783_297#_c_391_n N_A_c_699_n 2.39914e-19 $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_345 N_A_783_297#_c_393_n N_A_c_699_n 0.0185647f $X=7.262 $Y=0.945 $X2=0 $Y2=0
cc_346 N_A_783_297#_c_391_n A 0.016871f $X=7.12 $Y=0.85 $X2=0 $Y2=0
cc_347 N_A_783_297#_c_392_n A 0.00221618f $X=7.24 $Y=1.11 $X2=0 $Y2=0
cc_348 N_A_783_297#_c_386_n N_A_901_297#_M1006_s 8.58636e-19 $X=5.495 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_349 N_A_783_297#_c_400_n N_A_901_297#_c_738_n 0.0194501f $X=4.22 $Y=1.58
+ $X2=0 $Y2=0
cc_350 N_A_783_297#_c_386_n N_A_901_297#_c_738_n 0.0124002f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_351 N_A_783_297#_c_404_p N_A_901_297#_c_738_n 5.77119e-19 $X=4.305 $Y=0.85
+ $X2=0 $Y2=0
cc_352 N_A_783_297#_c_394_n N_A_901_297#_c_738_n 0.0604107f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_353 N_A_783_297#_c_397_n N_A_901_297#_c_746_n 0.00416703f $X=7.32 $Y=1.57
+ $X2=0 $Y2=0
cc_354 N_A_783_297#_c_390_n N_A_901_297#_c_740_n 0.00537182f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_355 N_A_783_297#_c_391_n N_A_901_297#_c_740_n 0.0052004f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_356 N_A_783_297#_c_393_n N_A_901_297#_c_740_n 0.00186387f $X=7.262 $Y=0.945
+ $X2=0 $Y2=0
cc_357 N_A_783_297#_M1016_g N_A_901_297#_c_758_n 0.00613906f $X=5.855 $Y=0.455
+ $X2=0 $Y2=0
cc_358 N_A_783_297#_c_385_n N_A_901_297#_c_758_n 3.69046e-19 $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_359 N_A_783_297#_c_386_n N_A_901_297#_c_758_n 0.0529767f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_360 N_A_783_297#_c_387_n N_A_901_297#_c_758_n 0.0955498f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_361 N_A_783_297#_c_388_n N_A_901_297#_c_758_n 0.026662f $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_362 N_A_783_297#_c_389_n N_A_901_297#_c_758_n 0.00310602f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_363 N_A_783_297#_c_390_n N_A_901_297#_c_758_n 0.0266136f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_783_297#_c_391_n N_A_901_297#_c_758_n 0.00475925f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_365 N_A_783_297#_c_393_n N_A_901_297#_c_758_n 0.00868614f $X=7.262 $Y=0.945
+ $X2=0 $Y2=0
cc_366 N_A_783_297#_c_386_n N_A_901_297#_c_742_n 0.0261258f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_367 N_A_783_297#_c_394_n N_A_901_297#_c_742_n 0.00683584f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_368 N_A_783_297#_c_386_n N_A_901_297#_c_743_n 0.00108548f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_369 N_A_783_297#_c_394_n N_A_901_297#_c_743_n 0.01151f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_370 N_A_783_297#_c_393_n N_A_901_297#_c_771_n 0.00156339f $X=7.262 $Y=0.945
+ $X2=0 $Y2=0
cc_371 N_A_783_297#_c_393_n N_A_901_297#_c_772_n 0.00805147f $X=7.262 $Y=0.945
+ $X2=0 $Y2=0
cc_372 N_A_783_297#_M1004_d N_VPWR_c_887_n 0.00367747f $X=3.915 $Y=1.485 $X2=0
+ $Y2=0
cc_373 N_A_783_297#_c_397_n N_VPWR_c_887_n 0.00650675f $X=7.32 $Y=1.57 $X2=0
+ $Y2=0
cc_374 N_A_783_297#_c_397_n N_VPWR_c_896_n 0.00434439f $X=7.32 $Y=1.57 $X2=0
+ $Y2=0
cc_375 N_A_783_297#_c_397_n N_VPWR_c_897_n 0.00129289f $X=7.32 $Y=1.57 $X2=0
+ $Y2=0
cc_376 N_A_783_297#_c_386_n N_A_351_325#_M1006_d 0.00134889f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_377 N_A_783_297#_c_388_n N_A_351_325#_M1006_d 5.4759e-19 $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_378 N_A_783_297#_c_389_n N_A_351_325#_M1006_d 0.00649965f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_379 N_A_783_297#_c_404_p N_A_351_325#_c_980_n 0.0023462f $X=4.305 $Y=0.85
+ $X2=0 $Y2=0
cc_380 N_A_783_297#_c_394_n N_A_351_325#_c_980_n 0.00358611f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_381 N_A_783_297#_c_400_n N_A_351_325#_c_981_n 0.0144171f $X=4.22 $Y=1.58
+ $X2=0 $Y2=0
cc_382 N_A_783_297#_c_394_n N_A_351_325#_c_981_n 0.00928178f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_383 N_A_783_297#_M1004_d N_A_351_325#_c_987_n 0.00767171f $X=3.915 $Y=1.485
+ $X2=0 $Y2=0
cc_384 N_A_783_297#_c_400_n N_A_351_325#_c_987_n 0.0315546f $X=4.22 $Y=1.58
+ $X2=0 $Y2=0
cc_385 N_A_783_297#_M1004_d N_A_351_325#_c_988_n 0.00313827f $X=3.915 $Y=1.485
+ $X2=0 $Y2=0
cc_386 N_A_783_297#_M1004_d N_A_351_325#_c_990_n 0.00318432f $X=3.915 $Y=1.485
+ $X2=0 $Y2=0
cc_387 N_A_783_297#_c_395_n N_A_351_325#_c_982_n 0.00131578f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_388 N_A_783_297#_c_383_n N_A_351_325#_c_982_n 6.52616e-19 $X=5.73 $Y=1.16
+ $X2=0 $Y2=0
cc_389 N_A_783_297#_c_384_n N_A_351_325#_c_982_n 3.9697e-19 $X=5.83 $Y=1.202
+ $X2=0 $Y2=0
cc_390 N_A_783_297#_c_385_n N_A_351_325#_c_982_n 0.0160828f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_391 N_A_783_297#_c_386_n N_A_351_325#_c_982_n 0.00616329f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_392 N_A_783_297#_c_388_n N_A_351_325#_c_982_n 0.00105141f $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_393 N_A_783_297#_c_389_n N_A_351_325#_c_982_n 0.00264545f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_394 N_A_783_297#_c_395_n N_A_351_325#_c_992_n 0.00258134f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_395 N_A_783_297#_c_397_n N_A_351_325#_c_992_n 0.00822576f $X=7.32 $Y=1.57
+ $X2=0 $Y2=0
cc_396 N_A_783_297#_M1016_g N_A_351_325#_c_1028_n 0.00223132f $X=5.855 $Y=0.455
+ $X2=0 $Y2=0
cc_397 N_A_783_297#_c_389_n N_A_351_325#_c_1028_n 0.00180873f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_398 N_A_783_297#_c_394_n N_A_351_325#_c_983_n 0.00616338f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_399 N_A_783_297#_c_383_n N_A_351_325#_c_984_n 2.22283e-19 $X=5.73 $Y=1.16
+ $X2=0 $Y2=0
cc_400 N_A_783_297#_c_385_n N_A_351_325#_c_984_n 0.00299453f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_401 N_A_783_297#_c_386_n N_A_351_325#_c_984_n 0.0171949f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_402 N_A_783_297#_c_388_n N_A_351_325#_c_984_n 0.00134696f $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_403 N_A_783_297#_c_389_n N_A_351_325#_c_984_n 0.0141636f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_404 N_A_783_297#_c_387_n N_A_375_49#_M1019_d 0.00140408f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_405 N_A_783_297#_c_390_n N_A_375_49#_M1019_d 0.00214439f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_406 N_A_783_297#_c_391_n N_A_375_49#_M1019_d 0.0050343f $X=7.12 $Y=0.85 $X2=0
+ $Y2=0
cc_407 N_A_783_297#_c_383_n N_A_375_49#_c_1136_n 0.00881942f $X=5.73 $Y=1.16
+ $X2=0 $Y2=0
cc_408 N_A_783_297#_c_385_n N_A_375_49#_c_1136_n 0.0271004f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_409 N_A_783_297#_c_386_n N_A_375_49#_c_1136_n 5.63647e-19 $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_410 N_A_783_297#_c_395_n N_A_375_49#_c_1173_n 0.00383389f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_411 N_A_783_297#_c_395_n N_A_375_49#_c_1137_n 0.0175777f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_412 N_A_783_297#_c_383_n N_A_375_49#_c_1137_n 7.42472e-19 $X=5.73 $Y=1.16
+ $X2=0 $Y2=0
cc_413 N_A_783_297#_c_384_n N_A_375_49#_c_1137_n 9.0109e-19 $X=5.83 $Y=1.202
+ $X2=0 $Y2=0
cc_414 N_A_783_297#_c_385_n N_A_375_49#_c_1137_n 0.00152864f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_415 N_A_783_297#_c_387_n N_A_375_49#_c_1137_n 0.00419686f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_416 N_A_783_297#_c_388_n N_A_375_49#_c_1137_n 6.55203e-19 $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_783_297#_c_395_n N_A_375_49#_c_1133_n 0.00139259f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_418 N_A_783_297#_M1016_g N_A_375_49#_c_1133_n 0.0164012f $X=5.855 $Y=0.455
+ $X2=0 $Y2=0
cc_419 N_A_783_297#_c_385_n N_A_375_49#_c_1133_n 0.0173003f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_420 N_A_783_297#_c_387_n N_A_375_49#_c_1133_n 0.0173494f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_421 N_A_783_297#_c_388_n N_A_375_49#_c_1133_n 0.00232583f $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_422 N_A_783_297#_c_389_n N_A_375_49#_c_1133_n 0.0185267f $X=5.64 $Y=0.85
+ $X2=0 $Y2=0
cc_423 N_A_783_297#_c_387_n N_A_375_49#_c_1186_n 0.00166303f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_424 N_A_783_297#_c_390_n N_A_375_49#_c_1187_n 3.55136e-19 $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_425 N_A_783_297#_c_391_n N_A_375_49#_c_1187_n 0.00528249f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_426 N_A_783_297#_c_393_n N_A_375_49#_c_1187_n 0.00335197f $X=7.262 $Y=0.945
+ $X2=0 $Y2=0
cc_427 N_A_783_297#_c_400_n N_A_375_49#_c_1139_n 0.0275977f $X=4.22 $Y=1.58
+ $X2=0 $Y2=0
cc_428 N_A_783_297#_c_385_n N_A_375_49#_c_1139_n 8.40027e-19 $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_429 N_A_783_297#_c_386_n N_A_375_49#_c_1139_n 0.0525103f $X=5.495 $Y=0.85
+ $X2=0 $Y2=0
cc_430 N_A_783_297#_c_404_p N_A_375_49#_c_1139_n 0.0124731f $X=4.305 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_783_297#_c_394_n N_A_375_49#_c_1139_n 0.00234688f $X=4.28 $Y=0.74
+ $X2=0 $Y2=0
cc_432 N_A_783_297#_c_395_n N_A_375_49#_c_1142_n 0.00348376f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_433 N_A_783_297#_c_383_n N_A_375_49#_c_1142_n 0.00431105f $X=5.73 $Y=1.16
+ $X2=0 $Y2=0
cc_434 N_A_783_297#_c_384_n N_A_375_49#_c_1142_n 2.0806e-19 $X=5.83 $Y=1.202
+ $X2=0 $Y2=0
cc_435 N_A_783_297#_c_385_n N_A_375_49#_c_1142_n 0.00243787f $X=5.62 $Y=0.995
+ $X2=0 $Y2=0
cc_436 N_A_783_297#_c_388_n N_A_375_49#_c_1142_n 0.015476f $X=5.785 $Y=0.85
+ $X2=0 $Y2=0
cc_437 N_A_783_297#_c_387_n N_A_1184_297#_M1016_d 0.00166227f $X=6.975 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_438 N_A_783_297#_c_395_n N_A_1184_297#_c_1268_n 0.00686704f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_439 N_A_783_297#_c_387_n N_A_1184_297#_c_1268_n 0.0181022f $X=6.975 $Y=0.85
+ $X2=0 $Y2=0
cc_440 N_A_783_297#_c_390_n N_A_1184_297#_c_1268_n 0.0020738f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_441 N_A_783_297#_c_391_n N_A_1184_297#_c_1268_n 0.00517339f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_783_297#_c_395_n N_A_1184_297#_c_1280_n 0.00431165f $X=5.83 $Y=1.41
+ $X2=0 $Y2=0
cc_443 N_A_783_297#_c_397_n N_A_1184_297#_c_1281_n 0.0165035f $X=7.32 $Y=1.57
+ $X2=0 $Y2=0
cc_444 N_A_783_297#_c_391_n N_A_1184_297#_c_1281_n 0.00161448f $X=7.12 $Y=0.85
+ $X2=0 $Y2=0
cc_445 N_A_783_297#_c_404_p N_VGND_c_1335_n 0.00371415f $X=4.305 $Y=0.85 $X2=0
+ $Y2=0
cc_446 N_A_783_297#_c_394_n N_VGND_c_1335_n 0.0242428f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_447 N_A_783_297#_M1016_g N_VGND_c_1340_n 0.00575161f $X=5.855 $Y=0.455 $X2=0
+ $Y2=0
cc_448 N_A_783_297#_c_389_n N_VGND_c_1340_n 0.00340751f $X=5.64 $Y=0.85 $X2=0
+ $Y2=0
cc_449 N_A_783_297#_c_391_n N_VGND_c_1340_n 0.00102193f $X=7.12 $Y=0.85 $X2=0
+ $Y2=0
cc_450 N_A_783_297#_c_393_n N_VGND_c_1340_n 0.00585385f $X=7.262 $Y=0.945 $X2=0
+ $Y2=0
cc_451 N_A_783_297#_c_394_n N_VGND_c_1340_n 0.0088551f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_452 N_A_783_297#_M1008_d N_VGND_c_1342_n 0.00198811f $X=4.145 $Y=0.235 $X2=0
+ $Y2=0
cc_453 N_A_783_297#_M1016_g N_VGND_c_1342_n 0.00668858f $X=5.855 $Y=0.455 $X2=0
+ $Y2=0
cc_454 N_A_783_297#_c_386_n N_VGND_c_1342_n 0.0112598f $X=5.495 $Y=0.85 $X2=0
+ $Y2=0
cc_455 N_A_783_297#_c_404_p N_VGND_c_1342_n 0.0148172f $X=4.305 $Y=0.85 $X2=0
+ $Y2=0
cc_456 N_A_783_297#_c_393_n N_VGND_c_1342_n 0.00635691f $X=7.262 $Y=0.945 $X2=0
+ $Y2=0
cc_457 N_A_783_297#_c_394_n N_VGND_c_1342_n 0.00448669f $X=4.28 $Y=0.74 $X2=0
+ $Y2=0
cc_458 N_B_c_567_n A 0.0014495f $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_459 N_B_c_570_n N_A_901_297#_c_738_n 0.003607f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_460 N_B_M1008_g N_A_901_297#_c_738_n 0.00120589f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_461 N_B_c_563_n N_A_901_297#_c_738_n 0.014573f $X=4.925 $Y=1.16 $X2=0 $Y2=0
cc_462 N_B_M1010_g N_A_901_297#_c_738_n 0.00424996f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_463 N_B_M1006_g N_A_901_297#_c_738_n 0.0035466f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_464 N_B_c_566_n N_A_901_297#_c_738_n 0.0011146f $X=5.025 $Y=1.16 $X2=0 $Y2=0
cc_465 B N_A_901_297#_c_746_n 0.008575f $X=7.035 $Y=1.445 $X2=0 $Y2=0
cc_466 N_B_M1006_g N_A_901_297#_c_758_n 0.00201366f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_467 N_B_c_569_n N_A_901_297#_c_758_n 0.0032563f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_468 N_B_M1008_g N_A_901_297#_c_742_n 4.212e-19 $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_469 N_B_M1006_g N_A_901_297#_c_742_n 9.17075e-19 $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_470 N_B_M1008_g N_A_901_297#_c_743_n 0.00491597f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_471 N_B_c_563_n N_A_901_297#_c_743_n 0.00309496f $X=4.925 $Y=1.16 $X2=0 $Y2=0
cc_472 N_B_c_570_n N_VPWR_c_889_n 0.0113699f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_473 N_B_c_570_n N_VPWR_c_887_n 0.00656627f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_474 N_B_c_573_n N_VPWR_c_887_n 0.0412005f $X=6.655 $Y=2.54 $X2=0 $Y2=0
cc_475 N_B_c_574_n N_VPWR_c_887_n 0.0071208f $X=5.125 $Y=2.54 $X2=0 $Y2=0
cc_476 N_B_c_570_n N_VPWR_c_896_n 0.00455828f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_477 N_B_c_574_n N_VPWR_c_896_n 0.0407088f $X=5.125 $Y=2.54 $X2=0 $Y2=0
cc_478 N_B_M1008_g N_A_351_325#_c_980_n 0.00316063f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_479 N_B_c_570_n N_A_351_325#_c_981_n 0.0127882f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_480 N_B_c_564_n N_A_351_325#_c_981_n 0.00535881f $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_481 N_B_c_570_n N_A_351_325#_c_987_n 0.0175458f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_482 N_B_c_570_n N_A_351_325#_c_988_n 0.00608631f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_483 N_B_M1010_g N_A_351_325#_c_988_n 8.94333e-19 $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_484 N_B_c_570_n N_A_351_325#_c_990_n 0.00366198f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_485 N_B_c_563_n N_A_351_325#_c_982_n 0.00354518f $X=4.925 $Y=1.16 $X2=0 $Y2=0
cc_486 N_B_M1010_g N_A_351_325#_c_982_n 0.0315935f $X=5.025 $Y=1.905 $X2=0 $Y2=0
cc_487 N_B_M1006_g N_A_351_325#_c_982_n 0.00651676f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_488 N_B_c_566_n N_A_351_325#_c_982_n 0.0105369f $X=5.025 $Y=1.16 $X2=0 $Y2=0
cc_489 N_B_M1010_g N_A_351_325#_c_992_n 0.00817171f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_490 N_B_c_573_n N_A_351_325#_c_992_n 0.0364604f $X=6.655 $Y=2.54 $X2=0 $Y2=0
cc_491 N_B_c_574_n N_A_351_325#_c_992_n 2.38151e-19 $X=5.125 $Y=2.54 $X2=0 $Y2=0
cc_492 N_B_M1011_g N_A_351_325#_c_992_n 0.0102069f $X=6.755 $Y=1.965 $X2=0 $Y2=0
cc_493 N_B_M1006_g N_A_351_325#_c_1028_n 5.73691e-19 $X=5.05 $Y=0.565 $X2=0
+ $Y2=0
cc_494 N_B_M1008_g N_A_351_325#_c_983_n 8.48623e-19 $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_495 N_B_c_564_n N_A_351_325#_c_983_n 0.0038653f $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_496 N_B_M1006_g N_A_351_325#_c_984_n 0.0136729f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_497 N_B_M1010_g N_A_351_325#_c_994_n 0.00716396f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_498 N_B_c_574_n N_A_351_325#_c_994_n 2.51585e-19 $X=5.125 $Y=2.54 $X2=0 $Y2=0
cc_499 N_B_c_564_n N_A_375_49#_c_1132_n 4.44674e-19 $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_500 N_B_M1010_g N_A_375_49#_c_1136_n 0.00145677f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_501 N_B_M1010_g N_A_375_49#_c_1173_n 0.00446449f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_502 N_B_c_569_n N_A_375_49#_c_1133_n 0.0026019f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_503 N_B_c_567_n N_A_375_49#_c_1186_n 0.0029291f $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_504 N_B_c_568_n N_A_375_49#_c_1186_n 4.30216e-19 $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_505 N_B_c_569_n N_A_375_49#_c_1186_n 0.00498906f $X=6.735 $Y=0.995 $X2=0
+ $Y2=0
cc_506 N_B_c_568_n N_A_375_49#_c_1187_n 0.00110831f $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_507 N_B_c_569_n N_A_375_49#_c_1208_n 0.00521263f $X=6.735 $Y=0.995 $X2=0
+ $Y2=0
cc_508 N_B_c_570_n N_A_375_49#_c_1139_n 0.00469456f $X=3.825 $Y=1.41 $X2=0 $Y2=0
cc_509 N_B_c_563_n N_A_375_49#_c_1139_n 0.00486395f $X=4.925 $Y=1.16 $X2=0 $Y2=0
cc_510 N_B_c_564_n N_A_375_49#_c_1139_n 2.58451e-19 $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_511 N_B_M1010_g N_A_375_49#_c_1139_n 0.00481446f $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_512 N_B_c_566_n N_A_375_49#_c_1139_n 2.29578e-19 $X=5.025 $Y=1.16 $X2=0 $Y2=0
cc_513 N_B_M1010_g N_A_375_49#_c_1142_n 4.48588e-19 $X=5.025 $Y=1.905 $X2=0
+ $Y2=0
cc_514 N_B_c_575_n N_A_1184_297#_c_1268_n 0.00160527f $X=6.755 $Y=1.47 $X2=0
+ $Y2=0
cc_515 N_B_M1011_g N_A_1184_297#_c_1268_n 0.00912353f $X=6.755 $Y=1.965 $X2=0
+ $Y2=0
cc_516 N_B_c_579_n N_A_1184_297#_c_1268_n 0.0142666f $X=6.735 $Y=1.445 $X2=0
+ $Y2=0
cc_517 N_B_c_567_n N_A_1184_297#_c_1268_n 0.0332296f $X=6.71 $Y=1.16 $X2=0 $Y2=0
cc_518 N_B_c_569_n N_A_1184_297#_c_1268_n 0.0105486f $X=6.735 $Y=0.995 $X2=0
+ $Y2=0
cc_519 N_B_M1011_g N_A_1184_297#_c_1281_n 0.011211f $X=6.755 $Y=1.965 $X2=0
+ $Y2=0
cc_520 N_B_c_579_n N_A_1184_297#_c_1281_n 0.00934779f $X=6.735 $Y=1.445 $X2=0
+ $Y2=0
cc_521 N_B_c_568_n N_A_1184_297#_c_1281_n 0.00114355f $X=6.71 $Y=1.16 $X2=0
+ $Y2=0
cc_522 B N_A_1184_297#_c_1281_n 0.0165342f $X=7.035 $Y=1.445 $X2=0 $Y2=0
cc_523 N_B_M1008_g N_VGND_c_1335_n 0.0190364f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_524 N_B_c_564_n N_VGND_c_1335_n 0.00541821f $X=4.145 $Y=1.16 $X2=0 $Y2=0
cc_525 N_B_M1008_g N_VGND_c_1340_n 0.00494995f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_526 N_B_M1006_g N_VGND_c_1340_n 0.00427876f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_527 N_B_c_569_n N_VGND_c_1340_n 0.00357877f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_528 N_B_M1008_g N_VGND_c_1342_n 0.00918586f $X=4.07 $Y=0.56 $X2=0 $Y2=0
cc_529 N_B_M1006_g N_VGND_c_1342_n 0.00718354f $X=5.05 $Y=0.565 $X2=0 $Y2=0
cc_530 N_B_c_569_n N_VGND_c_1342_n 0.00612424f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_531 N_A_c_698_n N_A_901_297#_c_736_n 0.0280559f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_532 A N_A_901_297#_c_736_n 0.00120954f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_533 N_A_c_699_n N_A_901_297#_c_737_n 0.0127509f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_534 N_A_c_698_n N_A_901_297#_c_746_n 0.0159729f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_535 A N_A_901_297#_c_746_n 0.0496316f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_536 N_A_c_698_n N_A_901_297#_c_739_n 5.76324e-19 $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_537 N_A_c_699_n N_A_901_297#_c_739_n 0.0126125f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_538 A N_A_901_297#_c_739_n 0.0305287f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_539 N_A_c_698_n N_A_901_297#_c_740_n 0.00444032f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_540 A N_A_901_297#_c_740_n 0.0219245f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_541 N_A_c_698_n N_A_901_297#_c_741_n 6.50193e-19 $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_542 N_A_c_699_n N_A_901_297#_c_741_n 0.00282528f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_543 A N_A_901_297#_c_741_n 0.0156105f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_544 N_A_c_698_n N_A_901_297#_c_748_n 0.0026346f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_545 A N_A_901_297#_c_771_n 0.00189901f $X=7.96 $Y=1.105 $X2=0 $Y2=0
cc_546 N_A_c_698_n N_VPWR_c_887_n 0.00449112f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_547 N_A_c_698_n N_VPWR_c_896_n 0.00365142f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_548 N_A_c_698_n N_VPWR_c_897_n 0.0154641f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_549 N_A_c_698_n N_A_351_325#_c_992_n 0.00151171f $X=7.875 $Y=1.41 $X2=0 $Y2=0
cc_550 N_A_c_698_n N_A_1184_297#_c_1281_n 0.0150455f $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_551 N_A_c_698_n N_A_1184_297#_c_1274_n 2.97458e-19 $X=7.875 $Y=1.41 $X2=0
+ $Y2=0
cc_552 N_A_c_699_n N_VGND_c_1336_n 0.00853835f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_553 N_A_c_699_n N_VGND_c_1340_n 0.00439206f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_554 N_A_c_699_n N_VGND_c_1342_n 0.00711209f $X=7.9 $Y=0.995 $X2=0 $Y2=0
cc_555 N_A_901_297#_c_746_n N_VPWR_M1014_d 0.0158767f $X=8.49 $Y=1.6 $X2=0 $Y2=0
cc_556 N_A_901_297#_c_736_n N_VPWR_c_892_n 0.00435494f $X=8.66 $Y=1.41 $X2=0
+ $Y2=0
cc_557 N_A_901_297#_M1005_d N_VPWR_c_887_n 0.00402227f $X=7.41 $Y=1.645 $X2=0
+ $Y2=0
cc_558 N_A_901_297#_c_736_n N_VPWR_c_887_n 0.00588068f $X=8.66 $Y=1.41 $X2=0
+ $Y2=0
cc_559 N_A_901_297#_c_736_n N_VPWR_c_897_n 0.0135348f $X=8.66 $Y=1.41 $X2=0
+ $Y2=0
cc_560 N_A_901_297#_c_758_n N_A_351_325#_M1006_d 0.00599198f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_561 N_A_901_297#_c_738_n N_A_351_325#_c_987_n 0.0132911f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_562 N_A_901_297#_c_738_n N_A_351_325#_c_988_n 0.00274773f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_563 N_A_901_297#_M1010_s N_A_351_325#_c_989_n 0.0102858f $X=4.505 $Y=1.485
+ $X2=0 $Y2=0
cc_564 N_A_901_297#_c_738_n N_A_351_325#_c_989_n 0.0128549f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_565 N_A_901_297#_c_738_n N_A_351_325#_c_982_n 0.0675972f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_566 N_A_901_297#_M1005_d N_A_351_325#_c_992_n 0.00265748f $X=7.41 $Y=1.645
+ $X2=0 $Y2=0
cc_567 N_A_901_297#_c_758_n N_A_351_325#_c_1028_n 0.0125715f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_568 N_A_901_297#_c_742_n N_A_351_325#_c_1028_n 0.0014251f $X=4.815 $Y=0.51
+ $X2=0 $Y2=0
cc_569 N_A_901_297#_c_743_n N_A_351_325#_c_1028_n 0.00331722f $X=4.67 $Y=0.51
+ $X2=0 $Y2=0
cc_570 N_A_901_297#_M1006_s N_A_351_325#_c_984_n 0.00152093f $X=4.665 $Y=0.245
+ $X2=0 $Y2=0
cc_571 N_A_901_297#_c_738_n N_A_351_325#_c_984_n 0.0123119f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_572 N_A_901_297#_c_758_n N_A_351_325#_c_984_n 0.00366657f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_573 N_A_901_297#_c_743_n N_A_351_325#_c_984_n 0.00172491f $X=4.67 $Y=0.51
+ $X2=0 $Y2=0
cc_574 N_A_901_297#_c_758_n N_A_375_49#_M1019_d 0.00419658f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_575 N_A_901_297#_c_758_n N_A_375_49#_c_1133_n 0.0147234f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_576 N_A_901_297#_c_758_n N_A_375_49#_c_1186_n 0.00610486f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_577 N_A_901_297#_c_758_n N_A_375_49#_c_1187_n 0.00980954f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_578 N_A_901_297#_c_771_n N_A_375_49#_c_1187_n 0.0012274f $X=7.63 $Y=0.51
+ $X2=0 $Y2=0
cc_579 N_A_901_297#_c_772_n N_A_375_49#_c_1187_n 0.00676871f $X=7.63 $Y=0.51
+ $X2=0 $Y2=0
cc_580 N_A_901_297#_c_758_n N_A_375_49#_c_1208_n 0.0119237f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_581 N_A_901_297#_M1010_s N_A_375_49#_c_1139_n 0.00802537f $X=4.505 $Y=1.485
+ $X2=0 $Y2=0
cc_582 N_A_901_297#_c_738_n N_A_375_49#_c_1139_n 0.0183124f $X=4.63 $Y=1.94
+ $X2=0 $Y2=0
cc_583 N_A_901_297#_c_758_n N_A_1184_297#_M1016_d 0.00653094f $X=7.485 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_584 N_A_901_297#_c_758_n N_A_1184_297#_c_1268_n 0.00162336f $X=7.485 $Y=0.51
+ $X2=0 $Y2=0
cc_585 N_A_901_297#_c_736_n N_A_1184_297#_c_1269_n 0.0195627f $X=8.66 $Y=1.41
+ $X2=0 $Y2=0
cc_586 N_A_901_297#_c_737_n N_A_1184_297#_c_1269_n 0.0097849f $X=8.685 $Y=0.995
+ $X2=0 $Y2=0
cc_587 N_A_901_297#_c_746_n N_A_1184_297#_c_1269_n 0.0112214f $X=8.49 $Y=1.6
+ $X2=0 $Y2=0
cc_588 N_A_901_297#_c_741_n N_A_1184_297#_c_1269_n 0.0381742f $X=8.575 $Y=1.325
+ $X2=0 $Y2=0
cc_589 N_A_901_297#_c_748_n N_A_1184_297#_c_1269_n 0.00830381f $X=8.575 $Y=1.495
+ $X2=0 $Y2=0
cc_590 N_A_901_297#_M1005_d N_A_1184_297#_c_1281_n 0.00774465f $X=7.41 $Y=1.645
+ $X2=0 $Y2=0
cc_591 N_A_901_297#_c_736_n N_A_1184_297#_c_1281_n 0.00346175f $X=8.66 $Y=1.41
+ $X2=0 $Y2=0
cc_592 N_A_901_297#_c_746_n N_A_1184_297#_c_1281_n 0.0539817f $X=8.49 $Y=1.6
+ $X2=0 $Y2=0
cc_593 N_A_901_297#_c_736_n N_A_1184_297#_c_1274_n 0.0129225f $X=8.66 $Y=1.41
+ $X2=0 $Y2=0
cc_594 N_A_901_297#_c_746_n N_A_1184_297#_c_1274_n 0.00653478f $X=8.49 $Y=1.6
+ $X2=0 $Y2=0
cc_595 N_A_901_297#_c_741_n N_A_1184_297#_c_1274_n 0.00278512f $X=8.575 $Y=1.325
+ $X2=0 $Y2=0
cc_596 N_A_901_297#_c_736_n N_A_1184_297#_c_1270_n 2.03932e-19 $X=8.66 $Y=1.41
+ $X2=0 $Y2=0
cc_597 N_A_901_297#_c_739_n N_VGND_M1009_d 0.00664804f $X=8.49 $Y=0.82 $X2=0
+ $Y2=0
cc_598 N_A_901_297#_c_741_n N_VGND_M1009_d 0.00108061f $X=8.575 $Y=1.325 $X2=0
+ $Y2=0
cc_599 N_A_901_297#_c_737_n N_VGND_c_1336_n 0.00767602f $X=8.685 $Y=0.995 $X2=0
+ $Y2=0
cc_600 N_A_901_297#_c_739_n N_VGND_c_1336_n 0.0344146f $X=8.49 $Y=0.82 $X2=0
+ $Y2=0
cc_601 N_A_901_297#_c_741_n N_VGND_c_1336_n 0.00164729f $X=8.575 $Y=1.325 $X2=0
+ $Y2=0
cc_602 N_A_901_297#_c_771_n N_VGND_c_1336_n 0.00124421f $X=7.63 $Y=0.51 $X2=0
+ $Y2=0
cc_603 N_A_901_297#_c_739_n N_VGND_c_1340_n 0.0027904f $X=8.49 $Y=0.82 $X2=0
+ $Y2=0
cc_604 N_A_901_297#_c_758_n N_VGND_c_1340_n 0.00574592f $X=7.485 $Y=0.51 $X2=0
+ $Y2=0
cc_605 N_A_901_297#_c_742_n N_VGND_c_1340_n 2.9688e-19 $X=4.815 $Y=0.51 $X2=0
+ $Y2=0
cc_606 N_A_901_297#_c_743_n N_VGND_c_1340_n 0.0250994f $X=4.67 $Y=0.51 $X2=0
+ $Y2=0
cc_607 N_A_901_297#_c_771_n N_VGND_c_1340_n 3.63685e-19 $X=7.63 $Y=0.51 $X2=0
+ $Y2=0
cc_608 N_A_901_297#_c_772_n N_VGND_c_1340_n 0.0149689f $X=7.63 $Y=0.51 $X2=0
+ $Y2=0
cc_609 N_A_901_297#_c_737_n N_VGND_c_1341_n 0.00536613f $X=8.685 $Y=0.995 $X2=0
+ $Y2=0
cc_610 N_A_901_297#_c_741_n N_VGND_c_1341_n 0.00182428f $X=8.575 $Y=1.325 $X2=0
+ $Y2=0
cc_611 N_A_901_297#_M1001_d N_VGND_c_1342_n 0.00244776f $X=7.42 $Y=0.235 $X2=0
+ $Y2=0
cc_612 N_A_901_297#_c_737_n N_VGND_c_1342_n 0.0108802f $X=8.685 $Y=0.995 $X2=0
+ $Y2=0
cc_613 N_A_901_297#_c_739_n N_VGND_c_1342_n 0.00734124f $X=8.49 $Y=0.82 $X2=0
+ $Y2=0
cc_614 N_A_901_297#_c_741_n N_VGND_c_1342_n 0.00405875f $X=8.575 $Y=1.325 $X2=0
+ $Y2=0
cc_615 N_A_901_297#_c_758_n N_VGND_c_1342_n 0.232931f $X=7.485 $Y=0.51 $X2=0
+ $Y2=0
cc_616 N_A_901_297#_c_742_n N_VGND_c_1342_n 0.028616f $X=4.815 $Y=0.51 $X2=0
+ $Y2=0
cc_617 N_A_901_297#_c_743_n N_VGND_c_1342_n 0.00392171f $X=4.67 $Y=0.51 $X2=0
+ $Y2=0
cc_618 N_A_901_297#_c_771_n N_VGND_c_1342_n 0.0285254f $X=7.63 $Y=0.51 $X2=0
+ $Y2=0
cc_619 N_A_901_297#_c_772_n N_VGND_c_1342_n 0.0036194f $X=7.63 $Y=0.51 $X2=0
+ $Y2=0
cc_620 N_X_c_869_n N_VPWR_c_888_n 0.0193871f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_621 N_X_c_869_n N_VPWR_c_890_n 0.0196165f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_622 N_X_M1000_s N_VPWR_c_887_n 0.00442207f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_623 N_X_c_869_n N_VPWR_c_887_n 0.0107063f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_624 N_X_c_866_n N_VGND_c_1334_n 0.0132437f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_625 N_X_c_866_n N_VGND_c_1339_n 0.0112745f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_626 N_X_M1012_s N_VGND_c_1342_n 0.00480511f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_627 N_X_c_866_n N_VGND_c_1342_n 0.00944103f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_628 N_VPWR_c_887_n N_A_351_325#_M1011_d 0.00241089f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_629 N_VPWR_c_889_n N_A_351_325#_c_985_n 0.00147971f $X=3.59 $Y=2.32 $X2=0
+ $Y2=0
cc_630 N_VPWR_c_891_n N_A_351_325#_c_985_n 0.012236f $X=3.425 $Y=2.72 $X2=0
+ $Y2=0
cc_631 N_VPWR_c_887_n N_A_351_325#_c_985_n 0.0223233f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_632 N_VPWR_M1004_s N_A_351_325#_c_981_n 0.00648603f $X=3.465 $Y=2.175 $X2=0
+ $Y2=0
cc_633 N_VPWR_M1004_s N_A_351_325#_c_987_n 0.00155527f $X=3.465 $Y=2.175 $X2=0
+ $Y2=0
cc_634 N_VPWR_c_889_n N_A_351_325#_c_987_n 0.00612755f $X=3.59 $Y=2.32 $X2=0
+ $Y2=0
cc_635 N_VPWR_c_887_n N_A_351_325#_c_987_n 0.0119497f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_636 N_VPWR_c_896_n N_A_351_325#_c_987_n 0.00666556f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_637 N_VPWR_c_889_n N_A_351_325#_c_988_n 0.00140976f $X=3.59 $Y=2.32 $X2=0
+ $Y2=0
cc_638 N_VPWR_c_887_n N_A_351_325#_c_989_n 0.0193106f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_639 N_VPWR_c_896_n N_A_351_325#_c_989_n 0.0300226f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_640 N_VPWR_c_889_n N_A_351_325#_c_990_n 0.00679194f $X=3.59 $Y=2.32 $X2=0
+ $Y2=0
cc_641 N_VPWR_c_887_n N_A_351_325#_c_990_n 0.00644598f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_642 N_VPWR_c_896_n N_A_351_325#_c_990_n 0.0105925f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_643 N_VPWR_c_887_n N_A_351_325#_c_992_n 0.0811181f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_644 N_VPWR_c_896_n N_A_351_325#_c_992_n 0.134682f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_645 N_VPWR_c_897_n N_A_351_325#_c_992_n 0.00713809f $X=8.595 $Y=2.54 $X2=0
+ $Y2=0
cc_646 N_VPWR_M1004_s N_A_351_325#_c_993_n 0.00233831f $X=3.465 $Y=2.175 $X2=0
+ $Y2=0
cc_647 N_VPWR_c_889_n N_A_351_325#_c_993_n 0.0144069f $X=3.59 $Y=2.32 $X2=0
+ $Y2=0
cc_648 N_VPWR_c_887_n N_A_351_325#_c_993_n 8.22076e-19 $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_649 N_VPWR_c_887_n N_A_351_325#_c_994_n 0.00587789f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_650 N_VPWR_c_896_n N_A_351_325#_c_994_n 0.0103509f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_651 N_VPWR_M1004_s N_A_375_49#_c_1139_n 0.00109947f $X=3.465 $Y=2.175 $X2=0
+ $Y2=0
cc_652 N_VPWR_c_887_n N_A_1184_297#_M1007_d 0.00259864f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_653 N_VPWR_c_892_n N_A_1184_297#_c_1272_n 0.0197624f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_654 N_VPWR_c_887_n N_A_1184_297#_c_1272_n 0.0111058f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_897_n N_A_1184_297#_c_1272_n 0.0126514f $X=8.595 $Y=2.54 $X2=0
+ $Y2=0
cc_656 N_VPWR_M1014_d N_A_1184_297#_c_1281_n 0.01324f $X=7.965 $Y=1.485 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_887_n N_A_1184_297#_c_1281_n 0.0167691f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_896_n N_A_1184_297#_c_1281_n 0.00725506f $X=7.915 $Y=2.54 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_897_n N_A_1184_297#_c_1281_n 0.0423107f $X=8.595 $Y=2.54 $X2=0
+ $Y2=0
cc_660 N_VPWR_c_892_n N_A_1184_297#_c_1274_n 0.0034505f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_887_n N_A_1184_297#_c_1274_n 0.00562459f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_662 N_A_351_325#_c_985_n N_A_375_49#_M1021_d 0.012215f $X=3.445 $Y=1.98 $X2=0
+ $Y2=0
cc_663 N_A_351_325#_c_992_n N_A_375_49#_M1010_d 0.00924946f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_664 N_A_351_325#_M1013_d N_A_375_49#_c_1144_n 0.0100433f $X=2.835 $Y=0.245
+ $X2=0 $Y2=0
cc_665 N_A_351_325#_c_979_n N_A_375_49#_c_1144_n 0.0200889f $X=3.335 $Y=0.37
+ $X2=0 $Y2=0
cc_666 N_A_351_325#_c_980_n N_A_375_49#_c_1144_n 0.0140571f $X=3.42 $Y=1.035
+ $X2=0 $Y2=0
cc_667 N_A_351_325#_M1013_d N_A_375_49#_c_1132_n 0.00270797f $X=2.835 $Y=0.245
+ $X2=0 $Y2=0
cc_668 N_A_351_325#_c_980_n N_A_375_49#_c_1132_n 0.0179157f $X=3.42 $Y=1.035
+ $X2=0 $Y2=0
cc_669 N_A_351_325#_c_981_n N_A_375_49#_c_1132_n 0.00902524f $X=3.53 $Y=1.895
+ $X2=0 $Y2=0
cc_670 N_A_351_325#_c_983_n N_A_375_49#_c_1132_n 0.0132103f $X=3.53 $Y=1.12
+ $X2=0 $Y2=0
cc_671 N_A_351_325#_c_982_n N_A_375_49#_c_1136_n 0.00870819f $X=4.97 $Y=2.275
+ $X2=0 $Y2=0
cc_672 N_A_351_325#_c_984_n N_A_375_49#_c_1136_n 2.53366e-19 $X=4.97 $Y=0.772
+ $X2=0 $Y2=0
cc_673 N_A_351_325#_c_982_n N_A_375_49#_c_1173_n 0.0255541f $X=4.97 $Y=2.275
+ $X2=0 $Y2=0
cc_674 N_A_351_325#_c_992_n N_A_375_49#_c_1173_n 0.0238103f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_675 N_A_351_325#_c_992_n N_A_375_49#_c_1137_n 0.0100462f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_676 N_A_351_325#_c_1028_n N_A_375_49#_c_1133_n 0.00253431f $X=5.26 $Y=0.545
+ $X2=0 $Y2=0
cc_677 N_A_351_325#_c_985_n N_A_375_49#_c_1139_n 0.00437461f $X=3.445 $Y=1.98
+ $X2=0 $Y2=0
cc_678 N_A_351_325#_c_981_n N_A_375_49#_c_1139_n 0.0161183f $X=3.53 $Y=1.895
+ $X2=0 $Y2=0
cc_679 N_A_351_325#_c_987_n N_A_375_49#_c_1139_n 0.01149f $X=4.19 $Y=1.98 $X2=0
+ $Y2=0
cc_680 N_A_351_325#_c_982_n N_A_375_49#_c_1139_n 0.0194408f $X=4.97 $Y=2.275
+ $X2=0 $Y2=0
cc_681 N_A_351_325#_c_983_n N_A_375_49#_c_1139_n 0.0052436f $X=3.53 $Y=1.12
+ $X2=0 $Y2=0
cc_682 N_A_351_325#_c_984_n N_A_375_49#_c_1139_n 8.86472e-19 $X=4.97 $Y=0.772
+ $X2=0 $Y2=0
cc_683 N_A_351_325#_c_985_n N_A_375_49#_c_1140_n 0.00415423f $X=3.445 $Y=1.98
+ $X2=0 $Y2=0
cc_684 N_A_351_325#_c_981_n N_A_375_49#_c_1140_n 0.00275249f $X=3.53 $Y=1.895
+ $X2=0 $Y2=0
cc_685 N_A_351_325#_c_985_n N_A_375_49#_c_1141_n 0.0251846f $X=3.445 $Y=1.98
+ $X2=0 $Y2=0
cc_686 N_A_351_325#_c_981_n N_A_375_49#_c_1141_n 0.0231767f $X=3.53 $Y=1.895
+ $X2=0 $Y2=0
cc_687 N_A_351_325#_c_982_n N_A_375_49#_c_1142_n 0.00127808f $X=4.97 $Y=2.275
+ $X2=0 $Y2=0
cc_688 N_A_351_325#_c_992_n N_A_1184_297#_M1018_d 0.00563686f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_689 N_A_351_325#_c_992_n N_A_1184_297#_c_1280_n 0.0129278f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_690 N_A_351_325#_M1011_d N_A_1184_297#_c_1281_n 0.00678674f $X=6.845 $Y=1.645
+ $X2=0 $Y2=0
cc_691 N_A_351_325#_c_992_n N_A_1184_297#_c_1281_n 0.0533312f $X=7.075 $Y=2.36
+ $X2=0 $Y2=0
cc_692 N_A_351_325#_c_979_n N_VGND_c_1335_n 0.0140424f $X=3.335 $Y=0.37 $X2=0
+ $Y2=0
cc_693 N_A_351_325#_c_980_n N_VGND_c_1335_n 0.0299545f $X=3.42 $Y=1.035 $X2=0
+ $Y2=0
cc_694 N_A_351_325#_c_979_n N_VGND_c_1337_n 0.0344776f $X=3.335 $Y=0.37 $X2=0
+ $Y2=0
cc_695 N_A_351_325#_c_1028_n N_VGND_c_1340_n 0.00800682f $X=5.26 $Y=0.545 $X2=0
+ $Y2=0
cc_696 N_A_351_325#_c_984_n N_VGND_c_1340_n 0.00283956f $X=4.97 $Y=0.772 $X2=0
+ $Y2=0
cc_697 N_A_351_325#_c_979_n N_VGND_c_1342_n 0.0232692f $X=3.335 $Y=0.37 $X2=0
+ $Y2=0
cc_698 N_A_351_325#_c_1028_n N_VGND_c_1342_n 0.0018012f $X=5.26 $Y=0.545 $X2=0
+ $Y2=0
cc_699 N_A_375_49#_c_1133_n N_A_1184_297#_M1016_d 0.00729398f $X=6.03 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_700 N_A_375_49#_c_1252_p N_A_1184_297#_M1016_d 0.0024562f $X=6.115 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_701 N_A_375_49#_c_1208_n N_A_1184_297#_M1016_d 0.0107136f $X=6.625 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_702 N_A_375_49#_c_1137_n N_A_1184_297#_M1018_d 0.00444096f $X=5.945 $Y=1.53
+ $X2=0 $Y2=0
cc_703 N_A_375_49#_c_1173_n N_A_1184_297#_c_1268_n 0.00453141f $X=5.46 $Y=1.62
+ $X2=0 $Y2=0
cc_704 N_A_375_49#_c_1137_n N_A_1184_297#_c_1268_n 0.013519f $X=5.945 $Y=1.53
+ $X2=0 $Y2=0
cc_705 N_A_375_49#_c_1133_n N_A_1184_297#_c_1268_n 0.062318f $X=6.03 $Y=1.445
+ $X2=0 $Y2=0
cc_706 N_A_375_49#_c_1208_n N_A_1184_297#_c_1268_n 0.0106102f $X=6.625 $Y=0.36
+ $X2=0 $Y2=0
cc_707 N_A_375_49#_c_1142_n N_A_1184_297#_c_1268_n 0.00130235f $X=5.64 $Y=1.53
+ $X2=0 $Y2=0
cc_708 N_A_375_49#_c_1139_n N_VGND_c_1335_n 0.00557009f $X=5.495 $Y=1.53 $X2=0
+ $Y2=0
cc_709 N_A_375_49#_c_1144_n N_VGND_c_1337_n 0.00321579f $X=2.995 $Y=0.71 $X2=0
+ $Y2=0
cc_710 N_A_375_49#_c_1252_p N_VGND_c_1340_n 0.0104913f $X=6.115 $Y=0.34 $X2=0
+ $Y2=0
cc_711 N_A_375_49#_c_1208_n N_VGND_c_1340_n 0.0617902f $X=6.625 $Y=0.36 $X2=0
+ $Y2=0
cc_712 N_A_375_49#_M1019_d N_VGND_c_1342_n 0.00226821f $X=6.725 $Y=0.245 $X2=0
+ $Y2=0
cc_713 N_A_375_49#_c_1252_p N_VGND_c_1342_n 0.00184693f $X=6.115 $Y=0.34 $X2=0
+ $Y2=0
cc_714 N_A_375_49#_c_1134_n N_VGND_c_1342_n 0.00750432f $X=2.225 $Y=0.765 $X2=0
+ $Y2=0
cc_715 N_A_375_49#_c_1208_n N_VGND_c_1342_n 0.00974346f $X=6.625 $Y=0.36 $X2=0
+ $Y2=0
cc_716 N_A_1184_297#_c_1270_n N_VGND_c_1341_n 0.0197576f $X=9.025 $Y=0.42 $X2=0
+ $Y2=0
cc_717 N_A_1184_297#_M1003_d N_VGND_c_1342_n 0.00399944f $X=8.76 $Y=0.235 $X2=0
+ $Y2=0
cc_718 N_A_1184_297#_c_1270_n N_VGND_c_1342_n 0.0113402f $X=9.025 $Y=0.42 $X2=0
+ $Y2=0
