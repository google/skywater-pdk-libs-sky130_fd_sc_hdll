# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dfstp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dfstp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.247200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.870000 1.005000 2.330000 1.625000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.540000 1.495000 10.485000 1.615000 ;
        RECT 9.540000 1.615000 10.015000 2.460000 ;
        RECT 9.685000 0.265000 10.015000 0.745000 ;
        RECT 9.685000 0.745000 10.485000 0.825000 ;
        RECT 9.750000 0.825000 10.485000 1.495000 ;
    END
  END Q
  PIN SET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 4.220000 0.735000 4.510000 0.780000 ;
        RECT 4.220000 0.780000 7.735000 0.920000 ;
        RECT 4.220000 0.920000 4.510000 0.965000 ;
        RECT 7.445000 0.735000 7.735000 0.780000 ;
        RECT 7.445000 0.920000 7.735000 0.965000 ;
    END
  END SET_B
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 10.580000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.555000  0.085000  1.885000 0.465000 ;
        RECT  3.910000  0.085000  4.370000 0.525000 ;
        RECT  5.140000  0.085000  5.530000 0.545000 ;
        RECT  7.320000  0.085000  8.030000 0.565000 ;
        RECT  9.070000  0.085000  9.450000 0.825000 ;
        RECT 10.185000  0.085000 10.450000 0.575000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 10.580000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.555000 2.135000  1.885000 2.635000 ;
        RECT  3.730000 2.255000  4.110000 2.635000 ;
        RECT  4.680000 2.255000  5.060000 2.635000 ;
        RECT  6.470000 2.255000  6.940000 2.635000 ;
        RECT  7.710000 1.945000  8.040000 2.635000 ;
        RECT  9.200000 1.495000  9.370000 2.635000 ;
        RECT 10.185000 1.785000 10.450000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.890000 0.805000 ;
      RECT 0.175000 1.795000 0.890000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.660000 0.805000 0.890000 1.795000 ;
      RECT 1.115000 0.345000 1.340000 2.465000 ;
      RECT 1.530000 0.635000 2.275000 0.825000 ;
      RECT 1.530000 0.825000 1.700000 1.795000 ;
      RECT 1.530000 1.795000 2.275000 1.965000 ;
      RECT 2.105000 0.305000 2.275000 0.635000 ;
      RECT 2.105000 1.965000 2.275000 2.465000 ;
      RECT 2.500000 0.705000 2.770000 1.575000 ;
      RECT 2.500000 1.575000 3.100000 1.955000 ;
      RECT 2.510000 2.250000 3.440000 2.420000 ;
      RECT 2.625000 0.265000 3.740000 0.465000 ;
      RECT 2.950000 0.645000 3.350000 1.015000 ;
      RECT 3.270000 1.230000 3.740000 1.235000 ;
      RECT 3.270000 1.235000 4.770000 1.405000 ;
      RECT 3.270000 1.405000 3.440000 2.250000 ;
      RECT 3.520000 0.465000 3.740000 1.230000 ;
      RECT 3.610000 1.575000 3.910000 1.835000 ;
      RECT 3.610000 1.835000 5.110000 2.085000 ;
      RECT 3.910000 0.735000 4.510000 1.065000 ;
      RECT 4.340000 2.085000 4.510000 2.375000 ;
      RECT 4.470000 1.405000 4.770000 1.565000 ;
      RECT 4.790000 0.295000 4.960000 0.725000 ;
      RECT 4.790000 0.725000 5.110000 1.065000 ;
      RECT 4.940000 1.065000 5.110000 1.835000 ;
      RECT 5.330000 0.725000 6.750000 0.895000 ;
      RECT 5.330000 0.895000 5.500000 1.655000 ;
      RECT 5.330000 1.655000 5.900000 1.965000 ;
      RECT 5.560000 2.165000 6.290000 2.415000 ;
      RECT 5.720000 1.065000 5.900000 1.475000 ;
      RECT 6.070000 1.235000 8.170000 1.405000 ;
      RECT 6.070000 1.405000 6.290000 1.915000 ;
      RECT 6.070000 1.915000 7.380000 2.085000 ;
      RECT 6.070000 2.085000 6.290000 2.165000 ;
      RECT 6.190000 0.305000 7.090000 0.475000 ;
      RECT 6.370000 0.895000 6.750000 1.015000 ;
      RECT 6.460000 1.575000 8.550000 1.745000 ;
      RECT 6.920000 0.475000 7.090000 1.235000 ;
      RECT 7.140000 2.085000 7.380000 2.375000 ;
      RECT 7.260000 0.735000 7.780000 1.005000 ;
      RECT 7.260000 1.005000 7.640000 1.065000 ;
      RECT 7.790000 1.175000 8.170000 1.235000 ;
      RECT 8.210000 0.350000 8.550000 0.680000 ;
      RECT 8.210000 1.745000 8.550000 1.765000 ;
      RECT 8.210000 1.765000 8.380000 2.375000 ;
      RECT 8.340000 0.680000 8.550000 1.575000 ;
      RECT 8.650000 1.915000 8.980000 2.425000 ;
      RECT 8.730000 0.345000 8.900000 0.995000 ;
      RECT 8.730000 0.995000 9.580000 1.325000 ;
      RECT 8.730000 1.325000 8.980000 1.915000 ;
    LAYER mcon ;
      RECT 0.665000 1.740000 0.835000 1.910000 ;
      RECT 1.165000 0.720000 1.335000 0.890000 ;
      RECT 2.645000 1.740000 2.815000 1.910000 ;
      RECT 3.155000 0.720000 3.325000 0.890000 ;
      RECT 4.280000 0.765000 4.450000 0.935000 ;
      RECT 5.705000 1.740000 5.875000 1.910000 ;
      RECT 5.725000 1.110000 5.895000 1.280000 ;
      RECT 7.505000 0.765000 7.675000 0.935000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 5.935000 1.940000 ;
      RECT 1.105000 0.690000 1.395000 0.780000 ;
      RECT 1.105000 0.780000 3.385000 0.920000 ;
      RECT 2.585000 1.710000 2.875000 1.800000 ;
      RECT 3.095000 0.690000 3.385000 0.780000 ;
      RECT 3.170000 0.920000 3.385000 1.120000 ;
      RECT 3.170000 1.120000 5.955000 1.260000 ;
      RECT 5.645000 1.710000 5.935000 1.800000 ;
      RECT 5.665000 1.080000 5.955000 1.120000 ;
      RECT 5.665000 1.260000 5.955000 1.310000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dfstp_2
