# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a22oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.675000 1.075000 6.285000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.510000 1.075000 8.535000 1.285000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.075000 4.440000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 2.095000 1.275000 ;
    END
  END B2
  PIN VGND
    ANTENNADIFFAREA  0.897000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.645000  0.085000 0.815000 0.555000 ;
        RECT 1.585000  0.085000 1.755000 0.555000 ;
        RECT 6.805000  0.085000 6.975000 0.555000 ;
        RECT 7.745000  0.085000 7.915000 0.555000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.160000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 4.885000 1.795000 5.135000 2.635000 ;
        RECT 5.825000 1.795000 6.075000 2.635000 ;
        RECT 6.765000 1.795000 7.015000 2.635000 ;
        RECT 7.705000 1.795000 7.955000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.024500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.645000 1.445000 3.675000 1.625000 ;
        RECT 0.645000 1.625000 0.855000 2.125000 ;
        RECT 1.545000 1.625000 1.795000 2.125000 ;
        RECT 2.395000 0.645000 6.115000 0.885000 ;
        RECT 2.395000 0.885000 2.695000 1.445000 ;
        RECT 2.485000 1.625000 2.735000 2.125000 ;
        RECT 3.425000 1.625000 3.675000 2.125000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.090000 1.455000 0.425000 2.295000 ;
      RECT 0.090000 2.295000 4.665000 2.465000 ;
      RECT 0.095000 0.255000 0.425000 0.725000 ;
      RECT 0.095000 0.725000 2.225000 0.905000 ;
      RECT 0.985000 0.255000 1.365000 0.725000 ;
      RECT 1.075000 1.795000 1.325000 2.295000 ;
      RECT 1.925000 0.255000 4.185000 0.475000 ;
      RECT 1.925000 0.475000 2.225000 0.725000 ;
      RECT 2.015000 1.795000 2.265000 2.295000 ;
      RECT 2.955000 1.795000 3.205000 2.295000 ;
      RECT 3.895000 1.455000 8.425000 1.625000 ;
      RECT 3.895000 1.625000 4.665000 2.295000 ;
      RECT 4.375000 0.255000 6.585000 0.475000 ;
      RECT 5.355000 1.625000 5.605000 2.465000 ;
      RECT 6.295000 1.625000 6.545000 2.465000 ;
      RECT 6.335000 0.475000 6.585000 0.725000 ;
      RECT 6.335000 0.725000 8.465000 0.905000 ;
      RECT 7.145000 0.255000 7.525000 0.725000 ;
      RECT 7.235000 1.625000 7.485000 2.465000 ;
      RECT 8.085000 0.255000 8.465000 0.725000 ;
      RECT 8.175000 1.625000 8.425000 2.465000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_4
