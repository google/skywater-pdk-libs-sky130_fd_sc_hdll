* NGSPICE file created from sky130_fd_sc_hdll__decap_12.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__decap_12 VGND VNB VPB VPWR
M1000 VPWR VGND VPWR VPB phighvt w=870000u l=4.73e+06u
+  ad=4.524e+11p pd=4.52e+06u as=0p ps=0u
M1001 VGND VPWR VGND VNB nshort w=550000u l=4.73e+06u
+  ad=2.86e+11p pd=3.24e+06u as=0p ps=0u
.ends

