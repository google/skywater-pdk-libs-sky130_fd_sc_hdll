* File: sky130_fd_sc_hdll__a211oi_1.pex.spice
* Created: Thu Aug 27 18:51:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%A2 1 3 4 6 7 8
r26 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.35
+ $Y=1.16 $X2=0.35 $Y2=1.16
r27 8 13 1.01686 $w=3.38e-07 $l=3e-08 $layer=LI1_cond $X=0.265 $Y=1.19 $X2=0.265
+ $Y2=1.16
r28 7 13 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.265 $Y=0.85
+ $X2=0.265 $Y2=1.16
r29 4 12 38.8967 $w=3.59e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.415 $Y2=1.16
r30 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r31 1 12 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.415 $Y2=1.16
r32 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%A1 1 3 4 6 7 8 9 10 18 27
r37 10 27 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.09 $Y=1.16 $X2=1.15
+ $Y2=1.16
r38 10 24 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=1.09 $Y=1.16
+ $X2=0.905 $Y2=1.16
r39 10 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.16 $X2=1.09 $Y2=1.16
r40 9 18 3.58108 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=1.16 $X2=0.755
+ $Y2=0.995
r41 9 24 3.25553 $w=3.3e-07 $l=1.5e-07 $layer=LI1_cond $X=0.755 $Y=1.16
+ $X2=0.905 $Y2=1.16
r42 8 18 5.57014 $w=2.98e-07 $l=1.45e-07 $layer=LI1_cond $X=0.755 $Y=0.85
+ $X2=0.755 $Y2=0.995
r43 7 8 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.755 $Y=0.51 $X2=0.755
+ $Y2=0.85
r44 4 16 47.8775 $w=2.99e-07 $l=2.79285e-07 $layer=POLY_cond $X=1 $Y=1.41
+ $X2=1.062 $Y2=1.16
r45 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.985
r46 1 16 38.5562 $w=2.99e-07 $l=2.03912e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=1.062 $Y2=1.16
r47 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%B1 1 3 4 6 7 8 9 10
r36 9 10 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=1.647 $Y=1.87
+ $X2=1.647 $Y2=2.21
r37 8 9 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=1.647 $Y=1.53
+ $X2=1.647 $Y2=1.87
r38 7 8 14.4544 $w=2.93e-07 $l=3.7e-07 $layer=LI1_cond $X=1.647 $Y=1.16
+ $X2=1.647 $Y2=1.53
r39 7 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.585
+ $Y=1.16 $X2=1.585 $Y2=1.16
r40 4 16 50.2707 $w=2.67e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.577 $Y2=1.16
r41 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.985
r42 1 16 38.9672 $w=2.67e-07 $l=1.95653e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.577 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995 $X2=1.51
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%C1 1 3 4 6 7 8
r25 7 8 14.9615 $w=2.83e-07 $l=3.7e-07 $layer=LI1_cond $X=2.122 $Y=1.16
+ $X2=2.122 $Y2=1.53
r26 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.065
+ $Y=1.16 $X2=2.065 $Y2=1.16
r27 4 12 47.4309 $w=3.07e-07 $l=2.81514e-07 $layer=POLY_cond $X=2.03 $Y=1.41
+ $X2=2.097 $Y2=1.16
r28 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.03 $Y=1.41 $X2=2.03
+ $Y2=1.985
r29 1 12 38.5336 $w=3.07e-07 $l=2.05925e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=2.097 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.005 $Y=0.995
+ $X2=2.005 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%A_27_297# 1 2 9 11 12 15
r21 13 15 7.49386 $w=1.83e-07 $l=1.25e-07 $layer=LI1_cond $X=1.237 $Y=1.725
+ $X2=1.237 $Y2=1.85
r22 11 13 6.82996 $w=2e-07 $l=1.38564e-07 $layer=LI1_cond $X=1.145 $Y=1.625
+ $X2=1.237 $Y2=1.725
r23 11 12 42.7 $w=1.98e-07 $l=7.7e-07 $layer=LI1_cond $X=1.145 $Y=1.625
+ $X2=0.375 $Y2=1.625
r24 7 12 6.92652 $w=2e-07 $l=1.67705e-07 $layer=LI1_cond $X=0.25 $Y=1.725
+ $X2=0.375 $Y2=1.625
r25 7 9 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.25 $Y=1.725
+ $X2=0.25 $Y2=1.85
r26 2 15 300 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.24 $Y2=1.85
r27 1 9 300 $w=1.7e-07 $l=4.31451e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%VPWR 1 6 8 10 20 21 24
r31 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r32 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 18 21 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r35 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r36 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 15 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=0.735 $Y2=2.72
r38 15 17 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 10 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.545 $Y=2.72
+ $X2=0.735 $Y2=2.72
r40 10 12 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.545 $Y=2.72
+ $X2=0.23 $Y2=2.72
r41 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r43 4 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=2.635
+ $X2=0.735 $Y2=2.72
r44 4 6 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=0.735 $Y=2.635
+ $X2=0.735 $Y2=2.02
r45 1 6 300 $w=1.7e-07 $l=6.07577e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.76 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%Y 1 2 3 12 14 15 18 20 22 23 24 25 36 39
+ 47 55 58
r43 52 55 3.12409 $w=6.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=2.12
+ $X2=2.53 $Y2=2.12
r44 36 39 1.87607 $w=2.13e-07 $l=3.5e-08 $layer=LI1_cond $X=2.542 $Y=0.815
+ $X2=2.542 $Y2=0.85
r45 25 58 0.0357038 $w=6.68e-07 $l=2e-09 $layer=LI1_cond $X=2.54 $Y=2.12
+ $X2=2.542 $Y2=2.12
r46 25 58 7.5304 $w=2.15e-07 $l=3.35e-07 $layer=LI1_cond $X=2.542 $Y=1.785
+ $X2=2.542 $Y2=2.12
r47 25 55 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=2.54 $Y=2.12 $X2=2.53
+ $Y2=2.12
r48 24 25 9.86223 $w=3.83e-07 $l=2.55e-07 $layer=LI1_cond $X=2.542 $Y=1.53
+ $X2=2.542 $Y2=1.785
r49 23 24 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=2.542 $Y=1.19
+ $X2=2.542 $Y2=1.53
r50 22 36 0.116746 $w=1.88e-07 $l=2e-09 $layer=LI1_cond $X=2.54 $Y=0.72
+ $X2=2.542 $Y2=0.72
r51 22 23 16.8846 $w=2.13e-07 $l=3.15e-07 $layer=LI1_cond $X=2.542 $Y=0.875
+ $X2=2.542 $Y2=1.19
r52 22 39 1.34005 $w=2.13e-07 $l=2.5e-08 $layer=LI1_cond $X=2.542 $Y=0.875
+ $X2=2.542 $Y2=0.85
r53 20 52 4.90928 $w=6.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.08 $Y=2.12
+ $X2=2.355 $Y2=2.12
r54 20 47 0.178519 $w=6.68e-07 $l=1e-08 $layer=LI1_cond $X=2.08 $Y=2.12 $X2=2.07
+ $Y2=2.12
r55 16 22 10.0986 $w=1.88e-07 $l=1.73e-07 $layer=LI1_cond $X=2.367 $Y=0.72
+ $X2=2.54 $Y2=0.72
r56 16 18 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.367 $Y=0.625
+ $X2=2.367 $Y2=0.53
r57 14 16 6.5378 $w=1.88e-07 $l=1.12e-07 $layer=LI1_cond $X=2.255 $Y=0.72
+ $X2=2.367 $Y2=0.72
r58 14 15 53.4115 $w=1.88e-07 $l=9.15e-07 $layer=LI1_cond $X=2.255 $Y=0.72
+ $X2=1.34 $Y2=0.72
r59 10 15 6.81807 $w=1.9e-07 $l=1.33641e-07 $layer=LI1_cond $X=1.247 $Y=0.625
+ $X2=1.34 $Y2=0.72
r60 10 12 5.69533 $w=1.83e-07 $l=9.5e-08 $layer=LI1_cond $X=1.247 $Y=0.625
+ $X2=1.247 $Y2=0.53
r61 3 52 600 $w=1.7e-07 $l=8.94818e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.485 $X2=2.355 $Y2=2.27
r62 3 52 600 $w=1.7e-07 $l=4.88569e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.485 $X2=2.355 $Y2=1.87
r63 2 18 182 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_NDIFF $count=1 $X=2.08
+ $Y=0.235 $X2=2.355 $Y2=0.53
r64 1 12 182 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.235 $X2=1.24 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_1%VGND 1 2 7 9 11 13 20 21 28
r38 28 31 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.74 $Y=0 $X2=1.74
+ $Y2=0.36
r39 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r40 21 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r41 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r42 18 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.74
+ $Y2=0
r43 18 20 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.53
+ $Y2=0
r44 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r45 16 17 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r46 14 24 4.90409 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r47 14 16 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r48 13 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=1.74
+ $Y2=0
r49 13 16 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=1.55 $Y=0 $X2=0.69
+ $Y2=0
r50 11 17 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r51 11 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r52 7 24 2.94706 $w=3.4e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.212 $Y2=0
r53 7 9 14.4055 $w=3.38e-07 $l=4.25e-07 $layer=LI1_cond $X=0.255 $Y=0.085
+ $X2=0.255 $Y2=0.51
r54 2 31 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.765 $Y2=0.36
r55 1 9 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

