* File: sky130_fd_sc_hdll__buf_6.pex.spice
* Created: Thu Aug 27 19:00:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_6%A 1 3 6 8 10 13 15 16 19 29 35
r49 29 30 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.225 $Y=1.217
+ $X2=1.25 $Y2=1.217
r50 27 29 22.1035 $w=3.38e-07 $l=1.55e-07 $layer=POLY_cond $X=1.07 $Y=1.217
+ $X2=1.225 $Y2=1.217
r51 25 27 41.355 $w=3.38e-07 $l=2.9e-07 $layer=POLY_cond $X=0.78 $Y=1.217
+ $X2=1.07 $Y2=1.217
r52 24 25 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=0.755 $Y=1.217
+ $X2=0.78 $Y2=1.217
r53 19 24 16.3496 $w=3.38e-07 $l=1.253e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.755 $Y2=1.217
r54 19 21 24.4391 $w=2.7e-07 $l=1.1e-07 $layer=POLY_cond $X=0.655 $Y=1.16
+ $X2=0.545 $Y2=1.16
r55 16 35 2.40092 $w=2.38e-07 $l=5e-08 $layer=LI1_cond $X=1.025 $Y=1.195
+ $X2=0.975 $Y2=1.195
r56 16 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.07
+ $Y=1.16 $X2=1.07 $Y2=1.16
r57 15 35 24.0092 $w=2.38e-07 $l=5e-07 $layer=LI1_cond $X=0.475 $Y=1.195
+ $X2=0.975 $Y2=1.195
r58 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.545
+ $Y=1.16 $X2=0.545 $Y2=1.16
r59 11 30 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.25 $Y=1.025
+ $X2=1.25 $Y2=1.217
r60 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.25 $Y=1.025
+ $X2=1.25 $Y2=0.56
r61 8 29 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.217
r62 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.985
r63 4 25 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.78 $Y=1.025
+ $X2=0.78 $Y2=1.217
r64 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.78 $Y=1.025
+ $X2=0.78 $Y2=0.56
r65 1 24 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.755 $Y2=1.217
r66 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.755 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_6%A_169_297# 1 2 9 11 13 16 18 20 23 25 27 30
+ 32 34 37 39 41 42 44 47 51 53 55 57 58 59 62 64 67 72 84
c151 84 0 1.46608e-19 $X=4.045 $Y=1.217
r152 84 85 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=4.045 $Y=1.217
+ $X2=4.07 $Y2=1.217
r153 83 84 69.9198 $w=3.24e-07 $l=4.7e-07 $layer=POLY_cond $X=3.575 $Y=1.217
+ $X2=4.045 $Y2=1.217
r154 82 83 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.55 $Y=1.217
+ $X2=3.575 $Y2=1.217
r155 81 82 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=3.105 $Y=1.217
+ $X2=3.55 $Y2=1.217
r156 80 81 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=3.08 $Y=1.217
+ $X2=3.105 $Y2=1.217
r157 79 80 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=2.635 $Y=1.217
+ $X2=3.08 $Y2=1.217
r158 78 79 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.61 $Y=1.217
+ $X2=2.635 $Y2=1.217
r159 77 78 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=2.165 $Y=1.217
+ $X2=2.61 $Y2=1.217
r160 76 77 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.14 $Y=1.217
+ $X2=2.165 $Y2=1.217
r161 73 74 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.67 $Y=1.217
+ $X2=1.695 $Y2=1.217
r162 68 76 56.5309 $w=3.24e-07 $l=3.8e-07 $layer=POLY_cond $X=1.76 $Y=1.217
+ $X2=2.14 $Y2=1.217
r163 68 74 9.66975 $w=3.24e-07 $l=6.5e-08 $layer=POLY_cond $X=1.76 $Y=1.217
+ $X2=1.695 $Y2=1.217
r164 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=1.16 $X2=1.76 $Y2=1.16
r165 65 72 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=1.16
+ $X2=1.54 $Y2=1.16
r166 65 67 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.625 $Y=1.16
+ $X2=1.76 $Y2=1.16
r167 63 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.245
+ $X2=1.54 $Y2=1.16
r168 63 64 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=1.54 $Y=1.245
+ $X2=1.54 $Y2=1.485
r169 62 72 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.54 $Y=1.075
+ $X2=1.54 $Y2=1.16
r170 61 62 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.54 $Y=0.905
+ $X2=1.54 $Y2=1.075
r171 60 71 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.155 $Y=1.57
+ $X2=0.965 $Y2=1.57
r172 59 64 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=1.57
+ $X2=1.54 $Y2=1.485
r173 59 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.455 $Y=1.57
+ $X2=1.155 $Y2=1.57
r174 57 61 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=0.82
+ $X2=1.54 $Y2=0.905
r175 57 58 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.455 $Y=0.82
+ $X2=1.155 $Y2=0.82
r176 53 71 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.965 $Y=1.655
+ $X2=0.965 $Y2=1.57
r177 53 55 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=0.965 $Y=1.655
+ $X2=0.965 $Y2=2.31
r178 49 58 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.965 $Y=0.735
+ $X2=1.155 $Y2=0.82
r179 49 51 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=0.965 $Y=0.735
+ $X2=0.965 $Y2=0.38
r180 45 85 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.07 $Y=1.025
+ $X2=4.07 $Y2=1.217
r181 45 47 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.07 $Y=1.025
+ $X2=4.07 $Y2=0.56
r182 42 84 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.217
r183 42 44 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.045 $Y=1.41
+ $X2=4.045 $Y2=1.985
r184 39 83 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.217
r185 39 41 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.575 $Y=1.41
+ $X2=3.575 $Y2=1.985
r186 35 82 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.55 $Y=1.025
+ $X2=3.55 $Y2=1.217
r187 35 37 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.55 $Y=1.025
+ $X2=3.55 $Y2=0.56
r188 32 81 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.217
r189 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.105 $Y=1.41
+ $X2=3.105 $Y2=1.985
r190 28 80 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.08 $Y=1.025
+ $X2=3.08 $Y2=1.217
r191 28 30 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.08 $Y=1.025
+ $X2=3.08 $Y2=0.56
r192 25 79 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.217
r193 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.635 $Y=1.41
+ $X2=2.635 $Y2=1.985
r194 21 78 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.61 $Y=1.025
+ $X2=2.61 $Y2=1.217
r195 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.61 $Y=1.025
+ $X2=2.61 $Y2=0.56
r196 18 77 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.217
r197 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.165 $Y=1.41
+ $X2=2.165 $Y2=1.985
r198 14 76 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.14 $Y=1.025
+ $X2=2.14 $Y2=1.217
r199 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.14 $Y=1.025
+ $X2=2.14 $Y2=0.56
r200 11 74 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.695 $Y=1.41
+ $X2=1.695 $Y2=1.217
r201 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.695 $Y=1.41
+ $X2=1.695 $Y2=1.985
r202 7 73 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.67 $Y=1.025
+ $X2=1.67 $Y2=1.217
r203 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.67 $Y=1.025
+ $X2=1.67 $Y2=0.56
r204 2 71 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.845
+ $Y=1.485 $X2=0.99 $Y2=1.63
r205 2 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.845
+ $Y=1.485 $X2=0.99 $Y2=2.31
r206 1 51 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.855
+ $Y=0.235 $X2=0.99 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_6%VPWR 1 2 3 4 5 18 24 28 32 34 36 41 42 44 45
+ 47 48 50 51 52 54 70 76
r82 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r83 73 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 70 75 5.10144 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=4.332 $Y2=2.72
r86 70 72 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=2.72
+ $X2=3.91 $Y2=2.72
r87 69 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r88 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r89 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r90 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r92 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r93 54 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 52 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 50 68 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.125 $Y=2.72
+ $X2=2.99 $Y2=2.72
r96 50 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=2.72
+ $X2=3.315 $Y2=2.72
r97 49 72 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.91 $Y2=2.72
r98 49 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.505 $Y=2.72
+ $X2=3.315 $Y2=2.72
r99 47 65 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 47 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.185 $Y=2.72
+ $X2=2.375 $Y2=2.72
r101 46 68 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.99 $Y2=2.72
r102 46 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.565 $Y=2.72
+ $X2=2.375 $Y2=2.72
r103 44 62 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.15 $Y2=2.72
r104 44 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.495 $Y2=2.72
r105 43 65 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=1.615 $Y=2.72
+ $X2=2.07 $Y2=2.72
r106 43 45 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.615 $Y=2.72
+ $X2=1.495 $Y2=2.72
r107 41 52 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.23 $Y2=2.72
r108 41 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.52 $Y2=2.72
r109 40 62 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=1.15 $Y2=2.72
r110 40 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.52 $Y2=2.72
r111 36 39 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.255 $Y=1.66
+ $X2=4.255 $Y2=2.34
r112 34 75 3.09525 $w=3.8e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.255 $Y=2.635
+ $X2=4.332 $Y2=2.72
r113 34 39 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.255 $Y=2.635
+ $X2=4.255 $Y2=2.34
r114 30 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=2.635
+ $X2=3.315 $Y2=2.72
r115 30 32 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.315 $Y=2.635
+ $X2=3.315 $Y2=2
r116 26 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=2.635
+ $X2=2.375 $Y2=2.72
r117 26 28 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.375 $Y=2.635
+ $X2=2.375 $Y2=2
r118 22 45 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.495 $Y=2.635
+ $X2=1.495 $Y2=2.72
r119 22 24 30.4917 $w=2.38e-07 $l=6.35e-07 $layer=LI1_cond $X=1.495 $Y=2.635
+ $X2=1.495 $Y2=2
r120 18 21 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.52 $Y=1.66
+ $X2=0.52 $Y2=2.34
r121 16 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=2.635
+ $X2=0.52 $Y2=2.72
r122 16 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.52 $Y=2.635
+ $X2=0.52 $Y2=2.34
r123 5 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.28 $Y2=2.34
r124 5 36 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.135
+ $Y=1.485 $X2=4.28 $Y2=1.66
r125 4 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.195
+ $Y=1.485 $X2=3.34 $Y2=2
r126 3 28 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.255
+ $Y=1.485 $X2=2.4 $Y2=2
r127 2 24 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.315
+ $Y=1.485 $X2=1.46 $Y2=2
r128 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.485 $X2=0.52 $Y2=2.34
r129 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.395
+ $Y=1.485 $X2=0.52 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_6%X 1 2 3 4 5 6 21 25 27 28 29 30 33 37 41 45
+ 47 55 59
r91 58 59 13.0318 $w=8.78e-07 $l=9.4e-07 $layer=LI1_cond $X=2.87 $Y=1.175
+ $X2=3.81 $Y2=1.175
r92 55 58 3.25795 $w=8.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.635 $Y=1.175
+ $X2=2.87 $Y2=1.175
r93 47 55 0.346591 $w=8.78e-07 $l=2.5e-08 $layer=LI1_cond $X=2.61 $Y=1.175
+ $X2=2.635 $Y2=1.175
r94 43 59 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=3.81 $Y=1.615
+ $X2=3.81 $Y2=1.175
r95 43 45 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.81 $Y=1.615
+ $X2=3.81 $Y2=1.755
r96 39 59 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=3.81 $Y=0.735
+ $X2=3.81 $Y2=1.175
r97 39 41 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.81 $Y=0.735
+ $X2=3.81 $Y2=0.56
r98 35 58 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=2.87 $Y=1.615
+ $X2=2.87 $Y2=1.175
r99 35 37 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=2.87 $Y=1.615
+ $X2=2.87 $Y2=1.755
r100 31 58 10.8514 $w=1.7e-07 $l=4.4e-07 $layer=LI1_cond $X=2.87 $Y=0.735
+ $X2=2.87 $Y2=1.175
r101 31 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.87 $Y=0.735
+ $X2=2.87 $Y2=0.56
r102 29 47 6.69542 $w=4.4e-07 $l=4.43875e-07 $layer=LI1_cond $X=2.41 $Y=1.53
+ $X2=2.61 $Y2=1.175
r103 29 30 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.41 $Y=1.53
+ $X2=2.015 $Y2=1.53
r104 27 47 6.69542 $w=4.4e-07 $l=4.43875e-07 $layer=LI1_cond $X=2.41 $Y=0.82
+ $X2=2.61 $Y2=1.175
r105 27 28 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=2.41 $Y=0.82
+ $X2=2.015 $Y2=0.82
r106 23 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.93 $Y=1.615
+ $X2=2.015 $Y2=1.53
r107 23 25 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.93 $Y=1.615
+ $X2=1.93 $Y2=1.755
r108 19 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.93 $Y=0.735
+ $X2=2.015 $Y2=0.82
r109 19 21 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.93 $Y=0.735
+ $X2=1.93 $Y2=0.56
r110 6 45 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.665
+ $Y=1.485 $X2=3.81 $Y2=1.755
r111 5 37 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.725
+ $Y=1.485 $X2=2.87 $Y2=1.755
r112 4 25 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.785
+ $Y=1.485 $X2=1.93 $Y2=1.755
r113 3 41 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=3.625
+ $Y=0.235 $X2=3.81 $Y2=0.56
r114 2 33 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=2.685
+ $Y=0.235 $X2=2.87 $Y2=0.56
r115 1 21 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=1.745
+ $Y=0.235 $X2=1.93 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_6%VGND 1 2 3 4 5 18 22 26 30 32 34 37 38 40 41
+ 43 44 46 47 48 50 66 72
c82 26 0 1.46608e-19 $X=2.4 $Y=0.4
r83 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r84 69 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r85 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r86 66 71 5.10144 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=4.332
+ $Y2=0
r87 66 68 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.065 $Y=0 $X2=3.91
+ $Y2=0
r88 65 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r89 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r90 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r91 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r93 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r94 50 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r95 48 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r96 46 64 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=2.99
+ $Y2=0
r97 46 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.125 $Y=0 $X2=3.315
+ $Y2=0
r98 45 68 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.91
+ $Y2=0
r99 45 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.315
+ $Y2=0
r100 43 61 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.185 $Y=0
+ $X2=2.07 $Y2=0
r101 43 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.185 $Y=0 $X2=2.375
+ $Y2=0
r102 42 64 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.565 $Y=0
+ $X2=2.99 $Y2=0
r103 42 44 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.375
+ $Y2=0
r104 40 58 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=0
+ $X2=1.15 $Y2=0
r105 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=0 $X2=1.46
+ $Y2=0
r106 39 61 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=1.545 $Y=0
+ $X2=2.07 $Y2=0
r107 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.545 $Y=0 $X2=1.46
+ $Y2=0
r108 37 48 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.23 $Y2=0
r109 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.435 $Y=0 $X2=0.52
+ $Y2=0
r110 36 58 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.605 $Y=0
+ $X2=1.15 $Y2=0
r111 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=0 $X2=0.52
+ $Y2=0
r112 32 71 3.09525 $w=3.8e-07 $l=1.17346e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.332 $Y2=0
r113 32 34 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=4.255 $Y=0.085
+ $X2=4.255 $Y2=0.38
r114 28 47 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0
r115 28 30 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.315 $Y=0.085
+ $X2=3.315 $Y2=0.4
r116 24 44 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0
r117 24 26 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.375 $Y=0.085
+ $X2=2.375 $Y2=0.4
r118 20 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.46 $Y=0.085
+ $X2=1.46 $Y2=0
r119 20 22 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.46 $Y=0.085
+ $X2=1.46 $Y2=0.4
r120 16 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0
r121 16 18 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0.4
r122 5 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.145
+ $Y=0.235 $X2=4.28 $Y2=0.38
r123 4 30 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.155
+ $Y=0.235 $X2=3.34 $Y2=0.4
r124 3 26 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.215
+ $Y=0.235 $X2=2.4 $Y2=0.4
r125 2 22 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=1.325
+ $Y=0.235 $X2=1.46 $Y2=0.4
r126 1 18 182 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=1 $X=0.395
+ $Y=0.235 $X2=0.52 $Y2=0.4
.ends

