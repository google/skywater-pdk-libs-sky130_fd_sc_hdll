* File: sky130_fd_sc_hdll__o22a_2.pex.spice
* Created: Wed Sep  2 08:45:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22A_2%A_83_21# 1 2 7 9 10 12 13 15 16 18 22 25 26
+ 27 28 30 32 34 36 42
c84 28 0 1.35542e-19 $X=2.075 $Y=0.77
r85 41 42 4.62192 $w=3.65e-07 $l=3.5e-08 $layer=POLY_cond $X=0.95 $Y=1.202
+ $X2=0.985 $Y2=1.202
r86 40 41 57.4438 $w=3.65e-07 $l=4.35e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.95 $Y2=1.202
r87 39 40 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r88 32 38 2.93335 $w=3.55e-07 $l=1.25e-07 $layer=LI1_cond $X=2.517 $Y=1.705
+ $X2=2.517 $Y2=1.58
r89 32 34 19.3156 $w=3.53e-07 $l=5.95e-07 $layer=LI1_cond $X=2.517 $Y=1.705
+ $X2=2.517 $Y2=2.3
r90 28 36 6.68437 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.77
+ $X2=1.95 $Y2=0.77
r91 28 30 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.77
+ $X2=2.2 $Y2=0.77
r92 26 38 4.15363 $w=2.5e-07 $l=1.77e-07 $layer=LI1_cond $X=2.34 $Y=1.58
+ $X2=2.517 $Y2=1.58
r93 26 27 45.4063 $w=2.48e-07 $l=9.85e-07 $layer=LI1_cond $X=2.34 $Y=1.58
+ $X2=1.355 $Y2=1.58
r94 25 36 36.6616 $w=1.78e-07 $l=5.95e-07 $layer=LI1_cond $X=1.355 $Y=0.805
+ $X2=1.95 $Y2=0.805
r95 23 42 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=1.235 $Y=1.202
+ $X2=0.985 $Y2=1.202
r96 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.235
+ $Y=1.16 $X2=1.235 $Y2=1.16
r97 20 27 6.84494 $w=2.5e-07 $l=1.92614e-07 $layer=LI1_cond $X=1.215 $Y=1.455
+ $X2=1.355 $Y2=1.58
r98 20 22 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.215 $Y=1.455
+ $X2=1.215 $Y2=1.16
r99 19 25 7.24404 $w=1.8e-07 $l=1.79444e-07 $layer=LI1_cond $X=1.215 $Y=0.895
+ $X2=1.355 $Y2=0.805
r100 19 22 10.9071 $w=2.78e-07 $l=2.65e-07 $layer=LI1_cond $X=1.215 $Y=0.895
+ $X2=1.215 $Y2=1.16
r101 16 42 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r102 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r103 13 41 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=1.202
r104 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.95 $Y=0.995
+ $X2=0.95 $Y2=0.56
r105 10 40 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r106 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r107 7 39 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r108 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
r109 2 38 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r110 2 34 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r111 1 30 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.2 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%B1 1 3 4 6 7 12
c31 7 0 1.46155e-19 $X=1.75 $Y=1.19
r32 12 13 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.965 $Y=1.202
+ $X2=1.99 $Y2=1.202
r33 10 12 31.6932 $w=3.65e-07 $l=2.4e-07 $layer=POLY_cond $X=1.725 $Y=1.202
+ $X2=1.965 $Y2=1.202
r34 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r35 4 13 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=1.202
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.99 $Y=0.995 $X2=1.99
+ $Y2=0.56
r37 1 12 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.202
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%B2 1 3 4 6 7 15
c33 1 0 2.70899e-19 $X=2.375 $Y=1.41
r34 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.16 $X2=2.41 $Y2=1.16
r35 7 15 7.76364 $w=1.98e-07 $l=1.4e-07 $layer=LI1_cond $X=2.215 $Y=1.175
+ $X2=2.355 $Y2=1.175
r36 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=2.41 $Y=0.995
+ $X2=2.435 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.41 $Y=0.995 $X2=2.41
+ $Y2=0.56
r38 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.435 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%A2 1 3 4 6 9 13
c36 13 0 1.7643e-19 $X=2.985 $Y=1.87
r37 12 13 25.3964 $w=2.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.04 $Y=1.275
+ $X2=3.04 $Y2=1.87
r38 9 12 4.46939 $w=3.78e-07 $l=1.15e-07 $layer=LI1_cond $X=2.985 $Y=1.16
+ $X2=2.985 $Y2=1.275
r39 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.96
+ $Y=1.16 $X2=2.96 $Y2=1.16
r40 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.07 $Y=0.995
+ $X2=2.975 $Y2=1.16
r41 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.07 $Y=0.995 $X2=3.07
+ $Y2=0.56
r42 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=3.045 $Y=1.41
+ $X2=2.975 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.045 $Y=1.41
+ $X2=3.045 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%A1 1 3 4 6 7 8 13
r23 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.54
+ $Y=1.16 $X2=3.54 $Y2=1.16
r24 7 8 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.525 $Y=1.19
+ $X2=3.525 $Y2=1.53
r25 7 13 0.960369 $w=3.58e-07 $l=3e-08 $layer=LI1_cond $X=3.525 $Y=1.19
+ $X2=3.525 $Y2=1.16
r26 4 12 38.7956 $w=3.51e-07 $l=1.83916e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.55 $Y2=1.16
r27 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995 $X2=3.51
+ $Y2=0.56
r28 1 12 45.736 $w=3.51e-07 $l=2.93684e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.55 $Y2=1.16
r29 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.455 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%VPWR 1 2 3 10 12 16 18 20 22 24 36 46 50
r46 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r47 40 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 40 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 39 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 36 39 11.3627 $w=7.98e-07 $l=7.6e-07 $layer=LI1_cond $X=1.495 $Y=1.96
+ $X2=1.495 $Y2=2.72
r52 33 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 31 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r54 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r56 28 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 25 39 10.2089 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=1.895 $Y=2.72 $X2=1.495
+ $Y2=2.72
r60 25 27 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 24 45 4.42303 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.855 $Y2=2.72
r62 24 30 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 22 50 0.00426813 $w=4.8e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=2.72
+ $X2=0.23 $Y2=2.72
r64 18 45 3.25908 $w=3.2e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.855 $Y2=2.72
r65 18 20 24.3093 $w=3.18e-07 $l=6.75e-07 $layer=LI1_cond $X=3.73 $Y=2.635
+ $X2=3.73 $Y2=1.96
r66 17 33 4.00981 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=2.72
+ $X2=0.182 $Y2=2.72
r67 16 39 10.2089 $w=1.7e-07 $l=4e-07 $layer=LI1_cond $X=1.095 $Y=2.72 $X2=1.495
+ $Y2=2.72
r68 16 17 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.365 $Y2=2.72
r69 12 15 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.62
+ $X2=0.24 $Y2=2.3
r70 10 33 3.13335 $w=2.5e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.182 $Y2=2.72
r71 10 15 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.3
r72 3 20 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.545
+ $Y=1.485 $X2=3.69 $Y2=1.96
r73 2 36 150 $w=1.7e-07 $l=8.6032e-07 $layer=licon1_PDIFF $count=4 $X=1.075
+ $Y=1.485 $X2=1.73 $Y2=1.96
r74 1 15 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r75 1 12 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%X 1 2 7 10
r17 10 13 47.2502 $w=2.48e-07 $l=1.025e-06 $layer=LI1_cond $X=0.73 $Y=0.595
+ $X2=0.73 $Y2=1.62
r18 7 17 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=0.73 $Y=2.21 $X2=0.73
+ $Y2=2.3
r19 7 13 27.1977 $w=2.48e-07 $l=5.9e-07 $layer=LI1_cond $X=0.73 $Y=2.21 $X2=0.73
+ $Y2=1.62
r20 2 17 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.3
r21 2 13 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.62
r22 1 10 182 $w=1.7e-07 $l=4.38862e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.74 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%VGND 1 2 3 10 12 14 18 22 25 26 27 37 38 44
+ 49
r56 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.23
+ $Y2=0
r57 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 41 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r59 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r60 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r61 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r62 32 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r63 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r64 31 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.99
+ $Y2=0
r65 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r66 29 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.215
+ $Y2=0
r67 29 31 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.61
+ $Y2=0
r68 27 49 0.00426813 $w=4.8e-07 $l=1.5e-08 $layer=MET1_cond $X=0.215 $Y=0
+ $X2=0.23 $Y2=0
r69 25 34 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.195 $Y=0 $X2=2.99
+ $Y2=0
r70 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.195 $Y=0 $X2=3.28
+ $Y2=0
r71 24 37 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.91
+ $Y2=0
r72 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.365 $Y=0 $X2=3.28
+ $Y2=0
r73 20 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0
r74 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.28 $Y=0.085
+ $X2=3.28 $Y2=0.36
r75 16 44 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0
r76 16 18 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0.38
r77 15 41 3.40825 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r78 14 44 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.215
+ $Y2=0
r79 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.355
+ $Y2=0
r80 10 41 3.40825 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.177 $Y2=0
r81 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r82 3 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.145
+ $Y=0.235 $X2=3.28 $Y2=0.36
r83 2 18 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.235 $X2=1.21 $Y2=0.38
r84 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_2%A_321_47# 1 2 3 10 14 15 16 20
c43 15 0 1.24744e-19 $X=2.76 $Y=0.695
r44 18 20 10.4924 $w=3.33e-07 $l=3.05e-07 $layer=LI1_cond $X=3.722 $Y=0.695
+ $X2=3.722 $Y2=0.39
r45 17 25 5.2341 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.93 $Y=0.78 $X2=2.76
+ $Y2=0.78
r46 16 18 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.555 $Y=0.78
+ $X2=3.722 $Y2=0.695
r47 16 17 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.555 $Y=0.78
+ $X2=2.93 $Y2=0.78
r48 15 25 2.61705 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.76 $Y=0.695
+ $X2=2.76 $Y2=0.78
r49 14 23 2.66241 $w=3.4e-07 $l=9e-08 $layer=LI1_cond $X=2.76 $Y=0.475 $X2=2.76
+ $Y2=0.385
r50 14 15 7.45698 $w=3.38e-07 $l=2.2e-07 $layer=LI1_cond $X=2.76 $Y=0.475
+ $X2=2.76 $Y2=0.695
r51 10 23 5.02899 $w=1.8e-07 $l=1.7e-07 $layer=LI1_cond $X=2.59 $Y=0.385
+ $X2=2.76 $Y2=0.385
r52 10 12 52.9899 $w=1.78e-07 $l=8.6e-07 $layer=LI1_cond $X=2.59 $Y=0.385
+ $X2=1.73 $Y2=0.385
r53 3 20 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.39
r54 2 25 182 $w=1.7e-07 $l=6.15366e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.755 $Y2=0.73
r55 2 23 182 $w=1.7e-07 $l=3.38748e-07 $layer=licon1_NDIFF $count=1 $X=2.485
+ $Y=0.235 $X2=2.755 $Y2=0.39
r56 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.73 $Y2=0.39
.ends

