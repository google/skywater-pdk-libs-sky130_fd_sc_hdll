* File: sky130_fd_sc_hdll__einvp_2.pxi.spice
* Created: Thu Aug 27 19:07:56 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVP_2%TE N_TE_M1008_g N_TE_c_67_n N_TE_c_68_n
+ N_TE_M1002_g N_TE_c_60_n N_TE_c_61_n N_TE_c_62_n N_TE_M1004_g N_TE_c_63_n
+ N_TE_c_64_n N_TE_M1005_g N_TE_c_65_n TE TE PM_SKY130_FD_SC_HDLL__EINVP_2%TE
x_PM_SKY130_FD_SC_HDLL__EINVP_2%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_115_n N_A_27_47#_M1001_g N_A_27_47#_c_116_n N_A_27_47#_c_117_n
+ N_A_27_47#_c_118_n N_A_27_47#_M1009_g N_A_27_47#_c_119_n N_A_27_47#_c_111_n
+ N_A_27_47#_c_120_n N_A_27_47#_c_121_n N_A_27_47#_c_112_n N_A_27_47#_c_113_n
+ N_A_27_47#_c_114_n PM_SKY130_FD_SC_HDLL__EINVP_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVP_2%A N_A_c_184_n N_A_M1000_g N_A_c_188_n
+ N_A_M1003_g N_A_c_189_n N_A_M1007_g N_A_c_185_n N_A_M1006_g A A A N_A_c_187_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%A
x_PM_SKY130_FD_SC_HDLL__EINVP_2%VPWR N_VPWR_M1002_d N_VPWR_M1001_d
+ N_VPWR_c_226_n N_VPWR_c_227_n N_VPWR_c_228_n VPWR N_VPWR_c_229_n
+ N_VPWR_c_230_n N_VPWR_c_225_n N_VPWR_c_232_n N_VPWR_c_233_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVP_2%A_235_309# N_A_235_309#_M1001_s
+ N_A_235_309#_M1009_s N_A_235_309#_M1007_d N_A_235_309#_c_272_n
+ N_A_235_309#_c_281_n N_A_235_309#_c_273_n N_A_235_309#_c_287_n
+ N_A_235_309#_c_274_n N_A_235_309#_c_307_n N_A_235_309#_c_275_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%A_235_309#
x_PM_SKY130_FD_SC_HDLL__EINVP_2%Z N_Z_M1000_d N_Z_M1003_s Z Z Z Z N_Z_c_315_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%Z
x_PM_SKY130_FD_SC_HDLL__EINVP_2%VGND N_VGND_M1008_d N_VGND_M1005_d
+ N_VGND_c_334_n VGND N_VGND_c_335_n N_VGND_c_336_n N_VGND_c_337_n
+ N_VGND_c_338_n N_VGND_c_339_n N_VGND_c_340_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%VGND
x_PM_SKY130_FD_SC_HDLL__EINVP_2%A_214_47# N_A_214_47#_M1004_s
+ N_A_214_47#_M1000_s N_A_214_47#_M1006_s N_A_214_47#_c_388_n
+ N_A_214_47#_c_384_n N_A_214_47#_c_390_n N_A_214_47#_c_385_n
+ N_A_214_47#_c_386_n N_A_214_47#_c_387_n
+ PM_SKY130_FD_SC_HDLL__EINVP_2%A_214_47#
cc_1 VNB N_TE_M1008_g 0.0346601f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_c_60_n 0.0199643f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.035
cc_3 VNB N_TE_c_61_n 0.040911f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.035
cc_4 VNB N_TE_c_62_n 0.0149371f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.96
cc_5 VNB N_TE_c_63_n 0.0251182f $X=-0.19 $Y=-0.24 $X2=1.39 $Y2=1.035
cc_6 VNB N_TE_c_64_n 0.0186925f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=0.96
cc_7 VNB N_TE_c_65_n 0.00649751f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.035
cc_8 VNB TE 0.0134128f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB N_A_27_47#_c_111_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=0.56
cc_10 VNB N_A_27_47#_c_112_n 0.00998586f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_11 VNB N_A_27_47#_c_113_n 0.00582006f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.142
cc_12 VNB N_A_27_47#_c_114_n 0.0313775f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_13 VNB N_A_c_184_n 0.0224159f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_14 VNB N_A_c_185_n 0.0196f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.035
cc_15 VNB A 0.021336f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.56
cc_16 VNB N_A_c_187_n 0.0635629f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_17 VNB N_VPWR_c_225_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_18 VNB N_VGND_c_334_n 0.00595067f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_19 VNB N_VGND_c_335_n 0.0143387f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.56
cc_20 VNB N_VGND_c_336_n 0.0139345f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=0.56
cc_21 VNB N_VGND_c_337_n 0.044959f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.142
cc_22 VNB N_VGND_c_338_n 0.205679f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.142
cc_23 VNB N_VGND_c_339_n 0.00604126f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_24 VNB N_VGND_c_340_n 0.00584155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_214_47#_c_384_n 0.00964742f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.56
cc_26 VNB N_A_214_47#_c_385_n 0.00333309f $X=-0.19 $Y=-0.24 $X2=1.465 $Y2=0.56
cc_27 VNB N_A_214_47#_c_386_n 0.0144618f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=1.035
cc_28 VNB N_A_214_47#_c_387_n 0.00191465f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_29 VPB N_TE_c_67_n 0.0260626f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_30 VPB N_TE_c_68_n 0.0324792f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_31 VPB N_TE_c_61_n 0.0103959f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.035
cc_32 VPB TE 0.0160339f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_27_47#_c_115_n 0.0195251f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_34 VPB N_A_27_47#_c_116_n 0.00851129f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.035
cc_35 VPB N_A_27_47#_c_117_n 0.0115354f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.035
cc_36 VPB N_A_27_47#_c_118_n 0.0173104f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.96
cc_37 VPB N_A_27_47#_c_119_n 0.00997866f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.035
cc_38 VPB N_A_27_47#_c_120_n 0.0198678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_121_n 0.0221716f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_40 VPB N_A_27_47#_c_113_n 0.011547f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.142
cc_41 VPB N_A_27_47#_c_114_n 0.0011297f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_42 VPB N_A_c_188_n 0.0171409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_c_189_n 0.0188133f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_44 VPB A 0.013525f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.56
cc_45 VPB N_A_c_187_n 0.0323965f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_46 VPB N_VPWR_c_226_n 0.00760933f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_47 VPB N_VPWR_c_227_n 0.0182895f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.035
cc_48 VPB N_VPWR_c_228_n 4.89148e-19 $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.035
cc_49 VPB N_VPWR_c_229_n 0.0150576f $X=-0.19 $Y=1.305 $X2=1.465 $Y2=0.56
cc_50 VPB N_VPWR_c_230_n 0.0436391f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.142
cc_51 VPB N_VPWR_c_225_n 0.0559585f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_52 VPB N_VPWR_c_232_n 0.00638089f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_53 VPB N_VPWR_c_233_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_235_309#_c_272_n 0.00798738f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=0.96
cc_55 VPB N_A_235_309#_c_273_n 0.00181253f $X=-0.19 $Y=1.305 $X2=1.39 $Y2=1.035
cc_56 VPB N_A_235_309#_c_274_n 0.00793407f $X=-0.19 $Y=1.305 $X2=0.995 $Y2=1.035
cc_57 VPB N_A_235_309#_c_275_n 0.0205972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 N_TE_c_63_n N_A_27_47#_c_117_n 0.00686273f $X=1.39 $Y=1.035 $X2=0 $Y2=0
cc_59 N_TE_c_68_n N_A_27_47#_c_120_n 0.00707894f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_60 N_TE_c_67_n N_A_27_47#_c_121_n 0.0146652f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_61 N_TE_c_68_n N_A_27_47#_c_121_n 0.0268362f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_62 N_TE_c_60_n N_A_27_47#_c_121_n 5.7676e-19 $X=0.92 $Y=1.035 $X2=0 $Y2=0
cc_63 N_TE_c_61_n N_A_27_47#_c_121_n 0.00264156f $X=0.595 $Y=1.035 $X2=0 $Y2=0
cc_64 TE N_A_27_47#_c_121_n 0.043173f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_65 N_TE_M1008_g N_A_27_47#_c_112_n 0.0245081f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_66 N_TE_c_60_n N_A_27_47#_c_112_n 0.0161511f $X=0.92 $Y=1.035 $X2=0 $Y2=0
cc_67 N_TE_c_61_n N_A_27_47#_c_112_n 0.0191449f $X=0.595 $Y=1.035 $X2=0 $Y2=0
cc_68 N_TE_c_62_n N_A_27_47#_c_112_n 0.00868069f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_69 N_TE_c_64_n N_A_27_47#_c_112_n 7.12865e-19 $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_70 N_TE_c_65_n N_A_27_47#_c_112_n 0.00171953f $X=0.995 $Y=1.035 $X2=0 $Y2=0
cc_71 TE N_A_27_47#_c_112_n 0.0471178f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_72 N_TE_c_63_n N_A_27_47#_c_113_n 0.0218309f $X=1.39 $Y=1.035 $X2=0 $Y2=0
cc_73 N_TE_c_65_n N_A_27_47#_c_113_n 0.0111081f $X=0.995 $Y=1.035 $X2=0 $Y2=0
cc_74 N_TE_c_63_n N_A_27_47#_c_114_n 0.00620476f $X=1.39 $Y=1.035 $X2=0 $Y2=0
cc_75 N_TE_c_68_n N_VPWR_c_226_n 0.0144429f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_76 N_TE_c_68_n N_VPWR_c_229_n 0.00427505f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_77 N_TE_c_68_n N_VPWR_c_225_n 0.0049402f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_78 N_TE_c_68_n N_A_235_309#_c_272_n 0.00550327f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_79 N_TE_c_67_n N_A_235_309#_c_273_n 6.88195e-19 $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_80 N_TE_c_63_n N_A_235_309#_c_273_n 0.00118725f $X=1.39 $Y=1.035 $X2=0 $Y2=0
cc_81 N_TE_c_62_n N_VGND_c_334_n 5.54177e-19 $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_82 N_TE_c_64_n N_VGND_c_334_n 0.0082289f $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_83 N_TE_M1008_g N_VGND_c_335_n 0.00342301f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_84 N_TE_c_62_n N_VGND_c_336_n 0.00565872f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_85 N_TE_c_64_n N_VGND_c_336_n 0.00341689f $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_86 N_TE_M1008_g N_VGND_c_338_n 0.00501518f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_87 N_TE_c_62_n N_VGND_c_338_n 0.00963525f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_88 N_TE_c_64_n N_VGND_c_338_n 0.00415805f $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_89 N_TE_M1008_g N_VGND_c_339_n 0.0128359f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_90 N_TE_c_60_n N_VGND_c_339_n 7.92531e-19 $X=0.92 $Y=1.035 $X2=0 $Y2=0
cc_91 N_TE_c_62_n N_VGND_c_339_n 0.00617076f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_92 N_TE_c_64_n N_VGND_c_339_n 5.38903e-19 $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_93 N_TE_c_62_n N_A_214_47#_c_388_n 0.00453937f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_94 N_TE_c_64_n N_A_214_47#_c_384_n 0.0125552f $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_95 N_TE_c_62_n N_A_214_47#_c_390_n 0.00122495f $X=0.995 $Y=0.96 $X2=0 $Y2=0
cc_96 N_TE_c_63_n N_A_214_47#_c_390_n 0.00289368f $X=1.39 $Y=1.035 $X2=0 $Y2=0
cc_97 N_TE_c_64_n N_A_214_47#_c_385_n 0.00305716f $X=1.465 $Y=0.96 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_118_n N_A_c_188_n 0.0181122f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_119_n N_A_c_188_n 0.00195253f $X=1.945 $Y=1.395 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_113_n N_A_c_187_n 0.00166709f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_114_n N_A_c_187_n 0.0120237f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_121_n N_VPWR_M1002_d 0.00270444f $X=0.712 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_27_47#_c_115_n N_VPWR_c_226_n 0.00290558f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_120_n N_VPWR_c_226_n 0.0263462f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_121_n N_VPWR_c_226_n 0.0276039f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_115_n N_VPWR_c_227_n 0.00622633f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_115_n N_VPWR_c_228_n 0.0128003f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_118_n N_VPWR_c_228_n 0.012625f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_120_n N_VPWR_c_229_n 0.0178308f $X=0.26 $Y=2.165 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_118_n N_VPWR_c_230_n 0.00622633f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_M1002_s N_VPWR_c_225_n 0.00252291f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_115_n N_VPWR_c_225_n 0.0116835f $X=1.535 $Y=1.47 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_118_n N_VPWR_c_225_n 0.0107403f $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_120_n N_VPWR_c_225_n 0.00986266f $X=0.26 $Y=2.165 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_c_121_n N_VPWR_c_225_n 0.00695765f $X=0.712 $Y=1.785 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_115_n N_A_235_309#_c_272_n 0.00651494f $X=1.535 $Y=1.47
+ $X2=0 $Y2=0
cc_117 N_A_27_47#_c_121_n N_A_235_309#_c_272_n 0.0162418f $X=0.712 $Y=1.785
+ $X2=0 $Y2=0
cc_118 N_A_27_47#_c_115_n N_A_235_309#_c_281_n 0.0184699f $X=1.535 $Y=1.47 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_116_n N_A_235_309#_c_281_n 0.00262074f $X=1.785 $Y=1.395
+ $X2=0 $Y2=0
cc_120 N_A_27_47#_c_118_n N_A_235_309#_c_281_n 0.0173569f $X=2.005 $Y=1.47 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_c_113_n N_A_235_309#_c_281_n 0.0360656f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_121_n N_A_235_309#_c_273_n 0.0127748f $X=0.712 $Y=1.785
+ $X2=0 $Y2=0
cc_123 N_A_27_47#_c_113_n N_A_235_309#_c_273_n 0.0167775f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A_27_47#_c_118_n N_A_235_309#_c_287_n 0.00489748f $X=2.005 $Y=1.47
+ $X2=0 $Y2=0
cc_125 N_A_27_47#_c_118_n N_Z_c_315_n 6.66076e-19 $X=2.005 $Y=1.47 $X2=0 $Y2=0
cc_126 N_A_27_47#_c_119_n N_Z_c_315_n 8.18929e-19 $X=1.945 $Y=1.395 $X2=0 $Y2=0
cc_127 N_A_27_47#_c_113_n N_Z_c_315_n 0.0102978f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_114_n N_Z_c_315_n 3.3604e-19 $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_112_n N_VGND_M1008_d 0.0035013f $X=0.925 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_27_47#_c_111_n N_VGND_c_335_n 0.0177719f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_112_n N_VGND_c_335_n 0.00273609f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_M1008_s N_VGND_c_338_n 0.00228937f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_111_n N_VGND_c_338_n 0.00989054f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_112_n N_VGND_c_338_n 0.00617642f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_112_n N_VGND_c_339_n 0.0270485f $X=0.925 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_117_n N_A_214_47#_c_384_n 8.32206e-19 $X=1.625 $Y=1.395
+ $X2=0 $Y2=0
cc_137 N_A_27_47#_c_113_n N_A_214_47#_c_384_n 0.0535561f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_c_114_n N_A_214_47#_c_384_n 0.00832597f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_112_n N_A_214_47#_c_390_n 0.0121615f $X=0.925 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_c_113_n N_A_214_47#_c_390_n 0.0155723f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_c_188_n N_VPWR_c_228_n 0.00107169f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_188_n N_VPWR_c_230_n 0.00429453f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_189_n N_VPWR_c_230_n 0.00429453f $X=3.095 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_188_n N_VPWR_c_225_n 0.00645807f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_189_n N_VPWR_c_225_n 0.00704999f $X=3.095 $Y=1.41 $X2=0 $Y2=0
cc_146 A N_A_235_309#_M1007_d 0.00461267f $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_147 N_A_c_188_n N_A_235_309#_c_281_n 0.00168697f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_188_n N_A_235_309#_c_287_n 0.00717311f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_188_n N_A_235_309#_c_274_n 0.0147259f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_189_n N_A_235_309#_c_274_n 0.0122476f $X=3.095 $Y=1.41 $X2=0 $Y2=0
cc_151 A N_A_235_309#_c_275_n 0.0257774f $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_152 N_A_c_187_n N_A_235_309#_c_275_n 0.0011073f $X=3.12 $Y=1.202 $X2=0 $Y2=0
cc_153 N_A_c_184_n N_Z_c_315_n 0.012153f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_188_n N_Z_c_315_n 0.0151788f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_189_n N_Z_c_315_n 0.0180386f $X=3.095 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_185_n N_Z_c_315_n 0.0121914f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_157 A N_Z_c_315_n 0.0613625f $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_158 N_A_c_187_n N_Z_c_315_n 0.0400277f $X=3.12 $Y=1.202 $X2=0 $Y2=0
cc_159 N_A_c_184_n N_VGND_c_334_n 0.0027212f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_c_184_n N_VGND_c_337_n 0.00357877f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_185_n N_VGND_c_337_n 0.00357877f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_184_n N_VGND_c_338_n 0.00689275f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_185_n N_VGND_c_338_n 0.00650683f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_164 A N_VGND_c_338_n 7.88603e-19 $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_165 A N_A_214_47#_M1006_s 0.00275832f $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A_c_184_n N_A_214_47#_c_386_n 0.0154277f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_185_n N_A_214_47#_c_386_n 0.011843f $X=3.12 $Y=0.995 $X2=0 $Y2=0
cc_168 A N_A_214_47#_c_386_n 0.0232068f $X=3.305 $Y=0.765 $X2=0 $Y2=0
cc_169 N_A_c_187_n N_A_214_47#_c_386_n 0.00173681f $X=3.12 $Y=1.202 $X2=0 $Y2=0
cc_170 N_VPWR_c_225_n N_A_235_309#_M1001_s 0.00425811f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_171 N_VPWR_c_225_n N_A_235_309#_M1009_s 0.00662844f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_172 N_VPWR_c_225_n N_A_235_309#_M1007_d 0.00217523f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_173 N_VPWR_c_226_n N_A_235_309#_c_272_n 0.0234767f $X=0.73 $Y=2.34 $X2=0
+ $Y2=0
cc_174 N_VPWR_c_227_n N_A_235_309#_c_272_n 0.0167762f $X=1.605 $Y=2.72 $X2=0
+ $Y2=0
cc_175 N_VPWR_c_228_n N_A_235_309#_c_272_n 0.0354158f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_176 N_VPWR_c_225_n N_A_235_309#_c_272_n 0.0091658f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_177 N_VPWR_M1001_d N_A_235_309#_c_281_n 0.0036863f $X=1.625 $Y=1.545 $X2=0
+ $Y2=0
cc_178 N_VPWR_c_228_n N_A_235_309#_c_281_n 0.0171295f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_228_n N_A_235_309#_c_287_n 0.0219309f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_230_n N_A_235_309#_c_274_n 0.0693025f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_c_225_n N_A_235_309#_c_274_n 0.0423961f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_228_n N_A_235_309#_c_307_n 0.0104344f $X=1.77 $Y=2.02 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_230_n N_A_235_309#_c_307_n 0.0119545f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_225_n N_A_235_309#_c_307_n 0.006547f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_185 N_VPWR_c_225_n N_Z_M1003_s 0.00232895f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_186 N_A_235_309#_c_274_n N_Z_M1003_s 0.00352392f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_187 N_A_235_309#_c_281_n N_Z_c_315_n 0.00948638f $X=2.185 $Y=1.64 $X2=0 $Y2=0
cc_188 N_A_235_309#_c_287_n N_Z_c_315_n 0.0199782f $X=2.27 $Y=1.96 $X2=0 $Y2=0
cc_189 N_A_235_309#_c_274_n N_Z_c_315_n 0.0231793f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_190 N_A_235_309#_c_275_n N_Z_c_315_n 0.0266244f $X=3.33 $Y=1.96 $X2=0 $Y2=0
cc_191 N_Z_M1000_d N_VGND_c_338_n 0.00297142f $X=2.675 $Y=0.235 $X2=1.92
+ $Y2=1.16
cc_192 N_Z_M1000_d N_A_214_47#_c_386_n 0.00503152f $X=2.675 $Y=0.235 $X2=0 $Y2=0
cc_193 N_Z_c_315_n N_A_214_47#_c_386_n 0.0235686f $X=2.86 $Y=0.76 $X2=0 $Y2=0
cc_194 N_VGND_c_338_n N_A_214_47#_M1004_s 0.00539683f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_195 N_VGND_c_338_n N_A_214_47#_M1000_s 0.00288008f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_338_n N_A_214_47#_M1006_s 0.00208521f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_197 N_VGND_c_336_n N_A_214_47#_c_388_n 0.0131946f $X=1.51 $Y=0 $X2=0 $Y2=0
cc_198 N_VGND_c_338_n N_A_214_47#_c_388_n 0.00739874f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_339_n N_A_214_47#_c_388_n 0.0143054f $X=0.69 $Y=0 $X2=0 $Y2=0
cc_200 N_VGND_M1005_d N_A_214_47#_c_384_n 0.00579475f $X=1.54 $Y=0.235 $X2=0
+ $Y2=0
cc_201 N_VGND_c_334_n N_A_214_47#_c_384_n 0.0238049f $X=1.695 $Y=0.38 $X2=0
+ $Y2=0
cc_202 N_VGND_c_336_n N_A_214_47#_c_384_n 0.00232396f $X=1.51 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_c_337_n N_A_214_47#_c_384_n 0.00453887f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_204 N_VGND_c_338_n N_A_214_47#_c_384_n 0.0130142f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_205 N_VGND_c_334_n N_A_214_47#_c_385_n 0.00372297f $X=1.695 $Y=0.38 $X2=0
+ $Y2=0
cc_206 N_VGND_c_337_n N_A_214_47#_c_386_n 0.0610419f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_338_n N_A_214_47#_c_386_n 0.0379531f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_334_n N_A_214_47#_c_387_n 0.0112643f $X=1.695 $Y=0.38 $X2=0
+ $Y2=0
cc_209 N_VGND_c_337_n N_A_214_47#_c_387_n 0.0230581f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_338_n N_A_214_47#_c_387_n 0.0128424f $X=3.45 $Y=0 $X2=0 $Y2=0
