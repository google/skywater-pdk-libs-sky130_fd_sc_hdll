* File: sky130_fd_sc_hdll__nand4b_2.pxi.spice
* Created: Wed Sep  2 08:38:45 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%A_N N_A_N_c_90_n N_A_N_c_91_n N_A_N_M1000_g
+ N_A_N_M1011_g A_N A_N N_A_N_c_89_n PM_SKY130_FD_SC_HDLL__NAND4B_2%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%A_27_47# N_A_27_47#_M1011_s N_A_27_47#_M1000_s
+ N_A_27_47#_c_127_n N_A_27_47#_M1009_g N_A_27_47#_c_118_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_128_n N_A_27_47#_M1016_g N_A_27_47#_c_119_n N_A_27_47#_M1014_g
+ N_A_27_47#_c_120_n N_A_27_47#_c_121_n N_A_27_47#_c_122_n N_A_27_47#_c_131_n
+ N_A_27_47#_c_123_n N_A_27_47#_c_124_n N_A_27_47#_c_125_n N_A_27_47#_c_126_n
+ N_A_27_47#_c_146_n PM_SKY130_FD_SC_HDLL__NAND4B_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%B N_B_c_207_n N_B_M1008_g N_B_c_211_n
+ N_B_M1001_g N_B_c_208_n N_B_M1010_g N_B_c_212_n N_B_M1006_g B B N_B_c_209_n
+ N_B_c_210_n B B PM_SKY130_FD_SC_HDLL__NAND4B_2%B
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%C N_C_c_260_n N_C_M1012_g N_C_c_256_n
+ N_C_M1005_g N_C_c_261_n N_C_M1017_g N_C_c_257_n N_C_M1015_g C C N_C_c_258_n C
+ C PM_SKY130_FD_SC_HDLL__NAND4B_2%C
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%D N_D_c_308_n N_D_M1003_g N_D_c_303_n
+ N_D_M1002_g N_D_c_309_n N_D_M1013_g N_D_c_304_n N_D_M1007_g N_D_c_305_n D D
+ N_D_c_307_n D D PM_SKY130_FD_SC_HDLL__NAND4B_2%D
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%VPWR N_VPWR_M1000_d N_VPWR_M1009_d
+ N_VPWR_M1016_d N_VPWR_M1006_d N_VPWR_M1017_d N_VPWR_M1013_d N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_356_n N_VPWR_c_357_n N_VPWR_c_358_n N_VPWR_c_359_n
+ N_VPWR_c_360_n N_VPWR_c_361_n VPWR N_VPWR_c_362_n N_VPWR_c_363_n
+ N_VPWR_c_364_n N_VPWR_c_365_n N_VPWR_c_348_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%Y N_Y_M1004_s N_Y_M1009_s N_Y_M1001_s
+ N_Y_M1012_s N_Y_M1003_s N_Y_c_445_n N_Y_c_440_n N_Y_c_449_n N_Y_c_441_n
+ N_Y_c_476_n N_Y_c_442_n N_Y_c_481_n N_Y_c_443_n N_Y_c_444_n Y Y Y N_Y_c_439_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%VGND N_VGND_M1011_d N_VGND_M1002_s
+ N_VGND_c_531_n N_VGND_c_532_n N_VGND_c_533_n VGND N_VGND_c_534_n
+ N_VGND_c_535_n N_VGND_c_536_n N_VGND_c_537_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_2%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%A_225_47# N_A_225_47#_M1004_d
+ N_A_225_47#_M1014_d N_A_225_47#_M1010_d N_A_225_47#_c_601_n
+ N_A_225_47#_c_602_n N_A_225_47#_c_611_n N_A_225_47#_c_603_n
+ N_A_225_47#_c_604_n PM_SKY130_FD_SC_HDLL__NAND4B_2%A_225_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%A_495_47# N_A_495_47#_M1008_s
+ N_A_495_47#_M1005_s N_A_495_47#_c_641_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_2%A_495_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_2%A_705_47# N_A_705_47#_M1005_d
+ N_A_705_47#_M1015_d N_A_705_47#_M1007_d N_A_705_47#_c_656_n
+ N_A_705_47#_c_667_n N_A_705_47#_c_657_n N_A_705_47#_c_658_n
+ N_A_705_47#_c_659_n PM_SKY130_FD_SC_HDLL__NAND4B_2%A_705_47#
cc_1 VNB N_A_N_M1011_g 0.043001f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.0134299f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_89_n 0.0395036f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_47#_c_118_n 0.0214729f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_27_47#_c_119_n 0.0166801f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_A_27_47#_c_120_n 0.0303277f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_7 VNB N_A_27_47#_c_121_n 0.0337477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_122_n 0.0147647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_123_n 0.0128299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_124_n 0.005642f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_125_n 6.40756e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_126_n 0.0166484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B_c_207_n 0.0164932f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_14 VNB N_B_c_208_n 0.0219752f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB N_B_c_209_n 0.0540351f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B_c_210_n 0.007669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C_c_256_n 0.0219752f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_18 VNB N_C_c_257_n 0.017682f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_19 VNB N_C_c_258_n 0.0457322f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=1.16
cc_20 VNB C 0.00770495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D_c_303_n 0.017682f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_22 VNB N_D_c_304_n 0.0219568f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_23 VNB N_D_c_305_n 0.0346998f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB D 0.00934205f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_25 VNB N_D_c_307_n 0.0347951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_348_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_Y_c_439_n 0.00101052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_531_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_532_n 0.0981619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_533_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_534_n 0.0143533f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_32 VNB N_VGND_c_535_n 0.0217464f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_536_n 0.310358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_537_n 0.0114568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_225_47#_c_601_n 0.00217944f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_36 VNB N_A_225_47#_c_602_n 0.00709211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_225_47#_c_603_n 0.00208278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_225_47#_c_604_n 0.00789203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_495_47#_c_641_n 0.0103416f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_40 VNB N_A_705_47#_c_656_n 0.00928571f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_41 VNB N_A_705_47#_c_657_n 0.0129041f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_42 VNB N_A_705_47#_c_658_n 0.0182049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_705_47#_c_659_n 0.00311367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_A_N_c_90_n 0.0476969f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_45 VPB N_A_N_c_91_n 0.0307843f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_46 VPB A_N 0.01652f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_47 VPB N_A_N_c_89_n 0.0103641f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_48 VPB N_A_27_47#_c_127_n 0.0191558f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_49 VPB N_A_27_47#_c_128_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_47#_c_120_n 0.0138206f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_51 VPB N_A_27_47#_c_121_n 0.021023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_131_n 0.0147827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_125_n 0.0198647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_B_c_211_n 0.0159796f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_55 VPB N_B_c_212_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_56 VPB N_B_c_209_n 0.0294897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_C_c_260_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_58 VPB N_C_c_261_n 0.0166564f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_59 VPB N_C_c_258_n 0.0263403f $X=-0.19 $Y=1.305 $X2=0.21 $Y2=1.16
cc_60 VPB N_D_c_308_n 0.0166564f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_61 VPB N_D_c_309_n 0.0209048f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_62 VPB N_D_c_305_n 0.0250596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_D_c_307_n 0.0109325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_349_n 0.0182684f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_65 VPB N_VPWR_c_350_n 0.00419147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_351_n 0.0115785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_352_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_353_n 0.0073282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_354_n 0.0052064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_355_n 0.0129627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_356_n 0.0455717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_357_n 0.0143307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_358_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_359_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_360_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_361_n 0.00497181f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_362_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_363_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_364_n 0.00842476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_365_n 0.012281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_348_n 0.0439966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_Y_c_440_n 0.00427918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_Y_c_441_n 0.0107683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_Y_c_442_n 0.00541418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_Y_c_443_n 0.00174301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_Y_c_444_n 0.00174301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 N_A_N_c_89_n N_A_27_47#_c_120_n 0.00900735f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_N_M1011_g N_A_27_47#_c_122_n 0.00425747f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_89 N_A_N_c_91_n N_A_27_47#_c_131_n 0.00449618f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_90 N_A_N_M1011_g N_A_27_47#_c_123_n 0.0141536f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_91 A_N N_A_27_47#_c_123_n 0.0174382f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_92 N_A_N_c_89_n N_A_27_47#_c_123_n 0.00596468f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_N_M1011_g N_A_27_47#_c_124_n 0.0123902f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_94 A_N N_A_27_47#_c_124_n 0.0056444f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_N_c_89_n N_A_27_47#_c_124_n 0.00253733f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_N_c_90_n N_A_27_47#_c_125_n 0.0274287f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_97 N_A_N_c_91_n N_A_27_47#_c_125_n 0.0198703f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_98 A_N N_A_27_47#_c_125_n 0.0407621f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_99 N_A_N_c_89_n N_A_27_47#_c_125_n 0.00494816f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_100 A_N N_A_27_47#_c_146_n 0.0132649f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A_N_c_89_n N_A_27_47#_c_146_n 0.0066797f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A_N_c_91_n N_VPWR_c_350_n 0.0126512f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_103 N_A_N_c_90_n N_VPWR_c_351_n 0.002358f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_104 N_A_N_c_91_n N_VPWR_c_351_n 0.00387233f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_105 N_A_N_c_91_n N_VPWR_c_357_n 0.00314304f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_106 N_A_N_c_91_n N_VPWR_c_348_n 0.00460683f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_107 N_A_N_M1011_g N_VGND_c_534_n 0.00198377f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_N_M1011_g N_VGND_c_536_n 0.00358947f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_N_M1011_g N_VGND_c_537_n 0.0123528f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_N_M1011_g N_A_225_47#_c_602_n 0.00438858f $X=0.52 $Y=0.445 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_119_n N_B_c_207_n 0.0223336f $X=1.98 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_27_47#_c_128_n N_B_c_211_n 0.0229911f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_121_n N_B_c_209_n 0.0223336f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_114 N_A_27_47#_c_121_n N_B_c_210_n 0.00210845f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_125_n N_VPWR_M1000_d 0.00107505f $X=0.61 $Y=1.915 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_27_47#_c_131_n N_VPWR_c_350_n 0.0169042f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_125_n N_VPWR_c_350_n 0.0108491f $X=0.61 $Y=1.915 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_127_n N_VPWR_c_351_n 0.00322167f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_27_47#_c_120_n N_VPWR_c_351_n 0.0062725f $X=1.385 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_125_n N_VPWR_c_351_n 0.0303972f $X=0.61 $Y=1.915 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_126_n N_VPWR_c_351_n 0.0177163f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_128_n N_VPWR_c_352_n 0.0052072f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_131_n N_VPWR_c_357_n 0.017116f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_125_n N_VPWR_c_357_n 0.00242775f $X=0.61 $Y=1.915 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_127_n N_VPWR_c_358_n 0.00597712f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_c_128_n N_VPWR_c_358_n 0.00673617f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_127_n N_VPWR_c_364_n 0.00606518f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_M1000_s N_VPWR_c_348_n 0.00239406f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_127_n N_VPWR_c_348_n 0.0112745f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_128_n N_VPWR_c_348_n 0.011869f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_131_n N_VPWR_c_348_n 0.00960198f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_125_n N_VPWR_c_348_n 0.00516589f $X=0.61 $Y=1.915 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_127_n N_Y_c_445_n 0.0121625f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_128_n N_Y_c_445_n 0.0106251f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_128_n N_Y_c_440_n 0.020382f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_121_n N_Y_c_440_n 4.93319e-19 $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_128_n N_Y_c_449_n 6.48386e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_127_n Y 0.00368288f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_128_n Y 8.77306e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_127_n N_Y_c_439_n 0.00199531f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_118_n N_Y_c_439_n 0.0105292f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_128_n N_Y_c_439_n 0.00103355f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_27_47#_c_119_n N_Y_c_439_n 0.00285271f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_121_n N_Y_c_439_n 0.0440368f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_126_n N_Y_c_439_n 0.0135488f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_123_n N_VGND_M1011_d 9.98338e-19 $X=0.61 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_27_47#_c_118_n N_VGND_c_532_n 0.00357877f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_119_n N_VGND_c_532_n 0.00357877f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_122_n N_VGND_c_534_n 0.017116f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_123_n N_VGND_c_534_n 0.00249162f $X=0.61 $Y=0.805 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1011_s N_VGND_c_536_n 0.00289329f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_118_n N_VGND_c_536_n 0.00668309f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_119_n N_VGND_c_536_n 0.00542415f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_122_n N_VGND_c_536_n 0.00960198f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_123_n N_VGND_c_536_n 0.00539505f $X=0.61 $Y=0.805 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_118_n N_VGND_c_537_n 0.00218593f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_122_n N_VGND_c_537_n 0.0161551f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_123_n N_VGND_c_537_n 0.0107888f $X=0.61 $Y=0.805 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_126_n N_VGND_c_537_n 0.00565372f $X=1.17 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_118_n N_A_225_47#_c_602_n 0.00456666f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_120_n N_A_225_47#_c_602_n 0.00634711f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_123_n N_A_225_47#_c_602_n 0.00848415f $X=0.61 $Y=0.805 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_124_n N_A_225_47#_c_602_n 0.00466249f $X=0.61 $Y=1.075 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_126_n N_A_225_47#_c_602_n 0.0199291f $X=1.17 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_118_n N_A_225_47#_c_611_n 0.0111679f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_119_n N_A_225_47#_c_611_n 0.0146117f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_120_n N_A_225_47#_c_611_n 0.00201482f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_121_n N_A_225_47#_c_611_n 4.68623e-19 $X=1.955 $Y=1.202
+ $X2=0 $Y2=0
cc_169 N_A_27_47#_c_119_n N_A_225_47#_c_603_n 7.54024e-19 $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_B_c_209_n N_C_c_258_n 0.0100132f $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_171 N_B_c_210_n N_C_c_258_n 7.3417e-19 $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_172 N_B_c_209_n C 8.19518e-19 $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_173 N_B_c_210_n C 0.0137573f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B_c_211_n N_VPWR_c_352_n 0.004751f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B_c_212_n N_VPWR_c_353_n 0.00817046f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_211_n N_VPWR_c_362_n 0.00597712f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B_c_212_n N_VPWR_c_362_n 0.00673617f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B_c_211_n N_VPWR_c_348_n 0.0100198f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_212_n N_VPWR_c_348_n 0.0131262f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_211_n N_Y_c_445_n 6.24674e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B_c_211_n N_Y_c_440_n 0.0113403f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B_c_209_n N_Y_c_440_n 3.10838e-19 $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_183 N_B_c_210_n N_Y_c_440_n 0.0212327f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B_c_211_n N_Y_c_449_n 0.0130707f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B_c_212_n N_Y_c_449_n 0.0153658f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_212_n N_Y_c_441_n 0.0179883f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_209_n N_Y_c_441_n 0.00709775f $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_188 N_B_c_210_n N_Y_c_441_n 0.0384032f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B_c_211_n N_Y_c_443_n 0.00292783f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_212_n N_Y_c_443_n 0.00116723f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_209_n N_Y_c_443_n 0.00786476f $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_192 N_B_c_210_n N_Y_c_443_n 0.0305798f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B_c_209_n N_Y_c_439_n 0.00125414f $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_194 N_B_c_210_n N_Y_c_439_n 0.0117738f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_195 N_B_c_207_n N_VGND_c_532_n 0.00411651f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B_c_208_n N_VGND_c_532_n 0.00357877f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_197 N_B_c_207_n N_VGND_c_536_n 0.00587071f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_198 N_B_c_208_n N_VGND_c_536_n 0.00672921f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B_c_210_n N_A_225_47#_c_603_n 0.00978542f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_207_n N_A_225_47#_c_604_n 0.0139704f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B_c_208_n N_A_225_47#_c_604_n 0.0117754f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B_c_209_n N_A_225_47#_c_604_n 0.0120291f $X=2.895 $Y=1.202 $X2=0 $Y2=0
cc_203 N_B_c_210_n N_A_225_47#_c_604_n 0.0756367f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_204 N_B_c_207_n N_A_495_47#_c_641_n 0.0028244f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_205 N_B_c_208_n N_A_495_47#_c_641_n 0.0112708f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_206 N_B_c_210_n N_A_495_47#_c_641_n 0.00175186f $X=3.115 $Y=1.16 $X2=0 $Y2=0
cc_207 N_B_c_208_n N_A_705_47#_c_656_n 4.99491e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_208 N_C_c_261_n N_D_c_308_n 0.0245765f $X=4.305 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_209 N_C_c_257_n N_D_c_303_n 0.0151684f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_210 N_C_c_258_n N_D_c_305_n 0.0276547f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_211 C N_D_c_305_n 0.00220274f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_212 C D 0.010601f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_213 N_C_c_260_n N_VPWR_c_353_n 0.0204445f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_214 N_C_c_261_n N_VPWR_c_354_n 0.00571162f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_215 N_C_c_260_n N_VPWR_c_360_n 0.00597712f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_216 N_C_c_261_n N_VPWR_c_360_n 0.00673617f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_217 N_C_c_260_n N_VPWR_c_348_n 0.0114039f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_218 N_C_c_261_n N_VPWR_c_348_n 0.0120675f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_219 N_C_c_260_n N_Y_c_441_n 0.0139912f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_220 N_C_c_258_n N_Y_c_441_n 2.7776e-19 $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_221 C N_Y_c_441_n 0.0181228f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_222 N_C_c_260_n N_Y_c_476_n 0.0178402f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_223 N_C_c_261_n N_Y_c_476_n 0.011049f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_224 N_C_c_261_n N_Y_c_442_n 0.0159401f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_225 N_C_c_258_n N_Y_c_442_n 0.00410828f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_226 C N_Y_c_442_n 0.0330941f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_227 N_C_c_261_n N_Y_c_481_n 6.27779e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_228 N_C_c_260_n N_Y_c_444_n 0.00292783f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_229 N_C_c_261_n N_Y_c_444_n 0.00116723f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_230 N_C_c_258_n N_Y_c_444_n 0.00787329f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_231 C N_Y_c_444_n 0.0305798f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_232 N_C_c_256_n N_VGND_c_532_n 0.00357877f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_233 N_C_c_257_n N_VGND_c_532_n 0.00425094f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_234 N_C_c_256_n N_VGND_c_536_n 0.00672921f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_235 N_C_c_257_n N_VGND_c_536_n 0.00625093f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_236 N_C_c_256_n N_A_225_47#_c_604_n 4.99491e-19 $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_237 N_C_c_256_n N_A_495_47#_c_641_n 0.0112708f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_238 N_C_c_256_n N_A_705_47#_c_656_n 0.0118634f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_239 N_C_c_257_n N_A_705_47#_c_656_n 0.0131204f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_240 N_C_c_258_n N_A_705_47#_c_656_n 0.0076395f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_241 C N_A_705_47#_c_656_n 0.0664799f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_242 N_C_c_258_n N_A_705_47#_c_659_n 0.00127974f $X=4.32 $Y=1.16 $X2=0 $Y2=0
cc_243 C N_A_705_47#_c_659_n 0.0151232f $X=4.365 $Y=1.19 $X2=0 $Y2=0
cc_244 N_D_c_308_n N_VPWR_c_354_n 0.00887722f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_245 N_D_c_309_n N_VPWR_c_356_n 0.0287414f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_246 D N_VPWR_c_356_n 0.02587f $X=5.65 $Y=1.105 $X2=0 $Y2=0
cc_247 N_D_c_307_n N_VPWR_c_356_n 0.00901782f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_248 N_D_c_308_n N_VPWR_c_363_n 0.00597712f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_249 N_D_c_309_n N_VPWR_c_363_n 0.00673617f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_250 N_D_c_308_n N_VPWR_c_348_n 0.0103045f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_251 N_D_c_309_n N_VPWR_c_348_n 0.0129848f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_252 N_D_c_308_n N_Y_c_476_n 6.74229e-19 $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_253 N_D_c_308_n N_Y_c_442_n 0.0190774f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_254 N_D_c_309_n N_Y_c_442_n 0.00747728f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_255 N_D_c_305_n N_Y_c_442_n 0.00859303f $X=5.485 $Y=1.16 $X2=0 $Y2=0
cc_256 D N_Y_c_442_n 0.0198871f $X=5.65 $Y=1.105 $X2=0 $Y2=0
cc_257 N_D_c_308_n N_Y_c_481_n 0.0151968f $X=4.865 $Y=1.41 $X2=0 $Y2=0
cc_258 N_D_c_309_n N_Y_c_481_n 0.0117384f $X=5.335 $Y=1.41 $X2=0 $Y2=0
cc_259 N_D_c_303_n N_VGND_c_531_n 0.00276126f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_260 N_D_c_304_n N_VGND_c_531_n 0.00376026f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_261 N_D_c_303_n N_VGND_c_532_n 0.00436487f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_262 N_D_c_304_n N_VGND_c_535_n 0.00422241f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_263 N_D_c_303_n N_VGND_c_536_n 0.00637915f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_264 N_D_c_304_n N_VGND_c_536_n 0.00698354f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_265 N_D_c_303_n N_A_705_47#_c_667_n 0.00469081f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_266 N_D_c_303_n N_A_705_47#_c_657_n 0.0155486f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_267 N_D_c_304_n N_A_705_47#_c_657_n 0.0105603f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_268 N_D_c_305_n N_A_705_47#_c_657_n 0.0054776f $X=5.485 $Y=1.16 $X2=0 $Y2=0
cc_269 D N_A_705_47#_c_657_n 0.0583175f $X=5.65 $Y=1.105 $X2=0 $Y2=0
cc_270 N_D_c_307_n N_A_705_47#_c_657_n 0.00778392f $X=5.695 $Y=1.16 $X2=0 $Y2=0
cc_271 N_D_c_303_n N_A_705_47#_c_658_n 6.77769e-19 $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_272 N_D_c_304_n N_A_705_47#_c_658_n 0.00693801f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_273 N_D_c_303_n N_A_705_47#_c_659_n 0.00172732f $X=4.94 $Y=0.995 $X2=0 $Y2=0
cc_274 N_D_c_305_n N_A_705_47#_c_659_n 0.00134197f $X=5.485 $Y=1.16 $X2=0 $Y2=0
cc_275 N_VPWR_c_348_n N_Y_M1009_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_276 N_VPWR_c_348_n N_Y_M1001_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_348_n N_Y_M1012_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_348_n N_Y_M1003_s 0.00231261f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_351_n N_Y_c_445_n 0.0452437f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_280 N_VPWR_c_352_n N_Y_c_445_n 0.0385613f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_281 N_VPWR_c_358_n N_Y_c_445_n 0.0223557f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_364_n N_Y_c_445_n 0.0175144f $X=1.15 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_348_n N_Y_c_445_n 0.0140101f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_M1016_d N_Y_c_440_n 0.00180012f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_285 N_VPWR_c_352_n N_Y_c_440_n 0.0139097f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_286 N_VPWR_c_352_n N_Y_c_449_n 0.0470327f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_287 N_VPWR_c_353_n N_Y_c_449_n 0.0426988f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_288 N_VPWR_c_362_n N_Y_c_449_n 0.0223557f $X=3.045 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_348_n N_Y_c_449_n 0.0140101f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_M1006_d N_Y_c_441_n 0.0107993f $X=2.985 $Y=1.485 $X2=0 $Y2=0
cc_291 N_VPWR_c_353_n N_Y_c_441_n 0.0528236f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_292 N_VPWR_c_353_n N_Y_c_476_n 0.0520395f $X=3.52 $Y=2 $X2=0 $Y2=0
cc_293 N_VPWR_c_354_n N_Y_c_476_n 0.0398033f $X=4.575 $Y=2 $X2=0 $Y2=0
cc_294 N_VPWR_c_360_n N_Y_c_476_n 0.0223557f $X=4.455 $Y=2.72 $X2=0 $Y2=0
cc_295 N_VPWR_c_348_n N_Y_c_476_n 0.0140101f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_296 N_VPWR_M1017_d N_Y_c_442_n 0.00296263f $X=4.395 $Y=1.485 $X2=0 $Y2=0
cc_297 N_VPWR_c_354_n N_Y_c_442_n 0.0213613f $X=4.575 $Y=2 $X2=0 $Y2=0
cc_298 N_VPWR_c_356_n N_Y_c_442_n 0.011627f $X=5.65 $Y=1.66 $X2=0 $Y2=0
cc_299 N_VPWR_c_354_n N_Y_c_481_n 0.0485357f $X=4.575 $Y=2 $X2=0 $Y2=0
cc_300 N_VPWR_c_356_n N_Y_c_481_n 0.0521605f $X=5.65 $Y=1.66 $X2=0 $Y2=0
cc_301 N_VPWR_c_363_n N_Y_c_481_n 0.0223557f $X=5.485 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_348_n N_Y_c_481_n 0.0140101f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_303 N_VPWR_c_351_n Y 0.0178254f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_304 N_Y_M1004_s N_VGND_c_536_n 0.00256987f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_305 N_Y_c_439_n N_A_225_47#_c_602_n 0.0207685f $X=1.72 $Y=0.72 $X2=0 $Y2=0
cc_306 N_Y_M1004_s N_A_225_47#_c_611_n 0.00399738f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_307 N_Y_c_439_n N_A_225_47#_c_611_n 0.0218008f $X=1.72 $Y=0.72 $X2=0 $Y2=0
cc_308 N_Y_c_440_n N_A_225_47#_c_603_n 0.00210886f $X=2.445 $Y=1.555 $X2=0 $Y2=0
cc_309 N_Y_c_439_n N_A_225_47#_c_603_n 0.00141443f $X=1.72 $Y=0.72 $X2=0 $Y2=0
cc_310 N_Y_c_441_n N_A_705_47#_c_656_n 0.00446358f $X=3.855 $Y=1.555 $X2=0 $Y2=0
cc_311 N_Y_c_442_n N_A_705_47#_c_657_n 0.00665764f $X=4.885 $Y=1.555 $X2=0 $Y2=0
cc_312 N_Y_c_442_n N_A_705_47#_c_659_n 0.00437829f $X=4.885 $Y=1.555 $X2=0 $Y2=0
cc_313 N_VGND_c_536_n N_A_225_47#_M1004_d 0.00250318f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_314 N_VGND_c_536_n N_A_225_47#_M1014_d 0.00235053f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_536_n N_A_225_47#_M1010_d 0.00251142f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_316 N_VGND_c_532_n N_A_225_47#_c_601_n 0.017577f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_536_n N_A_225_47#_c_601_n 0.00961661f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_c_537_n N_A_225_47#_c_601_n 0.0173456f $X=0.69 $Y=0 $X2=0 $Y2=0
cc_319 N_VGND_c_532_n N_A_225_47#_c_611_n 0.0538938f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_320 N_VGND_c_536_n N_A_225_47#_c_611_n 0.033904f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_532_n N_A_225_47#_c_604_n 0.00250396f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_536_n N_A_225_47#_c_604_n 0.00602355f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_536_n N_A_495_47#_M1008_s 0.00255381f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_324 N_VGND_c_536_n N_A_495_47#_M1005_s 0.00262311f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_325 N_VGND_c_532_n N_A_495_47#_c_641_n 0.108539f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_536_n N_A_495_47#_c_641_n 0.0671299f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_536_n N_A_705_47#_M1005_d 0.00251142f $X=5.75 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_328 N_VGND_c_536_n N_A_705_47#_M1015_d 0.00387859f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_329 N_VGND_c_536_n N_A_705_47#_M1007_d 0.00209319f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_330 N_VGND_c_532_n N_A_705_47#_c_656_n 0.0032051f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_331 N_VGND_c_536_n N_A_705_47#_c_656_n 0.00713708f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_332 N_VGND_c_532_n N_A_705_47#_c_667_n 0.0178751f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_333 N_VGND_c_536_n N_A_705_47#_c_667_n 0.00992425f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_334 N_VGND_M1002_s N_A_705_47#_c_657_n 0.0025045f $X=5.015 $Y=0.235 $X2=0
+ $Y2=0
cc_335 N_VGND_c_531_n N_A_705_47#_c_657_n 0.0127393f $X=5.15 $Y=0.38 $X2=0 $Y2=0
cc_336 N_VGND_c_532_n N_A_705_47#_c_657_n 0.00293397f $X=5.065 $Y=0 $X2=0 $Y2=0
cc_337 N_VGND_c_535_n N_A_705_47#_c_657_n 0.00273345f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_338 N_VGND_c_536_n N_A_705_47#_c_657_n 0.0120844f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_339 N_VGND_c_531_n N_A_705_47#_c_658_n 0.0175778f $X=5.15 $Y=0.38 $X2=0 $Y2=0
cc_340 N_VGND_c_535_n N_A_705_47#_c_658_n 0.0213324f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_341 N_VGND_c_536_n N_A_705_47#_c_658_n 0.0126042f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_342 N_VGND_c_532_n N_A_705_47#_c_659_n 7.60802e-19 $X=5.065 $Y=0 $X2=0 $Y2=0
cc_343 N_VGND_c_536_n N_A_705_47#_c_659_n 0.00117665f $X=5.75 $Y=0 $X2=0 $Y2=0
cc_344 N_A_225_47#_c_604_n N_A_495_47#_M1008_s 0.00214196f $X=3.13 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_345 N_A_225_47#_M1010_d N_A_495_47#_c_641_n 0.00632239f $X=2.945 $Y=0.235
+ $X2=0 $Y2=0
cc_346 N_A_225_47#_c_604_n N_A_495_47#_c_641_n 0.048335f $X=3.13 $Y=0.72 $X2=0
+ $Y2=0
cc_347 N_A_225_47#_c_604_n N_A_705_47#_c_656_n 0.0231991f $X=3.13 $Y=0.72 $X2=0
+ $Y2=0
cc_348 N_A_495_47#_c_641_n N_A_705_47#_M1005_d 0.00655451f $X=4.12 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_349 N_A_495_47#_M1005_s N_A_705_47#_c_656_n 0.00214196f $X=3.985 $Y=0.235
+ $X2=0 $Y2=0
cc_350 N_A_495_47#_c_641_n N_A_705_47#_c_656_n 0.0463395f $X=4.12 $Y=0.38 $X2=0
+ $Y2=0
