* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfstp_4 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q
X0 a_1663_329# a_693_369# a_1745_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X1 VGND a_693_369# a_877_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 a_27_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X3 a_119_47# SCE a_201_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 Q a_2447_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_2447_47# a_1745_329# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND a_2447_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR a_1075_413# a_1663_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X8 a_1075_413# a_877_369# a_1177_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_2067_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X10 VGND a_2447_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_201_47# a_349_21# a_27_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X12 a_2447_47# a_1745_329# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_211_369# D a_201_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X14 a_349_21# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X15 a_1075_413# a_693_369# a_1169_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X16 a_693_369# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND a_1745_329# a_1951_295# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_201_47# a_877_369# a_1075_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X19 a_349_21# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1229_21# a_1075_413# a_1467_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1169_413# a_1229_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X22 a_201_47# a_693_369# a_1075_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 Q a_2447_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR SCE a_211_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X25 a_1745_329# a_877_369# a_1891_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X26 VPWR a_1745_329# a_1951_295# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X27 VGND SCD a_119_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 VPWR a_2447_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VPWR a_693_369# a_877_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X30 VPWR a_1075_413# a_1229_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X31 a_295_47# a_349_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X32 a_1177_47# a_1229_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X33 a_1654_47# a_877_369# a_1745_329# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X34 a_1891_413# a_1951_295# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X35 a_693_369# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X36 a_201_47# D a_295_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X37 a_1229_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X38 a_1745_329# a_693_369# a_1995_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X39 VGND a_1075_413# a_1654_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X40 Q a_2447_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 a_1467_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 Q a_2447_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 VPWR SET_B a_1745_329# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X44 a_1995_47# a_1951_295# a_2067_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X45 VPWR a_2447_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
