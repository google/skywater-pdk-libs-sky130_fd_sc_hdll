* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__ebufn_2 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR A a_27_47# VPB phighvt w=640000u l=180000u
+  ad=5.254e+11p pd=4.53e+06u as=1.728e+11p ps=1.82e+06u
M1001 VGND a_224_47# a_412_47# VNB nshort w=650000u l=150000u
+  ad=3.54e+11p pd=3.53e+06u as=6.8575e+11p ps=6.01e+06u
M1002 a_224_47# TE_B VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1003 a_340_309# a_27_47# Z VPB phighvt w=1e+06u l=180000u
+  ad=1.3537e+12p pd=8.63e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_412_47# a_224_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_412_47# a_27_47# Z VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1006 a_224_47# TE_B VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_340_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR TE_B a_340_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Z a_27_47# a_340_309# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
M1011 Z a_27_47# a_412_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
