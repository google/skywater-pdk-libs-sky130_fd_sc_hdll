* File: sky130_fd_sc_hdll__conb_1.pex.spice
* Created: Wed Sep  2 08:27:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CONB_1%HI 1 3 5 6
r16 5 6 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.44 $Y=0.34
+ $X2=0.44 $Y2=0.34
r17 3 5 91.4009 $w=4.8e-07 $l=8.2e-07 $layer=POLY_cond $X=0.345 $Y=1.16
+ $X2=0.345 $Y2=0.34
r18 1 6 20.0113 $w=5.18e-07 $l=8.7e-07 $layer=LI1_cond $X=0.345 $Y=1.21
+ $X2=0.345 $Y2=0.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__CONB_1%VPWR 3 4 7 8 9 11 18 19
r18 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r19 9 19 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r20 9 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
r21 7 15 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.275 $Y=2.72 $X2=0.23
+ $Y2=2.72
r22 7 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.275 $Y=2.72 $X2=0.44
+ $Y2=2.72
r23 6 18 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 6 8 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.605 $Y=2.72 $X2=0.44
+ $Y2=2.72
r25 4 11 88.0569 $w=4.8e-07 $l=7.9e-07 $layer=POLY_cond $X=0.345 $Y=1.995
+ $X2=0.345 $Y2=1.205
r26 3 4 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.44 $Y=1.995
+ $X2=0.44 $Y2=1.995
r27 1 8 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.44 $Y=2.635 $X2=0.44
+ $Y2=2.72
r28 1 3 22.3504 $w=3.28e-07 $l=6.4e-07 $layer=LI1_cond $X=0.44 $Y=2.635 $X2=0.44
+ $Y2=1.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__CONB_1%VGND 1 3 4 6 8 11 18
r15 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r16 14 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r17 13 14 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r18 11 17 4.56849 $w=1.7e-07 $l=3.02e-07 $layer=LI1_cond $X=0.775 $Y=0 $X2=1.077
+ $Y2=0
r19 11 13 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0 $X2=0.69
+ $Y2=0
r20 6 14 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r21 4 8 93.6302 $w=4.8e-07 $l=8.4e-07 $layer=POLY_cond $X=1.035 $Y=0.32
+ $X2=1.035 $Y2=1.16
r22 3 4 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94 $Y=0.32
+ $X2=0.94 $Y2=0.32
r23 1 17 3.28266 $w=3.4e-07 $l=1.69245e-07 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=1.077 $Y2=0
r24 1 3 7.96542 $w=3.38e-07 $l=2.35e-07 $layer=LI1_cond $X=0.945 $Y=0.085
+ $X2=0.945 $Y2=0.32
.ends

.subckt PM_SKY130_FD_SC_HDLL__CONB_1%LO 1 3 5
r17 5 6 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.94 $Y=1.995
+ $X2=0.94 $Y2=1.995
r18 3 5 88.0569 $w=4.8e-07 $l=7.9e-07 $layer=POLY_cond $X=1.035 $Y=1.205
+ $X2=1.035 $Y2=1.995
r19 1 6 10.6957 $w=5.18e-07 $l=4.65e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=1.035 $Y2=1.995
.ends

