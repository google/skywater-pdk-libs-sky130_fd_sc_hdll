# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb8to1_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.915000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.525000 1.055000 6.345000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.535000 1.055000 7.355000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.965000 1.055000 12.785000 1.325000 ;
    END
  END D[3]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.975000 1.055000 13.795000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.405000 1.055000 19.225000 1.325000 ;
    END
  END D[5]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.415000 1.055000 20.235000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.845000 1.055000 25.665000 1.325000 ;
    END
  END D[7]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.790000 1.025000 3.125000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.315000 1.025000 3.650000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.230000 1.025000 9.565000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 9.755000 1.025000 10.090000 1.295000 ;
    END
  END S[3]
  PIN S[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.670000 1.025000 16.005000 1.295000 ;
    END
  END S[4]
  PIN S[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.195000 1.025000 16.530000 1.295000 ;
    END
  END S[5]
  PIN S[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.110000 1.025000 22.445000 1.295000 ;
    END
  END S[6]
  PIN S[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 22.635000 1.025000 22.970000 1.295000 ;
    END
  END S[7]
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  1.465000 1.755000  1.755000 1.800000 ;
        RECT  1.465000 1.800000 24.295000 1.940000 ;
        RECT  1.465000 1.940000  1.755000 1.985000 ;
        RECT  4.685000 1.755000  4.975000 1.800000 ;
        RECT  4.685000 1.940000  4.975000 1.985000 ;
        RECT  7.905000 1.755000  8.195000 1.800000 ;
        RECT  7.905000 1.940000  8.195000 1.985000 ;
        RECT 11.125000 1.755000 11.415000 1.800000 ;
        RECT 11.125000 1.940000 11.415000 1.985000 ;
        RECT 14.345000 1.755000 14.635000 1.800000 ;
        RECT 14.345000 1.940000 14.635000 1.985000 ;
        RECT 17.565000 1.755000 17.855000 1.800000 ;
        RECT 17.565000 1.940000 17.855000 1.985000 ;
        RECT 20.785000 1.755000 21.075000 1.800000 ;
        RECT 20.785000 1.940000 21.075000 1.985000 ;
        RECT 24.005000 1.755000 24.295000 1.800000 ;
        RECT 24.005000 1.940000 24.295000 1.985000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000 25.760000 2.805000 ;
      RECT  0.095000  1.495000  1.285000 1.665000 ;
      RECT  0.095000  1.665000  0.395000 2.210000 ;
      RECT  0.095000  2.210000  0.425000 2.465000 ;
      RECT  0.145000  0.255000  0.475000 0.715000 ;
      RECT  0.145000  0.715000  1.335000 0.885000 ;
      RECT  0.565000  1.835000  0.895000 2.105000 ;
      RECT  0.595000  2.105000  0.895000 2.635000 ;
      RECT  0.645000  0.085000  0.860000 0.545000 ;
      RECT  1.030000  0.255000  2.175000 0.425000 ;
      RECT  1.030000  0.425000  1.335000 0.715000 ;
      RECT  1.030000  0.885000  1.335000 0.925000 ;
      RECT  1.115000  1.665000  1.285000 2.295000 ;
      RECT  1.115000  2.295000  2.280000 2.465000 ;
      RECT  1.465000  1.755000  1.895000 2.125000 ;
      RECT  1.505000  0.595000  1.835000 0.885000 ;
      RECT  1.585000  0.885000  1.755000 1.755000 ;
      RECT  2.005000  0.425000  2.175000 0.770000 ;
      RECT  2.100000  1.205000  2.515000 1.305000 ;
      RECT  2.100000  1.305000  2.620000 1.465000 ;
      RECT  2.100000  1.465000  2.880000 1.475000 ;
      RECT  2.110000  1.645000  2.280000 2.295000 ;
      RECT  2.345000  0.585000  2.925000 0.755000 ;
      RECT  2.345000  0.755000  2.515000 1.205000 ;
      RECT  2.450000  1.475000  2.880000 1.635000 ;
      RECT  2.550000  1.635000  2.880000 2.465000 ;
      RECT  2.675000  0.330000  2.925000 0.585000 ;
      RECT  3.055000  1.465000  3.385000 2.635000 ;
      RECT  3.095000  0.085000  3.345000 0.660000 ;
      RECT  3.515000  0.330000  3.765000 0.585000 ;
      RECT  3.515000  0.585000  4.095000 0.755000 ;
      RECT  3.560000  1.465000  4.340000 1.475000 ;
      RECT  3.560000  1.475000  3.990000 1.635000 ;
      RECT  3.560000  1.635000  3.890000 2.465000 ;
      RECT  3.820000  1.305000  4.340000 1.465000 ;
      RECT  3.925000  0.755000  4.095000 1.205000 ;
      RECT  3.925000  1.205000  4.340000 1.305000 ;
      RECT  4.160000  1.645000  4.330000 2.295000 ;
      RECT  4.160000  2.295000  5.325000 2.465000 ;
      RECT  4.265000  0.255000  5.410000 0.425000 ;
      RECT  4.265000  0.425000  4.435000 0.770000 ;
      RECT  4.545000  1.755000  4.975000 2.125000 ;
      RECT  4.605000  0.595000  4.935000 0.885000 ;
      RECT  4.685000  0.885000  4.855000 1.755000 ;
      RECT  5.105000  0.425000  5.410000 0.715000 ;
      RECT  5.105000  0.715000  6.295000 0.885000 ;
      RECT  5.105000  0.885000  5.410000 0.925000 ;
      RECT  5.155000  1.495000  6.345000 1.665000 ;
      RECT  5.155000  1.665000  5.325000 2.295000 ;
      RECT  5.545000  1.835000  5.875000 2.105000 ;
      RECT  5.545000  2.105000  5.845000 2.635000 ;
      RECT  5.580000  0.085000  5.795000 0.545000 ;
      RECT  5.965000  0.255000  6.295000 0.715000 ;
      RECT  6.015000  2.210000  6.345000 2.465000 ;
      RECT  6.045000  1.665000  6.345000 2.210000 ;
      RECT  6.535000  1.495000  7.725000 1.665000 ;
      RECT  6.535000  1.665000  6.835000 2.210000 ;
      RECT  6.535000  2.210000  6.865000 2.465000 ;
      RECT  6.585000  0.255000  6.915000 0.715000 ;
      RECT  6.585000  0.715000  7.775000 0.885000 ;
      RECT  7.005000  1.835000  7.335000 2.105000 ;
      RECT  7.035000  2.105000  7.335000 2.635000 ;
      RECT  7.085000  0.085000  7.300000 0.545000 ;
      RECT  7.470000  0.255000  8.615000 0.425000 ;
      RECT  7.470000  0.425000  7.775000 0.715000 ;
      RECT  7.470000  0.885000  7.775000 0.925000 ;
      RECT  7.555000  1.665000  7.725000 2.295000 ;
      RECT  7.555000  2.295000  8.720000 2.465000 ;
      RECT  7.905000  1.755000  8.335000 2.125000 ;
      RECT  7.945000  0.595000  8.275000 0.885000 ;
      RECT  8.025000  0.885000  8.195000 1.755000 ;
      RECT  8.445000  0.425000  8.615000 0.770000 ;
      RECT  8.540000  1.205000  8.955000 1.305000 ;
      RECT  8.540000  1.305000  9.060000 1.465000 ;
      RECT  8.540000  1.465000  9.320000 1.475000 ;
      RECT  8.550000  1.645000  8.720000 2.295000 ;
      RECT  8.785000  0.585000  9.365000 0.755000 ;
      RECT  8.785000  0.755000  8.955000 1.205000 ;
      RECT  8.890000  1.475000  9.320000 1.635000 ;
      RECT  8.990000  1.635000  9.320000 2.465000 ;
      RECT  9.115000  0.330000  9.365000 0.585000 ;
      RECT  9.495000  1.465000  9.825000 2.635000 ;
      RECT  9.535000  0.085000  9.785000 0.660000 ;
      RECT  9.955000  0.330000 10.205000 0.585000 ;
      RECT  9.955000  0.585000 10.535000 0.755000 ;
      RECT 10.000000  1.465000 10.780000 1.475000 ;
      RECT 10.000000  1.475000 10.430000 1.635000 ;
      RECT 10.000000  1.635000 10.330000 2.465000 ;
      RECT 10.260000  1.305000 10.780000 1.465000 ;
      RECT 10.365000  0.755000 10.535000 1.205000 ;
      RECT 10.365000  1.205000 10.780000 1.305000 ;
      RECT 10.600000  1.645000 10.770000 2.295000 ;
      RECT 10.600000  2.295000 11.765000 2.465000 ;
      RECT 10.705000  0.255000 11.850000 0.425000 ;
      RECT 10.705000  0.425000 10.875000 0.770000 ;
      RECT 10.985000  1.755000 11.415000 2.125000 ;
      RECT 11.045000  0.595000 11.375000 0.885000 ;
      RECT 11.125000  0.885000 11.295000 1.755000 ;
      RECT 11.545000  0.425000 11.850000 0.715000 ;
      RECT 11.545000  0.715000 12.735000 0.885000 ;
      RECT 11.545000  0.885000 11.850000 0.925000 ;
      RECT 11.595000  1.495000 12.785000 1.665000 ;
      RECT 11.595000  1.665000 11.765000 2.295000 ;
      RECT 11.985000  1.835000 12.315000 2.105000 ;
      RECT 11.985000  2.105000 12.285000 2.635000 ;
      RECT 12.020000  0.085000 12.235000 0.545000 ;
      RECT 12.405000  0.255000 12.735000 0.715000 ;
      RECT 12.455000  2.210000 12.785000 2.465000 ;
      RECT 12.485000  1.665000 12.785000 2.210000 ;
      RECT 12.975000  1.495000 14.165000 1.665000 ;
      RECT 12.975000  1.665000 13.275000 2.210000 ;
      RECT 12.975000  2.210000 13.305000 2.465000 ;
      RECT 13.025000  0.255000 13.355000 0.715000 ;
      RECT 13.025000  0.715000 14.215000 0.885000 ;
      RECT 13.445000  1.835000 13.775000 2.105000 ;
      RECT 13.475000  2.105000 13.775000 2.635000 ;
      RECT 13.525000  0.085000 13.740000 0.545000 ;
      RECT 13.910000  0.255000 15.055000 0.425000 ;
      RECT 13.910000  0.425000 14.215000 0.715000 ;
      RECT 13.910000  0.885000 14.215000 0.925000 ;
      RECT 13.995000  1.665000 14.165000 2.295000 ;
      RECT 13.995000  2.295000 15.160000 2.465000 ;
      RECT 14.345000  1.755000 14.775000 2.125000 ;
      RECT 14.385000  0.595000 14.715000 0.885000 ;
      RECT 14.465000  0.885000 14.635000 1.755000 ;
      RECT 14.885000  0.425000 15.055000 0.770000 ;
      RECT 14.980000  1.205000 15.395000 1.305000 ;
      RECT 14.980000  1.305000 15.500000 1.465000 ;
      RECT 14.980000  1.465000 15.760000 1.475000 ;
      RECT 14.990000  1.645000 15.160000 2.295000 ;
      RECT 15.225000  0.585000 15.805000 0.755000 ;
      RECT 15.225000  0.755000 15.395000 1.205000 ;
      RECT 15.330000  1.475000 15.760000 1.635000 ;
      RECT 15.430000  1.635000 15.760000 2.465000 ;
      RECT 15.555000  0.330000 15.805000 0.585000 ;
      RECT 15.935000  1.465000 16.265000 2.635000 ;
      RECT 15.975000  0.085000 16.225000 0.660000 ;
      RECT 16.395000  0.330000 16.645000 0.585000 ;
      RECT 16.395000  0.585000 16.975000 0.755000 ;
      RECT 16.440000  1.465000 17.220000 1.475000 ;
      RECT 16.440000  1.475000 16.870000 1.635000 ;
      RECT 16.440000  1.635000 16.770000 2.465000 ;
      RECT 16.700000  1.305000 17.220000 1.465000 ;
      RECT 16.805000  0.755000 16.975000 1.205000 ;
      RECT 16.805000  1.205000 17.220000 1.305000 ;
      RECT 17.040000  1.645000 17.210000 2.295000 ;
      RECT 17.040000  2.295000 18.205000 2.465000 ;
      RECT 17.145000  0.255000 18.290000 0.425000 ;
      RECT 17.145000  0.425000 17.315000 0.770000 ;
      RECT 17.425000  1.755000 17.855000 2.125000 ;
      RECT 17.485000  0.595000 17.815000 0.885000 ;
      RECT 17.565000  0.885000 17.735000 1.755000 ;
      RECT 17.985000  0.425000 18.290000 0.715000 ;
      RECT 17.985000  0.715000 19.175000 0.885000 ;
      RECT 17.985000  0.885000 18.290000 0.925000 ;
      RECT 18.035000  1.495000 19.225000 1.665000 ;
      RECT 18.035000  1.665000 18.205000 2.295000 ;
      RECT 18.425000  1.835000 18.755000 2.105000 ;
      RECT 18.425000  2.105000 18.725000 2.635000 ;
      RECT 18.460000  0.085000 18.675000 0.545000 ;
      RECT 18.845000  0.255000 19.175000 0.715000 ;
      RECT 18.895000  2.210000 19.225000 2.465000 ;
      RECT 18.925000  1.665000 19.225000 2.210000 ;
      RECT 19.415000  1.495000 20.605000 1.665000 ;
      RECT 19.415000  1.665000 19.715000 2.210000 ;
      RECT 19.415000  2.210000 19.745000 2.465000 ;
      RECT 19.465000  0.255000 19.795000 0.715000 ;
      RECT 19.465000  0.715000 20.655000 0.885000 ;
      RECT 19.885000  1.835000 20.215000 2.105000 ;
      RECT 19.915000  2.105000 20.215000 2.635000 ;
      RECT 19.965000  0.085000 20.180000 0.545000 ;
      RECT 20.350000  0.255000 21.495000 0.425000 ;
      RECT 20.350000  0.425000 20.655000 0.715000 ;
      RECT 20.350000  0.885000 20.655000 0.925000 ;
      RECT 20.435000  1.665000 20.605000 2.295000 ;
      RECT 20.435000  2.295000 21.600000 2.465000 ;
      RECT 20.785000  1.755000 21.215000 2.125000 ;
      RECT 20.825000  0.595000 21.155000 0.885000 ;
      RECT 20.905000  0.885000 21.075000 1.755000 ;
      RECT 21.325000  0.425000 21.495000 0.770000 ;
      RECT 21.420000  1.205000 21.835000 1.305000 ;
      RECT 21.420000  1.305000 21.940000 1.465000 ;
      RECT 21.420000  1.465000 22.200000 1.475000 ;
      RECT 21.430000  1.645000 21.600000 2.295000 ;
      RECT 21.665000  0.585000 22.245000 0.755000 ;
      RECT 21.665000  0.755000 21.835000 1.205000 ;
      RECT 21.770000  1.475000 22.200000 1.635000 ;
      RECT 21.870000  1.635000 22.200000 2.465000 ;
      RECT 21.995000  0.330000 22.245000 0.585000 ;
      RECT 22.375000  1.465000 22.705000 2.635000 ;
      RECT 22.415000  0.085000 22.665000 0.660000 ;
      RECT 22.835000  0.330000 23.085000 0.585000 ;
      RECT 22.835000  0.585000 23.415000 0.755000 ;
      RECT 22.880000  1.465000 23.660000 1.475000 ;
      RECT 22.880000  1.475000 23.310000 1.635000 ;
      RECT 22.880000  1.635000 23.210000 2.465000 ;
      RECT 23.140000  1.305000 23.660000 1.465000 ;
      RECT 23.245000  0.755000 23.415000 1.205000 ;
      RECT 23.245000  1.205000 23.660000 1.305000 ;
      RECT 23.480000  1.645000 23.650000 2.295000 ;
      RECT 23.480000  2.295000 24.645000 2.465000 ;
      RECT 23.585000  0.255000 24.730000 0.425000 ;
      RECT 23.585000  0.425000 23.755000 0.770000 ;
      RECT 23.865000  1.755000 24.295000 2.125000 ;
      RECT 23.925000  0.595000 24.255000 0.885000 ;
      RECT 24.005000  0.885000 24.175000 1.755000 ;
      RECT 24.425000  0.425000 24.730000 0.715000 ;
      RECT 24.425000  0.715000 25.615000 0.885000 ;
      RECT 24.425000  0.885000 24.730000 0.925000 ;
      RECT 24.475000  1.495000 25.665000 1.665000 ;
      RECT 24.475000  1.665000 24.645000 2.295000 ;
      RECT 24.865000  1.835000 25.195000 2.105000 ;
      RECT 24.865000  2.105000 25.165000 2.635000 ;
      RECT 24.900000  0.085000 25.115000 0.545000 ;
      RECT 25.285000  0.255000 25.615000 0.715000 ;
      RECT 25.335000  2.210000 25.665000 2.465000 ;
      RECT 25.365000  1.665000 25.665000 2.210000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  1.785000  1.695000 1.955000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  1.785000  4.915000 1.955000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  1.785000  8.135000 1.955000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  1.785000 11.355000 1.955000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  1.785000 14.575000 1.955000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  1.785000 17.795000 1.955000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  1.785000 21.015000 1.955000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  1.785000 24.235000 1.955000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_2
END LIBRARY
