* File: sky130_fd_sc_hdll__or3b_1.spice
* Created: Wed Sep  2 08:48:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3b_1.pex.spice"
.subckt sky130_fd_sc_hdll__or3b_1  VNB VPB C_N B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_117_297#_M1006_d N_C_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_117_297#_M1002_g N_A_225_53#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_225_53#_M1000_d N_B_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.07665 AS=0.0567 PD=0.785 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_225_53#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0922822 AS=0.07665 PD=0.816449 PS=0.785 NRD=12.852 NRS=11.424 M=1 R=2.8
+ SA=75001.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1009 N_X_M1009_d N_A_225_53#_M1009_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.142818 PD=1.85 PS=1.26355 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_117_297#_M1003_d N_C_N_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1007 A_315_297# N_A_117_297#_M1007_g N_A_225_53#_M1007_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0504 AS=0.1134 PD=0.66 PS=1.38 NRD=30.4759 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1005 A_399_297# N_B_M1005_g A_315_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.07035
+ AS=0.0504 PD=0.755 PS=0.66 NRD=52.7566 NRS=30.4759 M=1 R=2.33333 SA=90000.6
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_399_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.07035 PD=0.804507 PS=0.755 NRD=76.83 NRS=52.7566 M=1
+ R=2.33333 SA=90001.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1008 N_X_M1008_d N_A_225_53#_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.285 AS=0.218803 PD=2.57 PS=1.91549 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_13 B B PROBETYPE=1
pX12_noxref noxref_14 A A PROBETYPE=1
c_66 VPB 0 2.17962e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__or3b_1.pxi.spice"
*
.ends
*
*
