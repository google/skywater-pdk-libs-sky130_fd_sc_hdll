* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or2_8 A B VGND VNB VPB VPWR X
X0 X a_123_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X a_123_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_123_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VPWR a_123_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 X a_123_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 X a_123_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND A a_123_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_123_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_123_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_123_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_123_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_123_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VGND a_123_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR a_123_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_123_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_123_47# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 X a_123_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND B a_123_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_123_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_27_297# B a_123_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR a_123_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 X a_123_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
