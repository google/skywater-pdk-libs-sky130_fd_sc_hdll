* File: sky130_fd_sc_hdll__and4b_2.spice
* Created: Wed Sep  2 08:23:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4b_2.pex.spice"
.subckt sky130_fd_sc_hdll__and4b_2  VNB VPB A_N B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1008 N_A_27_413#_M1008_d N_A_N_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 A_317_47# N_A_27_413#_M1010_g N_A_211_413#_M1010_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0546 AS=0.1092 PD=0.68 PS=1.36 NRD=21.42 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.7 A=0.063 P=1.14 MULT=1
MM1005 A_399_47# N_B_M1005_g A_317_47# VNB NSHORT L=0.15 W=0.42 AD=0.0945
+ AS=0.0546 PD=0.87 PS=0.68 NRD=48.564 NRS=21.42 M=1 R=2.8 SA=75000.6 SB=75002.3
+ A=0.063 P=1.14 MULT=1
MM1013 A_519_47# N_C_M1013_g A_399_47# VNB NSHORT L=0.15 W=0.42 AD=0.07245
+ AS=0.0945 PD=0.765 PS=0.87 NRD=33.564 NRS=48.564 M=1 R=2.8 SA=75001.2
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_D_M1002_g A_519_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0943822 AS=0.07245 PD=0.824299 PS=0.765 NRD=0 NRS=33.564 M=1 R=2.8
+ SA=75001.7 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1002_d N_A_211_413#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.146068 AS=0.115375 PD=1.2757 PS=1.005 NRD=23.076 NRS=5.532 M=1 R=4.33333
+ SA=75001.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_211_413#_M1012_g N_X_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.115375 PD=1.82 PS=1.005 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_N_M1001_g N_A_27_413#_M1001_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90003.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_211_413#_M1011_d N_A_27_413#_M1011_g N_VPWR_M1001_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.168 AS=0.0609 PD=1.22 PS=0.71 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.6 SB=90003.3 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_B_M1006_g N_A_211_413#_M1011_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0777 AS=0.168 PD=0.79 PS=1.22 NRD=39.8531 NRS=241.542 M=1 R=2.33333
+ SA=90001.6 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1009 N_A_211_413#_M1009_d N_C_M1009_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.06615 AS=0.0777 PD=0.735 PS=0.79 NRD=14.0658 NRS=2.3443 M=1 R=2.33333
+ SA=90002.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_D_M1000_g N_A_211_413#_M1009_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0914239 AS=0.06615 PD=0.810423 PS=0.735 NRD=39.8531 NRS=2.3443 M=1
+ R=2.33333 SA=90002.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_X_M1004_d N_A_211_413#_M1004_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.217676 PD=1.325 PS=1.92958 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1007 N_X_M1004_d N_A_211_413#_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.27 PD=1.325 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_16 C C PROBETYPE=1
pX16_noxref noxref_15 C C PROBETYPE=1
pX17_noxref noxref_17 X X PROBETYPE=1
pX18_noxref noxref_18 X X PROBETYPE=1
pX19_noxref noxref_19 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and4b_2.pxi.spice"
*
.ends
*
*
