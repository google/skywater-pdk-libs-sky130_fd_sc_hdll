# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__mux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__mux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.450000 0.995000 1.795000 1.615000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.965000 0.995000 2.585000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 0.995000 0.790000 1.325000 ;
        RECT 0.620000 0.635000 3.050000 0.805000 ;
        RECT 0.620000 0.805000 0.790000 0.995000 ;
        RECT 2.880000 0.805000 3.050000 0.995000 ;
        RECT 2.880000 0.995000 3.595000 1.325000 ;
    END
  END S
  PIN VGND
    ANTENNADIFFAREA  0.835250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.465000 ;
        RECT 3.615000  0.085000 3.995000 0.465000 ;
        RECT 4.555000  0.085000 4.935000 0.465000 ;
        RECT 5.495000  0.085000 5.875000 0.465000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.195000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.515000 1.835000 0.870000 2.635000 ;
        RECT 3.615000 2.255000 3.995000 2.635000 ;
        RECT 4.555000 1.915000 4.935000 2.635000 ;
        RECT 5.495000 1.915000 5.875000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.215000 0.255000 4.385000 0.635000 ;
        RECT 4.215000 0.635000 5.880000 0.805000 ;
        RECT 4.215000 1.575000 5.880000 1.745000 ;
        RECT 4.215000 1.745000 4.385000 2.465000 ;
        RECT 5.155000 0.255000 5.325000 0.635000 ;
        RECT 5.155000 1.745000 5.325000 2.465000 ;
        RECT 5.650000 0.805000 5.880000 1.575000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.090000 0.295000 0.345000 0.625000 ;
      RECT 0.090000 0.625000 0.260000 1.495000 ;
      RECT 0.090000 1.495000 1.180000 1.665000 ;
      RECT 0.090000 1.665000 0.345000 2.465000 ;
      RECT 0.960000 0.995000 1.180000 1.495000 ;
      RECT 1.040000 1.935000 1.440000 2.275000 ;
      RECT 1.040000 2.275000 2.970000 2.445000 ;
      RECT 1.630000 1.935000 3.445000 2.105000 ;
      RECT 2.075000 0.295000 3.430000 0.465000 ;
      RECT 2.130000 1.595000 3.985000 1.765000 ;
      RECT 3.260000 0.465000 3.430000 0.655000 ;
      RECT 3.260000 0.655000 3.985000 0.825000 ;
      RECT 3.275000 2.105000 3.445000 2.465000 ;
      RECT 3.815000 0.825000 3.985000 1.075000 ;
      RECT 3.815000 1.075000 5.430000 1.245000 ;
      RECT 3.815000 1.245000 3.985000 1.595000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__mux2_4
