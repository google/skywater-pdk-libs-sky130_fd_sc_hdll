* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor4_4 A B C D VGND VNB VPB VPWR Y
X0 a_497_297# C a_887_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_887_297# C a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_887_297# C a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_497_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_887_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 Y D a_887_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 Y D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_497_297# C a_887_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_27_297# B a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y D a_887_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_887_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_497_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_297# B a_497_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VGND D Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VGND C Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y C VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
