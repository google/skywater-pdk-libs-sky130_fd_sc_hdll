* File: sky130_fd_sc_hdll__dfrtp_1.spice
* Created: Wed Sep  2 08:28:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dfrtp_1.pex.spice"
.subckt sky130_fd_sc_hdll__dfrtp_1  VNB VPB CLK D RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1023 N_VGND_M1023_d N_CLK_M1023_g N_A_27_47#_M1023_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_211_363#_M1002_d N_A_27_47#_M1002_g N_VGND_M1023_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 N_A_436_413#_M1008_d N_D_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0720462 AS=0.1869 PD=0.807692 PS=1.73 NRD=0 NRS=45.708 M=1 R=2.8
+ SA=75000.4 SB=75005.4 A=0.063 P=1.14 MULT=1
MM1015 N_A_534_47#_M1015_d N_A_27_47#_M1015_g N_A_436_413#_M1008_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0702 AS=0.0617538 PD=0.75 PS=0.692308 NRD=16.656 NRS=16.656
+ M=1 R=2.4 SA=75000.8 SB=75005.8 A=0.054 P=1.02 MULT=1
MM1018 A_642_47# N_A_211_363#_M1018_g N_A_534_47#_M1015_d VNB NSHORT L=0.15
+ W=0.36 AD=0.126831 AS=0.0702 PD=1.00154 PS=0.75 NRD=99.096 NRS=19.992 M=1
+ R=2.4 SA=75001.4 SB=75005.2 A=0.054 P=1.02 MULT=1
MM1005 A_805_47# N_A_751_289#_M1005_g A_642_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.147969 PD=0.63 PS=1.16846 NRD=14.28 NRS=84.936 M=1 R=2.8
+ SA=75002 SB=75004 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_RESET_B_M1007_g A_805_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.127664 AS=0.0441 PD=0.990566 PS=0.63 NRD=47.136 NRS=14.28 M=1 R=2.8
+ SA=75002.3 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_751_289#_M1011_d N_A_534_47#_M1011_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.64 AD=0.127872 AS=0.194536 PD=1.2608 PS=1.50943 NRD=2.808 NRS=30.936 M=1
+ R=4.26667 SA=75002.1 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1014 N_A_1128_47#_M1014_d N_A_211_363#_M1014_g N_A_751_289#_M1011_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0711 AS=0.071928 PD=0.755 PS=0.7092 NRD=39.996 NRS=16.656
+ M=1 R=2.4 SA=75003.8 SB=75002.8 A=0.054 P=1.02 MULT=1
MM1019 A_1237_47# N_A_27_47#_M1019_g N_A_1128_47#_M1014_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0783692 AS=0.0711 PD=0.784615 PS=0.755 NRD=54.228 NRS=0 M=1 R=2.4
+ SA=75004.4 SB=75002.2 A=0.054 P=1.02 MULT=1
MM1009 N_VGND_M1009_d N_A_1323_21#_M1009_g A_1237_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.16695 AS=0.0914308 PD=1.215 PS=0.915385 NRD=1.428 NRS=46.476 M=1 R=2.8
+ SA=75004.3 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1020 A_1542_47# N_RESET_B_M1020_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.16695 PD=0.8 PS=1.215 NRD=38.568 NRS=145.704 M=1 R=2.8
+ SA=75005.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1021 N_A_1323_21#_M1021_d N_A_1128_47#_M1021_g A_1542_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0798 PD=1.36 PS=0.8 NRD=0 NRS=38.568 M=1 R=2.8
+ SA=75005.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_Q_M1003_d N_A_1323_21#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.2015 PD=1.86 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1025 N_A_211_363#_M1025_d N_A_27_47#_M1025_g N_VPWR_M1006_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1000 N_A_436_413#_M1000_d N_D_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0714 AS=0.1134 PD=0.76 PS=1.38 NRD=7.0329 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1026 N_A_534_47#_M1026_d N_A_211_363#_M1026_g N_A_436_413#_M1000_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07665 AS=0.0714 PD=0.785 PS=0.76 NRD=4.6886 NRS=21.0987 M=1
+ R=2.33333 SA=90000.7 SB=90002 A=0.0756 P=1.2 MULT=1
MM1004 N_A_649_413#_M1004_d N_A_27_47#_M1004_g N_A_534_47#_M1026_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1092 AS=0.07665 PD=0.94 PS=0.785 NRD=110.222 NRS=35.1645
+ M=1 R=2.33333 SA=90001.2 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_751_289#_M1010_g N_A_649_413#_M1004_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07455 AS=0.1092 PD=0.775 PS=0.94 NRD=32.8202 NRS=2.3443 M=1
+ R=2.33333 SA=90001.9 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1022 N_A_649_413#_M1022_d N_RESET_B_M1022_g N_VPWR_M1010_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.07455 PD=1.38 PS=0.775 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90002.5 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1016 N_A_751_289#_M1016_d N_A_534_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.1806 AS=0.2688 PD=1.60667 PS=2.32 NRD=5.8509 NRS=1.1623 M=1
+ R=4.66667 SA=90000.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1017 N_A_1128_47#_M1017_d N_A_27_47#_M1017_g N_A_751_289#_M1016_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0756 AS=0.0903 PD=0.78 PS=0.803333 NRD=7.0329 NRS=28.1316
+ M=1 R=2.33333 SA=90000.8 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1027 A_1330_413# N_A_211_363#_M1027_g N_A_1128_47#_M1017_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0483 AS=0.0756 PD=0.65 PS=0.78 NRD=28.1316 NRS=30.4759 M=1
+ R=2.33333 SA=90001.3 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1001 N_VPWR_M1001_d N_A_1323_21#_M1001_g A_1330_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1071 AS=0.0483 PD=0.93 PS=0.65 NRD=105.533 NRS=28.1316 M=1 R=2.33333
+ SA=90001.7 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1024 N_A_1323_21#_M1024_d N_RESET_B_M1024_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.063 AS=0.1071 PD=0.72 PS=0.93 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90002.4 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1013 N_VPWR_M1013_d N_A_1128_47#_M1013_g N_A_1323_21#_M1024_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1134 AS=0.063 PD=1.38 PS=0.72 NRD=2.3443 NRS=7.0329 M=1
+ R=2.33333 SA=90002.9 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1012 N_Q_M1012_d N_A_1323_21#_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.27 PD=2.58 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX28_noxref VNB VPB NWDIODE A=16.1142 P=23.29
c_186 VPB 0 2.7155e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__dfrtp_1.pxi.spice"
*
.ends
*
*
