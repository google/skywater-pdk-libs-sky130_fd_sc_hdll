* File: sky130_fd_sc_hdll__mux2_2.pxi.spice
* Created: Thu Aug 27 19:10:41 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2_2%A_79_21# N_A_79_21#_M1004_d N_A_79_21#_M1010_d
+ N_A_79_21#_c_77_n N_A_79_21#_M1006_g N_A_79_21#_c_84_n N_A_79_21#_M1000_g
+ N_A_79_21#_c_78_n N_A_79_21#_M1012_g N_A_79_21#_c_85_n N_A_79_21#_M1009_g
+ N_A_79_21#_c_86_n N_A_79_21#_c_79_n N_A_79_21#_c_155_p N_A_79_21#_c_87_n
+ N_A_79_21#_c_131_p N_A_79_21#_c_101_p N_A_79_21#_c_102_p N_A_79_21#_c_112_p
+ N_A_79_21#_c_80_n N_A_79_21#_c_93_p N_A_79_21#_c_81_n N_A_79_21#_c_82_n
+ N_A_79_21#_c_83_n PM_SKY130_FD_SC_HDLL__MUX2_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__MUX2_2%A_280_21# N_A_280_21#_M1013_d N_A_280_21#_M1001_d
+ N_A_280_21#_M1011_g N_A_280_21#_c_192_n N_A_280_21#_c_193_n
+ N_A_280_21#_M1008_g N_A_280_21#_c_189_n N_A_280_21#_c_190_n
+ N_A_280_21#_c_196_n N_A_280_21#_c_197_n N_A_280_21#_c_224_n
+ N_A_280_21#_c_191_n N_A_280_21#_c_199_n N_A_280_21#_c_200_n
+ PM_SKY130_FD_SC_HDLL__MUX2_2%A_280_21#
x_PM_SKY130_FD_SC_HDLL__MUX2_2%A0 N_A0_M1004_g N_A0_c_278_n N_A0_M1002_g
+ N_A0_c_279_n A0 A0 A0 A0 N_A0_c_282_n N_A0_c_283_n A0 A0
+ PM_SKY130_FD_SC_HDLL__MUX2_2%A0
x_PM_SKY130_FD_SC_HDLL__MUX2_2%A1 N_A1_M1007_g N_A1_c_334_n N_A1_c_340_n
+ N_A1_M1010_g N_A1_c_335_n N_A1_c_336_n A1 A1 N_A1_c_338_n
+ PM_SKY130_FD_SC_HDLL__MUX2_2%A1
x_PM_SKY130_FD_SC_HDLL__MUX2_2%S N_S_M1005_g N_S_c_385_n N_S_c_386_n N_S_M1003_g
+ N_S_c_387_n N_S_c_388_n N_S_M1001_g N_S_M1013_g S S S N_S_c_384_n
+ PM_SKY130_FD_SC_HDLL__MUX2_2%S
x_PM_SKY130_FD_SC_HDLL__MUX2_2%VPWR N_VPWR_M1000_d N_VPWR_M1009_d N_VPWR_M1003_d
+ N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n N_VPWR_c_434_n
+ N_VPWR_c_435_n N_VPWR_c_436_n VPWR N_VPWR_c_437_n N_VPWR_c_429_n
+ N_VPWR_c_439_n PM_SKY130_FD_SC_HDLL__MUX2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2_2%X N_X_M1006_s N_X_M1000_s N_X_c_490_n N_X_c_501_n
+ X X PM_SKY130_FD_SC_HDLL__MUX2_2%X
x_PM_SKY130_FD_SC_HDLL__MUX2_2%VGND N_VGND_M1006_d N_VGND_M1012_d N_VGND_M1005_d
+ N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n N_VGND_c_524_n
+ VGND N_VGND_c_525_n N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n
+ PM_SKY130_FD_SC_HDLL__MUX2_2%VGND
cc_1 VNB N_A_79_21#_c_77_n 0.0219887f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_78_n 0.0173392f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_79_21#_c_79_n 0.00292005f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.72
cc_4 VNB N_A_79_21#_c_80_n 0.00350755f $X=-0.19 $Y=-0.24 $X2=1.705 $Y2=0.43
cc_5 VNB N_A_79_21#_c_81_n 0.00306205f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.16
cc_6 VNB N_A_79_21#_c_82_n 0.00181439f $X=-0.19 $Y=-0.24 $X2=1.117 $Y2=0.995
cc_7 VNB N_A_79_21#_c_83_n 0.0554113f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_8 VNB N_A_280_21#_M1011_g 0.0298728f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_9 VNB N_A_280_21#_c_189_n 0.00100769f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_10 VNB N_A_280_21#_c_190_n 0.0253963f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.805
cc_11 VNB N_A_280_21#_c_191_n 0.0500924f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=2.34
cc_12 VNB N_A0_c_278_n 0.0085057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A0_c_279_n 4.2567e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_14 VNB A0 0.00814478f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB A0 0.00671156f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_16 VNB N_A0_c_282_n 0.0305507f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_17 VNB N_A0_c_283_n 0.0175405f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.995
cc_18 VNB N_A1_M1007_g 0.0225707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A1_c_334_n 0.01765f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A1_c_335_n 0.00877019f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_21 VNB N_A1_c_336_n 0.0358815f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_22 VNB A1 0.00298551f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_23 VNB N_A1_c_338_n 0.0051537f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.92
cc_24 VNB N_S_M1005_g 0.0332673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_S_M1013_g 0.033403f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_26 VNB S 0.00388431f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.805
cc_27 VNB N_S_c_384_n 0.0443155f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_429_n 0.193827f $X=-0.19 $Y=-0.24 $X2=1.117 $Y2=0.995
cc_29 VNB N_X_c_490_n 7.73293e-19 $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_30 VNB N_VGND_c_520_n 0.00997339f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_31 VNB N_VGND_c_521_n 0.0330966f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_32 VNB N_VGND_c_522_n 0.00491179f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_33 VNB N_VGND_c_523_n 0.0582511f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.805
cc_34 VNB N_VGND_c_524_n 0.00382076f $X=-0.19 $Y=-0.24 $X2=1.18 $Y2=0.995
cc_35 VNB N_VGND_c_525_n 0.0164934f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=0.72
cc_36 VNB N_VGND_c_526_n 0.0289273f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_527_n 0.249136f $X=-0.19 $Y=-0.24 $X2=1.117 $Y2=1.16
cc_38 VNB N_VGND_c_528_n 0.0090329f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=0.72
cc_39 VPB N_A_79_21#_c_84_n 0.0207574f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_40 VPB N_A_79_21#_c_85_n 0.0168411f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_41 VPB N_A_79_21#_c_86_n 0.00203598f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.835
cc_42 VPB N_A_79_21#_c_87_n 0.00333776f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.92
cc_43 VPB N_A_79_21#_c_81_n 0.00123844f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.16
cc_44 VPB N_A_79_21#_c_83_n 0.0278057f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_45 VPB N_A_280_21#_c_192_n 0.0241976f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_46 VPB N_A_280_21#_c_193_n 0.02689f $X=-0.19 $Y=1.305 $X2=0.94 $Y2=0.995
cc_47 VPB N_A_280_21#_c_189_n 0.00256734f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_48 VPB N_A_280_21#_c_190_n 0.00344177f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.805
cc_49 VPB N_A_280_21#_c_196_n 0.00501218f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=1.835
cc_50 VPB N_A_280_21#_c_197_n 0.0192783f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=0.72
cc_51 VPB N_A_280_21#_c_191_n 0.0278302f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=2.34
cc_52 VPB N_A_280_21#_c_199_n 0.0141757f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=0.43
cc_53 VPB N_A_280_21#_c_200_n 0.0284728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A0_c_278_n 0.0424629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A0_c_279_n 0.00825435f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_56 VPB A0 0.00611791f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_57 VPB N_A1_c_334_n 0.021982f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A1_c_340_n 0.0269075f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_59 VPB N_S_c_385_n 0.0174893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_S_c_386_n 0.0217648f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_61 VPB N_S_c_387_n 0.0205793f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_62 VPB N_S_c_388_n 0.0256439f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_63 VPB S 0.00348655f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.805
cc_64 VPB N_S_c_384_n 0.00490776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_430_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_66 VPB N_VPWR_c_431_n 0.0431474f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_67 VPB N_VPWR_c_432_n 0.0208473f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_68 VPB N_VPWR_c_433_n 0.00470153f $X=-0.19 $Y=1.305 $X2=1.18 $Y2=0.995
cc_69 VPB N_VPWR_c_434_n 0.00495385f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.72
cc_70 VPB N_VPWR_c_435_n 0.0540373f $X=-0.19 $Y=1.305 $X2=1.54 $Y2=2.005
cc_71 VPB N_VPWR_c_436_n 0.00420071f $X=-0.19 $Y=1.305 $X2=1.54 $Y2=2.255
cc_72 VPB N_VPWR_c_437_n 0.0270276f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.16
cc_73 VPB N_VPWR_c_429_n 0.0554144f $X=-0.19 $Y=1.305 $X2=1.117 $Y2=0.995
cc_74 VPB N_VPWR_c_439_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.202
cc_75 VPB N_X_c_490_n 0.00112597f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_76 N_A_79_21#_c_78_n N_A_280_21#_M1011_g 0.0185432f $X=0.94 $Y=0.995 $X2=0
+ $Y2=0
cc_77 N_A_79_21#_c_79_n N_A_280_21#_M1011_g 0.0108847f $X=1.535 $Y=0.72 $X2=0
+ $Y2=0
cc_78 N_A_79_21#_c_80_n N_A_280_21#_M1011_g 0.0107164f $X=1.705 $Y=0.43 $X2=0
+ $Y2=0
cc_79 N_A_79_21#_c_93_p N_A_280_21#_M1011_g 4.05547e-19 $X=2.165 $Y=0.43 $X2=0
+ $Y2=0
cc_80 N_A_79_21#_c_82_n N_A_280_21#_M1011_g 0.00257804f $X=1.117 $Y=0.995 $X2=0
+ $Y2=0
cc_81 N_A_79_21#_c_85_n N_A_280_21#_c_192_n 0.00967123f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_82 N_A_79_21#_c_86_n N_A_280_21#_c_192_n 0.00257804f $X=1.18 $Y=1.835 $X2=0
+ $Y2=0
cc_83 N_A_79_21#_c_83_n N_A_280_21#_c_192_n 0.00239585f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_84 N_A_79_21#_c_85_n N_A_280_21#_c_193_n 0.0205255f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_85 N_A_79_21#_c_86_n N_A_280_21#_c_193_n 6.85928e-19 $X=1.18 $Y=1.835 $X2=0
+ $Y2=0
cc_86 N_A_79_21#_c_87_n N_A_280_21#_c_193_n 0.0125829f $X=1.455 $Y=1.92 $X2=0
+ $Y2=0
cc_87 N_A_79_21#_c_101_p N_A_280_21#_c_193_n 0.00961653f $X=1.54 $Y=2.255 $X2=0
+ $Y2=0
cc_88 N_A_79_21#_c_102_p N_A_280_21#_c_193_n 0.008657f $X=1.625 $Y=2.34 $X2=0
+ $Y2=0
cc_89 N_A_79_21#_c_79_n N_A_280_21#_c_189_n 0.00672059f $X=1.535 $Y=0.72 $X2=0
+ $Y2=0
cc_90 N_A_79_21#_c_80_n N_A_280_21#_c_189_n 0.00922398f $X=1.705 $Y=0.43 $X2=0
+ $Y2=0
cc_91 N_A_79_21#_c_81_n N_A_280_21#_c_189_n 0.0374429f $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_79_21#_c_83_n N_A_280_21#_c_189_n 3.33026e-19 $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_80_n N_A_280_21#_c_190_n 0.00145753f $X=1.705 $Y=0.43 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_81_n N_A_280_21#_c_190_n 0.00257804f $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_83_n N_A_280_21#_c_190_n 0.0203215f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_86_n N_A_280_21#_c_196_n 0.00549775f $X=1.18 $Y=1.835 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_M1010_d N_A_280_21#_c_197_n 0.00227859f $X=2.55 $Y=1.845 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_112_p N_A_280_21#_c_197_n 0.0352098f $X=2.695 $Y=2.34 $X2=0
+ $Y2=0
cc_99 N_A_79_21#_c_87_n N_A_280_21#_c_224_n 0.00808719f $X=1.455 $Y=1.92 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_112_p N_A_280_21#_c_224_n 0.00894068f $X=2.695 $Y=2.34 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_86_n N_A_280_21#_c_199_n 0.0129412f $X=1.18 $Y=1.835 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_87_n N_A_280_21#_c_199_n 0.0143337f $X=1.455 $Y=1.92 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_112_p N_A_280_21#_c_199_n 0.00485029f $X=2.695 $Y=2.34 $X2=0
+ $Y2=0
cc_104 N_A_79_21#_c_112_p N_A0_c_278_n 0.00327688f $X=2.695 $Y=2.34 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_80_n A0 0.00254523f $X=1.705 $Y=0.43 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_93_p A0 0.0237984f $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_82_n A0 0.00496004f $X=1.117 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_93_p N_A0_c_282_n 7.44232e-19 $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_80_n N_A0_c_283_n 0.00425097f $X=1.705 $Y=0.43 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_93_p N_A0_c_283_n 0.0123074f $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_80_n N_A1_M1007_g 2.42031e-19 $X=1.705 $Y=0.43 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_112_p N_A1_c_340_n 0.0117722f $X=2.695 $Y=2.34 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_93_p A1 0.00529558f $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_112_p N_S_c_386_n 4.64095e-19 $X=2.695 $Y=2.34 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_86_n N_VPWR_M1009_d 0.00607726f $X=1.18 $Y=1.835 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_87_n N_VPWR_M1009_d 0.00334871f $X=1.455 $Y=1.92 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_131_p N_VPWR_M1009_d 0.00270618f $X=1.265 $Y=1.92 $X2=0
+ $Y2=0
cc_118 N_A_79_21#_c_84_n N_VPWR_c_431_n 0.00777278f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_84_n N_VPWR_c_432_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_85_n N_VPWR_c_432_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_85_n N_VPWR_c_433_n 0.00420128f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_79_21#_c_87_n N_VPWR_c_433_n 0.00144965f $X=1.455 $Y=1.92 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_131_p N_VPWR_c_433_n 0.0128103f $X=1.265 $Y=1.92 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_101_p N_VPWR_c_433_n 0.00558249f $X=1.54 $Y=2.255 $X2=0
+ $Y2=0
cc_125 N_A_79_21#_c_102_p N_VPWR_c_433_n 0.0133618f $X=1.625 $Y=2.34 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_87_n N_VPWR_c_435_n 0.00206015f $X=1.455 $Y=1.92 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_102_p N_VPWR_c_435_n 0.00821268f $X=1.625 $Y=2.34 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_c_112_p N_VPWR_c_435_n 0.0578461f $X=2.695 $Y=2.34 $X2=0 $Y2=0
cc_129 N_A_79_21#_M1010_d N_VPWR_c_429_n 0.00241975f $X=2.55 $Y=1.845 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_c_84_n N_VPWR_c_429_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_85_n N_VPWR_c_429_n 0.0126813f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_87_n N_VPWR_c_429_n 0.0044085f $X=1.455 $Y=1.92 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_131_p N_VPWR_c_429_n 0.00125604f $X=1.265 $Y=1.92 $X2=0
+ $Y2=0
cc_134 N_A_79_21#_c_102_p N_VPWR_c_429_n 0.00575824f $X=1.625 $Y=2.34 $X2=0
+ $Y2=0
cc_135 N_A_79_21#_c_112_p N_VPWR_c_429_n 0.0438553f $X=2.695 $Y=2.34 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_77_n N_X_c_490_n 0.0158841f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_84_n N_X_c_490_n 0.00703694f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_78_n N_X_c_490_n 0.00797783f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_85_n N_X_c_490_n 0.00170371f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_79_21#_c_86_n N_X_c_490_n 0.0113319f $X=1.18 $Y=1.835 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_155_p N_X_c_490_n 0.00921699f $X=1.265 $Y=0.72 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_81_n N_X_c_490_n 0.024279f $X=1.055 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_82_n N_X_c_490_n 0.00984496f $X=1.117 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_79_21#_c_83_n N_X_c_490_n 0.040921f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_145 N_A_79_21#_c_84_n N_X_c_501_n 0.00440365f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_79_21#_c_83_n N_X_c_501_n 0.00180397f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_147 N_A_79_21#_c_84_n X 0.0105729f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_79_21#_c_101_p X 0.00509128f $X=1.54 $Y=2.255 $X2=0 $Y2=0
cc_149 N_A_79_21#_c_112_p A_318_369# 0.020191f $X=2.695 $Y=2.34 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_79_21#_c_79_n N_VGND_M1012_d 0.00265709f $X=1.535 $Y=0.72 $X2=0 $Y2=0
cc_151 N_A_79_21#_c_155_p N_VGND_M1012_d 0.00469518f $X=1.265 $Y=0.72 $X2=0
+ $Y2=0
cc_152 N_A_79_21#_c_82_n N_VGND_M1012_d 0.00200923f $X=1.117 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_79_21#_c_77_n N_VGND_c_521_n 0.00318044f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_79_21#_c_79_n N_VGND_c_523_n 0.00255155f $X=1.535 $Y=0.72 $X2=0 $Y2=0
cc_155 N_A_79_21#_c_80_n N_VGND_c_523_n 0.00909399f $X=1.705 $Y=0.43 $X2=0 $Y2=0
cc_156 N_A_79_21#_c_93_p N_VGND_c_523_n 0.0303561f $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_77_n N_VGND_c_525_n 0.00541359f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_79_21#_c_78_n N_VGND_c_525_n 0.00468308f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_79_21#_M1004_d N_VGND_c_527_n 0.00513778f $X=2.03 $Y=0.235 $X2=0
+ $Y2=0
cc_160 N_A_79_21#_c_77_n N_VGND_c_527_n 0.0105827f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_79_21#_c_78_n N_VGND_c_527_n 0.00801881f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_79_21#_c_79_n N_VGND_c_527_n 0.00457575f $X=1.535 $Y=0.72 $X2=0 $Y2=0
cc_163 N_A_79_21#_c_155_p N_VGND_c_527_n 8.57032e-19 $X=1.265 $Y=0.72 $X2=0
+ $Y2=0
cc_164 N_A_79_21#_c_80_n N_VGND_c_527_n 0.00633526f $X=1.705 $Y=0.43 $X2=0 $Y2=0
cc_165 N_A_79_21#_c_93_p N_VGND_c_527_n 0.0197303f $X=2.165 $Y=0.43 $X2=0 $Y2=0
cc_166 N_A_79_21#_c_77_n N_VGND_c_528_n 4.73309e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_79_21#_c_78_n N_VGND_c_528_n 0.00761466f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_79_21#_c_79_n N_VGND_c_528_n 0.00591836f $X=1.535 $Y=0.72 $X2=0 $Y2=0
cc_169 N_A_79_21#_c_155_p N_VGND_c_528_n 0.0143265f $X=1.265 $Y=0.72 $X2=0 $Y2=0
cc_170 N_A_79_21#_c_81_n N_VGND_c_528_n 0.0024979f $X=1.055 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_79_21#_c_83_n N_VGND_c_528_n 6.12683e-19 $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_172 N_A_79_21#_c_80_n A_310_47# 0.00246712f $X=1.705 $Y=0.43 $X2=-0.19
+ $Y2=-0.24
cc_173 N_A_79_21#_c_93_p A_310_47# 0.00682357f $X=2.165 $Y=0.43 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_280_21#_c_197_n N_A0_c_278_n 0.0147834f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_175 N_A_280_21#_c_192_n N_A0_c_279_n 0.00153506f $X=1.5 $Y=1.67 $X2=0 $Y2=0
cc_176 N_A_280_21#_c_189_n N_A0_c_279_n 0.00981607f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_280_21#_c_190_n N_A0_c_279_n 4.92482e-19 $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_178 N_A_280_21#_c_197_n N_A0_c_279_n 0.0182718f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_179 N_A_280_21#_c_199_n N_A0_c_279_n 0.0156059f $X=1.88 $Y=1.58 $X2=0 $Y2=0
cc_180 N_A_280_21#_M1011_g A0 7.36251e-19 $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_181 N_A_280_21#_c_189_n A0 0.0154634f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_280_21#_c_190_n A0 0.00223847f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_280_21#_c_197_n A0 0.0503986f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_184 N_A_280_21#_c_189_n N_A0_c_282_n 3.39173e-19 $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_280_21#_c_190_n N_A0_c_282_n 0.00597f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_186 N_A_280_21#_c_199_n N_A0_c_282_n 0.00150231f $X=1.88 $Y=1.58 $X2=0 $Y2=0
cc_187 N_A_280_21#_M1011_g N_A0_c_283_n 0.0322139f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_280_21#_c_190_n N_A1_c_334_n 0.00219244f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_280_21#_c_196_n N_A1_c_334_n 0.00291318f $X=1.88 $Y=1.835 $X2=0 $Y2=0
cc_190 N_A_280_21#_c_199_n N_A1_c_334_n 0.00186037f $X=1.88 $Y=1.58 $X2=0 $Y2=0
cc_191 N_A_280_21#_c_196_n N_A1_c_340_n 0.00174455f $X=1.88 $Y=1.835 $X2=0 $Y2=0
cc_192 N_A_280_21#_c_197_n N_A1_c_340_n 0.0151681f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_193 N_A_280_21#_c_197_n N_S_c_386_n 0.0173758f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_194 N_A_280_21#_c_200_n N_S_c_386_n 8.56106e-19 $X=4.065 $Y=2 $X2=0 $Y2=0
cc_195 N_A_280_21#_c_197_n N_S_c_388_n 0.0126643f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_196 N_A_280_21#_c_191_n N_S_c_388_n 0.00259523f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_197 N_A_280_21#_c_200_n N_S_c_388_n 0.0127533f $X=4.065 $Y=2 $X2=0 $Y2=0
cc_198 N_A_280_21#_c_191_n N_S_M1013_g 0.0391993f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_199 N_A_280_21#_c_197_n S 0.0129203f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_200 N_A_280_21#_c_191_n S 0.033812f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_201 N_A_280_21#_c_197_n N_S_c_384_n 0.00226267f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_202 N_A_280_21#_c_197_n N_VPWR_M1003_d 0.00182309f $X=3.85 $Y=1.92 $X2=0
+ $Y2=0
cc_203 N_A_280_21#_c_193_n N_VPWR_c_433_n 0.00553176f $X=1.5 $Y=1.77 $X2=0 $Y2=0
cc_204 N_A_280_21#_c_197_n N_VPWR_c_434_n 0.0137405f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_205 N_A_280_21#_c_193_n N_VPWR_c_435_n 0.00460264f $X=1.5 $Y=1.77 $X2=0 $Y2=0
cc_206 N_A_280_21#_c_197_n N_VPWR_c_435_n 0.00756012f $X=3.85 $Y=1.92 $X2=0
+ $Y2=0
cc_207 N_A_280_21#_c_197_n N_VPWR_c_437_n 0.0020257f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_208 N_A_280_21#_c_200_n N_VPWR_c_437_n 0.0248195f $X=4.065 $Y=2 $X2=0 $Y2=0
cc_209 N_A_280_21#_M1001_d N_VPWR_c_429_n 0.00225715f $X=3.91 $Y=1.845 $X2=0
+ $Y2=0
cc_210 N_A_280_21#_c_193_n N_VPWR_c_429_n 0.00787179f $X=1.5 $Y=1.77 $X2=0 $Y2=0
cc_211 N_A_280_21#_c_197_n N_VPWR_c_429_n 0.0210048f $X=3.85 $Y=1.92 $X2=0 $Y2=0
cc_212 N_A_280_21#_c_200_n N_VPWR_c_429_n 0.0143976f $X=4.065 $Y=2 $X2=0 $Y2=0
cc_213 N_A_280_21#_c_197_n A_318_369# 0.00622228f $X=3.85 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_214 N_A_280_21#_c_224_n A_318_369# 0.0050135f $X=1.965 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_215 N_A_280_21#_c_197_n A_606_369# 0.00220509f $X=3.85 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_216 N_A_280_21#_c_191_n N_VGND_c_522_n 0.0164398f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_217 N_A_280_21#_M1011_g N_VGND_c_523_n 0.00420065f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_280_21#_c_191_n N_VGND_c_526_n 0.0174931f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_219 N_A_280_21#_M1013_d N_VGND_c_527_n 0.00447268f $X=3.92 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_A_280_21#_M1011_g N_VGND_c_527_n 0.00611525f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_280_21#_c_191_n N_VGND_c_527_n 0.00955092f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_222 N_A_280_21#_M1011_g N_VGND_c_528_n 0.00450023f $X=1.475 $Y=0.445 $X2=0
+ $Y2=0
cc_223 A0 N_A1_M1007_g 0.00860106f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_224 N_A0_c_282_n N_A1_M1007_g 0.0204296f $X=2.015 $Y=0.93 $X2=0 $Y2=0
cc_225 N_A0_c_283_n N_A1_M1007_g 0.0110449f $X=2.015 $Y=0.765 $X2=0 $Y2=0
cc_226 N_A0_c_278_n N_A1_c_334_n 0.0294622f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_227 A0 N_A1_c_334_n 0.0275759f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_228 N_A0_c_278_n N_A1_c_340_n 0.0231406f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_229 N_A0_c_278_n N_A1_c_335_n 6.8319e-19 $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_230 A0 N_A1_c_335_n 0.021522f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_231 A0 N_A1_c_335_n 0.0275376f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_232 N_A0_c_282_n N_A1_c_335_n 2.23372e-19 $X=2.015 $Y=0.93 $X2=0 $Y2=0
cc_233 N_A0_c_278_n N_A1_c_336_n 6.48195e-19 $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_234 A0 N_A1_c_336_n 0.00146939f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_235 A0 A1 3.28495e-19 $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A0_c_278_n N_A1_c_338_n 0.00130352f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_237 A0 N_A1_c_338_n 0.0178287f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_238 N_A0_c_278_n N_S_c_386_n 0.0498601f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_239 N_A0_c_278_n S 3.48231e-19 $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_240 A0 S 0.0192152f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_241 N_A0_c_278_n N_S_c_384_n 0.0306561f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_242 A0 N_S_c_384_n 0.00262612f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_243 N_A0_c_278_n N_VPWR_c_435_n 0.00519092f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_244 N_A0_c_278_n N_VPWR_c_429_n 0.00690099f $X=2.94 $Y=1.77 $X2=0 $Y2=0
cc_245 N_A0_c_283_n N_VGND_c_523_n 0.00359964f $X=2.015 $Y=0.765 $X2=0 $Y2=0
cc_246 A0 N_VGND_c_527_n 0.00241884f $X=1.985 $Y=0.765 $X2=0 $Y2=0
cc_247 N_A0_c_283_n N_VGND_c_527_n 0.00556941f $X=2.015 $Y=0.765 $X2=0 $Y2=0
cc_248 N_A1_c_336_n N_S_M1005_g 0.0053243f $X=2.615 $Y=0.94 $X2=0 $Y2=0
cc_249 A1 N_S_M1005_g 0.00991405f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_250 N_A1_c_338_n N_S_M1005_g 0.00383702f $X=2.972 $Y=0.775 $X2=0 $Y2=0
cc_251 N_A1_c_336_n S 2.05559e-19 $X=2.615 $Y=0.94 $X2=0 $Y2=0
cc_252 A1 S 9.82443e-19 $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_253 N_A1_c_338_n S 0.0181332f $X=2.972 $Y=0.775 $X2=0 $Y2=0
cc_254 N_A1_c_334_n N_S_c_384_n 0.0048084f $X=2.46 $Y=1.67 $X2=0 $Y2=0
cc_255 N_A1_c_340_n N_VPWR_c_435_n 0.00439333f $X=2.46 $Y=1.77 $X2=0 $Y2=0
cc_256 N_A1_c_340_n N_VPWR_c_429_n 0.00746349f $X=2.46 $Y=1.77 $X2=0 $Y2=0
cc_257 A1 N_VGND_c_522_n 0.00642214f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_258 N_A1_M1007_g N_VGND_c_523_n 0.00585385f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_259 A1 N_VGND_c_523_n 0.00685317f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_260 N_A1_M1007_g N_VGND_c_527_n 0.0122806f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_261 N_A1_c_335_n N_VGND_c_527_n 0.013115f $X=2.87 $Y=0.94 $X2=0 $Y2=0
cc_262 N_A1_c_336_n N_VGND_c_527_n 5.19133e-19 $X=2.615 $Y=0.94 $X2=0 $Y2=0
cc_263 A1 N_VGND_c_527_n 0.00711001f $X=2.905 $Y=0.425 $X2=0 $Y2=0
cc_264 A1 A_502_47# 0.011663f $X=2.905 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_265 N_S_c_386_n N_VPWR_c_434_n 0.00296873f $X=3.35 $Y=1.77 $X2=0 $Y2=0
cc_266 N_S_c_388_n N_VPWR_c_434_n 0.0028008f $X=3.82 $Y=1.77 $X2=0 $Y2=0
cc_267 N_S_c_386_n N_VPWR_c_435_n 0.00523784f $X=3.35 $Y=1.77 $X2=0 $Y2=0
cc_268 N_S_c_388_n N_VPWR_c_437_n 0.00493774f $X=3.82 $Y=1.77 $X2=0 $Y2=0
cc_269 N_S_c_386_n N_VPWR_c_429_n 0.00670171f $X=3.35 $Y=1.77 $X2=0 $Y2=0
cc_270 N_S_c_388_n N_VPWR_c_429_n 0.0076238f $X=3.82 $Y=1.77 $X2=0 $Y2=0
cc_271 N_S_M1005_g N_VGND_c_522_n 0.00726003f $X=3.325 $Y=0.445 $X2=0 $Y2=0
cc_272 N_S_M1013_g N_VGND_c_522_n 0.00451902f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_273 S N_VGND_c_522_n 0.00514911f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_274 N_S_c_384_n N_VGND_c_522_n 0.00504552f $X=3.845 $Y=1.16 $X2=0 $Y2=0
cc_275 N_S_M1005_g N_VGND_c_523_n 0.0054325f $X=3.325 $Y=0.445 $X2=0 $Y2=0
cc_276 S N_VGND_c_523_n 0.00197279f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_277 N_S_M1013_g N_VGND_c_526_n 0.00585385f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_278 N_S_M1005_g N_VGND_c_527_n 0.0109898f $X=3.325 $Y=0.445 $X2=0 $Y2=0
cc_279 N_S_M1013_g N_VGND_c_527_n 0.012005f $X=3.845 $Y=0.445 $X2=0 $Y2=0
cc_280 S N_VGND_c_527_n 0.00357008f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_281 N_VPWR_c_429_n N_X_M1000_s 0.00231261f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_431_n N_X_c_490_n 0.074106f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_283 N_VPWR_c_432_n X 0.0210575f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_433_n X 0.0177667f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_285 N_VPWR_c_429_n X 0.0133992f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_429_n A_318_369# 0.00640407f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_287 N_VPWR_c_429_n A_606_369# 0.00295606f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_288 N_VPWR_c_431_n N_VGND_c_521_n 0.00878083f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_289 N_X_c_490_n N_VGND_c_525_n 0.0178201f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_290 N_X_M1006_s N_VGND_c_527_n 0.00481003f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_291 N_X_c_490_n N_VGND_c_527_n 0.0106938f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_292 N_X_c_490_n N_VGND_c_528_n 0.0152614f $X=0.715 $Y=0.42 $X2=0 $Y2=0
cc_293 N_VGND_c_527_n A_310_47# 0.00264621f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_294 N_VGND_c_527_n A_502_47# 0.0144818f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
