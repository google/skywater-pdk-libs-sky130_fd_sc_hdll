* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__einvp_8 A TE VGND VNB VPB VPWR Z
X0 Z A a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_213_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Z A a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_27_47# a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X4 a_213_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_47# TE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 Z A a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_213_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Z A a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_27_47# a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X10 a_235_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_213_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_235_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X13 VGND TE a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 Z A a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_235_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_213_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_235_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X18 Z A a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND TE a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR a_27_47# a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X21 a_213_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND TE a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Z A a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 VPWR a_27_47# a_235_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X25 a_235_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 Z A a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_235_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X28 VGND TE a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# TE VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_213_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_235_309# A Z VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_235_309# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X33 a_213_47# A Z VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
