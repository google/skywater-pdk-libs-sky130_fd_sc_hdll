* File: sky130_fd_sc_hdll__nand3b_2.spice
* Created: Thu Aug 27 19:14:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand3b_2.pex.spice"
.subckt sky130_fd_sc_hdll__nand3b_2  VNB VPB A_N C B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* C	C
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1013 N_VGND_M1013_d N_A_N_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.102252 AS=0.1092 PD=0.859626 PS=1.36 NRD=32.136 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1013_d N_C_M1000_g N_A_228_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.158248 AS=0.12025 PD=1.33037 PS=1.02 NRD=10.152 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_C_M1007_g N_A_228_47#_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_448_47#_M1004_d N_B_M1004_g N_A_228_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_A_448_47#_M1005_d N_B_M1005_g N_A_228_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_A_27_47#_M1001_g N_A_448_47#_M1005_d VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_Y_M1001_d N_A_27_47#_M1010_g N_A_448_47#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_N_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.108165 AS=0.1134 PD=0.837042 PS=1.38 NRD=34.0022 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1002_d N_C_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.257535
+ AS=0.145 PD=1.99296 PS=1.29 NRD=12.7853 NRS=0.9653 M=1 R=5.55556 SA=90000.5
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_C_M1011_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.9
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1003_d N_B_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_27_47#_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_47#_M1009_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_35 VNB 0 9.80354e-20 $X=0.15 $Y=-0.085
*
.include "sky130_fd_sc_hdll__nand3b_2.pxi.spice"
*
.ends
*
*
