* File: sky130_fd_sc_hdll__sdfstp_4.pxi.spice
* Created: Wed Sep  2 08:51:58 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCD N_SCD_c_280_n N_SCD_c_284_n N_SCD_c_285_n
+ N_SCD_M1010_g N_SCD_c_281_n N_SCD_M1027_g SCD SCD
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCD
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCE N_SCE_M1037_g N_SCE_c_320_n N_SCE_c_321_n
+ N_SCE_M1039_g N_SCE_c_322_n N_SCE_c_323_n N_SCE_M1014_g N_SCE_M1007_g
+ N_SCE_c_315_n N_SCE_c_335_n N_SCE_c_360_p SCE N_SCE_c_316_n N_SCE_c_317_n
+ N_SCE_c_318_n N_SCE_c_319_n SCE PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCE
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%D N_D_c_423_n N_D_c_428_n N_D_M1041_g
+ N_D_M1035_g D D N_D_c_425_n N_D_c_426_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%D
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_349_21# N_A_349_21#_M1007_s
+ N_A_349_21#_M1014_s N_A_349_21#_M1001_g N_A_349_21#_c_478_n
+ N_A_349_21#_c_479_n N_A_349_21#_M1026_g N_A_349_21#_c_473_n
+ N_A_349_21#_c_474_n N_A_349_21#_c_475_n N_A_349_21#_c_476_n
+ N_A_349_21#_c_477_n N_A_349_21#_c_483_n N_A_349_21#_c_484_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_349_21#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%CLK N_CLK_M1044_g N_CLK_c_551_n N_CLK_M1021_g
+ N_CLK_c_552_n N_CLK_c_556_n N_CLK_c_557_n CLK N_CLK_c_553_n N_CLK_c_554_n
+ N_CLK_c_555_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%CLK
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_693_369# N_A_693_369#_M1021_s
+ N_A_693_369#_M1044_s N_A_693_369#_c_626_n N_A_693_369#_c_627_n
+ N_A_693_369#_M1031_g N_A_693_369#_c_609_n N_A_693_369#_M1018_g
+ N_A_693_369#_c_610_n N_A_693_369#_c_611_n N_A_693_369#_M1033_g
+ N_A_693_369#_c_628_n N_A_693_369#_M1042_g N_A_693_369#_c_629_n
+ N_A_693_369#_c_630_n N_A_693_369#_M1034_g N_A_693_369#_M1005_g
+ N_A_693_369#_c_613_n N_A_693_369#_c_642_n N_A_693_369#_c_614_n
+ N_A_693_369#_c_631_n N_A_693_369#_c_632_n N_A_693_369#_c_615_n
+ N_A_693_369#_c_616_n N_A_693_369#_c_707_p N_A_693_369#_c_617_n
+ N_A_693_369#_c_618_n N_A_693_369#_c_619_n N_A_693_369#_c_620_n
+ N_A_693_369#_c_621_n N_A_693_369#_c_622_n N_A_693_369#_c_623_n
+ N_A_693_369#_c_698_p N_A_693_369#_c_637_n N_A_693_369#_c_638_n
+ N_A_693_369#_c_639_n N_A_693_369#_c_640_n N_A_693_369#_c_751_p
+ N_A_693_369#_c_624_n N_A_693_369#_c_641_n N_A_693_369#_c_625_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_693_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_877_369# N_A_877_369#_M1018_d
+ N_A_877_369#_M1031_d N_A_877_369#_c_905_n N_A_877_369#_c_894_n
+ N_A_877_369#_c_906_n N_A_877_369#_c_907_n N_A_877_369#_c_908_n
+ N_A_877_369#_M1008_g N_A_877_369#_M1028_g N_A_877_369#_M1045_g
+ N_A_877_369#_c_910_n N_A_877_369#_M1006_g N_A_877_369#_c_897_n
+ N_A_877_369#_c_911_n N_A_877_369#_c_912_n N_A_877_369#_c_898_n
+ N_A_877_369#_c_899_n N_A_877_369#_c_900_n N_A_877_369#_c_901_n
+ N_A_877_369#_c_902_n N_A_877_369#_c_903_n N_A_877_369#_c_904_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_877_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1229_21# N_A_1229_21#_M1024_s
+ N_A_1229_21#_M1011_d N_A_1229_21#_M1019_g N_A_1229_21#_c_1078_n
+ N_A_1229_21#_c_1084_n N_A_1229_21#_M1043_g N_A_1229_21#_c_1085_n
+ N_A_1229_21#_c_1079_n N_A_1229_21#_c_1086_n N_A_1229_21#_c_1087_n
+ N_A_1229_21#_c_1080_n N_A_1229_21#_c_1140_p N_A_1229_21#_c_1081_n
+ N_A_1229_21#_c_1082_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1229_21#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1075_413# N_A_1075_413#_M1033_d
+ N_A_1075_413#_M1008_d N_A_1075_413#_c_1172_n N_A_1075_413#_c_1183_n
+ N_A_1075_413#_c_1184_n N_A_1075_413#_M1011_g N_A_1075_413#_c_1173_n
+ N_A_1075_413#_M1024_g N_A_1075_413#_M1023_g N_A_1075_413#_c_1185_n
+ N_A_1075_413#_c_1186_n N_A_1075_413#_M1032_g N_A_1075_413#_c_1174_n
+ N_A_1075_413#_c_1202_n N_A_1075_413#_c_1175_n N_A_1075_413#_c_1187_n
+ N_A_1075_413#_c_1176_n N_A_1075_413#_c_1177_n N_A_1075_413#_c_1178_n
+ N_A_1075_413#_c_1179_n N_A_1075_413#_c_1180_n N_A_1075_413#_c_1181_n
+ N_A_1075_413#_c_1182_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1075_413#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%SET_B N_SET_B_c_1329_n N_SET_B_c_1330_n
+ N_SET_B_M1000_g N_SET_B_M1017_g N_SET_B_c_1331_n N_SET_B_M1003_g
+ N_SET_B_M1015_g N_SET_B_c_1328_n N_SET_B_c_1334_n N_SET_B_c_1335_n
+ N_SET_B_c_1336_n N_SET_B_c_1337_n N_SET_B_c_1338_n SET_B N_SET_B_c_1339_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%SET_B
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1951_295# N_A_1951_295#_M1022_d
+ N_A_1951_295#_M1004_d N_A_1951_295#_c_1463_n N_A_1951_295#_c_1464_n
+ N_A_1951_295#_M1020_g N_A_1951_295#_c_1465_n N_A_1951_295#_c_1466_n
+ N_A_1951_295#_M1002_g N_A_1951_295#_c_1456_n N_A_1951_295#_c_1457_n
+ N_A_1951_295#_c_1458_n N_A_1951_295#_c_1459_n N_A_1951_295#_c_1469_n
+ N_A_1951_295#_c_1470_n N_A_1951_295#_c_1460_n N_A_1951_295#_c_1461_n
+ N_A_1951_295#_c_1462_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1951_295#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1745_329# N_A_1745_329#_M1045_d
+ N_A_1745_329#_M1034_d N_A_1745_329#_M1003_d N_A_1745_329#_M1022_g
+ N_A_1745_329#_c_1557_n N_A_1745_329#_M1004_g N_A_1745_329#_c_1558_n
+ N_A_1745_329#_c_1569_n N_A_1745_329#_M1040_g N_A_1745_329#_M1030_g
+ N_A_1745_329#_c_1560_n N_A_1745_329#_c_1561_n N_A_1745_329#_c_1562_n
+ N_A_1745_329#_c_1578_n N_A_1745_329#_c_1579_n N_A_1745_329#_c_1571_n
+ N_A_1745_329#_c_1563_n N_A_1745_329#_c_1564_n N_A_1745_329#_c_1565_n
+ N_A_1745_329#_c_1566_n N_A_1745_329#_c_1572_n N_A_1745_329#_c_1573_n
+ N_A_1745_329#_c_1574_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1745_329#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_2447_47# N_A_2447_47#_M1030_s
+ N_A_2447_47#_M1040_s N_A_2447_47#_c_1705_n N_A_2447_47#_M1012_g
+ N_A_2447_47#_c_1697_n N_A_2447_47#_M1009_g N_A_2447_47#_c_1706_n
+ N_A_2447_47#_M1016_g N_A_2447_47#_c_1698_n N_A_2447_47#_M1013_g
+ N_A_2447_47#_c_1707_n N_A_2447_47#_M1025_g N_A_2447_47#_c_1699_n
+ N_A_2447_47#_M1036_g N_A_2447_47#_c_1708_n N_A_2447_47#_M1029_g
+ N_A_2447_47#_c_1700_n N_A_2447_47#_M1038_g N_A_2447_47#_c_1701_n
+ N_A_2447_47#_c_1709_n N_A_2447_47#_c_1702_n N_A_2447_47#_c_1703_n
+ N_A_2447_47#_c_1704_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_2447_47#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_27_369# N_A_27_369#_M1010_s
+ N_A_27_369#_M1026_d N_A_27_369#_c_1796_n N_A_27_369#_c_1797_n
+ N_A_27_369#_c_1798_n N_A_27_369#_c_1813_n N_A_27_369#_c_1810_n
+ N_A_27_369#_c_1799_n PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_27_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%VPWR N_VPWR_M1010_d N_VPWR_M1014_d
+ N_VPWR_M1044_d N_VPWR_M1043_d N_VPWR_M1000_d N_VPWR_M1020_d N_VPWR_M1004_s
+ N_VPWR_M1040_d N_VPWR_M1016_s N_VPWR_M1029_s N_VPWR_c_1843_n N_VPWR_c_1844_n
+ N_VPWR_c_1845_n N_VPWR_c_1846_n N_VPWR_c_1847_n N_VPWR_c_1848_n
+ N_VPWR_c_1849_n N_VPWR_c_1850_n N_VPWR_c_1851_n N_VPWR_c_1852_n
+ N_VPWR_c_1853_n N_VPWR_c_1854_n N_VPWR_c_1855_n N_VPWR_c_1856_n
+ N_VPWR_c_1857_n VPWR N_VPWR_c_1858_n N_VPWR_c_1859_n N_VPWR_c_1860_n
+ N_VPWR_c_1861_n N_VPWR_c_1862_n N_VPWR_c_1863_n N_VPWR_c_1864_n
+ N_VPWR_c_1865_n N_VPWR_c_1866_n N_VPWR_c_1867_n N_VPWR_c_1868_n
+ N_VPWR_c_1869_n N_VPWR_c_1870_n N_VPWR_c_1871_n N_VPWR_c_1842_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_201_47# N_A_201_47#_M1037_d
+ N_A_201_47#_M1033_s N_A_201_47#_M1041_d N_A_201_47#_M1008_s
+ N_A_201_47#_c_2068_n N_A_201_47#_c_2057_n N_A_201_47#_c_2061_n
+ N_A_201_47#_c_2062_n N_A_201_47#_c_2071_n N_A_201_47#_c_2058_n
+ N_A_201_47#_c_2063_n N_A_201_47#_c_2064_n N_A_201_47#_c_2059_n
+ N_A_201_47#_c_2066_n N_A_201_47#_c_2060_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_201_47#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%Q N_Q_M1009_s N_Q_M1036_s N_Q_M1012_d
+ N_Q_M1025_d N_Q_c_2195_n N_Q_c_2197_n N_Q_c_2199_n N_Q_c_2193_n N_Q_c_2204_n
+ N_Q_c_2194_n N_Q_c_2210_n Q Q Q Q Q Q Q N_Q_c_2217_n Q N_Q_c_2218_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%Q
x_PM_SKY130_FD_SC_HDLL__SDFSTP_4%VGND N_VGND_M1027_s N_VGND_M1001_d
+ N_VGND_M1007_d N_VGND_M1021_d N_VGND_M1019_d N_VGND_M1017_d N_VGND_M1015_d
+ N_VGND_M1030_d N_VGND_M1013_d N_VGND_M1038_d N_VGND_c_2242_n N_VGND_c_2243_n
+ N_VGND_c_2244_n N_VGND_c_2245_n N_VGND_c_2246_n N_VGND_c_2247_n
+ N_VGND_c_2248_n N_VGND_c_2249_n N_VGND_c_2250_n N_VGND_c_2251_n
+ N_VGND_c_2252_n N_VGND_c_2253_n N_VGND_c_2254_n N_VGND_c_2255_n
+ N_VGND_c_2256_n VGND N_VGND_c_2257_n N_VGND_c_2258_n N_VGND_c_2259_n
+ N_VGND_c_2260_n N_VGND_c_2261_n N_VGND_c_2262_n N_VGND_c_2263_n
+ N_VGND_c_2264_n N_VGND_c_2265_n N_VGND_c_2266_n N_VGND_c_2267_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_4%VGND
cc_1 VNB N_SCD_c_280_n 0.0614876f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_2 VNB N_SCD_c_281_n 0.017667f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB SCD 0.0208496f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_SCE_M1037_g 0.0333651f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.77
cc_5 VNB N_SCE_M1007_g 0.0386452f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_6 VNB N_SCE_c_315_n 0.00641659f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_7 VNB N_SCE_c_316_n 0.0221836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_317_n 0.0327362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_318_n 0.00121258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_319_n 0.0063767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_c_423_n 0.00973242f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.62
cc_12 VNB D 0.00603948f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_13 VNB N_D_c_425_n 0.0284342f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_14 VNB N_D_c_426_n 0.0169241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_349_21#_M1001_g 0.030387f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_16 VNB N_A_349_21#_c_473_n 0.013066f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_17 VNB N_A_349_21#_c_474_n 0.00449025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_349_21#_c_475_n 0.0322814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_349_21#_c_476_n 0.0144986f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_20 VNB N_A_349_21#_c_477_n 0.00694339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_CLK_c_551_n 0.0175885f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_22 VNB N_CLK_c_552_n 0.0179572f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_23 VNB N_CLK_c_553_n 0.0169771f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_24 VNB N_CLK_c_554_n 0.016278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_CLK_c_555_n 0.0139632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_693_369#_c_609_n 0.0177594f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_27 VNB N_A_693_369#_c_610_n 0.0561083f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_28 VNB N_A_693_369#_c_611_n 0.0178231f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_29 VNB N_A_693_369#_M1005_g 0.0255213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_693_369#_c_613_n 0.0083546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_693_369#_c_614_n 0.00135304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_693_369#_c_615_n 0.00796372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_693_369#_c_616_n 0.0036336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_693_369#_c_617_n 0.00345628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_693_369#_c_618_n 0.0175281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_693_369#_c_619_n 0.00398691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_693_369#_c_620_n 0.028498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_693_369#_c_621_n 0.0104486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_693_369#_c_622_n 3.84112e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_693_369#_c_623_n 0.00472385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_693_369#_c_624_n 0.012173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_693_369#_c_625_n 0.0328018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_877_369#_c_894_n 0.0497739f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_44 VNB N_A_877_369#_M1028_g 0.0325688f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_45 VNB N_A_877_369#_M1045_g 0.0382341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_877_369#_c_897_n 0.00471247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_877_369#_c_898_n 0.0210013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_877_369#_c_899_n 5.03783e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_877_369#_c_900_n 0.00418782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_877_369#_c_901_n 0.00304349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_877_369#_c_902_n 0.00332697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_877_369#_c_903_n 0.00274772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_877_369#_c_904_n 0.017185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1229_21#_M1019_g 0.0191216f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_55 VNB N_A_1229_21#_c_1078_n 0.0139193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1229_21#_c_1079_n 0.0078726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1229_21#_c_1080_n 0.00452229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1229_21#_c_1081_n 0.0031057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1229_21#_c_1082_n 0.028204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1075_413#_c_1172_n 0.0139262f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_61 VNB N_A_1075_413#_c_1173_n 0.0164466f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.445
cc_62 VNB N_A_1075_413#_c_1174_n 0.0269257f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1075_413#_c_1175_n 0.0097997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1075_413#_c_1176_n 0.00369281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1075_413#_c_1177_n 0.0171906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1075_413#_c_1178_n 0.00204312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1075_413#_c_1179_n 0.00232092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1075_413#_c_1180_n 0.0249427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1075_413#_c_1181_n 0.0207836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1075_413#_c_1182_n 0.0196761f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_SET_B_M1017_g 0.0384509f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_72 VNB N_SET_B_M1015_g 0.0463357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_SET_B_c_1328_n 0.00805659f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_74 VNB N_A_1951_295#_M1002_g 0.0227251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1951_295#_c_1456_n 0.00746573f $X=-0.19 $Y=-0.24 $X2=0.255
+ $Y2=1.16
cc_76 VNB N_A_1951_295#_c_1457_n 0.0017077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1951_295#_c_1458_n 0.0316179f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_78 VNB N_A_1951_295#_c_1459_n 0.0108982f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1951_295#_c_1460_n 0.0122378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1951_295#_c_1461_n 0.00338281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1951_295#_c_1462_n 5.02844e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1745_329#_c_1557_n 0.00690736f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=0.765
cc_83 VNB N_A_1745_329#_c_1558_n 0.0328925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1745_329#_M1030_g 0.0312677f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_85 VNB N_A_1745_329#_c_1560_n 0.0170554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1745_329#_c_1561_n 0.0211706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1745_329#_c_1562_n 0.0031377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1745_329#_c_1563_n 0.00150402f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1745_329#_c_1564_n 0.00281159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1745_329#_c_1565_n 0.0100396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1745_329#_c_1566_n 0.0216888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2447_47#_c_1697_n 0.0176056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_2447_47#_c_1698_n 0.0169271f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_2447_47#_c_1699_n 0.0169253f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2447_47#_c_1700_n 0.0219834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_2447_47#_c_1701_n 0.00886299f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_A_2447_47#_c_1702_n 0.00563715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_2447_47#_c_1703_n 0.00180143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_A_2447_47#_c_1704_n 0.0970391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VPWR_c_1842_n 0.6303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_201_47#_c_2057_n 0.00432851f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_102 VNB N_A_201_47#_c_2058_n 0.00130739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_201_47#_c_2059_n 0.00392628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_201_47#_c_2060_n 0.00439899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_Q_c_2193_n 0.00106334f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_2242_n 0.0312931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2243_n 0.0352326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2244_n 0.00803967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2245_n 0.0164899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2246_n 0.00820979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2247_n 0.0027219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2248_n 0.00518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2249_n 0.00294656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2250_n 0.00570514f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2251_n 0.0113479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2252_n 0.0354721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2253_n 0.0146232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2254_n 0.00507625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2255_n 0.0214718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2256_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2257_n 0.0619169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2258_n 0.0698374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2259_n 0.031469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2260_n 0.0212612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2261_n 0.00506925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2262_n 0.00664466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2263_n 0.0167152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2264_n 0.0202344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2265_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2266_n 0.00625144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2267_n 0.700812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VPB N_SCD_c_280_n 0.00540609f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.325
cc_133 VPB N_SCD_c_284_n 0.0175267f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_134 VPB N_SCD_c_285_n 0.0494007f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_135 VPB SCD 0.0148037f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_136 VPB N_SCE_c_320_n 0.0133941f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_137 VPB N_SCE_c_321_n 0.0221672f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_138 VPB N_SCE_c_322_n 0.026286f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_139 VPB N_SCE_c_323_n 0.0343446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_SCE_c_316_n 0.0134821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_SCE_c_317_n 0.00642596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_SCE_c_318_n 0.00419291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_SCE_c_319_n 0.00484581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_D_c_423_n 0.0161429f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_145 VPB N_D_c_428_n 0.0222417f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_146 VPB D 0.0044569f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.695
cc_147 VPB N_A_349_21#_c_478_n 0.0220272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_349_21#_c_479_n 0.0251734f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_149 VPB N_A_349_21#_c_473_n 6.82321e-19 $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_150 VPB N_A_349_21#_c_474_n 0.0101942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_349_21#_c_475_n 0.0147247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_349_21#_c_483_n 0.00409949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_349_21#_c_484_n 0.0122482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_CLK_c_556_n 0.0121836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_CLK_c_557_n 0.040301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_CLK_c_553_n 0.0107275f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_157 VPB N_CLK_c_554_n 0.0204466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_693_369#_c_626_n 0.0149449f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_159 VPB N_A_693_369#_c_627_n 0.0251151f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.695
cc_160 VPB N_A_693_369#_c_628_n 0.0571336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_693_369#_c_629_n 0.0075279f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_693_369#_c_630_n 0.0208038f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_693_369#_c_631_n 0.0015983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_693_369#_c_632_n 0.00133399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_693_369#_c_617_n 0.00372107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_693_369#_c_618_n 0.0107422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_693_369#_c_619_n 0.00221239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_693_369#_c_620_n 0.00464409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_693_369#_c_637_n 0.00671353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_693_369#_c_638_n 3.87498e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_693_369#_c_639_n 0.00813324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_693_369#_c_640_n 0.0022021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_693_369#_c_641_n 0.00224736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_877_369#_c_905_n 0.0246271f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_175 VPB N_A_877_369#_c_906_n 0.0201586f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_176 VPB N_A_877_369#_c_907_n 0.0107019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_877_369#_c_908_n 0.0193133f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_178 VPB N_A_877_369#_M1045_g 0.0160839f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_877_369#_c_910_n 0.0701221f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.53
cc_180 VPB N_A_877_369#_c_911_n 0.004892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_877_369#_c_912_n 0.00997068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_A_877_369#_c_900_n 3.90977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_877_369#_c_901_n 0.00411878f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_877_369#_c_902_n 0.00122725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_877_369#_c_904_n 0.0170356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1229_21#_c_1078_n 0.0183639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_1229_21#_c_1084_n 0.064302f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_188 VPB N_A_1229_21#_c_1085_n 0.00179081f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_189 VPB N_A_1229_21#_c_1086_n 0.00606886f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.16
cc_190 VPB N_A_1229_21#_c_1087_n 7.95296e-19 $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_191 VPB N_A_1075_413#_c_1183_n 0.0317517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1075_413#_c_1184_n 0.0242898f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_193 VPB N_A_1075_413#_c_1185_n 0.0087284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1075_413#_c_1186_n 0.0214701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_A_1075_413#_c_1187_n 0.0165451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_A_1075_413#_c_1176_n 0.00646138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_A_1075_413#_c_1177_n 0.00210333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1075_413#_c_1178_n 0.0035338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1075_413#_c_1179_n 0.00131078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1075_413#_c_1180_n 0.00611954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1075_413#_c_1181_n 0.00983399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_1329_n 0.00905299f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_203 VPB N_SET_B_c_1330_n 0.0586682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_204 VPB N_SET_B_c_1331_n 0.0824845f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_SET_B_M1015_g 0.00888602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_SET_B_c_1328_n 0.00588959f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_207 VPB N_SET_B_c_1334_n 0.00856385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_1335_n 0.0140309f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.53
cc_209 VPB N_SET_B_c_1336_n 0.00241098f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_SET_B_c_1337_n 0.00604378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_SET_B_c_1338_n 0.00461355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_SET_B_c_1339_n 0.00985551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1951_295#_c_1463_n 0.0163304f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_214 VPB N_A_1951_295#_c_1464_n 0.0235005f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.695
cc_215 VPB N_A_1951_295#_c_1465_n 0.0295115f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1951_295#_c_1466_n 0.00792272f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_217 VPB N_A_1951_295#_c_1456_n 0.0123394f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_218 VPB N_A_1951_295#_c_1459_n 0.00760355f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1951_295#_c_1469_n 8.64549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1951_295#_c_1470_n 0.0187938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1745_329#_c_1557_n 0.0895167f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_222 VPB N_A_1745_329#_c_1558_n 0.0311166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1745_329#_c_1569_n 0.0192434f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_224 VPB N_A_1745_329#_c_1562_n 0.00623807f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1745_329#_c_1571_n 0.0150869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1745_329#_c_1572_n 0.00615721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_A_1745_329#_c_1573_n 0.00240612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1745_329#_c_1574_n 0.001738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_A_2447_47#_c_1705_n 0.0168351f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_230 VPB N_A_2447_47#_c_1706_n 0.0163246f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_231 VPB N_A_2447_47#_c_1707_n 0.0163246f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_232 VPB N_A_2447_47#_c_1708_n 0.0207521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_2447_47#_c_1709_n 0.0112297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_2447_47#_c_1702_n 0.00194757f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_2447_47#_c_1704_n 0.0604615f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_27_369#_c_1796_n 0.0170416f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_237 VPB N_A_27_369#_c_1797_n 0.00100316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_27_369#_c_1798_n 0.00945761f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_239 VPB N_A_27_369#_c_1799_n 0.00263317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1843_n 0.00252882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1844_n 0.00907525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1845_n 0.0164751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1846_n 0.0049533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1847_n 0.00925213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1848_n 0.00586716f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1849_n 0.0190443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1850_n 0.00567316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1851_n 0.00300019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1852_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1853_n 0.011322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1854_n 0.0453984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1855_n 0.0240535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1856_n 0.0214427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1857_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1858_n 0.0143786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1859_n 0.0512333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1860_n 0.0566134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1861_n 0.03085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1862_n 0.0257651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1863_n 0.0212612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1864_n 0.00464622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1865_n 0.00564769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1866_n 0.00547148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1867_n 0.0133607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1868_n 0.00644418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1869_n 0.00727646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1870_n 0.005797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1871_n 0.00628472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1842_n 0.0727137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_A_201_47#_c_2061_n 8.90825e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_A_201_47#_c_2062_n 0.00245242f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_272 VPB N_A_201_47#_c_2063_n 0.025058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_A_201_47#_c_2064_n 0.0031429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_A_201_47#_c_2059_n 0.00330318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_A_201_47#_c_2066_n 0.00776824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_A_201_47#_c_2060_n 0.00386251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_Q_c_2194_n 0.00154101f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 N_SCD_c_280_n N_SCE_M1037_g 0.00227875f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_279 N_SCD_c_281_n N_SCE_M1037_g 0.0377993f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_280 SCD N_SCE_M1037_g 3.82641e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_281 N_SCD_c_284_n N_SCE_c_320_n 0.00212959f $X=0.315 $Y=1.62 $X2=0 $Y2=0
cc_282 N_SCD_c_285_n N_SCE_c_320_n 0.00802922f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_283 SCD N_SCE_c_320_n 3.4065e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_284 N_SCD_c_285_n N_SCE_c_321_n 0.0232945f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_285 SCD N_SCE_c_335_n 0.00144346f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_286 N_SCD_c_280_n N_SCE_c_316_n 0.0152623f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_287 SCD N_SCE_c_316_n 3.22701e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_288 N_SCD_c_280_n N_SCE_c_319_n 0.0100034f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_289 N_SCD_c_285_n N_SCE_c_319_n 0.00381492f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_290 SCD N_SCE_c_319_n 0.0602867f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_291 N_SCD_c_285_n N_A_27_369#_c_1796_n 0.00843386f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_292 N_SCD_c_285_n N_A_27_369#_c_1797_n 0.0153318f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_293 N_SCD_c_280_n N_A_27_369#_c_1798_n 5.05332e-19 $X=0.315 $Y=1.325 $X2=0
+ $Y2=0
cc_294 N_SCD_c_285_n N_A_27_369#_c_1798_n 0.00332576f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_295 SCD N_A_27_369#_c_1798_n 0.0227399f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_296 N_SCD_c_285_n N_VPWR_c_1843_n 0.011563f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_297 N_SCD_c_285_n N_VPWR_c_1858_n 0.00317293f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_298 N_SCD_c_285_n N_VPWR_c_1842_n 0.0048112f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_299 N_SCD_c_281_n N_A_201_47#_c_2068_n 2.9719e-19 $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_300 N_SCD_c_280_n N_VGND_c_2243_n 0.00690102f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_301 N_SCD_c_281_n N_VGND_c_2243_n 0.0210021f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_302 SCD N_VGND_c_2243_n 0.0221805f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_303 SCD N_VGND_c_2267_n 9.88088e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_304 N_SCE_c_316_n N_D_c_423_n 0.0247422f $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_305 N_SCE_c_319_n N_D_c_423_n 4.55957e-19 $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_306 N_SCE_c_320_n N_D_c_428_n 0.016356f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_307 N_SCE_c_321_n N_D_c_428_n 0.0461727f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_308 N_SCE_M1037_g D 0.00355142f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_309 N_SCE_c_320_n D 0.00637589f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_310 N_SCE_c_321_n D 3.91386e-19 $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_311 N_SCE_c_315_n D 0.0313118f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_312 N_SCE_c_335_n D 0.00223888f $X=0.87 $Y=1.19 $X2=0 $Y2=0
cc_313 N_SCE_c_316_n D 0.00430657f $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_314 N_SCE_c_319_n D 0.0690236f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_315 N_SCE_M1037_g N_D_c_425_n 0.0192751f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_316 N_SCE_c_315_n N_D_c_425_n 0.00134139f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_317 N_SCE_c_319_n N_D_c_425_n 2.52791e-19 $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_318 N_SCE_M1037_g N_D_c_426_n 0.0134262f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_319 N_SCE_c_315_n N_A_349_21#_c_473_n 0.00480032f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_320 N_SCE_c_322_n N_A_349_21#_c_474_n 0.00674156f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_321 N_SCE_M1007_g N_A_349_21#_c_474_n 0.0025686f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_322 N_SCE_c_315_n N_A_349_21#_c_474_n 0.0173777f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_323 N_SCE_c_360_p N_A_349_21#_c_474_n 6.89964e-19 $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_324 N_SCE_c_317_n N_A_349_21#_c_474_n 0.00247942f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_325 N_SCE_c_318_n N_A_349_21#_c_474_n 0.0400811f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_326 N_SCE_c_315_n N_A_349_21#_c_475_n 0.0040858f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_327 N_SCE_c_317_n N_A_349_21#_c_475_n 0.0213661f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_328 N_SCE_c_318_n N_A_349_21#_c_475_n 7.19229e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_329 N_SCE_M1007_g N_A_349_21#_c_476_n 0.00827962f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_330 N_SCE_c_315_n N_A_349_21#_c_476_n 0.00905152f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_331 N_SCE_c_360_p N_A_349_21#_c_476_n 0.00104259f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_332 N_SCE_c_317_n N_A_349_21#_c_476_n 0.002964f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_333 N_SCE_c_318_n N_A_349_21#_c_476_n 0.00979853f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_SCE_M1007_g N_A_349_21#_c_477_n 0.00585491f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_335 N_SCE_c_323_n N_A_349_21#_c_484_n 0.00355437f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_336 N_SCE_c_317_n N_A_349_21#_c_484_n 4.82439e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_337 N_SCE_c_318_n N_A_349_21#_c_484_n 0.0105043f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_338 N_SCE_M1007_g N_CLK_c_552_n 0.00287881f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_339 N_SCE_c_322_n N_CLK_c_553_n 0.00124305f $X=2.835 $Y=1.67 $X2=0 $Y2=0
cc_340 N_SCE_c_317_n N_CLK_c_553_n 0.00331448f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_341 N_SCE_c_318_n N_CLK_c_553_n 3.6692e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_342 N_SCE_c_322_n N_CLK_c_554_n 0.00357902f $X=2.835 $Y=1.67 $X2=0 $Y2=0
cc_343 N_SCE_c_360_p N_CLK_c_554_n 0.00158915f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_344 N_SCE_c_317_n N_CLK_c_554_n 0.0033024f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_345 N_SCE_c_318_n N_CLK_c_554_n 0.0356601f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_346 N_SCE_c_317_n N_CLK_c_555_n 0.00287881f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_347 N_SCE_c_323_n N_A_693_369#_c_642_n 0.00347988f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_348 N_SCE_M1007_g N_A_693_369#_c_614_n 0.00346504f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_349 N_SCE_c_323_n N_A_693_369#_c_632_n 0.00464142f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_350 N_SCE_M1007_g N_A_693_369#_c_616_n 0.00350126f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_SCE_c_321_n N_A_27_369#_c_1797_n 0.0148547f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_352 N_SCE_c_315_n N_A_27_369#_c_1797_n 0.00494807f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_353 N_SCE_c_335_n N_A_27_369#_c_1797_n 0.00104089f $X=0.87 $Y=1.19 $X2=0
+ $Y2=0
cc_354 N_SCE_c_316_n N_A_27_369#_c_1797_n 7.84018e-19 $X=0.93 $Y=1.25 $X2=0
+ $Y2=0
cc_355 N_SCE_c_319_n N_A_27_369#_c_1797_n 0.0226263f $X=0.725 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_SCE_c_321_n N_A_27_369#_c_1810_n 0.00202367f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_357 N_SCE_c_321_n N_VPWR_c_1843_n 0.00296668f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_358 N_SCE_c_323_n N_VPWR_c_1844_n 0.0049892f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_359 N_SCE_c_321_n N_VPWR_c_1859_n 0.0052046f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_360 N_SCE_c_323_n N_VPWR_c_1859_n 0.00702461f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_361 N_SCE_c_321_n N_VPWR_c_1842_n 0.00671789f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_362 N_SCE_c_323_n N_VPWR_c_1842_n 0.0150885f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_363 N_SCE_M1037_g N_A_201_47#_c_2068_n 0.00782662f $X=0.93 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_SCE_c_315_n N_A_201_47#_c_2068_n 0.0112441f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_365 N_SCE_c_315_n N_A_201_47#_c_2071_n 0.00450485f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_366 N_SCE_c_322_n N_A_201_47#_c_2063_n 0.00811567f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_367 N_SCE_c_315_n N_A_201_47#_c_2063_n 0.0490896f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_SCE_c_360_p N_A_201_47#_c_2063_n 0.0249445f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_369 N_SCE_c_317_n N_A_201_47#_c_2063_n 4.55029e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_370 N_SCE_c_318_n N_A_201_47#_c_2063_n 0.0213105f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_371 N_SCE_c_315_n N_A_201_47#_c_2064_n 0.030535f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_372 N_SCE_c_315_n N_A_201_47#_c_2059_n 0.0185596f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_373 N_SCE_M1037_g N_VGND_c_2242_n 0.00456464f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_374 N_SCE_M1037_g N_VGND_c_2243_n 0.00569751f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_375 N_SCE_c_335_n N_VGND_c_2243_n 7.54179e-19 $X=0.87 $Y=1.19 $X2=0 $Y2=0
cc_376 N_SCE_c_316_n N_VGND_c_2243_n 3.94412e-19 $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_377 N_SCE_c_319_n N_VGND_c_2243_n 0.0152769f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_378 N_SCE_M1007_g N_VGND_c_2244_n 0.00178988f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_379 N_SCE_c_315_n N_VGND_c_2244_n 0.00127321f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_380 N_SCE_M1007_g N_VGND_c_2245_n 0.00486043f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_381 N_SCE_M1007_g N_VGND_c_2246_n 0.0100904f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_382 N_SCE_c_318_n N_VGND_c_2246_n 2.63385e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_383 N_SCE_M1037_g N_VGND_c_2267_n 0.00734604f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_384 N_SCE_M1007_g N_VGND_c_2267_n 0.00965187f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_385 N_SCE_c_319_n N_VGND_c_2267_n 0.00570024f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_386 D N_A_349_21#_M1001_g 3.18064e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_387 N_D_c_425_n N_A_349_21#_M1001_g 0.0203756f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_388 N_D_c_426_n N_A_349_21#_M1001_g 0.0310629f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_389 N_D_c_428_n N_A_349_21#_c_478_n 0.0157634f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_390 N_D_c_428_n N_A_349_21#_c_479_n 0.0234679f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_391 N_D_c_423_n N_A_349_21#_c_473_n 0.0157634f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_392 D N_A_349_21#_c_473_n 0.00160886f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_393 N_D_c_428_n N_A_27_369#_c_1797_n 0.00136438f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_394 D N_A_27_369#_c_1797_n 0.0137059f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_395 N_D_c_428_n N_A_27_369#_c_1813_n 0.00431987f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_396 N_D_c_428_n N_A_27_369#_c_1799_n 0.0135654f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_397 D N_A_27_369#_c_1799_n 0.00422562f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_398 N_D_c_428_n N_VPWR_c_1859_n 0.00429453f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_399 N_D_c_428_n N_VPWR_c_1842_n 0.0060009f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_400 D N_A_201_47#_c_2068_n 0.0313325f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_401 N_D_c_425_n N_A_201_47#_c_2068_n 0.00175893f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_402 N_D_c_426_n N_A_201_47#_c_2068_n 0.012197f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_403 N_D_c_428_n N_A_201_47#_c_2071_n 0.00519966f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_404 D N_A_201_47#_c_2071_n 0.00614145f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_405 D N_A_201_47#_c_2064_n 0.00778368f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_406 N_D_c_423_n N_A_201_47#_c_2059_n 0.00161643f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_407 N_D_c_428_n N_A_201_47#_c_2059_n 0.00355157f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_408 D N_A_201_47#_c_2059_n 0.0689424f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_409 N_D_c_425_n N_A_201_47#_c_2059_n 0.00193715f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_410 N_D_c_426_n N_A_201_47#_c_2059_n 0.00351003f $X=1.375 $Y=0.765 $X2=0
+ $Y2=0
cc_411 N_D_c_426_n N_VGND_c_2242_n 0.00357877f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_412 N_D_c_426_n N_VGND_c_2267_n 0.00539883f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_413 N_A_349_21#_c_484_n N_A_27_369#_M1026_d 0.00555261f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_414 N_A_349_21#_c_479_n N_A_27_369#_c_1799_n 0.011002f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_415 N_A_349_21#_c_483_n N_A_27_369#_c_1799_n 0.0148152f $X=2.595 $Y=1.927
+ $X2=0 $Y2=0
cc_416 N_A_349_21#_c_484_n N_A_27_369#_c_1799_n 0.0132953f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_417 N_A_349_21#_c_479_n N_VPWR_c_1859_n 0.00429453f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_418 N_A_349_21#_c_483_n N_VPWR_c_1859_n 0.0157393f $X=2.595 $Y=1.927 $X2=0
+ $Y2=0
cc_419 N_A_349_21#_c_484_n N_VPWR_c_1859_n 0.00432835f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_420 N_A_349_21#_M1014_s N_VPWR_c_1842_n 0.00304306f $X=2.475 $Y=1.845 $X2=0
+ $Y2=0
cc_421 N_A_349_21#_c_479_n N_VPWR_c_1842_n 0.00737353f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_422 N_A_349_21#_c_483_n N_VPWR_c_1842_n 0.00941222f $X=2.595 $Y=1.927 $X2=0
+ $Y2=0
cc_423 N_A_349_21#_c_484_n N_VPWR_c_1842_n 0.00699224f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_424 N_A_349_21#_M1001_g N_A_201_47#_c_2068_n 0.0106694f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_425 N_A_349_21#_c_477_n N_A_201_47#_c_2068_n 0.00154368f $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_426 N_A_349_21#_c_479_n N_A_201_47#_c_2071_n 0.00556528f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_427 N_A_349_21#_c_484_n N_A_201_47#_c_2071_n 0.0164794f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_428 N_A_349_21#_c_474_n N_A_201_47#_c_2063_n 0.0172766f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_429 N_A_349_21#_c_475_n N_A_201_47#_c_2063_n 0.00172463f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_430 N_A_349_21#_c_484_n N_A_201_47#_c_2063_n 0.0111897f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_431 N_A_349_21#_c_478_n N_A_201_47#_c_2064_n 0.00546081f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_432 N_A_349_21#_c_474_n N_A_201_47#_c_2064_n 0.00296292f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_433 N_A_349_21#_M1001_g N_A_201_47#_c_2059_n 0.00973696f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_434 N_A_349_21#_c_478_n N_A_201_47#_c_2059_n 0.0072174f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_435 N_A_349_21#_c_479_n N_A_201_47#_c_2059_n 0.00456775f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_436 N_A_349_21#_c_473_n N_A_201_47#_c_2059_n 0.00911472f $X=1.845 $Y=1.16
+ $X2=0 $Y2=0
cc_437 N_A_349_21#_c_474_n N_A_201_47#_c_2059_n 0.0488018f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_438 N_A_349_21#_c_476_n N_A_201_47#_c_2059_n 0.0125621f $X=2.59 $Y=0.715
+ $X2=0 $Y2=0
cc_439 N_A_349_21#_c_477_n N_A_201_47#_c_2059_n 0.00338006f $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_440 N_A_349_21#_c_484_n N_A_201_47#_c_2059_n 0.00494415f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_349_21#_M1001_g N_VGND_c_2242_n 0.00433573f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_442 N_A_349_21#_M1001_g N_VGND_c_2244_n 0.0105214f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_443 N_A_349_21#_c_475_n N_VGND_c_2244_n 0.00128608f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_444 N_A_349_21#_c_476_n N_VGND_c_2244_n 0.0174596f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_445 N_A_349_21#_c_477_n N_VGND_c_2244_n 0.0233257f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_446 N_A_349_21#_c_476_n N_VGND_c_2245_n 0.00268684f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_447 N_A_349_21#_c_477_n N_VGND_c_2245_n 0.0176923f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_448 N_A_349_21#_c_477_n N_VGND_c_2246_n 0.0190636f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_449 N_A_349_21#_M1007_s N_VGND_c_2267_n 0.00580108f $X=2.505 $Y=0.235 $X2=0
+ $Y2=0
cc_450 N_A_349_21#_M1001_g N_VGND_c_2267_n 0.00851845f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_451 N_A_349_21#_c_476_n N_VGND_c_2267_n 0.00551711f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_452 N_A_349_21#_c_477_n N_VGND_c_2267_n 0.00983733f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_453 N_CLK_c_556_n N_A_693_369#_c_626_n 0.0059319f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_454 N_CLK_c_557_n N_A_693_369#_c_626_n 0.00655864f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_455 N_CLK_c_554_n N_A_693_369#_c_626_n 3.04599e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_456 N_CLK_c_557_n N_A_693_369#_c_627_n 0.0222028f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_457 N_CLK_c_551_n N_A_693_369#_c_609_n 0.0116086f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_458 N_CLK_c_552_n N_A_693_369#_c_613_n 0.00767961f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_459 N_CLK_c_551_n N_A_693_369#_c_614_n 0.0056285f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_460 N_CLK_c_557_n N_A_693_369#_c_631_n 0.0161161f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_461 N_CLK_c_554_n N_A_693_369#_c_631_n 0.00934927f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_462 N_CLK_c_557_n N_A_693_369#_c_632_n 3.10042e-19 $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_463 N_CLK_c_553_n N_A_693_369#_c_632_n 5.4866e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_464 N_CLK_c_554_n N_A_693_369#_c_632_n 0.0133612f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_465 N_CLK_c_551_n N_A_693_369#_c_615_n 0.00401517f $X=3.88 $Y=0.73 $X2=0
+ $Y2=0
cc_466 N_CLK_c_552_n N_A_693_369#_c_615_n 0.00847863f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_467 N_CLK_c_554_n N_A_693_369#_c_615_n 0.00801255f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_468 N_CLK_c_555_n N_A_693_369#_c_615_n 0.00151794f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_469 N_CLK_c_552_n N_A_693_369#_c_616_n 0.00352145f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_470 N_CLK_c_553_n N_A_693_369#_c_616_n 8.54762e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_471 N_CLK_c_554_n N_A_693_369#_c_616_n 0.016187f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_472 N_CLK_c_555_n N_A_693_369#_c_616_n 5.61645e-19 $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_473 N_CLK_c_557_n N_A_693_369#_c_617_n 0.00461373f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_474 N_CLK_c_554_n N_A_693_369#_c_617_n 0.0379355f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_475 N_CLK_c_555_n N_A_693_369#_c_617_n 0.00572652f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_476 N_CLK_c_553_n N_A_693_369#_c_618_n 0.0164171f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_477 N_CLK_c_554_n N_A_693_369#_c_618_n 3.92042e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_478 N_CLK_c_555_n N_A_693_369#_c_624_n 0.0053784f $X=3.68 $Y=1.09 $X2=0 $Y2=0
cc_479 N_CLK_c_557_n N_VPWR_c_1844_n 0.00397623f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_480 N_CLK_c_554_n N_VPWR_c_1844_n 0.00278244f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_481 N_CLK_c_557_n N_VPWR_c_1845_n 0.00320592f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_482 N_CLK_c_557_n N_VPWR_c_1866_n 0.0111353f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_483 N_CLK_c_557_n N_VPWR_c_1842_n 0.00524235f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_484 N_CLK_c_556_n N_A_201_47#_c_2063_n 0.0011232f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_485 N_CLK_c_557_n N_A_201_47#_c_2063_n 0.00327618f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_486 N_CLK_c_554_n N_A_201_47#_c_2063_n 0.0533918f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_487 N_CLK_c_551_n N_VGND_c_2246_n 0.00207759f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_488 N_CLK_c_554_n N_VGND_c_2246_n 0.00829842f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_489 N_CLK_c_551_n N_VGND_c_2247_n 0.00817351f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_490 N_CLK_c_551_n N_VGND_c_2253_n 0.00348405f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_491 N_CLK_c_552_n N_VGND_c_2253_n 4.55781e-19 $X=3.88 $Y=0.805 $X2=0 $Y2=0
cc_492 N_CLK_c_551_n N_VGND_c_2267_n 0.00552264f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_493 N_A_693_369#_c_637_n N_A_877_369#_M1031_d 7.76593e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_494 N_A_693_369#_c_638_n N_A_877_369#_M1031_d 6.28941e-19 $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_495 N_A_693_369#_c_626_n N_A_877_369#_c_905_n 0.00683981f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_496 N_A_693_369#_c_627_n N_A_877_369#_c_905_n 0.0051976f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_497 N_A_693_369#_c_628_n N_A_877_369#_c_905_n 0.00286715f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_498 N_A_693_369#_c_637_n N_A_877_369#_c_905_n 0.00113464f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_499 N_A_693_369#_c_628_n N_A_877_369#_c_894_n 0.010354f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_500 N_A_693_369#_c_637_n N_A_877_369#_c_894_n 8.44234e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_501 N_A_693_369#_c_641_n N_A_877_369#_c_894_n 2.5741e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_502 N_A_693_369#_c_628_n N_A_877_369#_c_906_n 0.00899979f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_503 N_A_693_369#_c_637_n N_A_877_369#_c_906_n 0.00501369f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_504 N_A_693_369#_c_640_n N_A_877_369#_c_906_n 7.59275e-19 $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_505 N_A_693_369#_c_641_n N_A_877_369#_c_906_n 6.19475e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_506 N_A_693_369#_c_637_n N_A_877_369#_c_907_n 0.00175018f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_507 N_A_693_369#_c_628_n N_A_877_369#_c_908_n 0.0111876f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_508 N_A_693_369#_c_611_n N_A_877_369#_M1028_g 0.0150319f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_509 N_A_693_369#_c_629_n N_A_877_369#_M1045_g 0.00866971f $X=8.635 $Y=1.47
+ $X2=0 $Y2=0
cc_510 N_A_693_369#_c_630_n N_A_877_369#_M1045_g 0.00534181f $X=8.635 $Y=1.57
+ $X2=0 $Y2=0
cc_511 N_A_693_369#_M1005_g N_A_877_369#_M1045_g 0.0136211f $X=9.9 $Y=0.445
+ $X2=0 $Y2=0
cc_512 N_A_693_369#_c_619_n N_A_877_369#_M1045_g 0.00893179f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_513 N_A_693_369#_c_620_n N_A_877_369#_M1045_g 0.0206354f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_514 N_A_693_369#_c_621_n N_A_877_369#_M1045_g 0.0163585f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_515 N_A_693_369#_c_623_n N_A_877_369#_M1045_g 0.00133136f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_516 N_A_693_369#_c_625_n N_A_877_369#_M1045_g 0.00848925f $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_517 N_A_693_369#_c_630_n N_A_877_369#_c_910_n 0.0179968f $X=8.635 $Y=1.57
+ $X2=0 $Y2=0
cc_518 N_A_693_369#_c_621_n N_A_877_369#_c_910_n 0.00151205f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_519 N_A_693_369#_c_698_p N_A_877_369#_c_910_n 0.0033335f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_520 N_A_693_369#_c_609_n N_A_877_369#_c_897_n 0.00346646f $X=4.35 $Y=0.73
+ $X2=0 $Y2=0
cc_521 N_A_693_369#_c_610_n N_A_877_369#_c_897_n 0.015478f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_522 N_A_693_369#_c_615_n N_A_877_369#_c_897_n 0.0125458f $X=4.035 $Y=0.8
+ $X2=0 $Y2=0
cc_523 N_A_693_369#_c_617_n N_A_877_369#_c_897_n 0.0662039f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_524 N_A_693_369#_c_624_n N_A_877_369#_c_897_n 0.00343131f $X=4.235 $Y=1.09
+ $X2=0 $Y2=0
cc_525 N_A_693_369#_c_637_n N_A_877_369#_c_911_n 9.60456e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_526 N_A_693_369#_c_626_n N_A_877_369#_c_912_n 0.00343131f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_527 N_A_693_369#_c_627_n N_A_877_369#_c_912_n 0.00697298f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_528 N_A_693_369#_c_707_p N_A_877_369#_c_912_n 0.0109474f $X=4.165 $Y=1.83
+ $X2=0 $Y2=0
cc_529 N_A_693_369#_c_637_n N_A_877_369#_c_912_n 0.0215922f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_530 N_A_693_369#_c_638_n N_A_877_369#_c_912_n 0.00302262f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_531 N_A_693_369#_c_610_n N_A_877_369#_c_898_n 0.00209217f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_532 N_A_693_369#_c_619_n N_A_877_369#_c_898_n 0.0271596f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_533 N_A_693_369#_c_620_n N_A_877_369#_c_898_n 0.00288436f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_534 N_A_693_369#_c_621_n N_A_877_369#_c_898_n 0.0116627f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_535 N_A_693_369#_c_637_n N_A_877_369#_c_898_n 0.014567f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_536 N_A_693_369#_c_639_n N_A_877_369#_c_898_n 0.0618145f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_537 N_A_693_369#_c_640_n N_A_877_369#_c_898_n 0.0147711f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_538 N_A_693_369#_c_641_n N_A_877_369#_c_898_n 8.34727e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_539 N_A_693_369#_c_619_n N_A_877_369#_c_899_n 0.00222087f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_540 N_A_693_369#_c_621_n N_A_877_369#_c_899_n 0.0027091f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_541 N_A_693_369#_c_621_n N_A_877_369#_c_900_n 0.00293174f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_542 N_A_693_369#_c_623_n N_A_877_369#_c_900_n 0.00623523f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_543 N_A_693_369#_c_625_n N_A_877_369#_c_900_n 0.00392274f $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_544 N_A_693_369#_c_629_n N_A_877_369#_c_901_n 2.80207e-19 $X=8.635 $Y=1.47
+ $X2=0 $Y2=0
cc_545 N_A_693_369#_c_630_n N_A_877_369#_c_901_n 3.40634e-19 $X=8.635 $Y=1.57
+ $X2=0 $Y2=0
cc_546 N_A_693_369#_c_619_n N_A_877_369#_c_901_n 0.0260301f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_547 N_A_693_369#_c_620_n N_A_877_369#_c_901_n 4.25229e-19 $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_548 N_A_693_369#_c_621_n N_A_877_369#_c_901_n 0.0217551f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_549 N_A_693_369#_c_623_n N_A_877_369#_c_901_n 0.0118329f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_550 N_A_693_369#_c_698_p N_A_877_369#_c_901_n 0.0128627f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_551 N_A_693_369#_c_625_n N_A_877_369#_c_901_n 0.00143878f $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_552 N_A_693_369#_c_610_n N_A_877_369#_c_902_n 0.00266973f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_553 N_A_693_369#_c_618_n N_A_877_369#_c_902_n 0.00343131f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_554 N_A_693_369#_c_610_n N_A_877_369#_c_903_n 0.00247177f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_555 N_A_693_369#_c_617_n N_A_877_369#_c_903_n 0.00125608f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_556 N_A_693_369#_c_610_n N_A_877_369#_c_904_n 0.0528355f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_557 N_A_693_369#_c_617_n N_A_877_369#_c_904_n 2.72753e-19 $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_558 N_A_693_369#_c_618_n N_A_877_369#_c_904_n 0.0186987f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_559 N_A_693_369#_c_628_n N_A_1229_21#_c_1084_n 0.0334006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_560 N_A_693_369#_c_639_n N_A_1229_21#_c_1084_n 0.00848583f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_561 N_A_693_369#_c_639_n N_A_1229_21#_c_1085_n 0.0111901f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_562 N_A_693_369#_c_698_p N_A_1229_21#_c_1086_n 7.41551e-19 $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_563 N_A_693_369#_c_639_n N_A_1229_21#_c_1086_n 0.0287031f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_564 N_A_693_369#_c_639_n N_A_1229_21#_c_1087_n 0.0032337f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_565 N_A_693_369#_c_639_n N_A_1075_413#_c_1183_n 0.00384369f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_566 N_A_693_369#_c_639_n N_A_1075_413#_c_1184_n 7.54942e-19 $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_567 N_A_693_369#_c_629_n N_A_1075_413#_c_1185_n 0.0124551f $X=8.635 $Y=1.47
+ $X2=0 $Y2=0
cc_568 N_A_693_369#_c_619_n N_A_1075_413#_c_1185_n 0.001892f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_569 N_A_693_369#_c_630_n N_A_1075_413#_c_1186_n 0.0734562f $X=8.635 $Y=1.57
+ $X2=0 $Y2=0
cc_570 N_A_693_369#_c_619_n N_A_1075_413#_c_1186_n 7.14688e-19 $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_571 N_A_693_369#_c_698_p N_A_1075_413#_c_1186_n 0.0160277f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_572 N_A_693_369#_c_751_p N_A_1075_413#_c_1186_n 0.00203296f $X=8.295 $Y=1.87
+ $X2=0 $Y2=0
cc_573 N_A_693_369#_c_628_n N_A_1075_413#_c_1202_n 0.0154392f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_574 N_A_693_369#_c_637_n N_A_1075_413#_c_1202_n 0.00362812f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_575 N_A_693_369#_c_639_n N_A_1075_413#_c_1202_n 0.00492445f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_576 N_A_693_369#_c_640_n N_A_1075_413#_c_1202_n 0.00557824f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_577 N_A_693_369#_c_641_n N_A_1075_413#_c_1202_n 0.013294f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_578 N_A_693_369#_c_611_n N_A_1075_413#_c_1175_n 0.0028029f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_579 N_A_693_369#_c_628_n N_A_1075_413#_c_1187_n 0.00612006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_580 N_A_693_369#_c_639_n N_A_1075_413#_c_1187_n 0.0144347f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_581 N_A_693_369#_c_640_n N_A_1075_413#_c_1187_n 0.00314702f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_582 N_A_693_369#_c_641_n N_A_1075_413#_c_1187_n 0.0267088f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_583 N_A_693_369#_c_628_n N_A_1075_413#_c_1176_n 0.00266776f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_584 N_A_693_369#_c_637_n N_A_1075_413#_c_1176_n 0.00188086f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_585 N_A_693_369#_c_639_n N_A_1075_413#_c_1176_n 0.00794771f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_586 N_A_693_369#_c_640_n N_A_1075_413#_c_1176_n 0.00277252f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_587 N_A_693_369#_c_641_n N_A_1075_413#_c_1176_n 0.0162857f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_588 N_A_693_369#_c_619_n N_A_1075_413#_c_1177_n 0.0272879f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_589 N_A_693_369#_c_620_n N_A_1075_413#_c_1177_n 0.00195449f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_590 N_A_693_369#_c_698_p N_A_1075_413#_c_1177_n 0.0110153f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_591 N_A_693_369#_c_639_n N_A_1075_413#_c_1177_n 0.00254971f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_592 N_A_693_369#_c_639_n N_A_1075_413#_c_1178_n 0.00447966f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_593 N_A_693_369#_c_619_n N_A_1075_413#_c_1180_n 3.88379e-19 $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_594 N_A_693_369#_c_620_n N_A_1075_413#_c_1180_n 0.0124551f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_595 N_A_693_369#_c_698_p N_A_1075_413#_c_1180_n 0.00164261f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_596 N_A_693_369#_c_619_n N_A_1075_413#_c_1182_n 0.0022825f $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_597 N_A_693_369#_c_622_n N_A_1075_413#_c_1182_n 0.00403072f $X=8.885 $Y=0.812
+ $X2=0 $Y2=0
cc_598 N_A_693_369#_c_698_p N_SET_B_c_1330_n 0.00430764f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_599 N_A_693_369#_c_639_n N_SET_B_c_1330_n 0.00978683f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_600 N_A_693_369#_c_629_n N_SET_B_c_1335_n 5.55856e-19 $X=8.635 $Y=1.47 $X2=0
+ $Y2=0
cc_601 N_A_693_369#_c_630_n N_SET_B_c_1335_n 0.00106196f $X=8.635 $Y=1.57 $X2=0
+ $Y2=0
cc_602 N_A_693_369#_c_619_n N_SET_B_c_1335_n 0.024113f $X=8.67 $Y=1.16 $X2=0
+ $Y2=0
cc_603 N_A_693_369#_c_621_n N_SET_B_c_1335_n 0.00356101f $X=9.67 $Y=0.812 $X2=0
+ $Y2=0
cc_604 N_A_693_369#_c_623_n N_SET_B_c_1335_n 0.00179525f $X=9.79 $Y=1.09 $X2=0
+ $Y2=0
cc_605 N_A_693_369#_c_698_p N_SET_B_c_1335_n 0.0126888f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_606 N_A_693_369#_c_639_n N_SET_B_c_1335_n 0.0348253f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_607 N_A_693_369#_c_751_p N_SET_B_c_1335_n 0.0306606f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_608 N_A_693_369#_c_625_n N_SET_B_c_1335_n 3.78285e-19 $X=9.9 $Y=1.09 $X2=0
+ $Y2=0
cc_609 N_A_693_369#_c_639_n N_SET_B_c_1336_n 0.0304949f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_610 N_A_693_369#_c_623_n N_SET_B_c_1337_n 0.00770187f $X=9.79 $Y=1.09 $X2=0
+ $Y2=0
cc_611 N_A_693_369#_c_623_n N_SET_B_c_1338_n 0.0190534f $X=9.79 $Y=1.09 $X2=0
+ $Y2=0
cc_612 N_A_693_369#_c_625_n N_SET_B_c_1338_n 7.34482e-19 $X=9.9 $Y=1.09 $X2=0
+ $Y2=0
cc_613 N_A_693_369#_c_698_p N_SET_B_c_1339_n 0.00839482f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_614 N_A_693_369#_c_639_n N_SET_B_c_1339_n 0.011524f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_615 N_A_693_369#_c_623_n N_A_1951_295#_c_1466_n 2.4588e-19 $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_616 N_A_693_369#_c_625_n N_A_1951_295#_c_1466_n 0.0135231f $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_617 N_A_693_369#_M1005_g N_A_1951_295#_M1002_g 0.0366317f $X=9.9 $Y=0.445
+ $X2=0 $Y2=0
cc_618 N_A_693_369#_c_621_n N_A_1951_295#_M1002_g 0.00390523f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_619 N_A_693_369#_M1005_g N_A_1951_295#_c_1457_n 3.84849e-19 $X=9.9 $Y=0.445
+ $X2=0 $Y2=0
cc_620 N_A_693_369#_c_621_n N_A_1951_295#_c_1457_n 0.00348042f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_621 N_A_693_369#_c_623_n N_A_1951_295#_c_1457_n 0.018859f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_622 N_A_693_369#_c_623_n N_A_1951_295#_c_1458_n 0.00211266f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_623 N_A_693_369#_c_625_n N_A_1951_295#_c_1458_n 0.0366317f $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_624 N_A_693_369#_c_623_n N_A_1951_295#_c_1469_n 0.00422211f $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_625 N_A_693_369#_c_621_n N_A_1745_329#_M1045_d 0.0040046f $X=9.67 $Y=0.812
+ $X2=-0.19 $Y2=-0.24
cc_626 N_A_693_369#_c_619_n N_A_1745_329#_M1034_d 2.54843e-19 $X=8.67 $Y=1.16
+ $X2=0 $Y2=0
cc_627 N_A_693_369#_c_698_p N_A_1745_329#_M1034_d 0.00573907f $X=8.585 $Y=1.812
+ $X2=0 $Y2=0
cc_628 N_A_693_369#_c_630_n N_A_1745_329#_c_1578_n 0.00142794f $X=8.635 $Y=1.57
+ $X2=0 $Y2=0
cc_629 N_A_693_369#_M1005_g N_A_1745_329#_c_1579_n 0.0147933f $X=9.9 $Y=0.445
+ $X2=0 $Y2=0
cc_630 N_A_693_369#_c_621_n N_A_1745_329#_c_1579_n 0.0497339f $X=9.67 $Y=0.812
+ $X2=0 $Y2=0
cc_631 N_A_693_369#_c_625_n N_A_1745_329#_c_1579_n 6.4505e-19 $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_632 N_A_693_369#_c_623_n N_A_1745_329#_c_1573_n 7.54131e-19 $X=9.79 $Y=1.09
+ $X2=0 $Y2=0
cc_633 N_A_693_369#_c_625_n N_A_1745_329#_c_1573_n 3.84956e-19 $X=9.9 $Y=1.09
+ $X2=0 $Y2=0
cc_634 N_A_693_369#_c_631_n N_VPWR_M1044_d 7.92879e-19 $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_635 N_A_693_369#_c_707_p N_VPWR_M1044_d 0.00150754f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_636 N_A_693_369#_c_698_p N_VPWR_M1000_d 0.00927312f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_637 N_A_693_369#_c_642_n N_VPWR_c_1844_n 0.0102695f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_638 N_A_693_369#_c_642_n N_VPWR_c_1845_n 0.00603303f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_639 N_A_693_369#_c_631_n N_VPWR_c_1845_n 0.00195426f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_640 N_A_693_369#_c_751_p N_VPWR_c_1846_n 0.0039258f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_641 N_A_693_369#_c_698_p N_VPWR_c_1847_n 0.0381288f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_642 N_A_693_369#_c_639_n N_VPWR_c_1847_n 0.00793679f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_643 N_A_693_369#_c_627_n N_VPWR_c_1860_n 0.0055518f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_644 N_A_693_369#_c_628_n N_VPWR_c_1860_n 0.00429453f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_645 N_A_693_369#_c_707_p N_VPWR_c_1860_n 0.00103674f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_646 N_A_693_369#_c_627_n N_VPWR_c_1866_n 0.00815097f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_647 N_A_693_369#_c_642_n N_VPWR_c_1866_n 0.00373276f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_648 N_A_693_369#_c_631_n N_VPWR_c_1866_n 0.00632657f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_649 N_A_693_369#_c_707_p N_VPWR_c_1866_n 0.00632896f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_650 N_A_693_369#_c_638_n N_VPWR_c_1866_n 8.52709e-19 $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_651 N_A_693_369#_c_639_n N_VPWR_c_1867_n 0.00139085f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_652 N_A_693_369#_c_630_n N_VPWR_c_1868_n 0.0234092f $X=8.635 $Y=1.57 $X2=0
+ $Y2=0
cc_653 N_A_693_369#_c_698_p N_VPWR_c_1868_n 0.0110015f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_654 N_A_693_369#_M1044_s N_VPWR_c_1842_n 0.00400999f $X=3.465 $Y=1.845 $X2=0
+ $Y2=0
cc_655 N_A_693_369#_c_627_n N_VPWR_c_1842_n 0.00657032f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_656 N_A_693_369#_c_628_n N_VPWR_c_1842_n 0.00620168f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_657 N_A_693_369#_c_642_n N_VPWR_c_1842_n 0.00591039f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_658 N_A_693_369#_c_631_n N_VPWR_c_1842_n 0.004831f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_659 N_A_693_369#_c_707_p N_VPWR_c_1842_n 0.00153627f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_660 N_A_693_369#_c_698_p N_VPWR_c_1842_n 0.00693631f $X=8.585 $Y=1.812 $X2=0
+ $Y2=0
cc_661 N_A_693_369#_c_637_n N_VPWR_c_1842_n 0.0552922f $X=5.545 $Y=1.87 $X2=0
+ $Y2=0
cc_662 N_A_693_369#_c_638_n N_VPWR_c_1842_n 0.0167052f $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_663 N_A_693_369#_c_639_n N_VPWR_c_1842_n 0.103259f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_664 N_A_693_369#_c_640_n N_VPWR_c_1842_n 0.018311f $X=5.885 $Y=1.87 $X2=0
+ $Y2=0
cc_665 N_A_693_369#_c_751_p N_VPWR_c_1842_n 0.0168258f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_666 N_A_693_369#_c_611_n N_A_201_47#_c_2057_n 0.00439649f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_667 N_A_693_369#_c_628_n N_A_201_47#_c_2062_n 3.6876e-19 $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_668 N_A_693_369#_c_637_n N_A_201_47#_c_2062_n 0.0162746f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_669 N_A_693_369#_c_640_n N_A_201_47#_c_2062_n 0.00274259f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_670 N_A_693_369#_c_610_n N_A_201_47#_c_2058_n 0.0110036f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_671 N_A_693_369#_c_626_n N_A_201_47#_c_2063_n 0.00641873f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_672 N_A_693_369#_c_613_n N_A_201_47#_c_2063_n 0.00176142f $X=4.317 $Y=0.805
+ $X2=0 $Y2=0
cc_673 N_A_693_369#_c_631_n N_A_201_47#_c_2063_n 0.0099266f $X=4.035 $Y=1.915
+ $X2=0 $Y2=0
cc_674 N_A_693_369#_c_632_n N_A_201_47#_c_2063_n 0.00126159f $X=3.675 $Y=1.915
+ $X2=0 $Y2=0
cc_675 N_A_693_369#_c_615_n N_A_201_47#_c_2063_n 0.00714535f $X=4.035 $Y=0.8
+ $X2=0 $Y2=0
cc_676 N_A_693_369#_c_616_n N_A_201_47#_c_2063_n 7.07979e-19 $X=3.705 $Y=0.8
+ $X2=0 $Y2=0
cc_677 N_A_693_369#_c_617_n N_A_201_47#_c_2063_n 0.0221679f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_678 N_A_693_369#_c_637_n N_A_201_47#_c_2063_n 0.0423006f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_679 N_A_693_369#_c_638_n N_A_201_47#_c_2063_n 0.030156f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_680 N_A_693_369#_c_628_n N_A_201_47#_c_2066_n 0.00118188f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_681 N_A_693_369#_c_637_n N_A_201_47#_c_2066_n 0.0257219f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_682 N_A_693_369#_c_641_n N_A_201_47#_c_2066_n 0.00187515f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_683 N_A_693_369#_c_610_n N_A_201_47#_c_2060_n 0.0062731f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_684 N_A_693_369#_c_628_n N_A_201_47#_c_2060_n 0.00244962f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_685 N_A_693_369#_c_641_n N_A_201_47#_c_2060_n 0.0103278f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_686 N_A_693_369#_c_698_p A_1663_329# 0.00203785f $X=8.585 $Y=1.812 $X2=-0.19
+ $Y2=-0.24
cc_687 N_A_693_369#_c_751_p A_1663_329# 0.00166585f $X=8.295 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_688 N_A_693_369#_c_614_n N_VGND_c_2246_n 0.0239409f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_689 N_A_693_369#_c_609_n N_VGND_c_2247_n 0.00312892f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_690 N_A_693_369#_c_613_n N_VGND_c_2247_n 2.23286e-19 $X=4.317 $Y=0.805 $X2=0
+ $Y2=0
cc_691 N_A_693_369#_c_614_n N_VGND_c_2247_n 0.0176685f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_692 N_A_693_369#_c_615_n N_VGND_c_2247_n 0.0235008f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_693 N_A_693_369#_c_618_n N_VGND_c_2247_n 4.8449e-19 $X=4.21 $Y=1.255 $X2=0
+ $Y2=0
cc_694 N_A_693_369#_c_614_n N_VGND_c_2253_n 0.0127969f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_695 N_A_693_369#_c_615_n N_VGND_c_2253_n 0.00317989f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_696 N_A_693_369#_c_609_n N_VGND_c_2257_n 0.00565513f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_697 N_A_693_369#_c_610_n N_VGND_c_2257_n 0.00394222f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_698 N_A_693_369#_c_611_n N_VGND_c_2257_n 0.00585385f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_699 N_A_693_369#_c_615_n N_VGND_c_2257_n 6.403e-19 $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_700 N_A_693_369#_M1005_g N_VGND_c_2258_n 0.00362032f $X=9.9 $Y=0.445 $X2=0
+ $Y2=0
cc_701 N_A_693_369#_c_621_n N_VGND_c_2258_n 0.00468447f $X=9.67 $Y=0.812 $X2=0
+ $Y2=0
cc_702 N_A_693_369#_c_622_n N_VGND_c_2258_n 0.00486578f $X=8.885 $Y=0.812 $X2=0
+ $Y2=0
cc_703 N_A_693_369#_c_622_n N_VGND_c_2264_n 0.00757355f $X=8.885 $Y=0.812 $X2=0
+ $Y2=0
cc_704 N_A_693_369#_M1021_s N_VGND_c_2267_n 0.00388795f $X=3.495 $Y=0.235 $X2=0
+ $Y2=0
cc_705 N_A_693_369#_c_609_n N_VGND_c_2267_n 0.0113329f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_706 N_A_693_369#_c_610_n N_VGND_c_2267_n 0.00371212f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_707 N_A_693_369#_c_611_n N_VGND_c_2267_n 0.0121314f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_708 N_A_693_369#_M1005_g N_VGND_c_2267_n 0.00581448f $X=9.9 $Y=0.445 $X2=0
+ $Y2=0
cc_709 N_A_693_369#_c_614_n N_VGND_c_2267_n 0.00703355f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_710 N_A_693_369#_c_615_n N_VGND_c_2267_n 0.00765233f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_711 N_A_693_369#_c_621_n N_VGND_c_2267_n 0.010075f $X=9.67 $Y=0.812 $X2=0
+ $Y2=0
cc_712 N_A_693_369#_c_622_n N_VGND_c_2267_n 0.00847772f $X=8.885 $Y=0.812 $X2=0
+ $Y2=0
cc_713 N_A_693_369#_c_621_n A_1654_47# 0.00233778f $X=9.67 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_714 N_A_693_369#_c_622_n A_1654_47# 0.00945823f $X=8.885 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_715 N_A_877_369#_M1028_g N_A_1229_21#_M1019_g 0.0469974f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_716 N_A_877_369#_M1028_g N_A_1229_21#_c_1078_n 0.00658605f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_717 N_A_877_369#_c_898_n N_A_1229_21#_c_1078_n 0.0031108f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_718 N_A_877_369#_c_898_n N_A_1229_21#_c_1085_n 5.84337e-19 $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_719 N_A_877_369#_c_898_n N_A_1229_21#_c_1079_n 0.00911256f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_720 N_A_877_369#_M1028_g N_A_1229_21#_c_1081_n 0.00133724f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_721 N_A_877_369#_c_898_n N_A_1229_21#_c_1081_n 0.00983807f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_722 N_A_877_369#_c_898_n N_A_1229_21#_c_1082_n 0.00306049f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_723 N_A_877_369#_c_894_n N_A_1075_413#_c_1175_n 0.0141556f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_724 N_A_877_369#_M1028_g N_A_1075_413#_c_1175_n 0.0220882f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_725 N_A_877_369#_c_898_n N_A_1075_413#_c_1175_n 0.0327905f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_726 N_A_877_369#_c_898_n N_A_1075_413#_c_1187_n 3.47492e-19 $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_727 N_A_877_369#_c_894_n N_A_1075_413#_c_1176_n 0.00570521f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_728 N_A_877_369#_c_898_n N_A_1075_413#_c_1176_n 0.0218948f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_729 N_A_877_369#_c_904_n N_A_1075_413#_c_1176_n 3.61543e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_730 N_A_877_369#_c_898_n N_A_1075_413#_c_1177_n 0.0594233f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_731 N_A_877_369#_c_898_n N_A_1075_413#_c_1178_n 0.0189259f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_732 N_A_877_369#_c_898_n N_A_1075_413#_c_1179_n 0.0111401f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_733 N_A_877_369#_c_898_n N_A_1075_413#_c_1181_n 0.00146646f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_734 N_A_877_369#_M1045_g N_SET_B_c_1335_n 0.00172911f $X=9.14 $Y=0.555 $X2=0
+ $Y2=0
cc_735 N_A_877_369#_c_910_n N_SET_B_c_1335_n 0.00265142f $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_736 N_A_877_369#_c_898_n N_SET_B_c_1335_n 0.114413f $X=9.17 $Y=1.19 $X2=0
+ $Y2=0
cc_737 N_A_877_369#_c_899_n N_SET_B_c_1335_n 0.034199f $X=9.285 $Y=1.19 $X2=0
+ $Y2=0
cc_738 N_A_877_369#_c_901_n N_SET_B_c_1335_n 0.0188957f $X=9.365 $Y=1.19 $X2=0
+ $Y2=0
cc_739 N_A_877_369#_c_898_n N_SET_B_c_1336_n 0.0307796f $X=9.17 $Y=1.19 $X2=0
+ $Y2=0
cc_740 N_A_877_369#_c_910_n N_SET_B_c_1337_n 7.17593e-19 $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_741 N_A_877_369#_c_901_n N_SET_B_c_1337_n 0.00277925f $X=9.365 $Y=1.19 $X2=0
+ $Y2=0
cc_742 N_A_877_369#_M1045_g N_SET_B_c_1338_n 3.27076e-19 $X=9.14 $Y=0.555 $X2=0
+ $Y2=0
cc_743 N_A_877_369#_c_910_n N_SET_B_c_1338_n 8.85426e-19 $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_744 N_A_877_369#_c_901_n N_SET_B_c_1338_n 0.0163922f $X=9.365 $Y=1.19 $X2=0
+ $Y2=0
cc_745 N_A_877_369#_c_898_n N_SET_B_c_1339_n 0.00146727f $X=9.17 $Y=1.19 $X2=0
+ $Y2=0
cc_746 N_A_877_369#_c_901_n N_A_1951_295#_c_1463_n 0.00103803f $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_747 N_A_877_369#_c_910_n N_A_1951_295#_c_1464_n 0.0284644f $X=9.365 $Y=1.99
+ $X2=0 $Y2=0
cc_748 N_A_877_369#_M1045_g N_A_1951_295#_c_1466_n 0.00167318f $X=9.14 $Y=0.555
+ $X2=0 $Y2=0
cc_749 N_A_877_369#_c_910_n N_A_1951_295#_c_1466_n 0.0216246f $X=9.365 $Y=1.99
+ $X2=0 $Y2=0
cc_750 N_A_877_369#_c_901_n N_A_1951_295#_c_1466_n 5.0381e-19 $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_751 N_A_877_369#_c_900_n N_A_1951_295#_c_1456_n 0.00101096f $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_752 N_A_877_369#_c_901_n N_A_1951_295#_c_1456_n 0.00358367f $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_753 N_A_877_369#_c_910_n N_A_1745_329#_c_1578_n 0.0244065f $X=9.365 $Y=1.99
+ $X2=0 $Y2=0
cc_754 N_A_877_369#_c_901_n N_A_1745_329#_c_1578_n 0.016028f $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_755 N_A_877_369#_c_910_n N_A_1745_329#_c_1573_n 0.00479045f $X=9.365 $Y=1.99
+ $X2=0 $Y2=0
cc_756 N_A_877_369#_c_901_n N_A_1745_329#_c_1573_n 7.50645e-19 $X=9.365 $Y=1.19
+ $X2=0 $Y2=0
cc_757 N_A_877_369#_c_906_n N_VPWR_c_1860_n 4.12218e-19 $X=5.195 $Y=1.915 $X2=0
+ $Y2=0
cc_758 N_A_877_369#_c_907_n N_VPWR_c_1860_n 0.00206689f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_759 N_A_877_369#_c_908_n N_VPWR_c_1860_n 0.00702461f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_760 N_A_877_369#_c_911_n N_VPWR_c_1860_n 0.0242014f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_761 N_A_877_369#_c_910_n N_VPWR_c_1861_n 0.00430708f $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_762 N_A_877_369#_c_911_n N_VPWR_c_1866_n 0.0122663f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_763 N_A_877_369#_c_910_n N_VPWR_c_1868_n 0.0015408f $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_764 N_A_877_369#_M1031_d N_VPWR_c_1842_n 0.00224652f $X=4.385 $Y=1.845 $X2=0
+ $Y2=0
cc_765 N_A_877_369#_c_907_n N_VPWR_c_1842_n 0.00154765f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_766 N_A_877_369#_c_908_n N_VPWR_c_1842_n 0.00872443f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_767 N_A_877_369#_c_910_n N_VPWR_c_1842_n 0.00672267f $X=9.365 $Y=1.99 $X2=0
+ $Y2=0
cc_768 N_A_877_369#_c_911_n N_VPWR_c_1842_n 0.00627246f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_769 N_A_877_369#_c_897_n N_A_201_47#_c_2057_n 0.041221f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_770 N_A_877_369#_c_905_n N_A_201_47#_c_2061_n 0.00358193f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_771 N_A_877_369#_c_912_n N_A_201_47#_c_2061_n 0.0324615f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_772 N_A_877_369#_c_898_n N_A_201_47#_c_2061_n 6.11234e-19 $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_773 N_A_877_369#_c_905_n N_A_201_47#_c_2062_n 0.00244422f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_774 N_A_877_369#_c_906_n N_A_201_47#_c_2062_n 0.00940185f $X=5.195 $Y=1.915
+ $X2=0 $Y2=0
cc_775 N_A_877_369#_c_907_n N_A_201_47#_c_2062_n 0.00335679f $X=5.04 $Y=1.915
+ $X2=0 $Y2=0
cc_776 N_A_877_369#_c_908_n N_A_201_47#_c_2062_n 0.00398401f $X=5.285 $Y=1.99
+ $X2=0 $Y2=0
cc_777 N_A_877_369#_c_911_n N_A_201_47#_c_2062_n 0.0324615f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_778 N_A_877_369#_c_898_n N_A_201_47#_c_2058_n 0.00517494f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_779 N_A_877_369#_c_903_n N_A_201_47#_c_2058_n 3.91268e-19 $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_780 N_A_877_369#_c_904_n N_A_201_47#_c_2058_n 9.17329e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_781 N_A_877_369#_c_905_n N_A_201_47#_c_2063_n 0.00251435f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_782 N_A_877_369#_c_912_n N_A_201_47#_c_2063_n 0.0189338f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_783 N_A_877_369#_c_898_n N_A_201_47#_c_2063_n 0.00685911f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_784 N_A_877_369#_c_902_n N_A_201_47#_c_2063_n 0.0014563f $X=4.72 $Y=1.185
+ $X2=0 $Y2=0
cc_785 N_A_877_369#_c_903_n N_A_201_47#_c_2063_n 0.0250391f $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_786 N_A_877_369#_c_904_n N_A_201_47#_c_2063_n 8.40015e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_787 N_A_877_369#_c_905_n N_A_201_47#_c_2066_n 8.26579e-19 $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_788 N_A_877_369#_c_912_n N_A_201_47#_c_2066_n 0.00217539f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_789 N_A_877_369#_c_898_n N_A_201_47#_c_2066_n 0.0260799f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_790 N_A_877_369#_c_904_n N_A_201_47#_c_2066_n 5.52268e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_791 N_A_877_369#_c_905_n N_A_201_47#_c_2060_n 0.00416664f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_792 N_A_877_369#_c_894_n N_A_201_47#_c_2060_n 0.00791292f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_793 N_A_877_369#_M1028_g N_A_201_47#_c_2060_n 8.1098e-19 $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_794 N_A_877_369#_c_897_n N_A_201_47#_c_2060_n 0.0138333f $X=4.56 $Y=0.42
+ $X2=0 $Y2=0
cc_795 N_A_877_369#_c_912_n N_A_201_47#_c_2060_n 0.00871828f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_796 N_A_877_369#_c_898_n N_A_201_47#_c_2060_n 0.0126669f $X=9.17 $Y=1.19
+ $X2=0 $Y2=0
cc_797 N_A_877_369#_c_902_n N_A_201_47#_c_2060_n 0.0222258f $X=4.72 $Y=1.185
+ $X2=0 $Y2=0
cc_798 N_A_877_369#_c_903_n N_A_201_47#_c_2060_n 0.0023779f $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_799 N_A_877_369#_c_904_n N_A_201_47#_c_2060_n 0.00621958f $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_800 N_A_877_369#_M1028_g N_VGND_c_2257_n 0.00717785f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_801 N_A_877_369#_c_897_n N_VGND_c_2257_n 0.0144177f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_802 N_A_877_369#_M1045_g N_VGND_c_2258_n 0.00437171f $X=9.14 $Y=0.555 $X2=0
+ $Y2=0
cc_803 N_A_877_369#_M1045_g N_VGND_c_2264_n 0.0140162f $X=9.14 $Y=0.555 $X2=0
+ $Y2=0
cc_804 N_A_877_369#_c_898_n N_VGND_c_2264_n 0.00696859f $X=9.17 $Y=1.19 $X2=0
+ $Y2=0
cc_805 N_A_877_369#_M1018_d N_VGND_c_2267_n 0.00382094f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_806 N_A_877_369#_M1028_g N_VGND_c_2267_n 0.00537275f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_807 N_A_877_369#_M1045_g N_VGND_c_2267_n 0.00814253f $X=9.14 $Y=0.555 $X2=0
+ $Y2=0
cc_808 N_A_877_369#_c_897_n N_VGND_c_2267_n 0.00801045f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_809 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1172_n 5.62208e-19 $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_810 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1183_n 0.00632289f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_811 N_A_1229_21#_c_1084_n N_A_1075_413#_c_1183_n 0.0171889f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_812 N_A_1229_21#_c_1085_n N_A_1075_413#_c_1183_n 0.00183365f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_813 N_A_1229_21#_c_1084_n N_A_1075_413#_c_1184_n 0.0150522f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_814 N_A_1229_21#_c_1085_n N_A_1075_413#_c_1184_n 4.03149e-19 $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_815 N_A_1229_21#_c_1086_n N_A_1075_413#_c_1184_n 0.0160003f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_816 N_A_1229_21#_c_1079_n N_A_1075_413#_c_1173_n 0.00198418f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_817 N_A_1229_21#_c_1080_n N_A_1075_413#_c_1173_n 0.0077537f $X=6.95 $Y=0.51
+ $X2=0 $Y2=0
cc_818 N_A_1229_21#_M1019_g N_A_1075_413#_c_1174_n 8.49245e-19 $X=6.22 $Y=0.445
+ $X2=0 $Y2=0
cc_819 N_A_1229_21#_c_1079_n N_A_1075_413#_c_1174_n 0.00807215f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_820 N_A_1229_21#_c_1081_n N_A_1075_413#_c_1174_n 0.00110084f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_821 N_A_1229_21#_c_1082_n N_A_1075_413#_c_1174_n 0.00784562f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_822 N_A_1229_21#_M1019_g N_A_1075_413#_c_1175_n 0.00122809f $X=6.22 $Y=0.445
+ $X2=0 $Y2=0
cc_823 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1175_n 0.00261079f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_824 N_A_1229_21#_c_1081_n N_A_1075_413#_c_1175_n 0.0269973f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_825 N_A_1229_21#_c_1082_n N_A_1075_413#_c_1175_n 0.00113583f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_826 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1187_n 0.011517f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_827 N_A_1229_21#_c_1084_n N_A_1075_413#_c_1187_n 0.00116159f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_828 N_A_1229_21#_c_1085_n N_A_1075_413#_c_1187_n 0.0201747f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_829 N_A_1229_21#_c_1087_n N_A_1075_413#_c_1187_n 0.00880623f $X=6.595 $Y=2.02
+ $X2=0 $Y2=0
cc_830 N_A_1229_21#_c_1081_n N_A_1075_413#_c_1176_n 0.0192437f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_831 N_A_1229_21#_c_1082_n N_A_1075_413#_c_1176_n 0.0018579f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_832 N_A_1229_21#_c_1086_n N_A_1075_413#_c_1177_n 0.00267752f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_833 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1178_n 0.0152311f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_834 N_A_1229_21#_c_1084_n N_A_1075_413#_c_1178_n 0.00260846f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_835 N_A_1229_21#_c_1085_n N_A_1075_413#_c_1178_n 0.0109804f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_836 N_A_1229_21#_c_1079_n N_A_1075_413#_c_1178_n 0.00808722f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_837 N_A_1229_21#_c_1086_n N_A_1075_413#_c_1178_n 0.00696445f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_838 N_A_1229_21#_c_1082_n N_A_1075_413#_c_1178_n 5.30627e-19 $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_839 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1179_n 0.0017292f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_840 N_A_1229_21#_c_1079_n N_A_1075_413#_c_1179_n 0.0178097f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_841 N_A_1229_21#_c_1081_n N_A_1075_413#_c_1179_n 0.0020275f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_842 N_A_1229_21#_c_1082_n N_A_1075_413#_c_1179_n 0.00156611f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_843 N_A_1229_21#_c_1078_n N_A_1075_413#_c_1181_n 0.0115036f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_844 N_A_1229_21#_c_1079_n N_A_1075_413#_c_1181_n 0.00227132f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_845 N_A_1229_21#_c_1086_n N_A_1075_413#_c_1181_n 6.97279e-19 $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_846 N_A_1229_21#_c_1086_n N_SET_B_c_1330_n 0.00621496f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_847 N_A_1229_21#_c_1140_p N_SET_B_c_1330_n 0.00390541f $X=7.265 $Y=2.285
+ $X2=0 $Y2=0
cc_848 N_A_1229_21#_c_1085_n N_SET_B_c_1339_n 0.005781f $X=6.51 $Y=1.74 $X2=0
+ $Y2=0
cc_849 N_A_1229_21#_c_1086_n N_SET_B_c_1339_n 0.0157577f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_850 N_A_1229_21#_c_1086_n N_VPWR_M1043_d 0.00298622f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_851 N_A_1229_21#_c_1087_n N_VPWR_M1043_d 0.00153636f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_852 N_A_1229_21#_c_1086_n N_VPWR_c_1855_n 0.00479971f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_853 N_A_1229_21#_c_1140_p N_VPWR_c_1855_n 0.0165337f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_854 N_A_1229_21#_c_1084_n N_VPWR_c_1860_n 0.00743866f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_855 N_A_1229_21#_c_1084_n N_VPWR_c_1867_n 0.0056962f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_856 N_A_1229_21#_c_1086_n N_VPWR_c_1867_n 0.0164669f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_857 N_A_1229_21#_c_1087_n N_VPWR_c_1867_n 0.0102436f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_858 N_A_1229_21#_c_1140_p N_VPWR_c_1867_n 0.00867119f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_859 N_A_1229_21#_M1011_d N_VPWR_c_1842_n 0.00331536f $X=7.095 $Y=2.065 $X2=0
+ $Y2=0
cc_860 N_A_1229_21#_c_1084_n N_VPWR_c_1842_n 0.00849347f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_861 N_A_1229_21#_c_1086_n N_VPWR_c_1842_n 0.0042909f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_862 N_A_1229_21#_c_1087_n N_VPWR_c_1842_n 7.82982e-19 $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_863 N_A_1229_21#_c_1140_p N_VPWR_c_1842_n 0.00471488f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_864 N_A_1229_21#_c_1079_n N_VGND_M1019_d 8.64202e-19 $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_865 N_A_1229_21#_c_1081_n N_VGND_M1019_d 0.00133208f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_866 N_A_1229_21#_M1019_g N_VGND_c_2257_n 0.014377f $X=6.22 $Y=0.445 $X2=0
+ $Y2=0
cc_867 N_A_1229_21#_c_1079_n N_VGND_c_2257_n 0.00919218f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_868 N_A_1229_21#_c_1080_n N_VGND_c_2257_n 0.0164501f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_869 N_A_1229_21#_c_1081_n N_VGND_c_2257_n 0.0212099f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_870 N_A_1229_21#_c_1082_n N_VGND_c_2257_n 8.18098e-19 $X=6.31 $Y=0.93 $X2=0
+ $Y2=0
cc_871 N_A_1229_21#_c_1079_n N_VGND_c_2263_n 0.00346394f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_872 N_A_1229_21#_c_1080_n N_VGND_c_2263_n 0.0172232f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_873 N_A_1229_21#_c_1079_n N_VGND_c_2264_n 0.0118068f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_874 N_A_1229_21#_c_1080_n N_VGND_c_2264_n 0.0251021f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_875 N_A_1229_21#_M1024_s N_VGND_c_2267_n 0.00468266f $X=6.825 $Y=0.235 $X2=0
+ $Y2=0
cc_876 N_A_1229_21#_c_1079_n N_VGND_c_2267_n 0.00594673f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_877 N_A_1229_21#_c_1080_n N_VGND_c_2267_n 0.00949852f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_878 N_A_1229_21#_c_1081_n N_VGND_c_2267_n 0.00174322f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_879 N_A_1075_413#_c_1183_n N_SET_B_c_1329_n 0.0047982f $X=7.005 $Y=1.89 $X2=0
+ $Y2=0
cc_880 N_A_1075_413#_c_1185_n N_SET_B_c_1329_n 0.00304149f $X=8.225 $Y=1.47
+ $X2=0 $Y2=0
cc_881 N_A_1075_413#_c_1183_n N_SET_B_c_1330_n 0.0204443f $X=7.005 $Y=1.89 $X2=0
+ $Y2=0
cc_882 N_A_1075_413#_c_1184_n N_SET_B_c_1330_n 0.0108477f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_883 N_A_1075_413#_c_1186_n N_SET_B_c_1330_n 0.0262224f $X=8.225 $Y=1.57 $X2=0
+ $Y2=0
cc_884 N_A_1075_413#_c_1177_n N_SET_B_c_1330_n 7.94155e-19 $X=8.005 $Y=1.125
+ $X2=0 $Y2=0
cc_885 N_A_1075_413#_c_1172_n N_SET_B_M1017_g 0.00773331f $X=7.005 $Y=1.095
+ $X2=0 $Y2=0
cc_886 N_A_1075_413#_c_1173_n N_SET_B_M1017_g 0.0390147f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_887 N_A_1075_413#_c_1177_n N_SET_B_M1017_g 0.0118397f $X=8.005 $Y=1.125 $X2=0
+ $Y2=0
cc_888 N_A_1075_413#_c_1180_n N_SET_B_M1017_g 0.0214689f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_889 N_A_1075_413#_c_1182_n N_SET_B_M1017_g 0.0236625f $X=8.14 $Y=0.995 $X2=0
+ $Y2=0
cc_890 N_A_1075_413#_c_1185_n N_SET_B_c_1328_n 0.00161756f $X=8.225 $Y=1.47
+ $X2=0 $Y2=0
cc_891 N_A_1075_413#_c_1177_n N_SET_B_c_1328_n 0.00828332f $X=8.005 $Y=1.125
+ $X2=0 $Y2=0
cc_892 N_A_1075_413#_c_1179_n N_SET_B_c_1328_n 5.69298e-19 $X=6.975 $Y=1.185
+ $X2=0 $Y2=0
cc_893 N_A_1075_413#_c_1181_n N_SET_B_c_1328_n 0.0047982f $X=7.005 $Y=1.23 $X2=0
+ $Y2=0
cc_894 N_A_1075_413#_c_1185_n N_SET_B_c_1335_n 0.00138481f $X=8.225 $Y=1.47
+ $X2=0 $Y2=0
cc_895 N_A_1075_413#_c_1186_n N_SET_B_c_1335_n 0.00403144f $X=8.225 $Y=1.57
+ $X2=0 $Y2=0
cc_896 N_A_1075_413#_c_1177_n N_SET_B_c_1335_n 0.00966361f $X=8.005 $Y=1.125
+ $X2=0 $Y2=0
cc_897 N_A_1075_413#_c_1180_n N_SET_B_c_1335_n 7.77586e-19 $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_898 N_A_1075_413#_c_1183_n N_SET_B_c_1336_n 4.70557e-19 $X=7.005 $Y=1.89
+ $X2=0 $Y2=0
cc_899 N_A_1075_413#_c_1185_n N_SET_B_c_1336_n 6.48307e-19 $X=8.225 $Y=1.47
+ $X2=0 $Y2=0
cc_900 N_A_1075_413#_c_1186_n N_SET_B_c_1336_n 6.42433e-19 $X=8.225 $Y=1.57
+ $X2=0 $Y2=0
cc_901 N_A_1075_413#_c_1177_n N_SET_B_c_1336_n 0.00200562f $X=8.005 $Y=1.125
+ $X2=0 $Y2=0
cc_902 N_A_1075_413#_c_1183_n N_SET_B_c_1339_n 0.00646306f $X=7.005 $Y=1.89
+ $X2=0 $Y2=0
cc_903 N_A_1075_413#_c_1185_n N_SET_B_c_1339_n 0.00157368f $X=8.225 $Y=1.47
+ $X2=0 $Y2=0
cc_904 N_A_1075_413#_c_1186_n N_SET_B_c_1339_n 0.00172871f $X=8.225 $Y=1.57
+ $X2=0 $Y2=0
cc_905 N_A_1075_413#_c_1177_n N_SET_B_c_1339_n 0.0354578f $X=8.005 $Y=1.125
+ $X2=0 $Y2=0
cc_906 N_A_1075_413#_c_1186_n N_VPWR_c_1846_n 0.0264172f $X=8.225 $Y=1.57 $X2=0
+ $Y2=0
cc_907 N_A_1075_413#_c_1184_n N_VPWR_c_1855_n 0.00512994f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_908 N_A_1075_413#_c_1202_n N_VPWR_c_1860_n 0.0464661f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_909 N_A_1075_413#_c_1184_n N_VPWR_c_1867_n 0.00620668f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_910 N_A_1075_413#_M1008_d N_VPWR_c_1842_n 0.00231251f $X=5.375 $Y=2.065 $X2=0
+ $Y2=0
cc_911 N_A_1075_413#_c_1184_n N_VPWR_c_1842_n 0.00720657f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_912 N_A_1075_413#_c_1202_n N_VPWR_c_1842_n 0.012998f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_913 N_A_1075_413#_c_1175_n N_A_201_47#_c_2057_n 0.040178f $X=5.55 $Y=0.42
+ $X2=0 $Y2=0
cc_914 N_A_1075_413#_c_1176_n N_A_201_47#_c_2060_n 0.00906057f $X=6.205 $Y=1.31
+ $X2=0 $Y2=0
cc_915 N_A_1075_413#_c_1202_n A_1169_413# 0.00692155f $X=6.035 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_916 N_A_1075_413#_c_1187_n A_1169_413# 0.00130666f $X=6.12 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_917 N_A_1075_413#_c_1173_n N_VGND_c_2257_n 0.00172114f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_918 N_A_1075_413#_c_1175_n N_VGND_c_2257_n 0.0270576f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_919 N_A_1075_413#_c_1173_n N_VGND_c_2263_n 0.00271402f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_920 N_A_1075_413#_c_1174_n N_VGND_c_2263_n 0.00305109f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_921 N_A_1075_413#_c_1173_n N_VGND_c_2264_n 0.0187167f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_922 N_A_1075_413#_c_1174_n N_VGND_c_2264_n 0.00316742f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_923 N_A_1075_413#_c_1177_n N_VGND_c_2264_n 0.0870936f $X=8.005 $Y=1.125 $X2=0
+ $Y2=0
cc_924 N_A_1075_413#_c_1180_n N_VGND_c_2264_n 0.00108367f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_925 N_A_1075_413#_c_1182_n N_VGND_c_2264_n 0.0370231f $X=8.14 $Y=0.995 $X2=0
+ $Y2=0
cc_926 N_A_1075_413#_M1033_d N_VGND_c_2267_n 0.00428929f $X=5.415 $Y=0.235 $X2=0
+ $Y2=0
cc_927 N_A_1075_413#_c_1173_n N_VGND_c_2267_n 0.00630011f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_928 N_A_1075_413#_c_1174_n N_VGND_c_2267_n 0.00363714f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_929 N_A_1075_413#_c_1175_n N_VGND_c_2267_n 0.0155321f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_930 N_SET_B_c_1331_n N_A_1951_295#_c_1463_n 0.00779841f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_931 N_SET_B_c_1334_n N_A_1951_295#_c_1463_n 3.11511e-19 $X=10.78 $Y=1.63
+ $X2=0 $Y2=0
cc_932 N_SET_B_c_1338_n N_A_1951_295#_c_1463_n 0.00596497f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_933 N_SET_B_c_1331_n N_A_1951_295#_c_1464_n 0.0110556f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_934 N_SET_B_c_1334_n N_A_1951_295#_c_1465_n 0.0177936f $X=10.78 $Y=1.63 $X2=0
+ $Y2=0
cc_935 N_SET_B_c_1337_n N_A_1951_295#_c_1465_n 0.00171811f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_936 N_SET_B_c_1338_n N_A_1951_295#_c_1465_n 0.0048762f $X=9.875 $Y=1.53 $X2=0
+ $Y2=0
cc_937 N_SET_B_c_1338_n N_A_1951_295#_c_1466_n 0.00438471f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_938 N_SET_B_M1015_g N_A_1951_295#_M1002_g 0.0163085f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_939 N_SET_B_c_1331_n N_A_1951_295#_c_1456_n 0.0111834f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_940 N_SET_B_M1015_g N_A_1951_295#_c_1456_n 0.0079467f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_941 N_SET_B_c_1337_n N_A_1951_295#_c_1456_n 0.00162315f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_942 N_SET_B_c_1338_n N_A_1951_295#_c_1456_n 0.00166329f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_943 N_SET_B_M1015_g N_A_1951_295#_c_1457_n 0.00134295f $X=10.89 $Y=0.445
+ $X2=0 $Y2=0
cc_944 N_SET_B_c_1331_n N_A_1951_295#_c_1458_n 4.41093e-19 $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_945 N_SET_B_M1015_g N_A_1951_295#_c_1458_n 0.0133157f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_946 N_SET_B_c_1334_n N_A_1951_295#_c_1458_n 4.53365e-19 $X=10.78 $Y=1.63
+ $X2=0 $Y2=0
cc_947 N_SET_B_c_1331_n N_A_1951_295#_c_1459_n 0.00602516f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_948 N_SET_B_M1015_g N_A_1951_295#_c_1459_n 0.0113692f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_949 N_SET_B_c_1334_n N_A_1951_295#_c_1459_n 0.0353867f $X=10.78 $Y=1.63 $X2=0
+ $Y2=0
cc_950 N_SET_B_c_1334_n N_A_1951_295#_c_1469_n 0.0192836f $X=10.78 $Y=1.63 $X2=0
+ $Y2=0
cc_951 N_SET_B_c_1331_n N_A_1745_329#_c_1557_n 0.0181287f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_952 N_SET_B_c_1334_n N_A_1745_329#_c_1557_n 0.00239457f $X=10.78 $Y=1.63
+ $X2=0 $Y2=0
cc_953 N_SET_B_M1015_g N_A_1745_329#_c_1560_n 0.0182994f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_954 N_SET_B_M1015_g N_A_1745_329#_c_1561_n 0.0118803f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_955 N_SET_B_c_1335_n N_A_1745_329#_c_1578_n 0.0151371f $X=9.73 $Y=1.53 $X2=0
+ $Y2=0
cc_956 N_SET_B_M1015_g N_A_1745_329#_c_1579_n 0.010177f $X=10.89 $Y=0.445 $X2=0
+ $Y2=0
cc_957 N_SET_B_c_1331_n N_A_1745_329#_c_1571_n 0.0362752f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_958 N_SET_B_c_1334_n N_A_1745_329#_c_1571_n 0.0717923f $X=10.78 $Y=1.63 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1337_n N_A_1745_329#_c_1571_n 0.00136362f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_960 N_SET_B_c_1338_n N_A_1745_329#_c_1571_n 0.0133627f $X=9.875 $Y=1.53 $X2=0
+ $Y2=0
cc_961 N_SET_B_M1015_g N_A_1745_329#_c_1563_n 0.00837676f $X=10.89 $Y=0.445
+ $X2=0 $Y2=0
cc_962 N_SET_B_M1015_g N_A_1745_329#_c_1564_n 0.00528915f $X=10.89 $Y=0.445
+ $X2=0 $Y2=0
cc_963 N_SET_B_M1015_g N_A_1745_329#_c_1565_n 0.00603615f $X=10.89 $Y=0.445
+ $X2=0 $Y2=0
cc_964 N_SET_B_c_1331_n N_A_1745_329#_c_1566_n 0.0182994f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_965 N_SET_B_c_1331_n N_A_1745_329#_c_1572_n 5.50243e-19 $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_966 N_SET_B_c_1331_n N_A_1745_329#_c_1573_n 9.04123e-19 $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_967 N_SET_B_c_1335_n N_A_1745_329#_c_1573_n 0.00169667f $X=9.73 $Y=1.53 $X2=0
+ $Y2=0
cc_968 N_SET_B_c_1337_n N_A_1745_329#_c_1573_n 6.9852e-19 $X=9.875 $Y=1.53 $X2=0
+ $Y2=0
cc_969 N_SET_B_c_1338_n N_A_1745_329#_c_1573_n 0.00798024f $X=9.875 $Y=1.53
+ $X2=0 $Y2=0
cc_970 N_SET_B_c_1331_n N_A_1745_329#_c_1574_n 0.00268766f $X=10.565 $Y=1.99
+ $X2=0 $Y2=0
cc_971 N_SET_B_c_1334_n N_A_1745_329#_c_1574_n 0.00864864f $X=10.78 $Y=1.63
+ $X2=0 $Y2=0
cc_972 N_SET_B_c_1330_n N_VPWR_c_1847_n 0.00384082f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_973 N_SET_B_c_1331_n N_VPWR_c_1848_n 0.00533f $X=10.565 $Y=1.99 $X2=0 $Y2=0
cc_974 N_SET_B_c_1331_n N_VPWR_c_1849_n 0.00569972f $X=10.565 $Y=1.99 $X2=0
+ $Y2=0
cc_975 N_SET_B_c_1331_n N_VPWR_c_1850_n 0.00241392f $X=10.565 $Y=1.99 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1330_n N_VPWR_c_1855_n 0.00743866f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_977 N_SET_B_c_1335_n N_VPWR_c_1868_n 0.00119777f $X=9.73 $Y=1.53 $X2=0 $Y2=0
cc_978 N_SET_B_c_1330_n N_VPWR_c_1842_n 0.00869097f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_979 N_SET_B_c_1331_n N_VPWR_c_1842_n 0.00836421f $X=10.565 $Y=1.99 $X2=0
+ $Y2=0
cc_980 N_SET_B_M1015_g N_VGND_c_2248_n 0.0053804f $X=10.89 $Y=0.445 $X2=0 $Y2=0
cc_981 N_SET_B_M1015_g N_VGND_c_2258_n 0.00443798f $X=10.89 $Y=0.445 $X2=0 $Y2=0
cc_982 N_SET_B_M1017_g N_VGND_c_2264_n 0.0278746f $X=7.67 $Y=0.445 $X2=0 $Y2=0
cc_983 N_SET_B_c_1328_n N_VGND_c_2264_n 4.5828e-19 $X=7.62 $Y=1.365 $X2=0 $Y2=0
cc_984 N_SET_B_M1015_g N_VGND_c_2267_n 0.00656367f $X=10.89 $Y=0.445 $X2=0 $Y2=0
cc_985 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1557_n 0.0210784f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_986 N_A_1951_295#_c_1470_n N_A_1745_329#_c_1557_n 0.0278731f $X=11.84
+ $Y=2.285 $X2=0 $Y2=0
cc_987 N_A_1951_295#_c_1461_n N_A_1745_329#_c_1557_n 6.05607e-19 $X=11.84
+ $Y=0.42 $X2=0 $Y2=0
cc_988 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1558_n 0.0020184f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_989 N_A_1951_295#_c_1462_n N_A_1745_329#_c_1558_n 0.0180509f $X=11.885
+ $Y=1.28 $X2=0 $Y2=0
cc_990 N_A_1951_295#_c_1460_n N_A_1745_329#_M1030_g 6.78474e-19 $X=11.9 $Y=1.195
+ $X2=0 $Y2=0
cc_991 N_A_1951_295#_c_1461_n N_A_1745_329#_M1030_g 9.48411e-19 $X=11.84 $Y=0.42
+ $X2=0 $Y2=0
cc_992 N_A_1951_295#_c_1460_n N_A_1745_329#_c_1560_n 0.00150633f $X=11.9
+ $Y=1.195 $X2=0 $Y2=0
cc_993 N_A_1951_295#_c_1460_n N_A_1745_329#_c_1561_n 0.00693654f $X=11.9
+ $Y=1.195 $X2=0 $Y2=0
cc_994 N_A_1951_295#_c_1461_n N_A_1745_329#_c_1561_n 0.0082592f $X=11.84 $Y=0.42
+ $X2=0 $Y2=0
cc_995 N_A_1951_295#_c_1464_n N_A_1745_329#_c_1578_n 5.33833e-19 $X=9.855
+ $Y=1.99 $X2=0 $Y2=0
cc_996 N_A_1951_295#_M1002_g N_A_1745_329#_c_1579_n 0.0160958f $X=10.26 $Y=0.445
+ $X2=0 $Y2=0
cc_997 N_A_1951_295#_c_1457_n N_A_1745_329#_c_1579_n 0.0100001f $X=10.32 $Y=1.02
+ $X2=0 $Y2=0
cc_998 N_A_1951_295#_c_1458_n N_A_1745_329#_c_1579_n 0.00137429f $X=10.32
+ $Y=1.02 $X2=0 $Y2=0
cc_999 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1579_n 0.00662734f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1000 N_A_1951_295#_c_1464_n N_A_1745_329#_c_1571_n 0.0101951f $X=9.855
+ $Y=1.99 $X2=0 $Y2=0
cc_1001 N_A_1951_295#_c_1465_n N_A_1745_329#_c_1571_n 0.00233365f $X=10.185
+ $Y=1.55 $X2=0 $Y2=0
cc_1002 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1571_n 7.15895e-19 $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1003 N_A_1951_295#_M1002_g N_A_1745_329#_c_1563_n 0.0043272f $X=10.26
+ $Y=0.445 $X2=0 $Y2=0
cc_1004 N_A_1951_295#_M1002_g N_A_1745_329#_c_1564_n 0.00161591f $X=10.26
+ $Y=0.445 $X2=0 $Y2=0
cc_1005 N_A_1951_295#_c_1457_n N_A_1745_329#_c_1564_n 0.010594f $X=10.32 $Y=1.02
+ $X2=0 $Y2=0
cc_1006 N_A_1951_295#_c_1458_n N_A_1745_329#_c_1564_n 0.00125223f $X=10.32
+ $Y=1.02 $X2=0 $Y2=0
cc_1007 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1564_n 0.0154264f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1008 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1565_n 0.0492513f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1009 N_A_1951_295#_c_1460_n N_A_1745_329#_c_1565_n 0.0196589f $X=11.9
+ $Y=1.195 $X2=0 $Y2=0
cc_1010 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1566_n 0.0050268f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1011 N_A_1951_295#_c_1460_n N_A_1745_329#_c_1566_n 0.0067596f $X=11.9
+ $Y=1.195 $X2=0 $Y2=0
cc_1012 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1572_n 0.00650879f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1013 N_A_1951_295#_c_1464_n N_A_1745_329#_c_1573_n 0.01527f $X=9.855 $Y=1.99
+ $X2=0 $Y2=0
cc_1014 N_A_1951_295#_c_1459_n N_A_1745_329#_c_1574_n 0.0213588f $X=11.755
+ $Y=1.28 $X2=0 $Y2=0
cc_1015 N_A_1951_295#_c_1470_n N_A_1745_329#_c_1574_n 0.0360588f $X=11.84
+ $Y=2.285 $X2=0 $Y2=0
cc_1016 N_A_1951_295#_c_1461_n N_A_2447_47#_c_1701_n 0.0596014f $X=11.84 $Y=0.42
+ $X2=0 $Y2=0
cc_1017 N_A_1951_295#_c_1470_n N_A_2447_47#_c_1709_n 0.0883081f $X=11.84
+ $Y=2.285 $X2=0 $Y2=0
cc_1018 N_A_1951_295#_c_1462_n N_A_2447_47#_c_1709_n 0.0031876f $X=11.885
+ $Y=1.28 $X2=0 $Y2=0
cc_1019 N_A_1951_295#_c_1460_n N_A_2447_47#_c_1703_n 0.0172077f $X=11.9 $Y=1.195
+ $X2=0 $Y2=0
cc_1020 N_A_1951_295#_c_1462_n N_A_2447_47#_c_1703_n 0.0110951f $X=11.885
+ $Y=1.28 $X2=0 $Y2=0
cc_1021 N_A_1951_295#_c_1464_n N_VPWR_c_1848_n 0.00588614f $X=9.855 $Y=1.99
+ $X2=0 $Y2=0
cc_1022 N_A_1951_295#_c_1470_n N_VPWR_c_1850_n 0.0177194f $X=11.84 $Y=2.285
+ $X2=0 $Y2=0
cc_1023 N_A_1951_295#_c_1464_n N_VPWR_c_1861_n 0.00486131f $X=9.855 $Y=1.99
+ $X2=0 $Y2=0
cc_1024 N_A_1951_295#_c_1470_n N_VPWR_c_1862_n 0.0182101f $X=11.84 $Y=2.285
+ $X2=0 $Y2=0
cc_1025 N_A_1951_295#_M1004_d N_VPWR_c_1842_n 0.00404917f $X=11.695 $Y=2.065
+ $X2=0 $Y2=0
cc_1026 N_A_1951_295#_c_1464_n N_VPWR_c_1842_n 0.0071443f $X=9.855 $Y=1.99 $X2=0
+ $Y2=0
cc_1027 N_A_1951_295#_c_1470_n N_VPWR_c_1842_n 0.00993603f $X=11.84 $Y=2.285
+ $X2=0 $Y2=0
cc_1028 N_A_1951_295#_M1002_g N_VGND_c_2258_n 0.00362032f $X=10.26 $Y=0.445
+ $X2=0 $Y2=0
cc_1029 N_A_1951_295#_c_1461_n N_VGND_c_2259_n 0.0234496f $X=11.84 $Y=0.42 $X2=0
+ $Y2=0
cc_1030 N_A_1951_295#_M1022_d N_VGND_c_2267_n 0.00537869f $X=11.585 $Y=0.235
+ $X2=0 $Y2=0
cc_1031 N_A_1951_295#_M1002_g N_VGND_c_2267_n 0.00561157f $X=10.26 $Y=0.445
+ $X2=0 $Y2=0
cc_1032 N_A_1951_295#_c_1461_n N_VGND_c_2267_n 0.0129422f $X=11.84 $Y=0.42 $X2=0
+ $Y2=0
cc_1033 N_A_1745_329#_c_1569_n N_A_2447_47#_c_1705_n 0.00741781f $X=12.595
+ $Y=1.41 $X2=0 $Y2=0
cc_1034 N_A_1745_329#_M1030_g N_A_2447_47#_c_1697_n 0.0153146f $X=12.62 $Y=0.56
+ $X2=0 $Y2=0
cc_1035 N_A_1745_329#_M1030_g N_A_2447_47#_c_1701_n 0.0119139f $X=12.62 $Y=0.56
+ $X2=0 $Y2=0
cc_1036 N_A_1745_329#_c_1557_n N_A_2447_47#_c_1709_n 9.01204e-19 $X=11.605
+ $Y=1.99 $X2=0 $Y2=0
cc_1037 N_A_1745_329#_c_1558_n N_A_2447_47#_c_1709_n 0.00786815f $X=12.495
+ $Y=1.28 $X2=0 $Y2=0
cc_1038 N_A_1745_329#_c_1569_n N_A_2447_47#_c_1709_n 0.0117043f $X=12.595
+ $Y=1.41 $X2=0 $Y2=0
cc_1039 N_A_1745_329#_c_1562_n N_A_2447_47#_c_1709_n 0.00233005f $X=12.595
+ $Y=1.307 $X2=0 $Y2=0
cc_1040 N_A_1745_329#_c_1558_n N_A_2447_47#_c_1702_n 0.0026182f $X=12.495
+ $Y=1.28 $X2=0 $Y2=0
cc_1041 N_A_1745_329#_M1030_g N_A_2447_47#_c_1702_n 0.0136669f $X=12.62 $Y=0.56
+ $X2=0 $Y2=0
cc_1042 N_A_1745_329#_c_1562_n N_A_2447_47#_c_1702_n 0.0100836f $X=12.595
+ $Y=1.307 $X2=0 $Y2=0
cc_1043 N_A_1745_329#_c_1558_n N_A_2447_47#_c_1703_n 0.0109356f $X=12.495
+ $Y=1.28 $X2=0 $Y2=0
cc_1044 N_A_1745_329#_c_1566_n N_A_2447_47#_c_1703_n 2.95577e-19 $X=11.4 $Y=0.93
+ $X2=0 $Y2=0
cc_1045 N_A_1745_329#_M1030_g N_A_2447_47#_c_1704_n 0.021471f $X=12.62 $Y=0.56
+ $X2=0 $Y2=0
cc_1046 N_A_1745_329#_c_1562_n N_A_2447_47#_c_1704_n 0.00336889f $X=12.595
+ $Y=1.307 $X2=0 $Y2=0
cc_1047 N_A_1745_329#_c_1574_n N_VPWR_M1004_s 0.0028505f $X=11.37 $Y=1.69 $X2=0
+ $Y2=0
cc_1048 N_A_1745_329#_c_1571_n N_VPWR_c_1848_n 0.0285361f $X=10.61 $Y=1.98 $X2=0
+ $Y2=0
cc_1049 N_A_1745_329#_c_1573_n N_VPWR_c_1848_n 0.0138202f $X=9.755 $Y=1.98 $X2=0
+ $Y2=0
cc_1050 N_A_1745_329#_c_1571_n N_VPWR_c_1849_n 0.0263725f $X=10.61 $Y=1.98 $X2=0
+ $Y2=0
cc_1051 N_A_1745_329#_c_1572_n N_VPWR_c_1849_n 0.00332039f $X=11.205 $Y=1.98
+ $X2=0 $Y2=0
cc_1052 N_A_1745_329#_c_1557_n N_VPWR_c_1850_n 0.0135992f $X=11.605 $Y=1.99
+ $X2=0 $Y2=0
cc_1053 N_A_1745_329#_c_1571_n N_VPWR_c_1850_n 0.0169944f $X=10.61 $Y=1.98 $X2=0
+ $Y2=0
cc_1054 N_A_1745_329#_c_1574_n N_VPWR_c_1850_n 0.0284102f $X=11.37 $Y=1.69 $X2=0
+ $Y2=0
cc_1055 N_A_1745_329#_c_1569_n N_VPWR_c_1851_n 0.0220697f $X=12.595 $Y=1.41
+ $X2=0 $Y2=0
cc_1056 N_A_1745_329#_c_1578_n N_VPWR_c_1861_n 0.0435125f $X=9.67 $Y=2.292 $X2=0
+ $Y2=0
cc_1057 N_A_1745_329#_c_1571_n N_VPWR_c_1861_n 0.00364691f $X=10.61 $Y=1.98
+ $X2=0 $Y2=0
cc_1058 N_A_1745_329#_c_1573_n N_VPWR_c_1861_n 0.00927152f $X=9.755 $Y=1.98
+ $X2=0 $Y2=0
cc_1059 N_A_1745_329#_c_1557_n N_VPWR_c_1862_n 0.00448207f $X=11.605 $Y=1.99
+ $X2=0 $Y2=0
cc_1060 N_A_1745_329#_c_1569_n N_VPWR_c_1862_n 0.00427505f $X=12.595 $Y=1.41
+ $X2=0 $Y2=0
cc_1061 N_A_1745_329#_M1034_d N_VPWR_c_1842_n 0.00651684f $X=8.725 $Y=1.645
+ $X2=0 $Y2=0
cc_1062 N_A_1745_329#_M1003_d N_VPWR_c_1842_n 0.00259177f $X=10.655 $Y=2.065
+ $X2=0 $Y2=0
cc_1063 N_A_1745_329#_c_1557_n N_VPWR_c_1842_n 0.00895167f $X=11.605 $Y=1.99
+ $X2=0 $Y2=0
cc_1064 N_A_1745_329#_c_1569_n N_VPWR_c_1842_n 0.00861212f $X=12.595 $Y=1.41
+ $X2=0 $Y2=0
cc_1065 N_A_1745_329#_c_1578_n N_VPWR_c_1842_n 0.0268944f $X=9.67 $Y=2.292 $X2=0
+ $Y2=0
cc_1066 N_A_1745_329#_c_1571_n N_VPWR_c_1842_n 0.0263862f $X=10.61 $Y=1.98 $X2=0
+ $Y2=0
cc_1067 N_A_1745_329#_c_1572_n N_VPWR_c_1842_n 0.00529988f $X=11.205 $Y=1.98
+ $X2=0 $Y2=0
cc_1068 N_A_1745_329#_c_1573_n N_VPWR_c_1842_n 0.00608385f $X=9.755 $Y=1.98
+ $X2=0 $Y2=0
cc_1069 N_A_1745_329#_c_1574_n N_VPWR_c_1842_n 0.0017435f $X=11.37 $Y=1.69 $X2=0
+ $Y2=0
cc_1070 N_A_1745_329#_c_1578_n A_1891_413# 0.00509751f $X=9.67 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1071 N_A_1745_329#_c_1573_n A_1891_413# 0.00191133f $X=9.755 $Y=1.98
+ $X2=-0.19 $Y2=-0.24
cc_1072 N_A_1745_329#_c_1560_n N_VGND_c_2248_n 0.00383167f $X=11.425 $Y=0.925
+ $X2=0 $Y2=0
cc_1073 N_A_1745_329#_c_1561_n N_VGND_c_2248_n 0.00326191f $X=11.425 $Y=0.765
+ $X2=0 $Y2=0
cc_1074 N_A_1745_329#_c_1579_n N_VGND_c_2248_n 0.01594f $X=10.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1075 N_A_1745_329#_c_1565_n N_VGND_c_2248_n 0.0134367f $X=11.4 $Y=0.93 $X2=0
+ $Y2=0
cc_1076 N_A_1745_329#_M1030_g N_VGND_c_2249_n 0.0165842f $X=12.62 $Y=0.56 $X2=0
+ $Y2=0
cc_1077 N_A_1745_329#_c_1579_n N_VGND_c_2258_n 0.0875792f $X=10.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1078 N_A_1745_329#_M1030_g N_VGND_c_2259_n 0.00271402f $X=12.62 $Y=0.56 $X2=0
+ $Y2=0
cc_1079 N_A_1745_329#_c_1560_n N_VGND_c_2259_n 3.91476e-19 $X=11.425 $Y=0.925
+ $X2=0 $Y2=0
cc_1080 N_A_1745_329#_c_1561_n N_VGND_c_2259_n 0.00585385f $X=11.425 $Y=0.765
+ $X2=0 $Y2=0
cc_1081 N_A_1745_329#_M1045_d N_VGND_c_2267_n 0.00520375f $X=9.215 $Y=0.235
+ $X2=0 $Y2=0
cc_1082 N_A_1745_329#_M1030_g N_VGND_c_2267_n 0.00621952f $X=12.62 $Y=0.56 $X2=0
+ $Y2=0
cc_1083 N_A_1745_329#_c_1560_n N_VGND_c_2267_n 5.20533e-19 $X=11.425 $Y=0.925
+ $X2=0 $Y2=0
cc_1084 N_A_1745_329#_c_1561_n N_VGND_c_2267_n 0.00782368f $X=11.425 $Y=0.765
+ $X2=0 $Y2=0
cc_1085 N_A_1745_329#_c_1579_n N_VGND_c_2267_n 0.0595549f $X=10.71 $Y=0.41 $X2=0
+ $Y2=0
cc_1086 N_A_1745_329#_c_1565_n N_VGND_c_2267_n 0.0162134f $X=11.4 $Y=0.93 $X2=0
+ $Y2=0
cc_1087 N_A_1745_329#_c_1579_n A_1995_47# 0.00482916f $X=10.71 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1088 N_A_1745_329#_c_1579_n A_2067_47# 0.0111297f $X=10.71 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1089 N_A_1745_329#_c_1563_n A_2067_47# 0.0015298f $X=10.81 $Y=0.785 $X2=-0.19
+ $Y2=-0.24
cc_1090 N_A_2447_47#_c_1705_n N_VPWR_c_1851_n 0.00331097f $X=13.12 $Y=1.41 $X2=0
+ $Y2=0
cc_1091 N_A_2447_47#_c_1709_n N_VPWR_c_1851_n 0.0750937f $X=12.36 $Y=1.955 $X2=0
+ $Y2=0
cc_1092 N_A_2447_47#_c_1702_n N_VPWR_c_1851_n 0.0292881f $X=13.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1093 N_A_2447_47#_c_1704_n N_VPWR_c_1851_n 0.00251554f $X=14.58 $Y=1.202
+ $X2=0 $Y2=0
cc_1094 N_A_2447_47#_c_1706_n N_VPWR_c_1852_n 0.00608635f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1095 N_A_2447_47#_c_1707_n N_VPWR_c_1852_n 0.00575827f $X=14.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1096 N_A_2447_47#_c_1704_n N_VPWR_c_1852_n 0.00391367f $X=14.58 $Y=1.202
+ $X2=0 $Y2=0
cc_1097 N_A_2447_47#_c_1708_n N_VPWR_c_1854_n 0.00719044f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1098 N_A_2447_47#_c_1705_n N_VPWR_c_1856_n 0.00702461f $X=13.12 $Y=1.41 $X2=0
+ $Y2=0
cc_1099 N_A_2447_47#_c_1706_n N_VPWR_c_1856_n 0.0059915f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1100 N_A_2447_47#_c_1709_n N_VPWR_c_1862_n 0.0182101f $X=12.36 $Y=1.955 $X2=0
+ $Y2=0
cc_1101 N_A_2447_47#_c_1707_n N_VPWR_c_1863_n 0.00597712f $X=14.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1102 N_A_2447_47#_c_1708_n N_VPWR_c_1863_n 0.00521806f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1103 N_A_2447_47#_M1040_s N_VPWR_c_1842_n 0.00425811f $X=12.235 $Y=1.485
+ $X2=0 $Y2=0
cc_1104 N_A_2447_47#_c_1705_n N_VPWR_c_1842_n 0.0125663f $X=13.12 $Y=1.41 $X2=0
+ $Y2=0
cc_1105 N_A_2447_47#_c_1706_n N_VPWR_c_1842_n 0.0102479f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1106 N_A_2447_47#_c_1707_n N_VPWR_c_1842_n 0.0101168f $X=14.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1107 N_A_2447_47#_c_1708_n N_VPWR_c_1842_n 0.00923842f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1108 N_A_2447_47#_c_1709_n N_VPWR_c_1842_n 0.00993603f $X=12.36 $Y=1.955
+ $X2=0 $Y2=0
cc_1109 N_A_2447_47#_c_1698_n N_Q_c_2195_n 0.00505877f $X=13.615 $Y=0.995 $X2=0
+ $Y2=0
cc_1110 N_A_2447_47#_c_1699_n N_Q_c_2195_n 5.10522e-19 $X=14.135 $Y=0.995 $X2=0
+ $Y2=0
cc_1111 N_A_2447_47#_c_1706_n N_Q_c_2197_n 0.00416752f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1112 N_A_2447_47#_c_1704_n N_Q_c_2197_n 0.00315148f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1113 N_A_2447_47#_c_1706_n N_Q_c_2199_n 0.0169431f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1114 N_A_2447_47#_c_1697_n N_Q_c_2193_n 0.00397629f $X=13.145 $Y=0.995 $X2=0
+ $Y2=0
cc_1115 N_A_2447_47#_c_1698_n N_Q_c_2193_n 0.00431943f $X=13.615 $Y=0.995 $X2=0
+ $Y2=0
cc_1116 N_A_2447_47#_c_1702_n N_Q_c_2193_n 0.00369613f $X=13.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1117 N_A_2447_47#_c_1704_n N_Q_c_2193_n 0.00620199f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1118 N_A_2447_47#_c_1698_n N_Q_c_2204_n 0.00382124f $X=13.615 $Y=0.995 $X2=0
+ $Y2=0
cc_1119 N_A_2447_47#_c_1704_n N_Q_c_2204_n 0.00103509f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1120 N_A_2447_47#_c_1705_n N_Q_c_2194_n 0.00193705f $X=13.12 $Y=1.41 $X2=0
+ $Y2=0
cc_1121 N_A_2447_47#_c_1706_n N_Q_c_2194_n 0.00248354f $X=13.59 $Y=1.41 $X2=0
+ $Y2=0
cc_1122 N_A_2447_47#_c_1707_n N_Q_c_2194_n 5.49783e-19 $X=14.11 $Y=1.41 $X2=0
+ $Y2=0
cc_1123 N_A_2447_47#_c_1704_n N_Q_c_2194_n 0.00502225f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1124 N_A_2447_47#_c_1702_n N_Q_c_2210_n 0.0184883f $X=13.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1125 N_A_2447_47#_c_1704_n N_Q_c_2210_n 0.0136336f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1126 N_A_2447_47#_c_1704_n Q 0.0308047f $X=14.58 $Y=1.202 $X2=0 $Y2=0
cc_1127 N_A_2447_47#_c_1706_n Q 4.86048e-19 $X=13.59 $Y=1.41 $X2=0 $Y2=0
cc_1128 N_A_2447_47#_c_1707_n Q 0.0169696f $X=14.11 $Y=1.41 $X2=0 $Y2=0
cc_1129 N_A_2447_47#_c_1708_n Q 0.0236541f $X=14.58 $Y=1.41 $X2=0 $Y2=0
cc_1130 N_A_2447_47#_c_1704_n Q 0.00924318f $X=14.58 $Y=1.202 $X2=0 $Y2=0
cc_1131 N_A_2447_47#_c_1704_n N_Q_c_2217_n 0.0508509f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1132 N_A_2447_47#_c_1698_n N_Q_c_2218_n 5.26774e-19 $X=13.615 $Y=0.995 $X2=0
+ $Y2=0
cc_1133 N_A_2447_47#_c_1699_n N_Q_c_2218_n 0.0132952f $X=14.135 $Y=0.995 $X2=0
+ $Y2=0
cc_1134 N_A_2447_47#_c_1700_n N_Q_c_2218_n 0.0165529f $X=14.605 $Y=0.995 $X2=0
+ $Y2=0
cc_1135 N_A_2447_47#_c_1704_n N_Q_c_2218_n 0.0101075f $X=14.58 $Y=1.202 $X2=0
+ $Y2=0
cc_1136 N_A_2447_47#_c_1697_n N_VGND_c_2249_n 0.00631549f $X=13.145 $Y=0.995
+ $X2=0 $Y2=0
cc_1137 N_A_2447_47#_c_1701_n N_VGND_c_2249_n 0.0441275f $X=12.36 $Y=0.425 $X2=0
+ $Y2=0
cc_1138 N_A_2447_47#_c_1702_n N_VGND_c_2249_n 0.0310557f $X=13.04 $Y=1.16 $X2=0
+ $Y2=0
cc_1139 N_A_2447_47#_c_1704_n N_VGND_c_2249_n 0.00263742f $X=14.58 $Y=1.202
+ $X2=0 $Y2=0
cc_1140 N_A_2447_47#_c_1698_n N_VGND_c_2250_n 0.00522013f $X=13.615 $Y=0.995
+ $X2=0 $Y2=0
cc_1141 N_A_2447_47#_c_1699_n N_VGND_c_2250_n 0.00448853f $X=14.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1142 N_A_2447_47#_c_1704_n N_VGND_c_2250_n 0.00420888f $X=14.58 $Y=1.202
+ $X2=0 $Y2=0
cc_1143 N_A_2447_47#_c_1700_n N_VGND_c_2252_n 0.00631115f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1144 N_A_2447_47#_c_1697_n N_VGND_c_2255_n 0.00585385f $X=13.145 $Y=0.995
+ $X2=0 $Y2=0
cc_1145 N_A_2447_47#_c_1698_n N_VGND_c_2255_n 0.00542163f $X=13.615 $Y=0.995
+ $X2=0 $Y2=0
cc_1146 N_A_2447_47#_c_1701_n N_VGND_c_2259_n 0.0182101f $X=12.36 $Y=0.425 $X2=0
+ $Y2=0
cc_1147 N_A_2447_47#_c_1699_n N_VGND_c_2260_n 0.00465454f $X=14.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1148 N_A_2447_47#_c_1700_n N_VGND_c_2260_n 0.00465454f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1149 N_A_2447_47#_M1030_s N_VGND_c_2267_n 0.00600004f $X=12.235 $Y=0.235
+ $X2=0 $Y2=0
cc_1150 N_A_2447_47#_c_1697_n N_VGND_c_2267_n 0.0110943f $X=13.145 $Y=0.995
+ $X2=0 $Y2=0
cc_1151 N_A_2447_47#_c_1698_n N_VGND_c_2267_n 0.0100384f $X=13.615 $Y=0.995
+ $X2=0 $Y2=0
cc_1152 N_A_2447_47#_c_1699_n N_VGND_c_2267_n 0.00814434f $X=14.135 $Y=0.995
+ $X2=0 $Y2=0
cc_1153 N_A_2447_47#_c_1700_n N_VGND_c_2267_n 0.00894281f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1154 N_A_2447_47#_c_1701_n N_VGND_c_2267_n 0.00993603f $X=12.36 $Y=0.425
+ $X2=0 $Y2=0
cc_1155 N_A_27_369#_c_1797_n N_VPWR_M1010_d 0.00342966f $X=1.055 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_1156 N_A_27_369#_c_1796_n N_VPWR_c_1843_n 0.0205323f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1157 N_A_27_369#_c_1797_n N_VPWR_c_1843_n 0.0187115f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1158 N_A_27_369#_c_1796_n N_VPWR_c_1858_n 0.0180865f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1159 N_A_27_369#_c_1797_n N_VPWR_c_1858_n 0.00206566f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1160 N_A_27_369#_c_1797_n N_VPWR_c_1859_n 0.00290212f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1161 N_A_27_369#_c_1810_n N_VPWR_c_1859_n 0.00991509f $X=1.225 $Y=2.36 $X2=0
+ $Y2=0
cc_1162 N_A_27_369#_c_1799_n N_VPWR_c_1859_n 0.0582047f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1163 N_A_27_369#_M1010_s N_VPWR_c_1842_n 0.00244672f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1164 N_A_27_369#_M1026_d N_VPWR_c_1842_n 0.00217543f $X=1.935 $Y=1.845 $X2=0
+ $Y2=0
cc_1165 N_A_27_369#_c_1796_n N_VPWR_c_1842_n 0.00991202f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1166 N_A_27_369#_c_1797_n N_VPWR_c_1842_n 0.0103345f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1167 N_A_27_369#_c_1810_n N_VPWR_c_1842_n 0.00653118f $X=1.225 $Y=2.36 $X2=0
+ $Y2=0
cc_1168 N_A_27_369#_c_1799_n N_VPWR_c_1842_n 0.0364411f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1169 N_A_27_369#_c_1797_n A_211_369# 0.00274315f $X=1.055 $Y=1.935 $X2=-0.19
+ $Y2=1.305
cc_1170 N_A_27_369#_c_1813_n A_211_369# 0.00234118f $X=1.14 $Y=2.255 $X2=-0.19
+ $Y2=1.305
cc_1171 N_A_27_369#_c_1810_n A_211_369# 0.00110197f $X=1.225 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1172 N_A_27_369#_c_1799_n N_A_201_47#_M1041_d 0.0035404f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1173 N_A_27_369#_c_1797_n N_A_201_47#_c_2071_n 0.0151838f $X=1.055 $Y=1.935
+ $X2=0 $Y2=0
cc_1174 N_A_27_369#_c_1813_n N_A_201_47#_c_2071_n 0.00444947f $X=1.14 $Y=2.255
+ $X2=0 $Y2=0
cc_1175 N_A_27_369#_c_1799_n N_A_201_47#_c_2071_n 0.0229871f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1176 N_A_27_369#_c_1799_n N_A_201_47#_c_2064_n 0.00286705f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1177 N_VPWR_c_1842_n A_211_369# 0.00184693f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1178 N_VPWR_c_1842_n N_A_201_47#_M1041_d 0.00232895f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1179 N_VPWR_c_1842_n N_A_201_47#_M1008_s 0.0020949f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1180 N_VPWR_c_1860_n N_A_201_47#_c_2062_n 0.0135499f $X=6.445 $Y=2.72 $X2=0
+ $Y2=0
cc_1181 N_VPWR_c_1842_n N_A_201_47#_c_2062_n 0.00390749f $X=14.95 $Y=2.72 $X2=0
+ $Y2=0
cc_1182 N_VPWR_c_1844_n N_A_201_47#_c_2063_n 0.00826221f $X=3.07 $Y=2.34 $X2=0
+ $Y2=0
cc_1183 N_VPWR_c_1842_n A_1169_413# 0.00263276f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1184 N_VPWR_c_1846_n A_1663_329# 5.2056e-19 $X=8.425 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1185 N_VPWR_c_1868_n A_1663_329# 6.30678e-19 $X=8.765 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1186 N_VPWR_c_1842_n A_1891_413# 0.0024832f $X=14.95 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1187 N_VPWR_c_1842_n N_Q_M1012_d 0.0033595f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1188 N_VPWR_c_1842_n N_Q_M1025_d 0.00231261f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1189 N_VPWR_c_1852_n N_Q_c_2197_n 0.0577881f $X=13.875 $Y=1.66 $X2=0 $Y2=0
cc_1190 N_VPWR_c_1856_n N_Q_c_2199_n 0.0182467f $X=13.79 $Y=2.72 $X2=0 $Y2=0
cc_1191 N_VPWR_c_1842_n N_Q_c_2199_n 0.0121511f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1192 N_VPWR_c_1852_n Q 0.0737678f $X=13.875 $Y=1.66 $X2=0 $Y2=0
cc_1193 N_VPWR_c_1854_n Q 0.0766009f $X=14.865 $Y=1.66 $X2=0 $Y2=0
cc_1194 N_VPWR_c_1863_n Q 0.0291737f $X=14.78 $Y=2.72 $X2=0 $Y2=0
cc_1195 N_VPWR_c_1842_n Q 0.017404f $X=14.95 $Y=2.72 $X2=0 $Y2=0
cc_1196 N_VPWR_c_1852_n N_Q_c_2217_n 0.0136818f $X=13.875 $Y=1.66 $X2=0 $Y2=0
cc_1197 N_VPWR_c_1854_n N_VGND_c_2252_n 0.010033f $X=14.865 $Y=1.66 $X2=0 $Y2=0
cc_1198 N_A_201_47#_c_2068_n N_VGND_c_2242_n 0.0541179f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1199 N_A_201_47#_c_2068_n N_VGND_c_2243_n 0.0294921f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1200 N_A_201_47#_c_2068_n N_VGND_c_2244_n 0.0224969f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1201 N_A_201_47#_c_2057_n N_VGND_c_2257_n 0.0226408f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1202 N_A_201_47#_M1037_d N_VGND_c_2267_n 0.00255381f $X=1.005 $Y=0.235 $X2=0
+ $Y2=0
cc_1203 N_A_201_47#_M1033_s N_VGND_c_2267_n 0.0054218f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_1204 N_A_201_47#_c_2068_n N_VGND_c_2267_n 0.0334433f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1205 N_A_201_47#_c_2057_n N_VGND_c_2267_n 0.0123998f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1206 N_A_201_47#_c_2068_n A_295_47# 0.00393714f $X=1.655 $Y=0.425 $X2=-0.19
+ $Y2=-0.24
cc_1207 N_A_201_47#_c_2059_n A_295_47# 6.98288e-19 $X=1.76 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1208 N_Q_c_2195_n N_VGND_c_2250_n 0.0367673f $X=13.355 $Y=0.44 $X2=0 $Y2=0
cc_1209 N_Q_c_2217_n N_VGND_c_2250_n 0.0136816f $X=14.13 $Y=1.19 $X2=0 $Y2=0
cc_1210 N_Q_c_2218_n N_VGND_c_2250_n 0.0479113f $X=14.345 $Y=0.36 $X2=0 $Y2=0
cc_1211 N_Q_c_2218_n N_VGND_c_2252_n 0.049751f $X=14.345 $Y=0.36 $X2=0 $Y2=0
cc_1212 N_Q_c_2195_n N_VGND_c_2255_n 0.0174424f $X=13.355 $Y=0.44 $X2=0 $Y2=0
cc_1213 N_Q_c_2218_n N_VGND_c_2260_n 0.0292379f $X=14.345 $Y=0.36 $X2=0 $Y2=0
cc_1214 N_Q_M1009_s N_VGND_c_2267_n 0.00330789f $X=13.22 $Y=0.235 $X2=0 $Y2=0
cc_1215 N_Q_M1036_s N_VGND_c_2267_n 0.0025535f $X=14.21 $Y=0.235 $X2=0 $Y2=0
cc_1216 N_Q_c_2195_n N_VGND_c_2267_n 0.0123424f $X=13.355 $Y=0.44 $X2=0 $Y2=0
cc_1217 N_Q_c_2218_n N_VGND_c_2267_n 0.0175412f $X=14.345 $Y=0.36 $X2=0 $Y2=0
cc_1218 N_VGND_c_2243_n A_119_47# 0.00411471f $X=0.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1219 N_VGND_c_2267_n A_119_47# 0.00142631f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1220 N_VGND_c_2267_n A_295_47# 0.00216824f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1221 N_VGND_c_2257_n A_1177_47# 0.00329703f $X=6.06 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1222 N_VGND_c_2267_n A_1177_47# 0.00735224f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1223 N_VGND_c_2264_n A_1654_47# 0.0117508f $X=8.415 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1224 N_VGND_c_2267_n A_1654_47# 0.0135294f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1225 N_VGND_c_2267_n A_1995_47# 0.00169327f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1226 N_VGND_c_2267_n A_2067_47# 0.00389027f $X=14.95 $Y=0 $X2=-0.19 $Y2=-0.24
