* File: sky130_fd_sc_hdll__nand4bb_2.spice
* Created: Thu Aug 27 19:15:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4bb_2.pex.spice"
.subckt sky130_fd_sc_hdll__nand4bb_2  VNB VPB B_N A_N C D VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* D	D
* C	C
* A_N	A_N
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_B_N_M1012_g N_A_27_47#_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.9 A=0.063 P=1.14 MULT=1
MM1000 N_A_211_413#_M1000_d N_A_N_M1000_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1974 AS=0.0672 PD=1.78 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1003 N_A_361_47#_M1003_d N_A_211_413#_M1003_g N_Y_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_361_47#_M1004_d N_A_211_413#_M1004_g N_Y_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1015 N_A_361_47#_M1004_d N_A_27_47#_M1015_g N_A_641_47#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1018 N_A_361_47#_M1018_d N_A_27_47#_M1018_g N_A_641_47#_M1015_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_841_47#_M1011_d N_C_M1011_g N_A_641_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.104 PD=1.86 PS=0.97 NRD=2.76 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1019 N_A_841_47#_M1019_d N_C_M1019_g N_A_641_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_A_841_47#_M1019_d N_D_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_A_841_47#_M1008_d N_D_M1008_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_B_N_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1013 N_A_211_413#_M1013_d N_A_N_M1013_g N_VPWR_M1002_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.2016 AS=0.0609 PD=1.8 PS=0.71 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90000.4 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_211_413#_M1010_g N_Y_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_A_211_413#_M1014_g N_Y_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_A_27_47#_M1007_g N_VPWR_M1014_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003 A=0.18 P=2.36 MULT=1
MM1016 N_Y_M1007_d N_A_27_47#_M1016_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.39 PD=1.29 PS=1.78 NRD=0.9653 NRS=16.7253 M=1 R=5.55556
+ SA=90001.6 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_C_M1001_g N_VPWR_M1016_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.39 PD=1.29 PS=1.78 NRD=0.9653 NRS=10.8153 M=1 R=5.55556 SA=90002.5
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1001_d N_C_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1017_s N_D_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__nand4bb_2.pxi.spice"
*
.ends
*
*
