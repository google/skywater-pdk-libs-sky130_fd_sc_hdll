* NGSPICE file created from sky130_fd_sc_hdll__nor2b_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor2b_2 A B_N VGND VNB VPB VPWR Y
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=4.034e+11p pd=3.96e+06u as=8.5e+11p ps=7.7e+06u
M1001 a_27_297# a_271_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 VPWR B_N a_271_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.806e+11p ps=1.7e+06u
M1003 Y a_271_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y A VGND VNB nshort w=650000u l=150000u
+  ad=4.485e+11p pd=3.98e+06u as=6.8595e+11p ps=7.07e+06u
M1005 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_271_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Y a_271_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND B_N a_271_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.764e+11p ps=1.68e+06u
.ends

