* File: sky130_fd_sc_hdll__dlygate4sd1_1.pxi.spice
* Created: Thu Aug 27 19:06:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A N_A_M1007_g N_A_M1005_g A A N_A_c_68_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_27_47# N_A_27_47#_M1005_s
+ N_A_27_47#_M1007_s N_A_27_47#_M1004_g N_A_27_47#_M1000_g N_A_27_47#_c_106_n
+ N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_102_n N_A_27_47#_c_107_n
+ N_A_27_47#_c_108_n N_A_27_47#_c_103_n N_A_27_47#_c_110_n N_A_27_47#_c_104_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_213_47# N_A_213_47#_M1000_d
+ N_A_213_47#_M1004_d N_A_213_47#_c_177_n N_A_213_47#_M1002_g
+ N_A_213_47#_c_170_n N_A_213_47#_M1006_g N_A_213_47#_c_171_n
+ N_A_213_47#_c_172_n N_A_213_47#_c_173_n N_A_213_47#_c_174_n
+ N_A_213_47#_c_179_n N_A_213_47#_c_175_n N_A_213_47#_c_176_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_213_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_319_93# N_A_319_93#_M1006_s
+ N_A_319_93#_M1002_s N_A_319_93#_M1003_g N_A_319_93#_M1001_g
+ N_A_319_93#_c_239_n N_A_319_93#_c_233_n N_A_319_93#_c_240_n
+ N_A_319_93#_c_241_n N_A_319_93#_c_234_n N_A_319_93#_c_243_n
+ N_A_319_93#_c_235_n N_A_319_93#_c_236_n N_A_319_93#_c_237_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_319_93#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VPWR N_VPWR_M1007_d N_VPWR_M1002_d
+ N_VPWR_c_299_n N_VPWR_c_300_n N_VPWR_c_301_n N_VPWR_c_302_n VPWR
+ N_VPWR_c_303_n N_VPWR_c_304_n N_VPWR_c_298_n N_VPWR_c_306_n VPWR
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VPWR
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%X N_X_M1001_d N_X_M1003_d N_X_c_340_n
+ N_X_c_343_n N_X_c_341_n X X X PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%X
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VGND N_VGND_M1005_d N_VGND_M1006_d
+ N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n VGND
+ N_VGND_c_364_n N_VGND_c_365_n N_VGND_c_366_n N_VGND_c_367_n VGND
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VGND
cc_1 VNB N_A_M1005_g 0.0362104f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.0125899f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_A_c_68_n 0.0340348f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_47#_M1000_g 0.031984f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_5 VNB N_A_27_47#_c_100_n 0.0186036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_101_n 0.00873805f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.53
cc_7 VNB N_A_27_47#_c_102_n 0.00988907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_103_n 0.00521395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_104_n 0.026172f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_213_47#_c_170_n 0.0375794f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.445
cc_11 VNB N_A_213_47#_c_171_n 0.0105789f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_12 VNB N_A_213_47#_c_172_n 5.78778e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_213_47#_c_173_n 0.0100937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_213_47#_c_174_n 0.00414391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_213_47#_c_175_n 0.00212837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_213_47#_c_176_n 0.0403428f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_319_93#_c_233_n 0.00556952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_319_93#_c_234_n 0.00680248f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.53
cc_19 VNB N_A_319_93#_c_235_n 0.00798679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_319_93#_c_236_n 0.030671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_319_93#_c_237_n 0.0217033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_298_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_340_n 0.00558185f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.445
cc_24 VNB N_X_c_341_n 0.0219549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.0166789f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_26 VNB N_VGND_c_360_n 0.00493236f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_27 VNB N_VGND_c_361_n 0.00609109f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_28 VNB N_VGND_c_362_n 0.0343385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_363_n 0.00785847f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.16
cc_30 VNB N_VGND_c_364_n 0.0176957f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.16
cc_31 VNB N_VGND_c_365_n 0.0203986f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_366_n 0.193902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_367_n 0.00410458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_M1007_g 0.0644496f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=2.275
cc_35 VPB A 0.0179822f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_36 VPB N_A_c_68_n 0.00852761f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_37 VPB N_A_27_47#_M1004_g 0.0564089f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_38 VPB N_A_27_47#_c_106_n 0.0188411f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.16
cc_39 VPB N_A_27_47#_c_107_n 0.00971013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_108_n 0.012476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_103_n 6.81118e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_110_n 0.00337745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_104_n 0.00638495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_213_47#_c_177_n 0.0681786f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_45 VPB N_A_213_47#_c_172_n 0.0184675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_213_47#_c_179_n 0.00432408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_213_47#_c_176_n 0.0114838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_319_93#_M1003_g 0.0266947f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_49 VPB N_A_319_93#_c_239_n 0.00872646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_319_93#_c_240_n 0.00147342f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_319_93#_c_241_n 0.0031971f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_319_93#_c_234_n 2.3885e-19 $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.53
cc_53 VPB N_A_319_93#_c_243_n 0.00295275f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_319_93#_c_236_n 0.0080755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_299_n 0.00493236f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_56 VPB N_VPWR_c_300_n 0.00586751f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_57 VPB N_VPWR_c_301_n 0.0355964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_302_n 0.00709097f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.16
cc_59 VPB N_VPWR_c_303_n 0.0176016f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_60 VPB N_VPWR_c_304_n 0.0221506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_298_n 0.0597447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_306_n 0.00406576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_X_c_343_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_341_n 0.00896625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB X 0.0322452f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_66 N_A_M1007_g N_A_27_47#_M1004_g 0.0409596f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_67 A N_A_27_47#_M1004_g 8.58794e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_A_27_47#_M1000_g 0.0209556f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_69 N_A_M1007_g N_A_27_47#_c_106_n 0.0037728f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_70 N_A_M1005_g N_A_27_47#_c_100_n 0.00709694f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1005_g N_A_27_47#_c_101_n 0.013872f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_101_n 0.017067f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_c_68_n N_A_27_47#_c_101_n 0.00168708f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_74 A N_A_27_47#_c_102_n 0.0252593f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_75 N_A_c_68_n N_A_27_47#_c_102_n 0.00511105f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_M1007_g N_A_27_47#_c_107_n 0.0178074f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_77 A N_A_27_47#_c_107_n 0.017423f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_78 A N_A_27_47#_c_108_n 0.0271506f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A_c_68_n N_A_27_47#_c_108_n 8.59854e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_M1005_g N_A_27_47#_c_103_n 0.00366897f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_81 A N_A_27_47#_c_103_n 0.0232483f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A_c_68_n N_A_27_47#_c_103_n 8.544e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_M1007_g N_A_27_47#_c_110_n 0.00439862f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_84 A N_A_27_47#_c_110_n 0.0238071f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_85 A N_A_27_47#_c_104_n 8.94748e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_68_n N_A_27_47#_c_104_n 0.0213608f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_M1007_g N_VPWR_c_299_n 0.00304969f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_88 N_A_M1007_g N_VPWR_c_303_n 0.00523784f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_89 N_A_M1007_g N_VPWR_c_298_n 0.0077765f $X=0.505 $Y=2.275 $X2=0 $Y2=0
cc_90 N_A_M1005_g N_VGND_c_360_n 0.00308651f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_M1005_g N_VGND_c_364_n 0.00436487f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_92 N_A_M1005_g N_VGND_c_366_n 0.00697623f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_27_47#_M1000_g N_A_213_47#_c_171_n 0.0108753f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_103_n N_A_213_47#_c_171_n 0.0198042f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_104_n N_A_213_47#_c_171_n 7.01138e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_M1004_g N_A_213_47#_c_172_n 0.0195497f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_107_n N_A_213_47#_c_172_n 0.0113209f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_c_103_n N_A_213_47#_c_172_n 0.00371586f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_110_n N_A_213_47#_c_172_n 0.0212546f $X=0.86 $Y=1.785 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_104_n N_A_213_47#_c_172_n 4.37316e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_M1000_g N_A_213_47#_c_174_n 0.00657279f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_103_n N_A_213_47#_c_174_n 0.00294768f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_c_104_n N_A_213_47#_c_174_n 7.21452e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_M1004_g N_A_213_47#_c_179_n 0.00862725f $X=0.975 $Y=2.275
+ $X2=0 $Y2=0
cc_105 N_A_27_47#_c_103_n N_A_213_47#_c_175_n 0.0168575f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_104_n N_A_213_47#_c_175_n 0.00194717f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_104_n N_A_213_47#_c_176_n 0.00717325f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_M1004_g N_VPWR_c_299_n 0.00389952f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_107_n N_VPWR_c_299_n 0.0151692f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1004_g N_VPWR_c_301_n 0.0052151f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_107_n N_VPWR_c_301_n 0.0021103f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_112 N_A_27_47#_c_106_n N_VPWR_c_303_n 0.0199397f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_107_n N_VPWR_c_303_n 0.0031219f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_M1007_s N_VPWR_c_298_n 0.00242594f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_115 N_A_27_47#_M1004_g N_VPWR_c_298_n 0.00905583f $X=0.975 $Y=2.275 $X2=0
+ $Y2=0
cc_116 N_A_27_47#_c_106_n N_VPWR_c_298_n 0.0112839f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_107_n N_VPWR_c_298_n 0.00921336f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_118 N_A_27_47#_M1000_g N_VGND_c_360_n 0.0037144f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_101_n N_VGND_c_360_n 0.0115001f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_103_n N_VGND_c_360_n 0.00342769f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1000_g N_VGND_c_362_n 0.0043424f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_103_n N_VGND_c_362_n 0.00217856f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_123 N_A_27_47#_c_100_n N_VGND_c_364_n 0.0198425f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_101_n N_VGND_c_364_n 0.00312415f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_125 N_A_27_47#_M1005_s N_VGND_c_366_n 0.00281655f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_M1000_g N_VGND_c_366_n 0.00829313f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_100_n N_VGND_c_366_n 0.010877f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_101_n N_VGND_c_366_n 0.00573429f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_103_n N_VGND_c_366_n 0.00370966f $X=0.86 $Y=1.325 $X2=0
+ $Y2=0
cc_130 N_A_213_47#_c_177_n N_A_319_93#_M1003_g 0.0213988f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_131 N_A_213_47#_c_177_n N_A_319_93#_c_239_n 0.00932281f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_132 N_A_213_47#_c_172_n N_A_319_93#_c_239_n 0.029451f $X=1.335 $Y=2.175 $X2=0
+ $Y2=0
cc_133 N_A_213_47#_c_179_n N_A_319_93#_c_239_n 0.0191502f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_134 N_A_213_47#_c_170_n N_A_319_93#_c_233_n 0.0126703f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_135 N_A_213_47#_c_173_n N_A_319_93#_c_233_n 0.0112247f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_213_47#_c_176_n N_A_319_93#_c_233_n 0.0019749f $X=1.99 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_213_47#_c_177_n N_A_319_93#_c_240_n 0.0203668f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_138 N_A_213_47#_c_173_n N_A_319_93#_c_240_n 0.00712088f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_139 N_A_213_47#_c_176_n N_A_319_93#_c_240_n 9.73755e-19 $X=1.99 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_213_47#_c_172_n N_A_319_93#_c_241_n 0.012958f $X=1.335 $Y=2.175 $X2=0
+ $Y2=0
cc_141 N_A_213_47#_c_173_n N_A_319_93#_c_241_n 0.0120363f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_213_47#_c_176_n N_A_319_93#_c_241_n 0.00516661f $X=1.99 $Y=1.16 $X2=0
+ $Y2=0
cc_143 N_A_213_47#_c_170_n N_A_319_93#_c_234_n 0.00644328f $X=1.99 $Y=0.995
+ $X2=0 $Y2=0
cc_144 N_A_213_47#_c_173_n N_A_319_93#_c_234_n 0.00876131f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_213_47#_c_177_n N_A_319_93#_c_243_n 0.00492289f $X=1.975 $Y=1.325
+ $X2=0 $Y2=0
cc_146 N_A_213_47#_c_170_n N_A_319_93#_c_235_n 0.0103868f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_147 N_A_213_47#_c_171_n N_A_319_93#_c_235_n 0.0257191f $X=1.335 $Y=1.075
+ $X2=0 $Y2=0
cc_148 N_A_213_47#_c_173_n N_A_319_93#_c_235_n 0.0182754f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_149 N_A_213_47#_c_174_n N_A_319_93#_c_235_n 0.021598f $X=1.335 $Y=0.4 $X2=0
+ $Y2=0
cc_150 N_A_213_47#_c_176_n N_A_319_93#_c_235_n 0.00575864f $X=1.99 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_213_47#_c_176_n N_A_319_93#_c_236_n 0.00787314f $X=1.99 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_213_47#_c_170_n N_A_319_93#_c_237_n 0.0136124f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_213_47#_c_179_n N_VPWR_c_299_n 0.0222152f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_154 N_A_213_47#_c_177_n N_VPWR_c_300_n 0.0111922f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_155 N_A_213_47#_c_177_n N_VPWR_c_301_n 0.00702461f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_156 N_A_213_47#_c_179_n N_VPWR_c_301_n 0.026749f $X=1.335 $Y=2.32 $X2=0 $Y2=0
cc_157 N_A_213_47#_M1004_d N_VPWR_c_298_n 0.00209344f $X=1.065 $Y=2.065 $X2=0
+ $Y2=0
cc_158 N_A_213_47#_c_177_n N_VPWR_c_298_n 0.0145798f $X=1.975 $Y=1.325 $X2=0
+ $Y2=0
cc_159 N_A_213_47#_c_179_n N_VPWR_c_298_n 0.0159536f $X=1.335 $Y=2.32 $X2=0
+ $Y2=0
cc_160 N_A_213_47#_c_174_n N_VGND_c_360_n 0.0222153f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_161 N_A_213_47#_c_170_n N_VGND_c_361_n 0.00773202f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_213_47#_c_170_n N_VGND_c_362_n 0.00439206f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_213_47#_c_174_n N_VGND_c_362_n 0.0267806f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_164 N_A_213_47#_M1000_d N_VGND_c_366_n 0.00209344f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_165 N_A_213_47#_c_170_n N_VGND_c_366_n 0.00811115f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_A_213_47#_c_174_n N_VGND_c_366_n 0.0159581f $X=1.335 $Y=0.4 $X2=0 $Y2=0
cc_167 N_A_319_93#_c_240_n N_VPWR_M1002_d 0.0146765f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_168 N_A_319_93#_c_243_n N_VPWR_M1002_d 0.00179207f $X=2.505 $Y=1.575 $X2=0
+ $Y2=0
cc_169 N_A_319_93#_M1003_g N_VPWR_c_300_n 0.0105925f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_170 N_A_319_93#_c_239_n N_VPWR_c_300_n 0.0216036f $X=1.727 $Y=1.745 $X2=0
+ $Y2=0
cc_171 N_A_319_93#_c_240_n N_VPWR_c_300_n 0.030862f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_172 N_A_319_93#_c_239_n N_VPWR_c_301_n 0.0130885f $X=1.727 $Y=1.745 $X2=0
+ $Y2=0
cc_173 N_A_319_93#_M1003_g N_VPWR_c_304_n 0.00702461f $X=2.7 $Y=1.985 $X2=0
+ $Y2=0
cc_174 N_A_319_93#_M1003_g N_VPWR_c_298_n 0.0142556f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_175 N_A_319_93#_c_239_n N_VPWR_c_298_n 0.00844061f $X=1.727 $Y=1.745 $X2=0
+ $Y2=0
cc_176 N_A_319_93#_M1003_g N_X_c_343_n 0.0124445f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_177 N_A_319_93#_c_240_n N_X_c_343_n 0.0101894f $X=2.4 $Y=1.66 $X2=0 $Y2=0
cc_178 N_A_319_93#_M1003_g N_X_c_341_n 0.00371386f $X=2.7 $Y=1.985 $X2=0 $Y2=0
cc_179 N_A_319_93#_c_234_n N_X_c_341_n 0.0270787f $X=2.505 $Y=1.325 $X2=0 $Y2=0
cc_180 N_A_319_93#_c_243_n N_X_c_341_n 0.00770351f $X=2.505 $Y=1.575 $X2=0 $Y2=0
cc_181 N_A_319_93#_c_236_n N_X_c_341_n 0.00845268f $X=2.645 $Y=1.16 $X2=0 $Y2=0
cc_182 N_A_319_93#_c_237_n N_X_c_341_n 0.00368071f $X=2.685 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_319_93#_c_233_n N_VGND_M1006_d 0.00407602f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_184 N_A_319_93#_c_234_n N_VGND_M1006_d 0.00354068f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_185 N_A_319_93#_c_233_n N_VGND_c_361_n 0.0198976f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_186 N_A_319_93#_c_234_n N_VGND_c_361_n 0.0133517f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_187 N_A_319_93#_c_235_n N_VGND_c_361_n 0.0163002f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_188 N_A_319_93#_c_237_n N_VGND_c_361_n 0.00723006f $X=2.685 $Y=0.995 $X2=0
+ $Y2=0
cc_189 N_A_319_93#_c_233_n N_VGND_c_362_n 0.00338992f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_190 N_A_319_93#_c_235_n N_VGND_c_362_n 0.0159334f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_191 N_A_319_93#_c_234_n N_VGND_c_365_n 8.01519e-19 $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_192 N_A_319_93#_c_237_n N_VGND_c_365_n 0.00585385f $X=2.685 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_319_93#_c_233_n N_VGND_c_366_n 0.00822214f $X=2.4 $Y=0.82 $X2=0 $Y2=0
cc_194 N_A_319_93#_c_234_n N_VGND_c_366_n 0.0022347f $X=2.505 $Y=1.325 $X2=0
+ $Y2=0
cc_195 N_A_319_93#_c_235_n N_VGND_c_366_n 0.00857794f $X=1.72 $Y=0.74 $X2=0
+ $Y2=0
cc_196 N_A_319_93#_c_237_n N_VGND_c_366_n 0.0124757f $X=2.685 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_VPWR_c_298_n N_X_M1003_d 0.00472999f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_300_n X 0.0259609f $X=2.33 $Y=2 $X2=0 $Y2=0
cc_199 N_VPWR_c_304_n X 0.0182101f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_200 N_VPWR_c_298_n X 0.00993603f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_201 X N_VGND_c_365_n 0.0189908f $X=2.885 $Y=0.425 $X2=0 $Y2=0
cc_202 N_X_M1001_d N_VGND_c_366_n 0.00283025f $X=2.81 $Y=0.235 $X2=0 $Y2=0
cc_203 X N_VGND_c_366_n 0.0110704f $X=2.885 $Y=0.425 $X2=0 $Y2=0
