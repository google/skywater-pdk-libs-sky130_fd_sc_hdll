# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.470000 1.245000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.945000 2.125000 1.520000 2.465000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 0.305000 1.315000 0.750000 ;
        RECT 1.065000 0.750000 1.625000 1.245000 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA  0.509300 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 1.485000  0.085000 1.815000 0.580000 ;
        RECT 2.695000  0.085000 2.970000 0.745000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.410000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  0.832500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.085000 2.130000 0.765000 2.635000 ;
        RECT 0.525000 1.765000 0.905000 1.955000 ;
        RECT 0.525000 1.955000 0.765000 2.130000 ;
        RECT 1.705000 1.790000 1.920000 2.635000 ;
        RECT 2.790000 1.625000 3.050000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.511000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.255000 2.430000 0.715000 ;
        RECT 2.170000 1.795000 2.620000 2.465000 ;
        RECT 2.260000 0.715000 2.430000 0.925000 ;
        RECT 2.260000 0.925000 2.925000 1.445000 ;
        RECT 2.260000 1.445000 2.620000 1.795000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.100000 1.425000 2.040000 1.595000 ;
      RECT 0.100000 1.595000 0.355000 1.960000 ;
      RECT 0.105000 0.305000 0.895000 0.570000 ;
      RECT 0.690000 0.570000 0.895000 1.425000 ;
      RECT 1.180000 1.595000 1.480000 1.890000 ;
      RECT 1.810000 0.995000 2.040000 1.425000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_2
END LIBRARY
