* File: sky130_fd_sc_hdll__dfstp_1.spice
* Created: Wed Sep  2 08:28:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dfstp_1.pex.spice"
.subckt sky130_fd_sc_hdll__dfstp_1  VNB VPB CLK D SET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SET_B	SET_B
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1020 N_VGND_M1020_d N_CLK_M1020_g N_A_27_47#_M1020_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1001 N_A_211_363#_M1001_d N_A_27_47#_M1001_g N_VGND_M1020_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_A_409_329#_M1013_d N_D_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.64
+ AD=0.11968 AS=0.1984 PD=1.2352 PS=1.9 NRD=0 NRS=8.436 M=1 R=4.26667 SA=75000.2
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1002 N_A_506_47#_M1002_d N_A_27_47#_M1002_g N_A_409_329#_M1013_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.09 AS=0.06732 PD=0.86 PS=0.6948 NRD=39.996 NRS=16.656 M=1
+ R=2.4 SA=75000.7 SB=75002.4 A=0.054 P=1.02 MULT=1
MM1016 A_636_47# N_A_211_363#_M1016_g N_A_506_47#_M1002_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0618923 AS=0.09 PD=0.692308 PS=0.86 NRD=38.964 NRS=33.324 M=1
+ R=2.4 SA=75001.4 SB=75001.7 A=0.054 P=1.02 MULT=1
MM1022 N_VGND_M1022_d N_A_702_21#_M1022_g A_636_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0722077 PD=0.94 PS=0.807692 NRD=55.704 NRS=33.396 M=1 R=2.8
+ SA=75001.6 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1021 A_866_47# N_SET_B_M1021_g N_VGND_M1022_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.1092 PD=0.63 PS=0.94 NRD=14.28 NRS=12.852 M=1 R=2.8 SA=75002.3
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1025 N_A_702_21#_M1025_d N_A_506_47#_M1025_g A_866_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0441 PD=1.46 PS=0.63 NRD=12.852 NRS=14.28 M=1 R=2.8
+ SA=75002.6 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1015 A_1156_47# N_A_506_47#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0546 AS=0.1302 PD=0.68 PS=1.46 NRD=21.42 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1011 N_A_1126_413#_M1011_d N_A_211_363#_M1011_g A_1156_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.0798 AS=0.0546 PD=0.8 PS=0.68 NRD=7.14 NRS=21.42 M=1 R=2.8
+ SA=75000.6 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1004 A_1344_47# N_A_27_47#_M1004_g N_A_1126_413#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0441 AS=0.0798 PD=0.63 PS=0.8 NRD=14.28 NRS=21.42 M=1 R=2.8
+ SA=75001.2 SB=75001.6 A=0.063 P=1.14 MULT=1
MM1029 A_1416_47# N_A_1288_261#_M1029_g A_1344_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0441 AS=0.0441 PD=0.63 PS=0.63 NRD=14.28 NRS=14.28 M=1 R=2.8 SA=75001.5
+ SB=75001.3 A=0.063 P=1.14 MULT=1
MM1031 N_VGND_M1031_d N_SET_B_M1031_g A_1416_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.120487 AS=0.0441 PD=0.97125 PS=0.63 NRD=41.424 NRS=14.28 M=1 R=2.8
+ SA=75001.9 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1023 N_A_1288_261#_M1023_d N_A_1126_413#_M1023_g N_VGND_M1031_d VNB NSHORT
+ L=0.15 W=0.54 AD=0.1404 AS=0.154912 PD=1.6 PS=1.24875 NRD=0 NRS=32.22 M=1
+ R=3.6 SA=75002.1 SB=75000.2 A=0.081 P=1.38 MULT=1
MM1005 N_VGND_M1005_d N_A_1126_413#_M1005_g N_A_1738_47#_M1005_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0901822 AS=0.1302 PD=0.808598 PS=1.46 NRD=14.28 NRS=12.852
+ M=1 R=2.8 SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1009 N_Q_M1009_d N_A_1738_47#_M1009_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.19825 AS=0.139568 PD=1.91 PS=1.2514 NRD=7.38 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VPWR_M1006_d N_CLK_M1006_g N_A_27_47#_M1006_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1027 N_A_211_363#_M1027_d N_A_27_47#_M1027_g N_VPWR_M1006_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_A_409_329#_M1014_d N_D_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=0.84
+ AD=0.175 AS=0.2268 PD=1.59333 PS=2.22 NRD=1.1623 NRS=1.1623 M=1 R=4.66667
+ SA=90000.2 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1028 N_A_506_47#_M1028_d N_A_211_363#_M1028_g N_A_409_329#_M1014_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0609 AS=0.0875 PD=0.71 PS=0.796667 NRD=2.3443 NRS=32.8202
+ M=1 R=2.33333 SA=90000.7 SB=90004.2 A=0.0756 P=1.2 MULT=1
MM1019 A_610_413# N_A_27_47#_M1019_g N_A_506_47#_M1028_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0987 AS=0.0609 PD=0.89 PS=0.71 NRD=84.4145 NRS=2.3443 M=1
+ R=2.33333 SA=90001.2 SB=90003.8 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_A_702_21#_M1008_g A_610_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.084 AS=0.0987 PD=0.82 PS=0.89 NRD=25.7873 NRS=84.4145 M=1 R=2.33333
+ SA=90001.8 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1026 N_A_702_21#_M1026_d N_SET_B_M1026_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.084 PD=0.71 PS=0.82 NRD=2.3443 NRS=30.4759 M=1 R=2.33333
+ SA=90002.4 SB=90002.5 A=0.0756 P=1.2 MULT=1
MM1017 N_VPWR_M1017_d N_A_506_47#_M1017_g N_A_702_21#_M1026_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0609 AS=0.0609 PD=0.71 PS=0.71 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90002.9 SB=90002.1 A=0.0756 P=1.2 MULT=1
MM1012 A_1044_413# N_A_506_47#_M1012_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.0609 PD=0.65 PS=0.71 NRD=28.1316 NRS=2.3443 M=1 R=2.33333
+ SA=90003.4 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1030 N_A_1126_413#_M1030_d N_A_27_47#_M1030_g A_1044_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0861 AS=0.0483 PD=0.83 PS=0.65 NRD=2.3443 NRS=28.1316 M=1
+ R=2.33333 SA=90003.8 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1024 A_1244_413# N_A_211_363#_M1024_g N_A_1126_413#_M1030_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0483 AS=0.0861 PD=0.65 PS=0.83 NRD=28.1316 NRS=58.6272 M=1
+ R=2.33333 SA=90004.4 SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1288_261#_M1010_g A_1244_413# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.0483 PD=1.38 PS=0.65 NRD=2.3443 NRS=28.1316 M=1
+ R=2.33333 SA=90004.8 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_SET_B_M1000_g N_A_1126_413#_M1000_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0861 AS=0.1134 PD=0.793333 PS=1.38 NRD=30.4759 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1018 N_A_1288_261#_M1018_d N_A_1126_413#_M1018_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.2268 AS=0.1722 PD=2.22 PS=1.58667 NRD=1.1623 NRS=1.1623 M=1
+ R=4.66667 SA=90000.4 SB=90000.2 A=0.1512 P=2.04 MULT=1
MM1007 N_VPWR_M1007_d N_A_1126_413#_M1007_g N_A_1738_47#_M1007_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=18.4589 NRS=1.5366
+ M=1 R=3.55556 SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1003 N_Q_M1003_d N_A_1738_47#_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.32 AS=0.191707 PD=2.64 PS=1.64024 NRD=10.8153 NRS=0.9653 M=1 R=5.55556
+ SA=90000.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=16.8525 P=24.21
c_207 VPB 0 9.39049e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__dfstp_1.pxi.spice"
*
.ends
*
*
