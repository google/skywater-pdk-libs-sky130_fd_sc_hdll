* File: sky130_fd_sc_hdll__a21boi_1.pxi.spice
* Created: Wed Sep  2 08:16:45 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%B1_N N_B1_N_c_51_n N_B1_N_c_52_n N_B1_N_c_55_n
+ N_B1_N_M1000_g N_B1_N_c_53_n N_B1_N_M1002_g N_B1_N_c_56_n B1_N B1_N
+ N_B1_N_c_54_n PM_SKY130_FD_SC_HDLL__A21BOI_1%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%A_27_413# N_A_27_413#_M1002_s
+ N_A_27_413#_M1000_s N_A_27_413#_c_87_n N_A_27_413#_M1005_g N_A_27_413#_c_94_n
+ N_A_27_413#_M1007_g N_A_27_413#_c_89_n N_A_27_413#_c_96_n N_A_27_413#_c_97_n
+ N_A_27_413#_c_90_n N_A_27_413#_c_91_n N_A_27_413#_c_92_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_1%A_27_413#
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%A1 N_A1_c_153_n N_A1_M1001_g N_A1_c_154_n
+ N_A1_M1003_g A1 A1 A1 PM_SKY130_FD_SC_HDLL__A21BOI_1%A1
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%A2 N_A2_c_188_n N_A2_M1004_g N_A2_c_189_n
+ N_A2_M1006_g A2 A2 PM_SKY130_FD_SC_HDLL__A21BOI_1%A2
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_c_211_n N_VPWR_c_212_n N_VPWR_c_213_n N_VPWR_c_214_n VPWR
+ N_VPWR_c_215_n N_VPWR_c_216_n N_VPWR_c_210_n N_VPWR_c_218_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%Y N_Y_M1005_d N_Y_M1007_s Y Y Y Y Y N_Y_c_254_n
+ Y PM_SKY130_FD_SC_HDLL__A21BOI_1%Y
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%A_338_297# N_A_338_297#_M1007_d
+ N_A_338_297#_M1006_d N_A_338_297#_c_297_n N_A_338_297#_c_289_n
+ N_A_338_297#_c_291_n N_A_338_297#_c_294_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_1%A_338_297#
x_PM_SKY130_FD_SC_HDLL__A21BOI_1%VGND N_VGND_M1002_d N_VGND_M1004_d
+ N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n VGND N_VGND_c_308_n
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n
+ PM_SKY130_FD_SC_HDLL__A21BOI_1%VGND
cc_1 VNB N_B1_N_c_51_n 0.0379124f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_2 VNB N_B1_N_c_52_n 0.022461f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=0.83
cc_3 VNB N_B1_N_c_53_n 0.0204458f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.755
cc_4 VNB N_B1_N_c_54_n 0.0384937f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_5 VNB N_A_27_413#_c_87_n 0.0166923f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_6 VNB N_A_27_413#_M1005_g 0.0312382f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_7 VNB N_A_27_413#_c_89_n 0.0122703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_413#_c_90_n 0.00882695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_413#_c_91_n 0.0202329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_92_n 0.0109706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_153_n 0.0301118f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_12 VNB N_A1_c_154_n 0.0183511f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=2.275
cc_13 VNB A1 0.00211609f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_14 VNB N_A2_c_188_n 0.0225716f $X=-0.19 $Y=-0.24 $X2=0.79 $Y2=0.83
cc_15 VNB N_A2_c_189_n 0.0383657f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=2.275
cc_16 VNB A2 0.0142833f $X=-0.19 $Y=-0.24 $X2=0.865 $Y2=0.445
cc_17 VNB N_VPWR_c_210_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB Y 0.00222718f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_19 VNB N_Y_c_254_n 0.0082881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_305_n 0.00503731f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=0.905
cc_21 VNB N_VGND_c_306_n 0.0125968f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.815
cc_22 VNB N_VGND_c_307_n 0.0259848f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_23 VNB N_VGND_c_308_n 0.0302587f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_24 VNB N_VGND_c_309_n 0.0403496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_310_n 0.00442399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_311_n 0.188461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_B1_N_c_55_n 0.0214862f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.99
cc_28 VPB N_B1_N_c_56_n 0.0378059f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.815
cc_29 VPB N_B1_N_c_54_n 0.0488171f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_30 VPB N_A_27_413#_c_87_n 0.0160282f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_31 VPB N_A_27_413#_c_94_n 0.0193589f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_32 VPB N_A_27_413#_c_89_n 0.0116032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_413#_c_96_n 0.0173324f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_34 VPB N_A_27_413#_c_97_n 0.0133286f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.53
cc_35 VPB N_A_27_413#_c_90_n 0.00895493f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_413#_c_92_n 0.0303588f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A1_c_153_n 0.0275249f $X=-0.19 $Y=1.305 $X2=0.79 $Y2=0.83
cc_38 VPB A1 7.37302e-19 $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_39 VPB N_A2_c_189_n 0.0396543f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.275
cc_40 VPB A2 0.00815583f $X=-0.19 $Y=1.305 $X2=0.865 $Y2=0.445
cc_41 VPB N_VPWR_c_211_n 0.00624061f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=0.905
cc_42 VPB N_VPWR_c_212_n 0.00290346f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_43 VPB N_VPWR_c_213_n 0.0314344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_214_n 0.00583344f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_45 VPB N_VPWR_c_215_n 0.0148573f $X=-0.19 $Y=1.305 $X2=0.22 $Y2=1.16
cc_46 VPB N_VPWR_c_216_n 0.0239825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_210_n 0.0552916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_218_n 0.0056382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB Y 0.0140038f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=0.905
cc_50 VPB N_Y_c_254_n 0.0022423f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 N_B1_N_c_53_n N_A_27_413#_M1005_g 0.0125472f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_52 N_B1_N_c_55_n N_A_27_413#_c_96_n 0.00267678f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_53 N_B1_N_c_56_n N_A_27_413#_c_96_n 0.00251877f $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_54 N_B1_N_c_55_n N_A_27_413#_c_97_n 0.00449216f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_55 N_B1_N_c_56_n N_A_27_413#_c_97_n 0.0267787f $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_56 B1_N N_A_27_413#_c_97_n 0.0173893f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_57 N_B1_N_c_51_n N_A_27_413#_c_90_n 0.0243714f $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_58 N_B1_N_c_53_n N_A_27_413#_c_90_n 0.00124534f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_59 N_B1_N_c_56_n N_A_27_413#_c_90_n 0.00380052f $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_60 B1_N N_A_27_413#_c_90_n 0.0511021f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_61 N_B1_N_c_54_n N_A_27_413#_c_90_n 0.0109704f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B1_N_c_52_n N_A_27_413#_c_91_n 0.00669307f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_63 N_B1_N_c_53_n N_A_27_413#_c_91_n 0.0162503f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_64 N_B1_N_c_51_n N_A_27_413#_c_92_n 0.0152341f $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_65 B1_N N_A_27_413#_c_92_n 4.05914e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B1_N_c_54_n N_A_27_413#_c_92_n 0.0195991f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B1_N_c_55_n N_VPWR_c_211_n 0.0138923f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_68 N_B1_N_c_55_n N_VPWR_c_215_n 0.00333855f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_69 N_B1_N_c_56_n N_VPWR_c_215_n 3.30564e-19 $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_70 N_B1_N_c_55_n N_VPWR_c_210_n 0.00500193f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_71 N_B1_N_c_55_n Y 0.00456544f $X=0.5 $Y=1.99 $X2=0 $Y2=0
cc_72 N_B1_N_c_56_n Y 7.55401e-19 $X=0.24 $Y=1.815 $X2=0 $Y2=0
cc_73 N_B1_N_c_51_n Y 3.12237e-19 $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_74 N_B1_N_c_53_n N_VGND_c_305_n 0.00854696f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_75 N_B1_N_c_51_n N_VGND_c_308_n 6.22378e-19 $X=0.79 $Y=0.83 $X2=0 $Y2=0
cc_76 N_B1_N_c_52_n N_VGND_c_308_n 0.00533101f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_77 N_B1_N_c_53_n N_VGND_c_308_n 0.00489117f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_78 N_B1_N_c_52_n N_VGND_c_311_n 0.00698293f $X=0.375 $Y=0.83 $X2=0 $Y2=0
cc_79 N_B1_N_c_53_n N_VGND_c_311_n 0.0100926f $X=0.865 $Y=0.755 $X2=0 $Y2=0
cc_80 N_A_27_413#_M1005_g N_A1_c_153_n 0.00420089f $X=1.405 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_27_413#_c_94_n N_A1_c_153_n 0.0194733f $X=1.6 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_27_413#_c_89_n N_A1_c_153_n 0.0124387f $X=1.405 $Y=1.297 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_27_413#_M1005_g N_A1_c_154_n 0.0125058f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_84 N_A_27_413#_M1005_g A1 4.68875e-19 $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_85 N_A_27_413#_c_94_n N_VPWR_c_211_n 0.00324316f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_27_413#_c_97_n N_VPWR_c_211_n 0.0231213f $X=0.685 $Y=1.835 $X2=0 $Y2=0
cc_87 N_A_27_413#_c_92_n N_VPWR_c_211_n 0.00116902f $X=0.795 $Y=1.285 $X2=0
+ $Y2=0
cc_88 N_A_27_413#_c_94_n N_VPWR_c_212_n 0.00125863f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_27_413#_c_94_n N_VPWR_c_213_n 0.00681403f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_413#_c_96_n N_VPWR_c_215_n 0.014738f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_91 N_A_27_413#_c_97_n N_VPWR_c_215_n 0.00245093f $X=0.685 $Y=1.835 $X2=0
+ $Y2=0
cc_92 N_A_27_413#_M1000_s N_VPWR_c_210_n 0.00250649f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_93 N_A_27_413#_c_94_n N_VPWR_c_210_n 0.0135481f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_27_413#_c_96_n N_VPWR_c_210_n 0.00966027f $X=0.26 $Y=2.27 $X2=0 $Y2=0
cc_95 N_A_27_413#_c_97_n N_VPWR_c_210_n 0.00529104f $X=0.685 $Y=1.835 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_87_n Y 0.00882756f $X=1.33 $Y=1.285 $X2=0 $Y2=0
cc_97 N_A_27_413#_c_94_n Y 0.0349271f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_27_413#_c_89_n Y 0.0074768f $X=1.405 $Y=1.297 $X2=0 $Y2=0
cc_99 N_A_27_413#_c_97_n Y 0.0131166f $X=0.685 $Y=1.835 $X2=0 $Y2=0
cc_100 N_A_27_413#_c_90_n Y 0.0348863f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_101 N_A_27_413#_c_92_n Y 0.00257784f $X=0.795 $Y=1.285 $X2=0 $Y2=0
cc_102 N_A_27_413#_M1005_g Y 0.0171385f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_27_413#_c_89_n Y 0.00118864f $X=1.405 $Y=1.297 $X2=0 $Y2=0
cc_104 N_A_27_413#_c_90_n Y 0.00546706f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_105 N_A_27_413#_c_87_n N_Y_c_254_n 0.0118189f $X=1.33 $Y=1.285 $X2=0 $Y2=0
cc_106 N_A_27_413#_M1005_g N_Y_c_254_n 0.0118905f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_107 N_A_27_413#_c_89_n N_Y_c_254_n 0.0188273f $X=1.405 $Y=1.297 $X2=0 $Y2=0
cc_108 N_A_27_413#_c_90_n N_Y_c_254_n 0.0214345f $X=0.77 $Y=1.44 $X2=0 $Y2=0
cc_109 N_A_27_413#_c_87_n N_VGND_c_305_n 0.00248136f $X=1.33 $Y=1.285 $X2=0
+ $Y2=0
cc_110 N_A_27_413#_M1005_g N_VGND_c_305_n 0.005221f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_111 N_A_27_413#_c_91_n N_VGND_c_305_n 0.0463141f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_112 N_A_27_413#_c_91_n N_VGND_c_308_n 0.0300406f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_113 N_A_27_413#_M1005_g N_VGND_c_309_n 0.00526721f $X=1.405 $Y=0.56 $X2=0
+ $Y2=0
cc_114 N_A_27_413#_M1002_s N_VGND_c_311_n 0.00296656f $X=0.425 $Y=0.235 $X2=0
+ $Y2=0
cc_115 N_A_27_413#_M1005_g N_VGND_c_311_n 0.010104f $X=1.405 $Y=0.56 $X2=0 $Y2=0
cc_116 N_A_27_413#_c_91_n N_VGND_c_311_n 0.0183483f $X=0.55 $Y=0.45 $X2=0 $Y2=0
cc_117 N_A1_c_154_n N_A2_c_188_n 0.0238718f $X=2.095 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_118 A1 N_A2_c_188_n 0.00689065f $X=2.025 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_119 N_A1_c_153_n N_A2_c_189_n 0.0372727f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_120 A1 N_A2_c_189_n 0.00164319f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_121 N_A1_c_153_n A2 0.00122266f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_122 A1 A2 0.0130641f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_123 N_A1_c_153_n N_VPWR_c_212_n 0.0153018f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_153_n N_VPWR_c_213_n 0.00447018f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_153_n N_VPWR_c_210_n 0.00768581f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A1_c_153_n Y 0.00118657f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A1_c_153_n Y 4.73303e-19 $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A1_c_154_n Y 0.00510974f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_129 A1 Y 0.0291297f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_130 N_A1_c_153_n N_Y_c_254_n 0.00254172f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_131 A1 N_Y_c_254_n 0.0215548f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_132 N_A1_c_153_n N_A_338_297#_c_289_n 0.0174281f $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_133 A1 N_A_338_297#_c_289_n 0.0168779f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_134 N_A1_c_153_n N_A_338_297#_c_291_n 5.98561e-19 $X=2.08 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_154_n N_VGND_c_307_n 0.00189125f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_136 A1 N_VGND_c_307_n 0.0151956f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_137 N_A1_c_154_n N_VGND_c_309_n 0.00381508f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_138 A1 N_VGND_c_309_n 0.008037f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_139 N_A1_c_154_n N_VGND_c_311_n 0.00627634f $X=2.095 $Y=0.995 $X2=0 $Y2=0
cc_140 A1 N_VGND_c_311_n 0.00838783f $X=2.025 $Y=0.425 $X2=0 $Y2=0
cc_141 A1 A_434_47# 0.00732205f $X=2.025 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_142 N_A2_c_189_n N_VPWR_c_212_n 0.00984323f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A2_c_189_n N_VPWR_c_216_n 0.00702461f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_189_n N_VPWR_c_210_n 0.0139495f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_189_n N_A_338_297#_c_289_n 0.0243113f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_146 A2 N_A_338_297#_c_289_n 0.0253498f $X=2.865 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A2_c_189_n N_A_338_297#_c_294_n 0.00691099f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A2_c_188_n N_VGND_c_307_n 0.0157822f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_189_n N_VGND_c_307_n 0.00717335f $X=2.68 $Y=1.41 $X2=0 $Y2=0
cc_150 A2 N_VGND_c_307_n 0.0260817f $X=2.865 $Y=1.105 $X2=0 $Y2=0
cc_151 N_A2_c_188_n N_VGND_c_309_n 0.00525069f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_188_n N_VGND_c_311_n 0.00923482f $X=2.655 $Y=0.995 $X2=0 $Y2=0
cc_153 N_VPWR_c_210_n N_Y_M1007_s 0.00263814f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_154 N_VPWR_c_211_n Y 0.0241189f $X=0.74 $Y=2.34 $X2=0 $Y2=0
cc_155 N_VPWR_c_213_n Y 0.0285397f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_210_n Y 0.0174906f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_210_n N_A_338_297#_M1007_d 0.00621398f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_158 N_VPWR_c_210_n N_A_338_297#_M1006_d 0.00589812f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_213_n N_A_338_297#_c_297_n 0.0123577f $X=2.105 $Y=2.72 $X2=0
+ $Y2=0
cc_160 N_VPWR_c_210_n N_A_338_297#_c_297_n 0.0071952f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_161 N_VPWR_M1001_d N_A_338_297#_c_289_n 0.0169214f $X=2.17 $Y=1.485 $X2=0
+ $Y2=0
cc_162 N_VPWR_c_212_n N_A_338_297#_c_289_n 0.0249236f $X=2.32 $Y=2.02 $X2=0
+ $Y2=0
cc_163 N_VPWR_c_212_n N_A_338_297#_c_294_n 0.0249674f $X=2.32 $Y=2.02 $X2=0
+ $Y2=0
cc_164 N_VPWR_c_216_n N_A_338_297#_c_294_n 0.0111013f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_165 N_VPWR_c_210_n N_A_338_297#_c_294_n 0.00643939f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_166 N_Y_c_254_n N_A_338_297#_c_291_n 0.00280418f $X=1.61 $Y=1.045 $X2=0 $Y2=0
cc_167 Y N_VGND_c_305_n 0.042544f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_168 N_Y_c_254_n N_VGND_c_305_n 0.0156069f $X=1.61 $Y=1.045 $X2=0 $Y2=0
cc_169 Y N_VGND_c_309_n 0.0203957f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_170 N_Y_M1005_d N_VGND_c_311_n 0.0115745f $X=1.48 $Y=0.235 $X2=0 $Y2=0
cc_171 Y N_VGND_c_311_n 0.0127759f $X=1.53 $Y=0.425 $X2=0 $Y2=0
cc_172 N_VGND_c_311_n A_434_47# 0.0151758f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
