* File: sky130_fd_sc_hdll__or2b_1.pxi.spice
* Created: Thu Aug 27 19:23:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2B_1%B_N N_B_N_c_58_n N_B_N_M1002_g N_B_N_M1000_g B_N
+ N_B_N_c_57_n B_N PM_SKY130_FD_SC_HDLL__OR2B_1%B_N
x_PM_SKY130_FD_SC_HDLL__OR2B_1%A_27_53# N_A_27_53#_M1000_s N_A_27_53#_M1002_d
+ N_A_27_53#_M1006_g N_A_27_53#_c_84_n N_A_27_53#_M1003_g N_A_27_53#_c_85_n
+ N_A_27_53#_c_86_n N_A_27_53#_c_87_n N_A_27_53#_c_91_n N_A_27_53#_c_88_n
+ N_A_27_53#_c_89_n PM_SKY130_FD_SC_HDLL__OR2B_1%A_27_53#
x_PM_SKY130_FD_SC_HDLL__OR2B_1%A N_A_c_135_n N_A_c_133_n N_A_M1005_g N_A_M1004_g
+ N_A_c_138_n A N_A_c_140_n A PM_SKY130_FD_SC_HDLL__OR2B_1%A
x_PM_SKY130_FD_SC_HDLL__OR2B_1%A_229_297# N_A_229_297#_M1006_d
+ N_A_229_297#_M1003_s N_A_229_297#_c_180_n N_A_229_297#_M1007_g
+ N_A_229_297#_c_181_n N_A_229_297#_M1001_g N_A_229_297#_c_191_n
+ N_A_229_297#_c_229_p N_A_229_297#_c_182_n N_A_229_297#_c_183_n
+ N_A_229_297#_c_187_n N_A_229_297#_c_188_n N_A_229_297#_c_184_n
+ N_A_229_297#_c_185_n PM_SKY130_FD_SC_HDLL__OR2B_1%A_229_297#
x_PM_SKY130_FD_SC_HDLL__OR2B_1%VPWR N_VPWR_M1002_s N_VPWR_M1005_d N_VPWR_c_240_n
+ N_VPWR_c_241_n N_VPWR_c_242_n VPWR N_VPWR_c_243_n N_VPWR_c_244_n
+ N_VPWR_c_239_n N_VPWR_c_246_n PM_SKY130_FD_SC_HDLL__OR2B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2B_1%X N_X_M1001_d N_X_M1007_d N_X_c_272_n N_X_c_274_n
+ N_X_c_273_n X N_X_c_276_n PM_SKY130_FD_SC_HDLL__OR2B_1%X
x_PM_SKY130_FD_SC_HDLL__OR2B_1%VGND N_VGND_M1000_d N_VGND_M1004_d VGND
+ N_VGND_c_290_n N_VGND_c_291_n N_VGND_c_292_n N_VGND_c_293_n N_VGND_c_294_n
+ N_VGND_c_295_n PM_SKY130_FD_SC_HDLL__OR2B_1%VGND
cc_1 VNB N_B_N_M1000_g 0.0401282f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB B_N 0.0092769f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_B_N_c_57_n 0.0431049f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_27_53#_M1006_g 0.0342798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_53#_c_84_n 0.0385104f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_6 VNB N_A_27_53#_c_85_n 0.0205152f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_A_27_53#_c_86_n 0.00342105f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_8 VNB N_A_27_53#_c_87_n 0.00940306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_88_n 0.00460073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_53#_c_89_n 0.0132332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_133_n 0.0106012f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_12 VNB N_A_M1004_g 0.0347972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_229_297#_c_180_n 0.0265082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_229_297#_c_181_n 0.0209378f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_15 VNB N_A_229_297#_c_182_n 0.00237161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_229_297#_c_183_n 0.00445587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_229_297#_c_184_n 0.00390081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_229_297#_c_185_n 0.00183865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_239_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_272_n 0.0193786f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_21 VNB N_X_c_273_n 0.0307968f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_22 VNB N_VGND_c_290_n 0.0147625f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_23 VNB N_VGND_c_291_n 0.0259761f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_24 VNB N_VGND_c_292_n 0.193254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_293_n 0.018858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_294_n 0.0227524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_295_n 0.0102714f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_B_N_c_58_n 0.0238148f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_29 VPB B_N 8.85293e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_30 VPB N_B_N_c_57_n 0.0190244f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_31 VPB N_A_27_53#_c_84_n 0.0334901f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_32 VPB N_A_27_53#_c_91_n 0.00464761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_53#_c_88_n 0.00639441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_53#_c_89_n 0.00350361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_c_135_n 0.0365664f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_A_c_133_n 0.006635f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_37 VPB N_A_M1005_g 0.0117887f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_38 VPB N_A_c_138_n 0.0290475f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_39 VPB A 0.0284548f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_40 VPB N_A_c_140_n 0.0372853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_229_297#_c_180_n 0.0326577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_229_297#_c_187_n 0.00156472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_229_297#_c_188_n 0.008297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_229_297#_c_184_n 2.03541e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_240_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_241_n 0.0554415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_242_n 0.0121493f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_48 VPB N_VPWR_c_243_n 0.0436263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_244_n 0.0254436f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_239_n 0.0677334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_246_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_274_n 0.0118171f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_53 VPB N_X_c_273_n 0.0111555f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_54 VPB N_X_c_276_n 0.0374223f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.2
cc_55 N_B_N_c_57_n N_A_27_53#_c_84_n 0.00528959f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_56 N_B_N_M1000_g N_A_27_53#_c_85_n 0.00300084f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_57 N_B_N_M1000_g N_A_27_53#_c_86_n 0.0187886f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_58 B_N N_A_27_53#_c_86_n 3.30304e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_59 N_B_N_c_57_n N_A_27_53#_c_86_n 0.00104773f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_60 B_N N_A_27_53#_c_87_n 0.0255233f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_61 N_B_N_c_57_n N_A_27_53#_c_87_n 0.00800665f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_62 N_B_N_c_58_n N_A_27_53#_c_91_n 0.00630275f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B_N_c_57_n N_A_27_53#_c_91_n 0.00650453f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_64 N_B_N_M1000_g N_A_27_53#_c_89_n 0.00807875f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_65 B_N N_A_27_53#_c_89_n 0.0159063f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_66 N_B_N_c_58_n A 0.00227571f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_B_N_c_57_n A 2.63734e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_68 N_B_N_c_58_n N_A_229_297#_c_188_n 0.00166948f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B_N_c_58_n N_VPWR_c_241_n 0.00874982f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 B_N N_VPWR_c_241_n 0.0206483f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_B_N_c_57_n N_VPWR_c_241_n 0.00545118f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_72 N_B_N_c_58_n N_VPWR_c_243_n 0.00298464f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_B_N_c_58_n N_VPWR_c_239_n 0.0037574f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B_N_M1000_g N_VGND_c_292_n 0.00754515f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_75 N_B_N_M1000_g N_VGND_c_293_n 0.00413798f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_76 N_B_N_M1000_g N_VGND_c_294_n 0.00505351f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_77 N_A_27_53#_c_84_n N_A_c_135_n 0.010421f $X=1.505 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_27_53#_c_84_n N_A_c_133_n 0.0183953f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_27_53#_c_88_n N_A_c_133_n 8.05573e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_27_53#_c_84_n N_A_M1005_g 0.0358735f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_53#_M1006_g N_A_M1004_g 0.0181421f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_82 N_A_27_53#_c_84_n N_A_M1004_g 0.00719371f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_27_53#_c_88_n N_A_M1004_g 5.70471e-19 $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_53#_c_84_n A 0.00205903f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_27_53#_c_91_n A 0.0124285f $X=0.73 $Y=1.62 $X2=0 $Y2=0
cc_86 N_A_27_53#_c_84_n N_A_229_297#_c_191_n 0.0126327f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_87 N_A_27_53#_M1006_g N_A_229_297#_c_183_n 0.00459933f $X=1.47 $Y=0.475 $X2=0
+ $Y2=0
cc_88 N_A_27_53#_c_84_n N_A_229_297#_c_183_n 3.06238e-19 $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_89 N_A_27_53#_c_84_n N_A_229_297#_c_188_n 0.0155597f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_90 N_A_27_53#_c_91_n N_A_229_297#_c_188_n 0.0253576f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_91 N_A_27_53#_c_88_n N_A_229_297#_c_188_n 0.0267679f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_27_53#_c_91_n N_VPWR_c_241_n 0.0192276f $X=0.73 $Y=1.62 $X2=0 $Y2=0
cc_93 N_A_27_53#_M1006_g N_VGND_c_290_n 0.00555245f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_94 N_A_27_53#_M1006_g N_VGND_c_292_n 0.0114814f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_85_n N_VGND_c_292_n 0.0117861f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_27_53#_c_86_n N_VGND_c_292_n 0.0050353f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_97 N_A_27_53#_c_89_n N_VGND_c_292_n 0.00105248f $X=0.77 $Y=0.82 $X2=0 $Y2=0
cc_98 N_A_27_53#_c_85_n N_VGND_c_293_n 0.0192939f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_99 N_A_27_53#_c_86_n N_VGND_c_293_n 0.00299761f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_27_53#_M1006_g N_VGND_c_294_n 0.00352149f $X=1.47 $Y=0.475 $X2=0
+ $Y2=0
cc_101 N_A_27_53#_c_84_n N_VGND_c_294_n 0.004553f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_27_53#_c_88_n N_VGND_c_294_n 0.0194332f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_103 N_A_27_53#_c_89_n N_VGND_c_294_n 0.0214575f $X=0.77 $Y=0.82 $X2=0 $Y2=0
cc_104 N_A_27_53#_M1006_g N_VGND_c_295_n 5.8523e-19 $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_105 N_A_c_133_n N_A_229_297#_c_180_n 0.00272261f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_A_229_297#_c_180_n 0.016126f $X=1.915 $Y=1.695 $X2=0 $Y2=0
cc_107 N_A_M1004_g N_A_229_297#_c_180_n 0.0198015f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_108 N_A_M1004_g N_A_229_297#_c_181_n 0.0175751f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_109 N_A_c_135_n N_A_229_297#_c_191_n 7.85782e-19 $X=1.815 $Y=2.34 $X2=0 $Y2=0
cc_110 N_A_M1005_g N_A_229_297#_c_191_n 0.0195895f $X=1.915 $Y=1.695 $X2=0 $Y2=0
cc_111 A N_A_229_297#_c_191_n 0.0127859f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_112 N_A_c_133_n N_A_229_297#_c_182_n 0.00127717f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_M1004_g N_A_229_297#_c_182_n 0.0133141f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_114 N_A_M1005_g N_A_229_297#_c_187_n 0.00173315f $X=1.915 $Y=1.695 $X2=0
+ $Y2=0
cc_115 N_A_c_135_n N_A_229_297#_c_188_n 9.83498e-19 $X=1.815 $Y=2.34 $X2=0 $Y2=0
cc_116 N_A_M1005_g N_A_229_297#_c_188_n 0.00115522f $X=1.915 $Y=1.695 $X2=0
+ $Y2=0
cc_117 A N_A_229_297#_c_188_n 0.0344364f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_118 N_A_c_140_n N_A_229_297#_c_188_n 0.00119166f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_119 N_A_c_133_n N_A_229_297#_c_184_n 0.0060279f $X=1.915 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_M1004_g N_A_229_297#_c_185_n 0.0060279f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_121 A N_VPWR_c_241_n 0.0258572f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_122 N_A_c_140_n N_VPWR_c_241_n 9.23051e-19 $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_123 N_A_M1005_g N_VPWR_c_242_n 0.00443253f $X=1.915 $Y=1.695 $X2=0 $Y2=0
cc_124 N_A_c_138_n N_VPWR_c_242_n 0.00487993f $X=1.915 $Y=2.34 $X2=0 $Y2=0
cc_125 A N_VPWR_c_242_n 0.0216404f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_126 A N_VPWR_c_243_n 0.0637422f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_127 N_A_c_140_n N_VPWR_c_243_n 0.0240252f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_128 A N_VPWR_c_239_n 0.0469078f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_129 N_A_c_140_n N_VPWR_c_239_n 0.0331114f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_130 N_A_M1004_g N_VGND_c_290_n 0.00188229f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_131 N_A_M1004_g N_VGND_c_292_n 0.00261357f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_132 N_A_M1004_g N_VGND_c_295_n 0.0100787f $X=1.94 $Y=0.475 $X2=0 $Y2=0
cc_133 N_A_229_297#_c_191_n N_VPWR_M1005_d 0.00563715f $X=2.215 $Y=1.58 $X2=0
+ $Y2=0
cc_134 N_A_229_297#_c_180_n N_VPWR_c_242_n 0.00522717f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_229_297#_c_191_n N_VPWR_c_242_n 0.0204259f $X=2.215 $Y=1.58 $X2=0
+ $Y2=0
cc_136 N_A_229_297#_c_188_n N_VPWR_c_242_n 0.00230358f $X=1.25 $Y=1.58 $X2=0
+ $Y2=0
cc_137 N_A_229_297#_c_180_n N_VPWR_c_244_n 0.00702461f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_229_297#_c_180_n N_VPWR_c_239_n 0.0148945f $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_229_297#_c_191_n A_319_297# 0.003951f $X=2.215 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_229_297#_c_180_n N_X_c_274_n 0.0129488f $X=2.455 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_229_297#_c_191_n N_X_c_274_n 0.0118073f $X=2.215 $Y=1.58 $X2=0 $Y2=0
cc_142 N_A_229_297#_c_180_n N_X_c_273_n 0.00189669f $X=2.455 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_229_297#_c_181_n N_X_c_273_n 0.0148863f $X=2.48 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_229_297#_c_187_n N_X_c_273_n 0.00803295f $X=2.3 $Y=1.495 $X2=0 $Y2=0
cc_145 N_A_229_297#_c_184_n N_X_c_273_n 0.018793f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_229_297#_c_185_n N_X_c_273_n 0.00717901f $X=2.33 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_229_297#_c_182_n N_VGND_M1004_d 0.00670822f $X=2.215 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_229_297#_c_185_n N_VGND_M1004_d 6.98847e-19 $X=2.33 $Y=0.995 $X2=0
+ $Y2=0
cc_149 N_A_229_297#_c_229_p N_VGND_c_290_n 0.00861358f $X=1.68 $Y=0.47 $X2=0
+ $Y2=0
cc_150 N_A_229_297#_c_182_n N_VGND_c_290_n 0.00232988f $X=2.215 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_229_297#_c_181_n N_VGND_c_291_n 0.00585385f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_229_297#_c_181_n N_VGND_c_292_n 0.012382f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_229_297#_c_229_p N_VGND_c_292_n 0.00625722f $X=1.68 $Y=0.47 $X2=0
+ $Y2=0
cc_154 N_A_229_297#_c_182_n N_VGND_c_292_n 0.00689417f $X=2.215 $Y=0.74 $X2=0
+ $Y2=0
cc_155 N_A_229_297#_c_180_n N_VGND_c_295_n 5.00515e-19 $X=2.455 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_229_297#_c_181_n N_VGND_c_295_n 0.00498808f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_157 N_A_229_297#_c_229_p N_VGND_c_295_n 0.0135697f $X=1.68 $Y=0.47 $X2=0
+ $Y2=0
cc_158 N_A_229_297#_c_182_n N_VGND_c_295_n 0.0278587f $X=2.215 $Y=0.74 $X2=0
+ $Y2=0
cc_159 N_VPWR_c_239_n N_X_M1007_d 0.00438284f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_244_n N_X_c_276_n 0.0343278f $X=2.345 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_239_n N_X_c_276_n 0.0186012f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_162 N_X_c_272_n N_VGND_c_291_n 0.0166207f $X=2.69 $Y=0.59 $X2=0 $Y2=0
cc_163 N_X_M1001_d N_VGND_c_292_n 0.00414673f $X=2.555 $Y=0.235 $X2=0 $Y2=0
cc_164 N_X_c_272_n N_VGND_c_292_n 0.0168832f $X=2.69 $Y=0.59 $X2=0 $Y2=0
