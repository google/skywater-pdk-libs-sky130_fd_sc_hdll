* File: sky130_fd_sc_hdll__a32oi_2.spice
* Created: Wed Sep  2 08:21:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32oi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a32oi_2  VNB VPB B2 B1 A1 A2 A3 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1002 N_A_27_47#_M1002_d N_B2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1014 N_A_27_47#_M1014_d N_B2_M1014_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_27_47#_M1014_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1015 N_Y_M1004_d N_B1_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_507_47#_M1011_d N_A1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1012 N_A_507_47#_M1012_d N_A1_M1012_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.08775 PD=0.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.6
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1008 N_A_507_47#_M1012_d N_A2_M1008_g N_A_757_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1016 N_A_507_47#_M1016_d N_A2_M1016_g N_A_757_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A3_M1006_g N_A_757_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26975 AS=0.1365 PD=2.13 PS=1.07 NRD=27.684 NRS=3.684 M=1 R=4.33333
+ SA=75000.3 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A3_M1019_g N_A_757_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.1365 PD=1.82 PS=1.07 NRD=0 NRS=22.152 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_297#_M1001_d N_B2_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90005.6 A=0.18 P=2.36 MULT=1
MM1007 N_A_27_297#_M1007_d N_B2_M1007_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90005.2 A=0.18 P=2.36 MULT=1
MM1013 N_A_27_297#_M1007_d N_B1_M1013_g N_Y_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90004.7 A=0.18 P=2.36 MULT=1
MM1018 N_A_27_297#_M1018_d N_B1_M1018_g N_Y_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1018_d N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.355 PD=1.29 PS=1.71 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90002.1 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_27_297#_M1010_d N_A1_M1010_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.355 PD=1.29 PS=1.71 NRD=0.9653 NRS=9.8303 M=1 R=5.55556
+ SA=90002.9 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_27_297#_M1010_d VPB PHIGHVT L=0.18 W=1
+ AD=0.315 AS=0.145 PD=1.63 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.4 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1000_d N_A2_M1017_g N_A_27_297#_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.315 AS=0.15 PD=1.63 PS=1.3 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1005 N_A_27_297#_M1017_s N_A3_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.37 PD=1.3 PS=1.74 NRD=2.9353 NRS=6.8753 M=1 R=5.55556 SA=90004.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_A_27_297#_M1009_d N_A3_M1009_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.37 PD=2.54 PS=1.74 NRD=0.9653 NRS=6.8753 M=1 R=5.55556 SA=90005.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9541 P=16.86
c_72 VPB 0 4.0732e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__a32oi_2.pxi.spice"
*
.ends
*
*
