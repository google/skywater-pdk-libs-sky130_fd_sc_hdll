* File: sky130_fd_sc_hdll__nand3_1.pex.spice
* Created: Wed Sep  2 08:37:33 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%C 1 3 4 6 7 8 14
r29 14 15 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 12 14 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r32 7 8 16.239 $w=2.18e-07 $l=3.1e-07 $layer=LI1_cond $X=0.22 $Y=0.85 $X2=0.22
+ $Y2=1.16
r33 4 15 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r35 1 14 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%B 1 3 4 6 7 8
r33 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r34 8 13 0.934413 $w=3.68e-07 $l=3e-08 $layer=LI1_cond $X=1.1 $Y=1.19 $X2=1.1
+ $Y2=1.16
r35 7 13 9.6556 $w=3.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.1 $Y=0.85 $X2=1.1
+ $Y2=1.16
r36 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1.025 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r38 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1.025 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%A 1 3 4 6 7 13
r26 7 13 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=1.625 $Y=1.16
+ $X2=1.615 $Y2=1.16
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.705
+ $Y=1.16 $X2=1.705 $Y2=1.16
r28 4 10 44.9511 $w=3.94e-07 $l=3.04959e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.617 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
r30 1 10 39.4698 $w=3.94e-07 $l=2.26892e-07 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.617 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%VPWR 1 2 7 9 13 17 19 23 24 30
r31 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r32 24 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r33 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 21 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.23 $Y2=2.72
r35 21 23 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=2.07 $Y2=2.72
r36 19 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 19 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r38 15 30 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r39 15 17 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2
r40 14 27 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r41 13 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.23 $Y2=2.72
r42 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r43 9 12 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r44 7 27 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r45 7 12 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r46 2 17 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r47 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r48 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%Y 1 2 3 12 14 16 18 20 22 24 27 31
r60 31 35 2.88588 $w=3.4e-07 $l=1.15e-07 $layer=LI1_cond $X=0.63 $Y=0.425
+ $X2=0.745 $Y2=0.425
r61 31 35 0.237268 $w=3.38e-07 $l=7e-09 $layer=LI1_cond $X=0.752 $Y=0.425
+ $X2=0.745 $Y2=0.425
r62 27 31 25.8622 $w=3.38e-07 $l=7.63e-07 $layer=LI1_cond $X=1.515 $Y=0.425
+ $X2=0.752 $Y2=0.425
r63 26 27 1.386 $w=3.4e-07 $l=1.9e-07 $layer=LI1_cond $X=1.705 $Y=0.425
+ $X2=1.515 $Y2=0.425
r64 24 26 1.36474 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=1.705 $Y=0.38
+ $X2=1.705 $Y2=0.425
r65 20 31 28.1625 $w=3.83e-07 $l=9e-07 $layer=LI1_cond $X=0.63 $Y=1.495 $X2=0.63
+ $Y2=0.595
r66 20 22 3.10218 $w=3.05e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.63 $Y=1.495
+ $X2=0.705 $Y2=1.58
r67 16 30 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=1.58
r68 16 18 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.705 $Y=1.665
+ $X2=1.705 $Y2=2.34
r69 15 22 3.51065 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r70 14 30 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.515 $Y=1.58
+ $X2=1.705 $Y2=1.58
r71 14 15 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.515 $Y=1.58
+ $X2=0.895 $Y2=1.58
r72 10 22 3.10218 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.58
r73 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r74 3 30 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.485 $X2=1.73 $Y2=1.66
r75 3 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.585
+ $Y=1.485 $X2=1.73 $Y2=2.34
r76 2 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r77 2 12 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r78 1 24 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.545
+ $Y=0.235 $X2=1.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3_1%VGND 1 4 6 8 15 16
r25 15 16 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r26 13 16 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r27 12 15 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r28 12 13 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r29 10 19 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r30 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r31 8 13 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r32 8 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r33 4 19 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r34 4 6 14.688 $w=2.53e-07 $l=3.25e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.41
r35 1 6 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.41
.ends

