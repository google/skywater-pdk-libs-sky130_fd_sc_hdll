* File: sky130_fd_sc_hdll__or3_4.pxi.spice
* Created: Thu Aug 27 19:24:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3_4%C N_C_c_80_n N_C_M1005_g N_C_c_77_n N_C_M1010_g C
+ N_C_c_79_n PM_SKY130_FD_SC_HDLL__OR3_4%C
x_PM_SKY130_FD_SC_HDLL__OR3_4%B N_B_c_105_n N_B_M1000_g N_B_c_106_n N_B_M1001_g
+ N_B_c_107_n N_B_c_108_n B B PM_SKY130_FD_SC_HDLL__OR3_4%B
x_PM_SKY130_FD_SC_HDLL__OR3_4%A N_A_c_143_n N_A_M1003_g N_A_c_144_n N_A_M1012_g
+ A A PM_SKY130_FD_SC_HDLL__OR3_4%A
x_PM_SKY130_FD_SC_HDLL__OR3_4%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1001_d
+ N_A_27_47#_M1005_s N_A_27_47#_c_193_n N_A_27_47#_M1002_g N_A_27_47#_c_179_n
+ N_A_27_47#_M1006_g N_A_27_47#_c_194_n N_A_27_47#_M1004_g N_A_27_47#_c_180_n
+ N_A_27_47#_M1007_g N_A_27_47#_c_195_n N_A_27_47#_M1009_g N_A_27_47#_c_181_n
+ N_A_27_47#_M1008_g N_A_27_47#_c_196_n N_A_27_47#_M1013_g N_A_27_47#_c_182_n
+ N_A_27_47#_M1011_g N_A_27_47#_c_183_n N_A_27_47#_c_197_n N_A_27_47#_c_198_n
+ N_A_27_47#_c_184_n N_A_27_47#_c_185_n N_A_27_47#_c_209_n N_A_27_47#_c_210_n
+ N_A_27_47#_c_226_n N_A_27_47#_c_186_n N_A_27_47#_c_230_n N_A_27_47#_c_219_n
+ N_A_27_47#_c_187_n N_A_27_47#_c_188_n N_A_27_47#_c_189_n N_A_27_47#_c_190_n
+ N_A_27_47#_c_191_n N_A_27_47#_c_192_n PM_SKY130_FD_SC_HDLL__OR3_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__OR3_4%VPWR N_VPWR_M1012_d N_VPWR_M1004_d N_VPWR_M1013_d
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n VPWR N_VPWR_c_352_n N_VPWR_c_353_n
+ N_VPWR_c_344_n N_VPWR_c_355_n PM_SKY130_FD_SC_HDLL__OR3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3_4%X N_X_M1006_s N_X_M1008_s N_X_M1002_s N_X_M1009_s
+ N_X_c_410_n N_X_c_446_n N_X_c_405_n N_X_c_406_n N_X_c_399_n N_X_c_400_n
+ N_X_c_428_n N_X_c_450_n N_X_c_407_n N_X_c_401_n N_X_c_402_n N_X_c_408_n X
+ N_X_c_404_n PM_SKY130_FD_SC_HDLL__OR3_4%X
x_PM_SKY130_FD_SC_HDLL__OR3_4%VGND N_VGND_M1010_d N_VGND_M1003_d N_VGND_M1007_d
+ N_VGND_M1011_d N_VGND_c_475_n N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n
+ N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n VGND N_VGND_c_482_n
+ N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n VGND
+ PM_SKY130_FD_SC_HDLL__OR3_4%VGND
cc_1 VNB N_C_c_77_n 0.022163f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB C 0.00894111f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C_c_79_n 0.0375026f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_c_105_n 0.0219213f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_c_106_n 0.0166804f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B_c_107_n 0.00213548f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_B_c_108_n 0.00168216f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_8 VNB N_A_c_143_n 0.0200373f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_A_c_144_n 0.0250547f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB A 0.00454573f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_179_n 0.0196226f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_12 VNB N_A_27_47#_c_180_n 0.016746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_181_n 0.0167612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_182_n 0.0197218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_183_n 0.0187495f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_184_n 0.0027452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_185_n 0.00984759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_186_n 0.00529957f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_187_n 0.00298992f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_188_n 3.90207e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_189_n 0.0015776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_190_n 0.00311049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_191_n 0.00113699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_192_n 0.0978134f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VPWR_c_344_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_399_n 0.00264486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_400_n 0.0023255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_401_n 0.00241217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_402_n 0.0023255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.0232136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_404_n 0.0111589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_475_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_476_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_477_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_478_n 0.0201421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_479_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_480_n 0.0195143f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_481_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_482_n 0.0149319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_483_n 0.242064f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_484_n 0.0219024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_485_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_486_n 0.0211525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VPB N_C_c_80_n 0.0212409f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_45 VPB C 0.00107117f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_46 VPB N_C_c_79_n 0.0165525f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_47 VPB N_B_c_105_n 0.0286264f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_48 VPB N_B_c_108_n 3.9349e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_49 VPB B 0.00308784f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_50 VPB N_A_c_144_n 0.0308007f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_51 VPB A 0.00194607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_193_n 0.0191527f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_53 VPB N_A_27_47#_c_194_n 0.0158902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_195_n 0.0158728f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_196_n 0.0192069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_197_n 0.00760212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_198_n 0.031746f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_188_n 0.00364539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_192_n 0.05671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_345_n 0.0077057f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_61 VPB N_VPWR_c_346_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_347_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_348_n 0.0208333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_349_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_350_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_351_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_352_n 0.0401334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_353_n 0.014713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_344_n 0.0518293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_355_n 0.0134384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_X_c_405_n 0.00202512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_X_c_406_n 0.0019944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_407_n 0.016631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_X_c_408_n 0.00158256f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB X 0.00835245f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 N_C_c_80_n N_B_c_105_n 0.0465224f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_77 N_C_c_79_n N_B_c_105_n 0.0255995f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_78 N_C_c_77_n N_B_c_106_n 0.0213001f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_79 C N_B_c_107_n 0.019637f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_80 N_C_c_79_n N_B_c_107_n 0.00225961f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_81 N_C_c_80_n B 0.00482378f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_C_c_79_n B 0.00230592f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_83 N_C_c_80_n N_A_27_47#_c_197_n 4.66918e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_84 N_C_c_80_n N_A_27_47#_c_198_n 0.0110053f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 C N_A_27_47#_c_198_n 0.0249698f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_86 N_C_c_79_n N_A_27_47#_c_198_n 0.00614661f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_87 N_C_c_77_n N_A_27_47#_c_184_n 0.0156229f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_88 N_C_c_79_n N_A_27_47#_c_184_n 8.91444e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_89 C N_A_27_47#_c_185_n 0.0281891f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_90 N_C_c_79_n N_A_27_47#_c_185_n 0.00777596f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_91 N_C_c_80_n N_A_27_47#_c_209_n 0.0129415f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_C_c_77_n N_A_27_47#_c_210_n 5.82315e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_93 N_C_c_80_n N_VPWR_c_352_n 0.00429425f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_C_c_80_n N_VPWR_c_344_n 0.00700259f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C_c_77_n N_VGND_c_475_n 0.00276126f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_96 N_C_c_77_n N_VGND_c_483_n 0.00703099f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_97 N_C_c_77_n N_VGND_c_484_n 0.00437852f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B_c_106_n N_A_c_143_n 0.0124239f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_99 N_B_c_105_n N_A_c_144_n 0.0758548f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_108_n N_A_c_144_n 8.7243e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B_c_105_n A 8.22176e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_108_n A 0.0224512f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_103 N_B_c_105_n N_A_27_47#_c_198_n 8.73858e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_105_n N_A_27_47#_c_184_n 0.00289838f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B_c_106_n N_A_27_47#_c_184_n 0.00616748f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_107_n N_A_27_47#_c_184_n 0.019812f $X=0.83 $Y=1.2 $X2=0 $Y2=0
cc_107 N_B_c_108_n N_A_27_47#_c_184_n 0.011123f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_108 N_B_c_105_n N_A_27_47#_c_209_n 0.0164077f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_109 B N_A_27_47#_c_209_n 0.00979454f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_110 N_B_c_106_n N_A_27_47#_c_210_n 0.00850899f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_c_105_n N_A_27_47#_c_219_n 5.45826e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_108_n N_A_27_47#_c_219_n 0.00403579f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B_c_105_n N_A_27_47#_c_190_n 0.00153559f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_106_n N_A_27_47#_c_190_n 0.00269873f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B_c_108_n N_A_27_47#_c_190_n 0.0137766f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_116 B A_117_297# 0.00751942f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_117 N_B_c_105_n N_VPWR_c_352_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B_c_105_n N_VPWR_c_344_n 0.00615826f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B_c_106_n N_VGND_c_475_n 0.00359159f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B_c_106_n N_VGND_c_483_n 0.00573353f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_106_n N_VGND_c_485_n 0.00396605f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_144_n N_A_27_47#_c_209_n 0.00434133f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_143_n N_A_27_47#_c_210_n 0.011462f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A_c_144_n N_A_27_47#_c_226_n 0.0189401f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_143_n N_A_27_47#_c_186_n 0.0109318f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_144_n N_A_27_47#_c_186_n 0.00487325f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_127 A N_A_27_47#_c_186_n 0.03606f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_128 N_A_c_144_n N_A_27_47#_c_230_n 0.0187681f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_129 A N_A_27_47#_c_230_n 0.0332549f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_130 N_A_c_144_n N_A_27_47#_c_219_n 0.00225738f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_131 A N_A_27_47#_c_219_n 0.00232727f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_132 N_A_c_143_n N_A_27_47#_c_187_n 0.0021454f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_144_n N_A_27_47#_c_187_n 0.00150782f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_144_n N_A_27_47#_c_188_n 0.00455986f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_135 A N_A_27_47#_c_188_n 0.00661024f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_136 N_A_c_143_n N_A_27_47#_c_190_n 0.00112787f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_137 A N_A_27_47#_c_190_n 0.00320352f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_138 N_A_c_144_n N_A_27_47#_c_191_n 4.82199e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_139 A N_A_27_47#_c_191_n 0.0155295f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_140 N_A_c_144_n N_A_27_47#_c_192_n 0.0101395f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_141 A N_A_27_47#_c_192_n 9.33627e-19 $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_142 N_A_c_144_n N_VPWR_c_345_n 0.0211587f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_144_n N_VPWR_c_352_n 0.00672099f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_144_n N_VPWR_c_344_n 0.0132832f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_143_n N_VGND_c_483_n 0.00719234f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_143_n N_VGND_c_485_n 0.00423334f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_143_n N_VGND_c_486_n 0.00618046f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_209_n A_117_297# 0.00385499f $X=1.1 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_27_47#_c_209_n A_211_297# 0.00172119f $X=1.1 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_27_47#_c_226_n A_211_297# 0.0013201f $X=1.232 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A_27_47#_c_219_n A_211_297# 0.0033751f $X=1.365 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_27_47#_c_230_n N_VPWR_M1012_d 0.0193483f $X=2.02 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_27_47#_c_188_n N_VPWR_M1012_d 2.36704e-19 $X=2.13 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_27_47#_c_193_n N_VPWR_c_345_n 0.00875484f $X=2.435 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_209_n N_VPWR_c_345_n 0.0121434f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_226_n N_VPWR_c_345_n 0.0306024f $X=1.232 $Y=2.295 $X2=0
+ $Y2=0
cc_157 N_A_27_47#_c_230_n N_VPWR_c_345_n 0.0550186f $X=2.02 $Y=1.58 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_189_n N_VPWR_c_345_n 0.00129928f $X=3.725 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_192_n N_VPWR_c_345_n 0.00158942f $X=3.845 $Y=1.202 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_194_n N_VPWR_c_346_n 0.00300743f $X=2.905 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_195_n N_VPWR_c_346_n 0.00300743f $X=3.375 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_196_n N_VPWR_c_347_n 0.00479105f $X=3.845 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_193_n N_VPWR_c_348_n 0.00702461f $X=2.435 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_194_n N_VPWR_c_348_n 0.00702461f $X=2.905 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_195_n N_VPWR_c_350_n 0.00702461f $X=3.375 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_196_n N_VPWR_c_350_n 0.00702461f $X=3.845 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_27_47#_c_197_n N_VPWR_c_352_n 0.0219164f $X=0.255 $Y=2.295 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_209_n N_VPWR_c_352_n 0.0538421f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_169 N_A_27_47#_M1005_s N_VPWR_c_344_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_170 N_A_27_47#_c_193_n N_VPWR_c_344_n 0.0137919f $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_194_n N_VPWR_c_344_n 0.0124092f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_195_n N_VPWR_c_344_n 0.0124092f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_196_n N_VPWR_c_344_n 0.0134885f $X=3.845 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_197_n N_VPWR_c_344_n 0.0129301f $X=0.255 $Y=2.295 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_209_n N_VPWR_c_344_n 0.0337013f $X=1.1 $Y=2.38 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_179_n N_X_c_410_n 0.0132627f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_186_n N_X_c_410_n 6.63905e-19 $X=2.02 $Y=0.815 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_194_n N_X_c_405_n 0.015887f $X=2.905 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_195_n N_X_c_405_n 0.0159694f $X=3.375 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_189_n N_X_c_405_n 0.0422526f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_192_n N_X_c_405_n 0.00888237f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_193_n N_X_c_406_n 4.68563e-19 $X=2.435 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_188_n N_X_c_406_n 0.00247314f $X=2.13 $Y=1.495 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_189_n N_X_c_406_n 0.0178591f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_192_n N_X_c_406_n 0.00678113f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_180_n N_X_c_399_n 0.0107068f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_181_n N_X_c_399_n 0.0060427f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_189_n N_X_c_399_n 0.0391606f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_192_n N_X_c_399_n 0.00345061f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_179_n N_X_c_400_n 0.00403483f $X=2.46 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_186_n N_X_c_400_n 0.0124162f $X=2.02 $Y=0.815 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_189_n N_X_c_400_n 0.030144f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_192_n N_X_c_400_n 0.00358132f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_180_n N_X_c_428_n 6.12918e-19 $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_181_n N_X_c_428_n 0.00862393f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_196_n N_X_c_407_n 0.0177141f $X=3.845 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_189_n N_X_c_407_n 0.0125781f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_192_n N_X_c_407_n 9.07829e-19 $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_182_n N_X_c_401_n 0.0122646f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_189_n N_X_c_401_n 0.0115602f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_181_n N_X_c_402_n 0.00266207f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_189_n N_X_c_402_n 0.030144f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_192_n N_X_c_402_n 0.00358132f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_189_n N_X_c_408_n 0.0178591f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_192_n N_X_c_408_n 0.00678113f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_206 N_A_27_47#_c_196_n X 0.00127652f $X=3.845 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_182_n X 0.00691871f $X=3.87 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_189_n X 0.0141296f $X=3.725 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_192_n X 0.00809906f $X=3.845 $Y=1.202 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_184_n N_VGND_M1010_d 0.00251047f $X=0.985 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_211 N_A_27_47#_c_186_n N_VGND_M1003_d 0.0128665f $X=2.02 $Y=0.815 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_184_n N_VGND_c_475_n 0.0127273f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_210_n N_VGND_c_475_n 0.0223967f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_180_n N_VGND_c_476_n 0.00276126f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_181_n N_VGND_c_476_n 0.0037534f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_182_n N_VGND_c_477_n 0.00438629f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_179_n N_VGND_c_478_n 0.00466554f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_180_n N_VGND_c_478_n 0.00439206f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_181_n N_VGND_c_480_n 0.00398337f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_182_n N_VGND_c_480_n 0.00439206f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_M1010_s N_VGND_c_483_n 0.00258952f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1001_d N_VGND_c_483_n 0.00215201f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_179_n N_VGND_c_483_n 0.00922919f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_180_n N_VGND_c_483_n 0.00616524f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_181_n N_VGND_c_483_n 0.0058274f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_182_n N_VGND_c_483_n 0.00716551f $X=3.87 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_183_n N_VGND_c_483_n 0.0130015f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_184_n N_VGND_c_483_n 0.00977515f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_229 N_A_27_47#_c_210_n N_VGND_c_483_n 0.0139016f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_186_n N_VGND_c_483_n 0.00780437f $X=2.02 $Y=0.815 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_183_n N_VGND_c_484_n 0.0225107f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_184_n N_VGND_c_484_n 0.00254521f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_233 N_A_27_47#_c_184_n N_VGND_c_485_n 0.00199443f $X=0.985 $Y=0.815 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_210_n N_VGND_c_485_n 0.0222529f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_186_n N_VGND_c_485_n 0.00266636f $X=2.02 $Y=0.815 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_179_n N_VGND_c_486_n 0.00612723f $X=2.46 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_210_n N_VGND_c_486_n 0.0204879f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_186_n N_VGND_c_486_n 0.0528905f $X=2.02 $Y=0.815 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_189_n N_VGND_c_486_n 0.00146636f $X=3.725 $Y=1.16 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_c_192_n N_VGND_c_486_n 0.00173974f $X=3.845 $Y=1.202 $X2=0
+ $Y2=0
cc_241 A_117_297# N_VPWR_c_344_n 0.00232895f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_242 A_211_297# N_VPWR_c_344_n 0.00232871f $X=1.055 $Y=1.485 $X2=1.1 $Y2=2.38
cc_243 N_VPWR_c_344_n N_X_M1002_s 0.00370124f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_244 N_VPWR_c_344_n N_X_M1009_s 0.00370124f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_348_n N_X_c_446_n 0.0149311f $X=3.015 $Y=2.72 $X2=0 $Y2=0
cc_246 N_VPWR_c_344_n N_X_c_446_n 0.00955092f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_247 N_VPWR_M1004_d N_X_c_405_n 0.00191634f $X=2.995 $Y=1.485 $X2=0 $Y2=0
cc_248 N_VPWR_c_346_n N_X_c_405_n 0.0137198f $X=3.14 $Y=1.96 $X2=0 $Y2=0
cc_249 N_VPWR_c_350_n N_X_c_450_n 0.0149311f $X=3.955 $Y=2.72 $X2=0 $Y2=0
cc_250 N_VPWR_c_344_n N_X_c_450_n 0.00955092f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_251 N_VPWR_M1013_d N_X_c_407_n 0.00826072f $X=3.935 $Y=1.485 $X2=0 $Y2=0
cc_252 N_VPWR_c_347_n N_X_c_407_n 0.0172399f $X=4.08 $Y=1.96 $X2=0 $Y2=0
cc_253 N_X_c_399_n N_VGND_M1007_d 0.00255557f $X=3.395 $Y=0.82 $X2=0 $Y2=0
cc_254 N_X_c_401_n N_VGND_M1011_d 0.00119049f $X=4.115 $Y=0.82 $X2=0 $Y2=0
cc_255 N_X_c_404_n N_VGND_M1011_d 0.00359674f $X=4.285 $Y=0.905 $X2=0 $Y2=0
cc_256 N_X_c_399_n N_VGND_c_476_n 0.012101f $X=3.395 $Y=0.82 $X2=0 $Y2=0
cc_257 N_X_c_428_n N_VGND_c_476_n 0.0216501f $X=3.61 $Y=0.39 $X2=0 $Y2=0
cc_258 N_X_c_401_n N_VGND_c_477_n 0.00840877f $X=4.115 $Y=0.82 $X2=0 $Y2=0
cc_259 N_X_c_404_n N_VGND_c_477_n 0.00404097f $X=4.285 $Y=0.905 $X2=0 $Y2=0
cc_260 N_X_c_410_n N_VGND_c_478_n 0.0216696f $X=2.67 $Y=0.39 $X2=0 $Y2=0
cc_261 N_X_c_399_n N_VGND_c_478_n 0.00248202f $X=3.395 $Y=0.82 $X2=0 $Y2=0
cc_262 N_X_c_399_n N_VGND_c_480_n 0.00194552f $X=3.395 $Y=0.82 $X2=0 $Y2=0
cc_263 N_X_c_428_n N_VGND_c_480_n 0.0216696f $X=3.61 $Y=0.39 $X2=0 $Y2=0
cc_264 N_X_c_401_n N_VGND_c_480_n 0.00248202f $X=4.115 $Y=0.82 $X2=0 $Y2=0
cc_265 N_X_c_404_n N_VGND_c_482_n 0.00474764f $X=4.285 $Y=0.905 $X2=0 $Y2=0
cc_266 N_X_M1006_s N_VGND_c_483_n 0.00264648f $X=2.535 $Y=0.235 $X2=0 $Y2=0
cc_267 N_X_M1008_s N_VGND_c_483_n 0.00264648f $X=3.475 $Y=0.235 $X2=0 $Y2=0
cc_268 N_X_c_410_n N_VGND_c_483_n 0.0140292f $X=2.67 $Y=0.39 $X2=0 $Y2=0
cc_269 N_X_c_399_n N_VGND_c_483_n 0.0096764f $X=3.395 $Y=0.82 $X2=0 $Y2=0
cc_270 N_X_c_428_n N_VGND_c_483_n 0.0140292f $X=3.61 $Y=0.39 $X2=0 $Y2=0
cc_271 N_X_c_401_n N_VGND_c_483_n 0.00538201f $X=4.115 $Y=0.82 $X2=0 $Y2=0
cc_272 N_X_c_404_n N_VGND_c_483_n 0.00836179f $X=4.285 $Y=0.905 $X2=0 $Y2=0
cc_273 N_X_c_410_n N_VGND_c_486_n 0.0241592f $X=2.67 $Y=0.39 $X2=0 $Y2=0
