* File: sky130_fd_sc_hdll__a32o_1.pxi.spice
* Created: Wed Sep  2 08:20:34 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32O_1%A_93_21# N_A_93_21#_M1003_d N_A_93_21#_M1002_d
+ N_A_93_21#_c_60_n N_A_93_21#_M1005_g N_A_93_21#_c_61_n N_A_93_21#_M1001_g
+ N_A_93_21#_c_65_n N_A_93_21#_c_69_p N_A_93_21#_c_112_p N_A_93_21#_c_70_p
+ N_A_93_21#_c_116_p N_A_93_21#_c_75_p N_A_93_21#_c_76_p N_A_93_21#_c_71_p
+ N_A_93_21#_c_101_p N_A_93_21#_c_62_n N_A_93_21#_c_63_n
+ PM_SKY130_FD_SC_HDLL__A32O_1%A_93_21#
x_PM_SKY130_FD_SC_HDLL__A32O_1%A3 N_A3_c_157_n N_A3_M1009_g N_A3_c_158_n
+ N_A3_M1000_g A3 A3 PM_SKY130_FD_SC_HDLL__A32O_1%A3
x_PM_SKY130_FD_SC_HDLL__A32O_1%A2 N_A2_c_191_n N_A2_M1004_g N_A2_c_192_n
+ N_A2_M1007_g A2 A2 PM_SKY130_FD_SC_HDLL__A32O_1%A2
x_PM_SKY130_FD_SC_HDLL__A32O_1%A1 N_A1_c_226_n N_A1_M1008_g N_A1_c_227_n
+ N_A1_M1003_g A1 A1 N_A1_c_229_n PM_SKY130_FD_SC_HDLL__A32O_1%A1
x_PM_SKY130_FD_SC_HDLL__A32O_1%B1 N_B1_c_259_n N_B1_M1002_g N_B1_c_260_n
+ N_B1_M1006_g B1 B1 PM_SKY130_FD_SC_HDLL__A32O_1%B1
x_PM_SKY130_FD_SC_HDLL__A32O_1%B2 N_B2_c_291_n N_B2_M1011_g N_B2_c_292_n
+ N_B2_M1010_g N_B2_c_293_n B2 B2 N_B2_c_294_n PM_SKY130_FD_SC_HDLL__A32O_1%B2
x_PM_SKY130_FD_SC_HDLL__A32O_1%X N_X_M1005_s N_X_M1001_s X X X X X X X
+ N_X_c_321_n X PM_SKY130_FD_SC_HDLL__A32O_1%X
x_PM_SKY130_FD_SC_HDLL__A32O_1%VPWR N_VPWR_M1001_d N_VPWR_M1007_d N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_341_n N_VPWR_c_342_n VPWR N_VPWR_c_343_n
+ N_VPWR_c_344_n N_VPWR_c_338_n N_VPWR_c_346_n PM_SKY130_FD_SC_HDLL__A32O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A32O_1%A_268_297# N_A_268_297#_M1009_d
+ N_A_268_297#_M1008_d N_A_268_297#_M1010_d N_A_268_297#_c_391_n
+ N_A_268_297#_c_409_n N_A_268_297#_c_392_n N_A_268_297#_c_393_n
+ N_A_268_297#_c_387_n N_A_268_297#_c_418_n N_A_268_297#_c_388_n
+ PM_SKY130_FD_SC_HDLL__A32O_1%A_268_297#
x_PM_SKY130_FD_SC_HDLL__A32O_1%VGND N_VGND_M1005_d N_VGND_M1011_d N_VGND_c_420_n
+ N_VGND_c_421_n N_VGND_c_422_n VGND N_VGND_c_423_n N_VGND_c_424_n
+ N_VGND_c_425_n N_VGND_c_426_n PM_SKY130_FD_SC_HDLL__A32O_1%VGND
cc_1 VNB N_A_93_21#_c_60_n 0.0214698f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB N_A_93_21#_c_61_n 0.0278773f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.41
cc_3 VNB N_A_93_21#_c_62_n 0.00285601f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_4 VNB N_A_93_21#_c_63_n 0.00204748f $X=-0.19 $Y=-0.24 $X2=0.707 $Y2=0.995
cc_5 VNB N_A3_c_157_n 0.0271101f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0.235
cc_6 VNB N_A3_c_158_n 0.0191663f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB A3 0.00284997f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_8 VNB N_A2_c_191_n 0.0175079f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0.235
cc_9 VNB N_A2_c_192_n 0.0237946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A2 0.00401345f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_11 VNB N_A1_c_226_n 0.0252664f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0.235
cc_12 VNB N_A1_c_227_n 0.0193357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A1 4.61796e-19 $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_14 VNB N_A1_c_229_n 0.00421814f $X=-0.19 $Y=-0.24 $X2=0.76 $Y2=0.825
cc_15 VNB N_B1_c_259_n 0.0251324f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0.235
cc_16 VNB N_B1_c_260_n 0.0169386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB B1 0.00273498f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_18 VNB N_B2_c_291_n 0.0207468f $X=-0.19 $Y=-0.24 $X2=2.53 $Y2=0.235
cc_19 VNB N_B2_c_292_n 0.0287521f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B2_c_293_n 8.57664e-19 $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_21 VNB N_B2_c_294_n 0.0208583f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=0.74
cc_22 VNB X 0.0341419f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_23 VNB N_X_c_321_n 0.0104776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_338_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0.707 $Y2=0.995
cc_25 VNB N_VGND_c_420_n 0.00315146f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.56
cc_26 VNB N_VGND_c_421_n 0.0164311f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.985
cc_27 VNB N_VGND_c_422_n 0.025814f $X=-0.19 $Y=-0.24 $X2=0.76 $Y2=0.825
cc_28 VNB N_VGND_c_423_n 0.0171616f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=0.74
cc_29 VNB N_VGND_c_424_n 0.062984f $X=-0.19 $Y=-0.24 $X2=1.23 $Y2=0.655
cc_30 VNB N_VGND_c_425_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0.707 $Y2=1.16
cc_31 VNB N_VGND_c_426_n 0.225558f $X=-0.19 $Y=-0.24 $X2=0.707 $Y2=1.325
cc_32 VPB N_A_93_21#_c_61_n 0.0327672f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.41
cc_33 VPB N_A_93_21#_c_65_n 0.00284944f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=1.495
cc_34 VPB N_A_93_21#_c_62_n 4.93889e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_35 VPB N_A3_c_157_n 0.0299156f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=0.235
cc_36 VPB A3 0.00104734f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_37 VPB N_A2_c_192_n 0.0289498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB A2 0.00220454f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_39 VPB N_A1_c_226_n 0.0294497f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=0.235
cc_40 VPB N_A1_c_229_n 0.00202173f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=0.825
cc_41 VPB N_B1_c_259_n 0.0279228f $X=-0.19 $Y=1.305 $X2=2.53 $Y2=0.235
cc_42 VPB B1 0.00105015f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_43 VPB N_B2_c_292_n 0.0323824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_B2_c_293_n 0.00126766f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_45 VPB B2 0.019644f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=0.825
cc_46 VPB N_B2_c_294_n 8.73081e-19 $X=-0.19 $Y=1.305 $X2=1.145 $Y2=0.74
cc_47 VPB X 0.025687f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_48 VPB X 0.0065071f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.985
cc_49 VPB X 0.0136697f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.985
cc_50 VPB N_VPWR_c_339_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_51 VPB N_VPWR_c_340_n 0.00564356f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=0.825
cc_52 VPB N_VPWR_c_341_n 0.0223171f $X=-0.19 $Y=1.305 $X2=0.76 $Y2=1.495
cc_53 VPB N_VPWR_c_342_n 0.00632158f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=0.74
cc_54 VPB N_VPWR_c_343_n 0.0241764f $X=-0.19 $Y=1.305 $X2=2.745 $Y2=0.4
cc_55 VPB N_VPWR_c_344_n 0.0475383f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.16
cc_56 VPB N_VPWR_c_338_n 0.0505846f $X=-0.19 $Y=1.305 $X2=0.707 $Y2=0.995
cc_57 VPB N_VPWR_c_346_n 0.00631679f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_268_297#_c_387_n 0.00759475f $X=-0.19 $Y=1.305 $X2=0.845 $Y2=0.74
cc_59 VPB N_A_268_297#_c_388_n 0.019434f $X=-0.19 $Y=1.305 $X2=1.23 $Y2=0.655
cc_60 N_A_93_21#_c_61_n N_A3_c_157_n 0.0362026f $X=0.565 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_61 N_A_93_21#_c_65_n N_A3_c_157_n 0.00326099f $X=0.76 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A_93_21#_c_69_p N_A3_c_157_n 0.00275737f $X=1.145 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_63 N_A_93_21#_c_70_p N_A3_c_157_n 0.0222711f $X=3.155 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_93_21#_c_71_p N_A3_c_157_n 0.0016757f $X=2.745 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_93_21#_c_62_n N_A3_c_157_n 9.02808e-19 $X=0.655 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_93_21#_c_60_n N_A3_c_158_n 0.00899518f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_93_21#_c_69_p N_A3_c_158_n 0.00710672f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_68 N_A_93_21#_c_75_p N_A3_c_158_n 0.00560289f $X=1.23 $Y=0.655 $X2=0 $Y2=0
cc_69 N_A_93_21#_c_76_p N_A3_c_158_n 0.00425099f $X=1.315 $Y=0.4 $X2=0 $Y2=0
cc_70 N_A_93_21#_c_71_p N_A3_c_158_n 0.00589174f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_71 N_A_93_21#_c_63_n N_A3_c_158_n 0.0030684f $X=0.707 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_93_21#_c_61_n A3 0.00105576f $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_73 N_A_93_21#_c_69_p A3 0.0210144f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_93_21#_c_70_p A3 0.022465f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A_93_21#_c_71_p A3 0.00115107f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_76 N_A_93_21#_c_62_n A3 0.0271209f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_93_21#_c_69_p N_A2_c_191_n 2.00732e-19 $X=1.145 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_93_21#_c_75_p N_A2_c_191_n 9.22582e-19 $X=1.23 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_93_21#_c_71_p N_A2_c_191_n 0.0113566f $X=2.745 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_93_21#_c_70_p N_A2_c_192_n 0.0155584f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_93_21#_c_71_p N_A2_c_192_n 0.00168277f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_82 N_A_93_21#_c_69_p A2 0.0113525f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_93_21#_c_70_p A2 0.029267f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_84 N_A_93_21#_c_71_p A2 0.0219141f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_85 N_A_93_21#_c_70_p N_A1_c_226_n 0.0157465f $X=3.155 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_93_21#_c_71_p N_A1_c_226_n 0.00178923f $X=2.745 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_93_21#_c_71_p N_A1_c_227_n 0.0118757f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_88 N_A_93_21#_M1003_d A1 0.0028545f $X=2.53 $Y=0.235 $X2=0 $Y2=0
cc_89 N_A_93_21#_c_71_p A1 0.0158347f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_90 N_A_93_21#_c_70_p N_A1_c_229_n 0.0271881f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_93_21#_c_71_p N_A1_c_229_n 0.00356529f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_92 N_A_93_21#_c_70_p N_B1_c_259_n 0.0161052f $X=3.155 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_93_21#_c_71_p N_B1_c_259_n 2.06151e-19 $X=2.745 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_93_21#_c_101_p N_B1_c_259_n 0.00558198f $X=3.24 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_93_21#_c_71_p N_B1_c_260_n 0.00272261f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_96 N_A_93_21#_M1003_d B1 0.00387504f $X=2.53 $Y=0.235 $X2=0 $Y2=0
cc_97 N_A_93_21#_c_70_p B1 0.019323f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_98 N_A_93_21#_c_71_p B1 0.00555891f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_99 N_A_93_21#_c_70_p N_B2_c_292_n 0.00322653f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_100 N_A_93_21#_c_101_p N_B2_c_292_n 0.00449951f $X=3.24 $Y=1.96 $X2=0 $Y2=0
cc_101 N_A_93_21#_c_70_p B2 0.00472671f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_93_21#_c_60_n X 0.021481f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_93_21#_c_61_n X 0.0142768f $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_93_21#_c_65_n X 0.00801843f $X=0.76 $Y=1.495 $X2=0 $Y2=0
cc_105 N_A_93_21#_c_112_p X 0.00866435f $X=0.845 $Y=0.74 $X2=0 $Y2=0
cc_106 N_A_93_21#_c_62_n X 0.0204748f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_93_21#_c_63_n X 0.00809463f $X=0.707 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_93_21#_c_70_p N_VPWR_M1001_d 0.00958444f $X=3.155 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_109 N_A_93_21#_c_116_p N_VPWR_M1001_d 0.00311522f $X=0.845 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_110 N_A_93_21#_c_70_p N_VPWR_M1007_d 0.0146872f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_111 N_A_93_21#_c_61_n N_VPWR_c_339_n 0.0123596f $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_93_21#_c_70_p N_VPWR_c_339_n 0.0169675f $X=3.155 $Y=1.58 $X2=0 $Y2=0
cc_113 N_A_93_21#_c_116_p N_VPWR_c_339_n 0.0106842f $X=0.845 $Y=1.58 $X2=0 $Y2=0
cc_114 N_A_93_21#_c_61_n N_VPWR_c_341_n 0.00702461f $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_93_21#_M1002_d N_VPWR_c_338_n 0.00240926f $X=3.09 $Y=1.485 $X2=0
+ $Y2=0
cc_116 N_A_93_21#_c_61_n N_VPWR_c_338_n 0.0141659f $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_93_21#_c_70_p N_A_268_297#_M1009_d 0.00686999f $X=3.155 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_118 N_A_93_21#_c_70_p N_A_268_297#_M1008_d 0.0111156f $X=3.155 $Y=1.58 $X2=0
+ $Y2=0
cc_119 N_A_93_21#_c_70_p N_A_268_297#_c_391_n 0.0162181f $X=3.155 $Y=1.58 $X2=0
+ $Y2=0
cc_120 N_A_93_21#_c_70_p N_A_268_297#_c_392_n 0.0426634f $X=3.155 $Y=1.58 $X2=0
+ $Y2=0
cc_121 N_A_93_21#_c_70_p N_A_268_297#_c_393_n 0.0189669f $X=3.155 $Y=1.58 $X2=0
+ $Y2=0
cc_122 N_A_93_21#_M1002_d N_A_268_297#_c_387_n 0.00403964f $X=3.09 $Y=1.485
+ $X2=0 $Y2=0
cc_123 N_A_93_21#_c_70_p N_A_268_297#_c_387_n 0.00431302f $X=3.155 $Y=1.58 $X2=0
+ $Y2=0
cc_124 N_A_93_21#_c_101_p N_A_268_297#_c_387_n 0.0127257f $X=3.24 $Y=1.96 $X2=0
+ $Y2=0
cc_125 N_A_93_21#_c_101_p N_A_268_297#_c_388_n 0.0159059f $X=3.24 $Y=1.96 $X2=0
+ $Y2=0
cc_126 N_A_93_21#_c_69_p N_VGND_M1005_d 0.0110651f $X=1.145 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_93_21#_c_112_p N_VGND_M1005_d 0.0051458f $X=0.845 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_128 N_A_93_21#_c_75_p N_VGND_M1005_d 0.00265633f $X=1.23 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_129 N_A_93_21#_c_76_p N_VGND_M1005_d 0.00199936f $X=1.315 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_93_21#_c_63_n N_VGND_M1005_d 0.00144856f $X=0.707 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_93_21#_c_60_n N_VGND_c_420_n 0.0103776f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_93_21#_c_61_n N_VGND_c_420_n 5.9868e-19 $X=0.565 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_93_21#_c_69_p N_VGND_c_420_n 0.00986995f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_93_21#_c_112_p N_VGND_c_420_n 0.014416f $X=0.845 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_93_21#_c_76_p N_VGND_c_420_n 0.0146233f $X=1.315 $Y=0.4 $X2=0 $Y2=0
cc_136 N_A_93_21#_c_62_n N_VGND_c_420_n 0.00157277f $X=0.655 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_93_21#_c_71_p N_VGND_c_422_n 0.0052136f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_138 N_A_93_21#_c_60_n N_VGND_c_423_n 0.00505556f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_93_21#_c_69_p N_VGND_c_424_n 0.00283163f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_140 N_A_93_21#_c_76_p N_VGND_c_424_n 0.0069528f $X=1.315 $Y=0.4 $X2=0 $Y2=0
cc_141 N_A_93_21#_c_71_p N_VGND_c_424_n 0.0669684f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_142 N_A_93_21#_M1003_d N_VGND_c_426_n 0.00446095f $X=2.53 $Y=0.235 $X2=0
+ $Y2=0
cc_143 N_A_93_21#_c_60_n N_VGND_c_426_n 0.00963589f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_93_21#_c_69_p N_VGND_c_426_n 0.0053278f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_93_21#_c_112_p N_VGND_c_426_n 8.26975e-19 $X=0.845 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_93_21#_c_76_p N_VGND_c_426_n 0.00588979f $X=1.315 $Y=0.4 $X2=0 $Y2=0
cc_147 N_A_93_21#_c_71_p N_VGND_c_426_n 0.0554977f $X=2.745 $Y=0.4 $X2=0 $Y2=0
cc_148 N_A_93_21#_c_71_p A_276_47# 0.00568658f $X=2.745 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_93_21#_c_71_p A_366_47# 0.01753f $X=2.745 $Y=0.4 $X2=-0.19 $Y2=-0.24
cc_150 N_A3_c_158_n N_A2_c_191_n 0.0365601f $X=1.305 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A3_c_157_n N_A2_c_192_n 0.0430721f $X=1.25 $Y=1.41 $X2=0 $Y2=0
cc_152 A3 N_A2_c_192_n 2.57201e-19 $X=1.12 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A3_c_157_n A2 0.00247386f $X=1.25 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A3_c_158_n A2 0.0055162f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_155 A3 A2 0.0266717f $X=1.12 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A3_c_157_n N_VPWR_c_339_n 0.01119f $X=1.25 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A3_c_157_n N_VPWR_c_343_n 0.00702461f $X=1.25 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A3_c_157_n N_VPWR_c_338_n 0.0133143f $X=1.25 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A3_c_158_n N_VGND_c_420_n 0.00477504f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A3_c_158_n N_VGND_c_424_n 0.00370003f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A3_c_158_n N_VGND_c_426_n 0.00608187f $X=1.305 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_192_n N_A1_c_226_n 0.0530506f $X=1.78 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_163 A2 N_A1_c_226_n 0.00109533f $X=1.585 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_164 N_A2_c_191_n N_A1_c_227_n 0.017921f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_165 A2 N_A1_c_227_n 0.00235163f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_166 N_A2_c_191_n A1 3.00622e-19 $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_167 A2 A1 0.0112236f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_168 N_A2_c_192_n N_A1_c_229_n 0.00109563f $X=1.78 $Y=1.41 $X2=0 $Y2=0
cc_169 A2 N_A1_c_229_n 0.0181324f $X=1.585 $Y=0.765 $X2=0 $Y2=0
cc_170 N_A2_c_192_n N_VPWR_c_340_n 0.00653952f $X=1.78 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A2_c_192_n N_VPWR_c_343_n 0.00517074f $X=1.78 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A2_c_192_n N_VPWR_c_338_n 0.0074085f $X=1.78 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A2_c_192_n N_A_268_297#_c_392_n 0.0127248f $X=1.78 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_191_n N_VGND_c_424_n 0.00370116f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_c_191_n N_VGND_c_426_n 0.00598773f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_176 A2 A_276_47# 0.0033096f $X=1.585 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_177 A2 A_366_47# 0.00381643f $X=1.585 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_178 N_A1_c_226_n N_B1_c_259_n 0.0422794f $X=2.43 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_179 N_A1_c_229_n N_B1_c_259_n 0.00119392f $X=2.345 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A1_c_227_n N_B1_c_260_n 0.0207598f $X=2.455 $Y=0.995 $X2=0 $Y2=0
cc_181 A1 N_B1_c_260_n 8.57919e-19 $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_182 N_A1_c_227_n B1 0.00192735f $X=2.455 $Y=0.995 $X2=0 $Y2=0
cc_183 A1 B1 0.0540782f $X=2.44 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A1_c_226_n N_VPWR_c_340_n 0.00642273f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A1_c_226_n N_VPWR_c_344_n 0.00517074f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A1_c_226_n N_VPWR_c_338_n 0.00749122f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A1_c_226_n N_A_268_297#_c_392_n 0.0127248f $X=2.43 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A1_c_227_n N_VGND_c_424_n 0.00370116f $X=2.455 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_227_n N_VGND_c_426_n 0.00636922f $X=2.455 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_260_n N_B2_c_291_n 0.037167f $X=3.095 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_191 B1 N_B2_c_291_n 0.0027437f $X=2.89 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_192 N_B1_c_259_n N_B2_c_292_n 0.0748219f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B1_c_259_n N_B2_c_293_n 0.00107771f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_194 B1 N_B2_c_293_n 0.0165339f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_195 N_B1_c_259_n N_VPWR_c_344_n 0.00429453f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B1_c_259_n N_VPWR_c_338_n 0.00640989f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_259_n N_A_268_297#_c_387_n 0.0138137f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B1_c_260_n N_VGND_c_422_n 0.0032765f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_199 B1 N_VGND_c_422_n 0.00584599f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_200 N_B1_c_260_n N_VGND_c_424_n 0.00466229f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_201 B1 N_VGND_c_424_n 0.0034258f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_202 N_B1_c_260_n N_VGND_c_426_n 0.00746504f $X=3.095 $Y=0.995 $X2=0 $Y2=0
cc_203 B1 N_VGND_c_426_n 0.00620946f $X=2.89 $Y=0.765 $X2=0 $Y2=0
cc_204 N_B2_c_292_n N_VPWR_c_344_n 0.00429453f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B2_c_292_n N_VPWR_c_338_n 0.00714844f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_206 B2 N_A_268_297#_M1010_d 0.00264558f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_207 N_B2_c_292_n N_A_268_297#_c_387_n 0.0143719f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B2_c_292_n N_A_268_297#_c_388_n 0.00122211f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B2_c_293_n N_A_268_297#_c_388_n 0.00613441f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_210 B2 N_A_268_297#_c_388_n 0.00899927f $X=3.825 $Y=1.445 $X2=0 $Y2=0
cc_211 N_B2_c_291_n N_VGND_c_422_n 0.0159154f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B2_c_292_n N_VGND_c_422_n 0.00390066f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B2_c_293_n N_VGND_c_422_n 0.0193969f $X=3.79 $Y=1.16 $X2=0 $Y2=0
cc_214 N_B2_c_294_n N_VGND_c_422_n 0.00798179f $X=3.91 $Y=1.325 $X2=0 $Y2=0
cc_215 N_B2_c_291_n N_VGND_c_424_n 0.00486043f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B2_c_291_n N_VGND_c_426_n 0.00814024f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_217 X N_VPWR_c_339_n 0.00345753f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_218 X N_VPWR_c_341_n 0.0184261f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_219 N_X_M1001_s N_VPWR_c_338_n 0.00455261f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_220 X N_VPWR_c_338_n 0.0125459f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_221 N_X_c_321_n N_VGND_c_423_n 0.0175601f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_222 N_X_M1005_s N_VGND_c_426_n 0.00412857f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_223 N_X_c_321_n N_VGND_c_426_n 0.012458f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_224 N_VPWR_c_338_n N_A_268_297#_M1009_d 0.00336199f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_225 N_VPWR_c_338_n N_A_268_297#_M1008_d 0.0032252f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_226 N_VPWR_c_338_n N_A_268_297#_M1010_d 0.00221622f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_227 N_VPWR_c_343_n N_A_268_297#_c_409_n 0.018092f $X=1.94 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_c_338_n N_A_268_297#_c_409_n 0.0108535f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_229 N_VPWR_M1007_d N_A_268_297#_c_392_n 0.00885533f $X=1.87 $Y=1.485 $X2=0
+ $Y2=0
cc_230 N_VPWR_c_340_n N_A_268_297#_c_392_n 0.025328f $X=2.105 $Y=2.34 $X2=0
+ $Y2=0
cc_231 N_VPWR_c_343_n N_A_268_297#_c_392_n 0.00386992f $X=1.94 $Y=2.72 $X2=0
+ $Y2=0
cc_232 N_VPWR_c_344_n N_A_268_297#_c_392_n 0.00360543f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_VPWR_c_338_n N_A_268_297#_c_392_n 0.0154596f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_344_n N_A_268_297#_c_387_n 0.059987f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_338_n N_A_268_297#_c_387_n 0.0366007f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_344_n N_A_268_297#_c_418_n 0.0211241f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_338_n N_A_268_297#_c_418_n 0.0126619f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VGND_c_426_n A_276_47# 0.00246016f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_239 N_VGND_c_426_n A_366_47# 0.00454223f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
cc_240 N_VGND_c_426_n A_634_47# 0.00897657f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
