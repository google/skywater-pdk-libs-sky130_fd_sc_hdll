* File: sky130_fd_sc_hdll__mux2_1.spice
* Created: Thu Aug 27 19:10:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2_1.pex.spice"
.subckt sky130_fd_sc_hdll__mux2_1  VNB VPB S A1 A0 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_A_79_21#_M1010_g N_X_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.178537 AS=0.169 PD=1.43364 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1000 A_245_47# N_S_M1000_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42 AD=0.0756
+ AS=0.115363 PD=0.78 PS=0.926355 NRD=35.712 NRS=58.56 M=1 R=2.8 SA=75000.9
+ SB=75003 A=0.063 P=1.14 MULT=1
MM1004 N_A_79_21#_M1004_d N_A1_M1004_g A_245_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.0756 PD=1.03 PS=0.78 NRD=0 NRS=35.712 M=1 R=2.8 SA=75001.4
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 A_499_47# N_A0_M1007_g N_A_79_21#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1659 AS=0.1281 PD=1.21 PS=1.03 NRD=97.14 NRS=95.712 M=1 R=2.8 SA=75002.1
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_657_21#_M1001_g A_499_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0903 AS=0.1659 PD=0.85 PS=1.21 NRD=30 NRS=97.14 M=1 R=2.8 SA=75003.1
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_657_21#_M1008_d N_S_M1008_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0903 PD=1.36 PS=0.85 NRD=0 NRS=12.852 M=1 R=2.8 SA=75003.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_VPWR_M1005_d N_A_79_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.24338 AS=0.27 PD=2.04225 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1009 A_243_374# N_S_M1009_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.08715 AS=0.10222 PD=0.835 PS=0.857746 NRD=71.511 NRS=78.5636 M=1
+ R=2.33333 SA=90000.8 SB=90003 A=0.0756 P=1.2 MULT=1
MM1002 N_A_79_21#_M1002_d N_A0_M1002_g A_243_374# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.22575 AS=0.08715 PD=1.495 PS=0.835 NRD=28.1316 NRS=71.511 M=1 R=2.33333
+ SA=90001.4 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1003 A_613_374# N_A1_M1003_g N_A_79_21#_M1002_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.22575 PD=0.65 PS=1.495 NRD=28.1316 NRS=98.4803 M=1 R=2.33333
+ SA=90002.7 SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_657_21#_M1006_g A_613_374# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0735 AS=0.0483 PD=0.77 PS=0.65 NRD=25.7873 NRS=28.1316 M=1 R=2.33333
+ SA=90003.1 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_A_657_21#_M1011_d N_S_M1011_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1218 AS=0.0735 PD=1.42 PS=0.77 NRD=2.3443 NRS=7.0329 M=1 R=2.33333
+ SA=90003.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX13_noxref noxref_15 A0 A0 PROBETYPE=1
c_35 VNB 0 1.9931e-19 $X=0.42 $Y=-0.085
*
.include "sky130_fd_sc_hdll__mux2_1.pxi.spice"
*
.ends
*
*
