* File: sky130_fd_sc_hdll__or4b_1.spice
* Created: Thu Aug 27 19:25:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4b_1.pex.spice"
.subckt sky130_fd_sc_hdll__or4b_1  VNB VPB D_N C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1000 N_A_117_297#_M1000_d N_D_N_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_225_297#_M1001_d N_A_117_297#_M1001_g N_VGND_M1001_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.07455 AS=0.1302 PD=0.775 PS=1.46 NRD=7.14 NRS=12.852 M=1
+ R=2.8 SA=75000.2 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_225_297#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0609 AS=0.07455 PD=0.71 PS=0.775 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.7
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1006 N_A_225_297#_M1006_d N_B_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0735 AS=0.0609 PD=0.77 PS=0.71 NRD=7.14 NRS=4.284 M=1 R=2.8 SA=75001.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_M1003_g N_A_225_297#_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.0735 PD=0.816449 PS=0.77 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_225_297#_M1002_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17875 AS=0.143516 PD=1.85 PS=1.26355 NRD=0 NRS=11.988 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_117_297#_M1004_d N_D_N_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1009 A_315_297# N_A_117_297#_M1009_g N_A_225_297#_M1009_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.06825 AS=0.1134 PD=0.745 PS=1.38 NRD=50.4123 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1010 A_416_297# N_C_M1010_g A_315_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0546
+ AS=0.06825 PD=0.68 PS=0.745 NRD=35.1645 NRS=50.4123 M=1 R=2.33333 SA=90000.7
+ SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1005 A_504_297# N_B_M1005_g A_416_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0672
+ AS=0.0546 PD=0.74 PS=0.68 NRD=49.25 NRS=35.1645 M=1 R=2.33333 SA=90001.1
+ SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_504_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0672 PD=0.804507 PS=0.74 NRD=76.83 NRS=49.25 M=1 R=2.33333
+ SA=90001.6 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1011 N_X_M1011_d N_A_225_297#_M1011_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.285 AS=0.218803 PD=2.57 PS=1.91549 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90001 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_15 B B PROBETYPE=1
pX14_noxref noxref_16 B B PROBETYPE=1
pX15_noxref noxref_17 C C PROBETYPE=1
pX16_noxref noxref_18 C C PROBETYPE=1
pX17_noxref noxref_19 B B PROBETYPE=1
c_70 VPB 0 2.02209e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or4b_1.pxi.spice"
*
.ends
*
*
