* File: sky130_fd_sc_hdll__nand4_2.pex.spice
* Created: Wed Sep  2 08:38:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%D 3 5 8 10 12 15 17 18 21 26
c46 18 0 1.26238e-19 $X=0.695 $Y=1.19
c47 15 0 8.56806e-20 $X=0.99 $Y=0.56
r48 26 27 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=0.99 $Y2=1.217
r49 24 26 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=0.73 $Y=1.217
+ $X2=0.965 $Y2=1.217
r50 22 24 29.9467 $w=3.38e-07 $l=2.1e-07 $layer=POLY_cond $X=0.52 $Y=1.217
+ $X2=0.73 $Y2=1.217
r51 21 22 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.52 $Y2=1.217
r52 18 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=1.16 $X2=0.73 $Y2=1.16
r53 17 18 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r54 13 27 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.217
r55 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r56 10 26 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r57 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r58 6 22 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.217
r59 6 8 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r60 3 21 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r61 3 5 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%C 3 5 7 8 10 13 15 16 24
c48 24 0 1.26238e-19 $X=1.905 $Y=1.217
c49 16 0 1.89496e-19 $X=1.765 $Y=1.19
c50 3 0 1.79953e-19 $X=1.41 $Y=0.56
r51 24 25 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r52 22 24 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=1.67 $Y=1.217
+ $X2=1.905 $Y2=1.217
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r54 20 22 33.5118 $w=3.38e-07 $l=2.35e-07 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.67 $Y2=1.217
r55 19 20 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.217
+ $X2=1.435 $Y2=1.217
r56 16 23 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=1.765 $Y=1.175
+ $X2=1.67 $Y2=1.175
r57 15 23 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=1.255 $Y=1.175
+ $X2=1.67 $Y2=1.175
r58 11 25 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r59 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r60 8 24 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r61 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r62 5 20 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r63 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r64 1 19 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.217
r65 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%B 1 3 4 6 9 13 15 19 20 21 30
c52 21 0 1.68817e-19 $X=3.295 $Y=1.19
c53 15 0 1.89496e-19 $X=3.105 $Y=1.16
r54 26 30 22.1818 $w=1.98e-07 $l=4e-07 $layer=LI1_cond $X=3.19 $Y=1.175 $X2=2.79
+ $Y2=1.175
r55 25 26 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.19
+ $Y=1.16 $X2=3.19 $Y2=1.16
r56 21 26 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=3.295 $Y=1.175
+ $X2=3.19 $Y2=1.175
r57 20 30 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.785 $Y=1.175
+ $X2=2.79 $Y2=1.175
r58 19 25 47.7673 $w=2.7e-07 $l=2.15e-07 $layer=POLY_cond $X=3.405 $Y=1.16
+ $X2=3.19 $Y2=1.16
r59 17 18 0.713018 $w=3.38e-07 $l=5e-09 $layer=POLY_cond $X=3.005 $Y=1.217
+ $X2=3.01 $Y2=1.217
r60 16 17 67.0237 $w=3.38e-07 $l=4.7e-07 $layer=POLY_cond $X=2.535 $Y=1.217
+ $X2=3.005 $Y2=1.217
r61 15 25 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=3.105 $Y=1.16
+ $X2=3.19 $Y2=1.16
r62 15 18 15.6366 $w=3.38e-07 $l=1.20167e-07 $layer=POLY_cond $X=3.105 $Y=1.16
+ $X2=3.01 $Y2=1.217
r63 11 19 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=3.48 $Y=1.025
+ $X2=3.405 $Y2=1.16
r64 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.48 $Y=1.025
+ $X2=3.48 $Y2=0.56
r65 7 18 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=3.01 $Y2=1.217
r66 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.01 $Y=1.025
+ $X2=3.01 $Y2=0.56
r67 4 17 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.217
r68 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.985
r69 1 16 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.535 $Y=1.41
+ $X2=2.535 $Y2=1.217
r70 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.535 $Y=1.41
+ $X2=2.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%A 3 5 7 10 12 14 15 20 23 28
c40 15 0 1.68817e-19 $X=4.495 $Y=1.165
r41 23 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.78
+ $Y=1.16 $X2=4.78 $Y2=1.16
r42 20 28 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=4.82 $Y=1.175 $X2=4.78
+ $Y2=1.175
r43 18 19 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=4.37 $Y=1.217
+ $X2=4.395 $Y2=1.217
r44 17 18 63.4586 $w=3.38e-07 $l=4.45e-07 $layer=POLY_cond $X=3.925 $Y=1.217
+ $X2=4.37 $Y2=1.217
r45 16 17 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=3.9 $Y=1.217
+ $X2=3.925 $Y2=1.217
r46 15 23 61.0581 $w=2.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.495 $Y=1.165
+ $X2=4.78 $Y2=1.165
r47 15 19 15.8222 $w=3.38e-07 $l=1.23288e-07 $layer=POLY_cond $X=4.495 $Y=1.165
+ $X2=4.395 $Y2=1.217
r48 12 19 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.217
r49 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.985
r50 8 18 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=1.217
r51 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.37 $Y=1.025
+ $X2=4.37 $Y2=0.56
r52 5 17 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.217
r53 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.985
r54 1 16 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.9 $Y=1.025 $X2=3.9
+ $Y2=1.217
r55 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.9 $Y=1.025 $X2=3.9
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%VPWR 1 2 3 4 5 16 18 22 26 28 32 36 38 40
+ 44 46 51 60 63 66 70
r74 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r75 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r76 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r77 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r78 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r79 55 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r80 55 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r82 52 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.485 $Y2=2.72
r83 52 54 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=4.37 $Y2=2.72
r84 51 69 4.59886 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.802 $Y2=2.72
r85 51 54 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.545 $Y=2.72
+ $X2=4.37 $Y2=2.72
r86 50 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r87 50 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r88 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r89 47 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.22 $Y2=2.72
r90 47 49 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.385 $Y=2.72
+ $X2=2.99 $Y2=2.72
r91 46 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.485 $Y2=2.72
r92 46 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=2.99 $Y2=2.72
r93 44 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 44 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 40 43 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=4.71 $Y=1.66
+ $X2=4.71 $Y2=2.34
r96 38 69 3.16731 $w=3.3e-07 $l=1.27609e-07 $layer=LI1_cond $X=4.71 $Y=2.635
+ $X2=4.802 $Y2=2.72
r97 38 43 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.71 $Y=2.635
+ $X2=4.71 $Y2=2.34
r98 34 66 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=2.635
+ $X2=3.485 $Y2=2.72
r99 34 36 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=3.485 $Y=2.635
+ $X2=3.485 $Y2=2
r100 30 63 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.635
+ $X2=2.22 $Y2=2.72
r101 30 32 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.22 $Y=2.635
+ $X2=2.22 $Y2=2
r102 29 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r103 28 63 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.22 $Y2=2.72
r104 28 29 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r105 24 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r106 24 26 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r107 23 57 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r108 22 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r109 22 23 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r110 18 21 30.7318 $w=2.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.217 $Y=1.66
+ $X2=0.217 $Y2=2.34
r111 16 57 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.172 $Y2=2.72
r112 16 21 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=2.635
+ $X2=0.217 $Y2=2.34
r113 5 43 400 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.485 $X2=4.71 $Y2=2.34
r114 5 40 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=4.485 $Y=1.485
+ $X2=4.71 $Y2=1.66
r115 4 36 300 $w=1.7e-07 $l=6.73201e-07 $layer=licon1_PDIFF $count=2 $X=3.095
+ $Y=1.485 $X2=3.46 $Y2=2
r116 3 32 300 $w=1.7e-07 $l=6.17333e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.22 $Y2=2
r117 2 26 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r118 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r119 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%Y 1 2 3 4 5 16 18 20 24 26 30 34 38 43 44
+ 45 46 47 56
c98 47 0 1.77658e-19 $X=3.8 $Y=1.53
r99 69 70 1.74479 $w=6.03e-07 $l=5e-09 $layer=LI1_cond $X=4.022 $Y=1.66
+ $X2=4.022 $Y2=1.665
r100 54 56 17.0247 $w=2.18e-07 $l=3.25e-07 $layer=LI1_cond $X=2.935 $Y=1.555
+ $X2=3.26 $Y2=1.555
r101 47 69 2.07584 $w=6.03e-07 $l=1.05e-07 $layer=LI1_cond $X=4.022 $Y=1.555
+ $X2=4.022 $Y2=1.66
r102 46 47 6.72176 $w=6.03e-07 $l=3.4e-07 $layer=LI1_cond $X=4.022 $Y=1.19
+ $X2=4.022 $Y2=1.53
r103 46 64 4.31488 $w=6.03e-07 $l=1.35e-07 $layer=LI1_cond $X=4.022 $Y=1.19
+ $X2=4.022 $Y2=1.055
r104 45 47 14.7305 $w=3.88e-07 $l=4.25e-07 $layer=LI1_cond $X=3.295 $Y=1.555
+ $X2=3.72 $Y2=1.555
r105 45 56 1.83343 $w=2.18e-07 $l=3.5e-08 $layer=LI1_cond $X=3.295 $Y=1.555
+ $X2=3.26 $Y2=1.555
r106 44 54 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.745 $Y=1.555
+ $X2=2.935 $Y2=1.555
r107 38 70 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.135 $Y=2.34
+ $X2=4.135 $Y2=1.665
r108 34 64 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.135 $Y=0.72
+ $X2=4.135 $Y2=1.055
r109 28 44 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=2.745 $Y=1.665
+ $X2=2.745 $Y2=1.555
r110 28 30 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.745 $Y=1.665
+ $X2=2.745 $Y2=2.34
r111 27 43 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.555
+ $X2=1.645 $Y2=1.555
r112 26 44 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=2.555 $Y=1.555
+ $X2=2.745 $Y2=1.555
r113 26 27 37.7163 $w=2.18e-07 $l=7.2e-07 $layer=LI1_cond $X=2.555 $Y=1.555
+ $X2=1.835 $Y2=1.555
r114 22 43 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=1.555
r115 22 24 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.645 $Y=1.665
+ $X2=1.645 $Y2=2.34
r116 21 41 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.555
+ $X2=0.705 $Y2=1.555
r117 20 43 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=1.645 $Y2=1.555
r118 20 21 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.555
+ $X2=0.895 $Y2=1.555
r119 16 41 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=1.555
r120 16 18 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.705 $Y=1.665
+ $X2=0.705 $Y2=2.34
r121 5 69 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.485 $X2=4.16 $Y2=1.66
r122 5 38 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.485 $X2=4.16 $Y2=2.34
r123 4 44 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=1.485 $X2=2.77 $Y2=1.66
r124 4 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=1.485 $X2=2.77 $Y2=2.34
r125 3 43 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r126 3 24 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r127 2 41 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r128 2 18 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r129 1 34 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.235 $X2=4.16 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%A_27_47# 1 2 3 12 14 15 16 19 22
c41 14 0 1.79953e-19 $X=0.985 $Y=0.82
r42 20 25 4.17428 $w=2.1e-07 $l=1.5e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=1.135 $Y2=0.36
r43 20 22 46.2121 $w=2.08e-07 $l=8.75e-07 $layer=LI1_cond $X=1.285 $Y=0.36
+ $X2=2.16 $Y2=0.36
r44 17 19 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.135 $Y=0.735
+ $X2=1.135 $Y2=0.72
r45 16 25 2.92199 $w=3e-07 $l=1.05e-07 $layer=LI1_cond $X=1.135 $Y=0.465
+ $X2=1.135 $Y2=0.36
r46 16 19 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=1.135 $Y=0.465
+ $X2=1.135 $Y2=0.72
r47 14 17 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=1.135 $Y2=0.735
r48 14 15 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.82
+ $X2=0.425 $Y2=0.82
r49 10 15 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.425 $Y2=0.82
r50 10 12 12.2125 $w=3.33e-07 $l=3.55e-07 $layer=LI1_cond $X=0.257 $Y=0.735
+ $X2=0.257 $Y2=0.38
r51 3 22 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.16 $Y2=0.38
r52 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r53 2 19 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.72
r54 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%VGND 1 8 10 17 18 21
r54 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r55 17 18 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r56 15 18 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r57 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r58 14 17 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r59 14 15 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r60 12 21 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r61 12 14 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r62 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r63 6 21 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0
r64 6 8 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085 $X2=0.73
+ $Y2=0.38
r65 1 8 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%A_297_47# 1 2 11
c23 11 0 2.63339e-19 $X=3.22 $Y=0.72
r24 8 11 66.1588 $w=2.68e-07 $l=1.55e-06 $layer=LI1_cond $X=1.67 $Y=0.77
+ $X2=3.22 $Y2=0.77
r25 2 11 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.72
r26 1 8 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND4_2%A_511_47# 1 2 3 10 16 18 20 22 25
r34 20 27 2.82476 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=4.71 $Y=0.465
+ $X2=4.71 $Y2=0.36
r35 20 22 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.71 $Y=0.465
+ $X2=4.71 $Y2=0.72
r36 19 25 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.775 $Y=0.36 $X2=3.69
+ $Y2=0.36
r37 18 27 4.43891 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=4.545 $Y=0.36
+ $X2=4.71 $Y2=0.36
r38 18 19 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=4.545 $Y=0.36
+ $X2=3.775 $Y2=0.36
r39 14 25 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=3.69 $Y=0.465
+ $X2=3.69 $Y2=0.36
r40 14 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.69 $Y=0.465
+ $X2=3.69 $Y2=0.72
r41 10 25 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.605 $Y=0.36 $X2=3.69
+ $Y2=0.36
r42 10 12 46.2121 $w=2.08e-07 $l=8.75e-07 $layer=LI1_cond $X=3.605 $Y=0.36
+ $X2=2.73 $Y2=0.36
r43 3 27 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.71 $Y2=0.38
r44 3 22 182 $w=1.7e-07 $l=6.03117e-07 $layer=licon1_NDIFF $count=1 $X=4.445
+ $Y=0.235 $X2=4.71 $Y2=0.72
r45 2 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.69 $Y2=0.38
r46 2 16 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.555
+ $Y=0.235 $X2=3.69 $Y2=0.72
r47 1 12 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.73 $Y2=0.38
.ends

