* File: sky130_fd_sc_hdll__o211ai_2.pxi.spice
* Created: Wed Sep  2 08:42:47 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211AI_2%C1 N_C1_c_68_n N_C1_M1003_g N_C1_c_64_n
+ N_C1_M1007_g N_C1_c_69_n N_C1_M1014_g N_C1_c_65_n N_C1_M1013_g C1 N_C1_c_66_n
+ N_C1_c_67_n PM_SKY130_FD_SC_HDLL__O211AI_2%C1
x_PM_SKY130_FD_SC_HDLL__O211AI_2%B1 N_B1_c_109_n N_B1_M1006_g N_B1_c_105_n
+ N_B1_M1000_g N_B1_c_110_n N_B1_M1015_g N_B1_c_106_n N_B1_M1002_g B1
+ N_B1_c_107_n N_B1_c_108_n B1 PM_SKY130_FD_SC_HDLL__O211AI_2%B1
x_PM_SKY130_FD_SC_HDLL__O211AI_2%A2 N_A2_c_158_n N_A2_M1001_g N_A2_c_154_n
+ N_A2_M1004_g N_A2_c_159_n N_A2_M1008_g N_A2_c_155_n N_A2_M1011_g A2
+ N_A2_c_156_n N_A2_c_157_n A2 PM_SKY130_FD_SC_HDLL__O211AI_2%A2
x_PM_SKY130_FD_SC_HDLL__O211AI_2%A1 N_A1_c_202_n N_A1_M1005_g N_A1_c_197_n
+ N_A1_M1009_g N_A1_c_203_n N_A1_M1012_g N_A1_c_198_n N_A1_M1010_g N_A1_c_199_n
+ A1 N_A1_c_201_n PM_SKY130_FD_SC_HDLL__O211AI_2%A1
x_PM_SKY130_FD_SC_HDLL__O211AI_2%VPWR N_VPWR_M1003_d N_VPWR_M1014_d
+ N_VPWR_M1015_d N_VPWR_M1005_d N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n
+ N_VPWR_c_243_n N_VPWR_c_244_n N_VPWR_c_245_n N_VPWR_c_246_n VPWR
+ N_VPWR_c_247_n N_VPWR_c_248_n N_VPWR_c_249_n N_VPWR_c_239_n N_VPWR_c_251_n
+ N_VPWR_c_252_n PM_SKY130_FD_SC_HDLL__O211AI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O211AI_2%Y N_Y_M1007_s N_Y_M1003_s N_Y_M1006_s
+ N_Y_M1001_d N_Y_c_310_n N_Y_c_311_n N_Y_c_343_n N_Y_c_309_n N_Y_c_312_n
+ N_Y_c_325_n N_Y_c_332_n Y N_Y_c_308_n PM_SKY130_FD_SC_HDLL__O211AI_2%Y
x_PM_SKY130_FD_SC_HDLL__O211AI_2%A_527_297# N_A_527_297#_M1001_s
+ N_A_527_297#_M1008_s N_A_527_297#_M1012_s N_A_527_297#_c_361_n
+ N_A_527_297#_c_358_n N_A_527_297#_c_363_n N_A_527_297#_c_359_n
+ N_A_527_297#_c_360_n PM_SKY130_FD_SC_HDLL__O211AI_2%A_527_297#
x_PM_SKY130_FD_SC_HDLL__O211AI_2%A_27_47# N_A_27_47#_M1007_d N_A_27_47#_M1013_d
+ N_A_27_47#_M1002_s N_A_27_47#_c_387_n N_A_27_47#_c_388_n N_A_27_47#_c_389_n
+ N_A_27_47#_c_412_p PM_SKY130_FD_SC_HDLL__O211AI_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O211AI_2%A_316_47# N_A_316_47#_M1000_d
+ N_A_316_47#_M1004_d N_A_316_47#_M1009_d N_A_316_47#_c_419_n
+ N_A_316_47#_c_431_n PM_SKY130_FD_SC_HDLL__O211AI_2%A_316_47#
x_PM_SKY130_FD_SC_HDLL__O211AI_2%VGND N_VGND_M1004_s N_VGND_M1011_s
+ N_VGND_M1010_s N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n N_VGND_c_454_n
+ N_VGND_c_455_n VGND N_VGND_c_456_n N_VGND_c_457_n N_VGND_c_458_n
+ PM_SKY130_FD_SC_HDLL__O211AI_2%VGND
cc_1 VNB N_C1_c_64_n 0.0220124f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_2 VNB N_C1_c_65_n 0.0173165f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_3 VNB N_C1_c_66_n 0.0161079f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_4 VNB N_C1_c_67_n 0.0619731f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_5 VNB N_B1_c_105_n 0.0173594f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_6 VNB N_B1_c_106_n 0.0225567f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_7 VNB N_B1_c_107_n 0.00675983f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_8 VNB N_B1_c_108_n 0.0466204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A2_c_154_n 0.0227798f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_10 VNB N_A2_c_155_n 0.0168231f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_11 VNB N_A2_c_156_n 0.00707185f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.202
cc_12 VNB N_A2_c_157_n 0.043948f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_13 VNB N_A1_c_197_n 0.0171812f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_14 VNB N_A1_c_198_n 0.0194093f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_15 VNB N_A1_c_199_n 0.00197161f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_16 VNB A1 0.0304127f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_17 VNB N_A1_c_201_n 0.0424259f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VPWR_c_239_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_308_n 0.00104662f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_387_n 0.00871655f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_21 VNB N_A_27_47#_c_388_n 0.00232037f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_22 VNB N_A_27_47#_c_389_n 0.00238482f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.202
cc_23 VNB N_A_316_47#_c_419_n 0.0149027f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.995
cc_24 VNB N_VGND_c_451_n 0.00718344f $X=-0.19 $Y=-0.24 $X2=1.025 $Y2=0.56
cc_25 VNB N_VGND_c_452_n 0.0618103f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.202
cc_26 VNB N_VGND_c_453_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_27 VNB N_VGND_c_454_n 0.00781369f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_28 VNB N_VGND_c_455_n 0.0153474f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_29 VNB N_VGND_c_456_n 0.0147729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_457_n 0.0255559f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_458_n 0.262598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_C1_c_68_n 0.0188939f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_33 VPB N_C1_c_69_n 0.0158156f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_34 VPB N_C1_c_66_n 0.0273111f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_35 VPB N_C1_c_67_n 0.0317635f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.202
cc_36 VPB N_B1_c_109_n 0.0164153f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_37 VPB N_B1_c_110_n 0.0200756f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_38 VPB N_B1_c_107_n 0.00673895f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_39 VPB N_B1_c_108_n 0.0243823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A2_c_158_n 0.0211704f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_41 VPB N_A2_c_159_n 0.0166059f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_42 VPB N_A2_c_156_n 0.00780287f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.202
cc_43 VPB N_A2_c_157_n 0.023657f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.202
cc_44 VPB N_A1_c_202_n 0.0161826f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_45 VPB N_A1_c_203_n 0.0210264f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.41
cc_46 VPB N_A1_c_201_n 0.0242013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_240_n 0.0107363f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.445
cc_48 VPB N_VPWR_c_241_n 0.0165871f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.202
cc_49 VPB N_VPWR_c_242_n 3.36964e-19 $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.202
cc_50 VPB N_VPWR_c_243_n 0.00962827f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_244_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_245_n 0.0386828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_246_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_247_n 0.0165388f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_248_n 0.0145309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_249_n 0.0207856f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_239_n 0.0587379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_251_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_252_n 0.00583344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_Y_c_309_n 0.0214284f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_527_297#_c_358_n 0.00759381f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_62 VPB N_A_527_297#_c_359_n 0.0292274f $X=-0.19 $Y=1.305 $X2=1 $Y2=1.202
cc_63 VPB N_A_527_297#_c_360_n 0.00429005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 N_C1_c_69_n N_B1_c_109_n 0.0219165f $X=1 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_65 N_C1_c_65_n N_B1_c_105_n 0.0096399f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_66 N_C1_c_67_n N_B1_c_107_n 0.00277095f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_67 N_C1_c_67_n N_B1_c_108_n 0.0266003f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_68 N_C1_c_66_n N_VPWR_M1003_d 0.00796434f $X=0.24 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_69 N_C1_c_66_n N_VPWR_c_240_n 4.72765e-19 $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_70 N_C1_c_68_n N_VPWR_c_241_n 0.003211f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_71 N_C1_c_66_n N_VPWR_c_241_n 0.0190991f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_72 N_C1_c_68_n N_VPWR_c_242_n 6.9258e-19 $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C1_c_69_n N_VPWR_c_242_n 0.0141023f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C1_c_68_n N_VPWR_c_247_n 0.00605302f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C1_c_69_n N_VPWR_c_247_n 0.00447018f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_76 N_C1_c_68_n N_VPWR_c_239_n 0.0111262f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_77 N_C1_c_69_n N_VPWR_c_239_n 0.00766229f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_78 N_C1_c_66_n N_VPWR_c_239_n 0.00201653f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C1_c_68_n N_Y_c_310_n 0.0187821f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_80 N_C1_c_69_n N_Y_c_311_n 0.0173162f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_81 N_C1_c_68_n N_Y_c_312_n 0.00349845f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_82 N_C1_c_69_n N_Y_c_312_n 0.00198297f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_83 N_C1_c_68_n N_Y_c_308_n 0.00344488f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_84 N_C1_c_64_n N_Y_c_308_n 0.017999f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_85 N_C1_c_69_n N_Y_c_308_n 0.00402639f $X=1 $Y=1.41 $X2=0 $Y2=0
cc_86 N_C1_c_65_n N_Y_c_308_n 0.00314807f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_87 N_C1_c_66_n N_Y_c_308_n 0.0394462f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C1_c_67_n N_Y_c_308_n 0.0357707f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_89 N_C1_c_64_n N_A_27_47#_c_387_n 0.0110269f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_c_65_n N_A_27_47#_c_387_n 0.0131648f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_91 N_C1_c_66_n N_A_27_47#_c_387_n 0.00888263f $X=0.24 $Y=1.16 $X2=0 $Y2=0
cc_92 N_C1_c_67_n N_A_27_47#_c_387_n 0.00385336f $X=1 $Y=1.202 $X2=0 $Y2=0
cc_93 N_C1_c_64_n N_VGND_c_452_n 0.00357877f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_94 N_C1_c_65_n N_VGND_c_452_n 0.00357877f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_95 N_C1_c_64_n N_VGND_c_458_n 0.00640069f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_96 N_C1_c_65_n N_VGND_c_458_n 0.0055497f $X=1.025 $Y=0.995 $X2=0 $Y2=0
cc_97 N_B1_c_107_n N_A2_c_156_n 0.0130201f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_98 N_B1_c_108_n N_A2_c_156_n 0.00147293f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_99 N_B1_c_107_n N_A2_c_157_n 0.00155656f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_100 N_B1_c_109_n N_VPWR_c_242_n 0.0104414f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B1_c_110_n N_VPWR_c_242_n 5.87114e-19 $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B1_c_109_n N_VPWR_c_243_n 6.23977e-19 $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B1_c_110_n N_VPWR_c_243_n 0.0149753f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B1_c_109_n N_VPWR_c_248_n 0.00642146f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B1_c_110_n N_VPWR_c_248_n 0.00447018f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B1_c_109_n N_VPWR_c_239_n 0.0107337f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_VPWR_c_239_n 0.00766229f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B1_c_109_n N_Y_c_311_n 0.0163127f $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B1_c_107_n N_Y_c_311_n 0.0257426f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_110 N_B1_c_108_n N_Y_c_311_n 3.43217e-19 $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_111 N_B1_c_110_n N_Y_c_309_n 0.0168398f $X=1.96 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B1_c_107_n N_Y_c_309_n 0.0246095f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_113 N_B1_c_107_n N_Y_c_325_n 0.0157997f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_108_n N_Y_c_325_n 0.0013343f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_115 N_B1_c_109_n N_Y_c_308_n 5.88217e-19 $X=1.48 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B1_c_107_n N_Y_c_308_n 0.016464f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_c_108_n N_Y_c_308_n 8.77378e-19 $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_118 N_B1_c_105_n N_A_27_47#_c_388_n 0.00473388f $X=1.505 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B1_c_107_n N_A_27_47#_c_388_n 0.00967171f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B1_c_108_n N_A_27_47#_c_388_n 6.09178e-19 $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_121 N_B1_c_105_n N_A_27_47#_c_389_n 0.0101363f $X=1.505 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B1_c_106_n N_A_27_47#_c_389_n 0.00910135f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B1_c_107_n N_A_27_47#_c_389_n 0.00360235f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_124 N_B1_c_108_n N_A_27_47#_c_389_n 0.00157298f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_125 N_B1_c_105_n N_A_316_47#_c_419_n 0.0050364f $X=1.505 $Y=0.995 $X2=0 $Y2=0
cc_126 N_B1_c_106_n N_A_316_47#_c_419_n 0.01238f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B1_c_107_n N_A_316_47#_c_419_n 0.0363906f $X=1.835 $Y=1.16 $X2=0 $Y2=0
cc_128 N_B1_c_108_n N_A_316_47#_c_419_n 0.00357425f $X=1.96 $Y=1.202 $X2=0 $Y2=0
cc_129 N_B1_c_106_n N_VGND_c_451_n 0.00219146f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B1_c_105_n N_VGND_c_452_n 0.00357877f $X=1.505 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_c_106_n N_VGND_c_452_n 0.00357877f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B1_c_105_n N_VGND_c_458_n 0.0055497f $X=1.505 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B1_c_106_n N_VGND_c_458_n 0.00670797f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A2_c_159_n N_A1_c_202_n 0.0183326f $X=3.48 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_135 N_A2_c_155_n N_A1_c_197_n 0.0244776f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A2_c_156_n N_A1_c_199_n 0.0203733f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A2_c_157_n N_A1_c_199_n 7.6318e-19 $X=3.48 $Y=1.202 $X2=0 $Y2=0
cc_138 N_A2_c_156_n N_A1_c_201_n 0.00237275f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A2_c_157_n N_A1_c_201_n 0.024989f $X=3.48 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A2_c_158_n N_VPWR_c_243_n 0.0055638f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A2_c_159_n N_VPWR_c_244_n 0.00108143f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_158_n N_VPWR_c_245_n 0.00429453f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A2_c_159_n N_VPWR_c_245_n 0.00429453f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_158_n N_VPWR_c_239_n 0.0073737f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_159_n N_VPWR_c_239_n 0.00614026f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_158_n N_Y_c_309_n 0.0105713f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A2_c_156_n N_Y_c_309_n 0.0229267f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A2_c_158_n N_Y_c_332_n 0.0176943f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A2_c_159_n N_Y_c_332_n 0.00700328f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A2_c_156_n N_Y_c_332_n 0.0248542f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A2_c_157_n N_Y_c_332_n 0.00171303f $X=3.48 $Y=1.202 $X2=0 $Y2=0
cc_152 N_A2_c_158_n N_A_527_297#_c_361_n 0.0104438f $X=3 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A2_c_159_n N_A_527_297#_c_361_n 0.0139438f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_156_n N_A_527_297#_c_363_n 7.66876e-19 $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A2_c_154_n N_A_316_47#_c_419_n 0.0137547f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A2_c_155_n N_A_316_47#_c_419_n 0.0137174f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A2_c_156_n N_A_316_47#_c_419_n 0.0509228f $X=3.42 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A2_c_157_n N_A_316_47#_c_419_n 0.00416996f $X=3.48 $Y=1.202 $X2=0 $Y2=0
cc_159 N_A2_c_154_n N_VGND_c_451_n 0.00332888f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_154_n N_VGND_c_454_n 0.00119077f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_155_n N_VGND_c_454_n 0.011111f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_154_n N_VGND_c_455_n 0.00425094f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_155_n N_VGND_c_455_n 0.00198377f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_154_n N_VGND_c_458_n 0.00719146f $X=3.025 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A2_c_155_n N_VGND_c_458_n 0.00285026f $X=3.53 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_202_n N_VPWR_c_244_n 0.0156078f $X=3.96 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A1_c_203_n N_VPWR_c_244_n 0.0127915f $X=4.44 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A1_c_202_n N_VPWR_c_245_n 0.00447018f $X=3.96 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A1_c_203_n N_VPWR_c_249_n 0.00642146f $X=4.44 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A1_c_202_n N_VPWR_c_239_n 0.00768581f $X=3.96 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A1_c_203_n N_VPWR_c_239_n 0.0117169f $X=4.44 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A1_c_202_n N_A_527_297#_c_358_n 0.0148511f $X=3.96 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A1_c_203_n N_A_527_297#_c_358_n 0.0188f $X=4.44 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A1_c_199_n N_A_527_297#_c_358_n 0.0313358f $X=4.465 $Y=1.185 $X2=0
+ $Y2=0
cc_175 A1 N_A_527_297#_c_358_n 0.0245103f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_176 N_A1_c_201_n N_A_527_297#_c_358_n 0.00646734f $X=4.44 $Y=1.202 $X2=0
+ $Y2=0
cc_177 N_A1_c_199_n N_A_527_297#_c_363_n 6.04866e-19 $X=4.465 $Y=1.185 $X2=0
+ $Y2=0
cc_178 N_A1_c_197_n N_A_316_47#_c_419_n 0.0113482f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A1_c_199_n N_A_316_47#_c_419_n 0.0139644f $X=4.465 $Y=1.185 $X2=0 $Y2=0
cc_180 N_A1_c_201_n N_A_316_47#_c_419_n 0.0017792f $X=4.44 $Y=1.202 $X2=0 $Y2=0
cc_181 N_A1_c_199_n N_A_316_47#_c_431_n 0.0109257f $X=4.465 $Y=1.185 $X2=0 $Y2=0
cc_182 A1 N_A_316_47#_c_431_n 0.00610165f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_183 N_A1_c_201_n N_A_316_47#_c_431_n 0.00348404f $X=4.44 $Y=1.202 $X2=0 $Y2=0
cc_184 A1 N_VGND_M1010_s 0.00438531f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_185 N_A1_c_197_n N_VGND_c_454_n 0.00167049f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A1_c_197_n N_VGND_c_456_n 0.00425094f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A1_c_198_n N_VGND_c_456_n 0.00271402f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A1_c_197_n N_VGND_c_457_n 0.00118155f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A1_c_198_n N_VGND_c_457_n 0.0125297f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_190 A1 N_VGND_c_457_n 0.0170368f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_191 N_A1_c_197_n N_VGND_c_458_n 0.00587843f $X=3.985 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A1_c_198_n N_VGND_c_458_n 0.00509204f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_193 A1 N_VGND_c_458_n 0.00336628f $X=4.685 $Y=0.765 $X2=0 $Y2=0
cc_194 N_VPWR_c_239_n N_Y_M1003_s 0.00430227f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_195 N_VPWR_c_239_n N_Y_M1006_s 0.00621163f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_196 N_VPWR_c_239_n N_Y_M1001_d 0.00240926f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_197 N_VPWR_c_247_n N_Y_c_310_n 0.0194684f $X=1.025 $Y=2.72 $X2=0 $Y2=0
cc_198 N_VPWR_c_239_n N_Y_c_310_n 0.0114913f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_199 N_VPWR_M1014_d N_Y_c_311_n 0.00477701f $X=1.09 $Y=1.485 $X2=0 $Y2=0
cc_200 N_VPWR_c_242_n N_Y_c_311_n 0.0182017f $X=1.24 $Y=2 $X2=0 $Y2=0
cc_201 N_VPWR_c_248_n N_Y_c_343_n 0.0131506f $X=1.985 $Y=2.72 $X2=0 $Y2=0
cc_202 N_VPWR_c_239_n N_Y_c_343_n 0.00722976f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_203 N_VPWR_M1015_d N_Y_c_309_n 0.00889266f $X=2.05 $Y=1.485 $X2=0 $Y2=0
cc_204 N_VPWR_c_243_n N_Y_c_309_n 0.0224717f $X=2.2 $Y=2 $X2=0 $Y2=0
cc_205 N_VPWR_c_243_n N_Y_c_332_n 0.00533309f $X=2.2 $Y=2 $X2=0 $Y2=0
cc_206 N_VPWR_c_239_n N_A_527_297#_M1001_s 0.00220818f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_207 N_VPWR_c_239_n N_A_527_297#_M1008_s 0.00426761f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_239_n N_A_527_297#_M1012_s 0.00412552f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_245_n N_A_527_297#_c_361_n 0.055006f $X=3.985 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_239_n N_A_527_297#_c_361_n 0.0341944f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_M1005_d N_A_527_297#_c_358_n 0.00374937f $X=4.05 $Y=1.485 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_244_n N_A_527_297#_c_358_n 0.0209901f $X=4.2 $Y=1.95 $X2=0 $Y2=0
cc_213 N_VPWR_c_249_n N_A_527_297#_c_359_n 0.0181615f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_214 N_VPWR_c_239_n N_A_527_297#_c_359_n 0.00993081f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_215 N_VPWR_c_243_n N_A_527_297#_c_360_n 0.0244369f $X=2.2 $Y=2 $X2=0 $Y2=0
cc_216 N_VPWR_c_245_n N_A_527_297#_c_360_n 0.0173659f $X=3.985 $Y=2.72 $X2=0
+ $Y2=0
cc_217 N_VPWR_c_239_n N_A_527_297#_c_360_n 0.00977772f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_218 N_Y_c_309_n N_A_527_297#_M1001_s 0.00768619f $X=3.025 $Y=1.625 $X2=-0.19
+ $Y2=-0.24
cc_219 N_Y_M1001_d N_A_527_297#_c_361_n 0.00372414f $X=3.09 $Y=1.485 $X2=0 $Y2=0
cc_220 N_Y_c_309_n N_A_527_297#_c_361_n 0.00278684f $X=3.025 $Y=1.625 $X2=0
+ $Y2=0
cc_221 N_Y_c_332_n N_A_527_297#_c_361_n 0.0194343f $X=3.24 $Y=1.7 $X2=0 $Y2=0
cc_222 N_Y_c_309_n N_A_527_297#_c_360_n 0.0108975f $X=3.025 $Y=1.625 $X2=0 $Y2=0
cc_223 N_Y_M1007_s N_A_27_47#_c_387_n 0.00445202f $X=0.62 $Y=0.235 $X2=0 $Y2=0
cc_224 N_Y_c_308_n N_A_27_47#_c_387_n 0.017214f $X=0.76 $Y=0.76 $X2=0 $Y2=0
cc_225 N_Y_c_311_n N_A_27_47#_c_388_n 0.00214885f $X=1.625 $Y=1.625 $X2=0 $Y2=0
cc_226 N_Y_c_308_n N_A_27_47#_c_388_n 2.69592e-19 $X=0.76 $Y=0.76 $X2=0 $Y2=0
cc_227 N_Y_M1007_s N_VGND_c_458_n 0.00265018f $X=0.62 $Y=0.235 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_389_n N_A_316_47#_M1000_d 0.00419293f $X=2.2 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_229 N_A_27_47#_M1002_s N_A_316_47#_c_419_n 0.00998507f $X=2.06 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_27_47#_c_388_n N_A_316_47#_c_419_n 0.0164761f $X=1.24 $Y=0.705 $X2=0
+ $Y2=0
cc_231 N_A_27_47#_c_389_n N_A_316_47#_c_419_n 0.0479183f $X=2.2 $Y=0.36 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_c_389_n N_VGND_c_451_n 0.013521f $X=2.2 $Y=0.36 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_387_n N_VGND_c_452_n 0.060302f $X=1.145 $Y=0.35 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_389_n N_VGND_c_452_n 0.0589721f $X=2.2 $Y=0.36 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_412_p N_VGND_c_452_n 0.0128805f $X=1.24 $Y=0.36 $X2=0 $Y2=0
cc_236 N_A_27_47#_M1007_d N_VGND_c_458_n 0.00270836f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_M1013_d N_VGND_c_458_n 0.00263394f $X=1.1 $Y=0.235 $X2=0 $Y2=0
cc_238 N_A_27_47#_M1002_s N_VGND_c_458_n 0.00229841f $X=2.06 $Y=0.235 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_c_387_n N_VGND_c_458_n 0.0376909f $X=1.145 $Y=0.35 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_389_n N_VGND_c_458_n 0.0370265f $X=2.2 $Y=0.36 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_412_p N_VGND_c_458_n 0.00730424f $X=1.24 $Y=0.36 $X2=0 $Y2=0
cc_242 N_A_316_47#_c_419_n N_VGND_M1004_s 0.00966312f $X=4.105 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_316_47#_c_419_n N_VGND_M1011_s 0.00819164f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_244 N_A_316_47#_c_419_n N_VGND_c_451_n 0.0208531f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_245 N_A_316_47#_c_419_n N_VGND_c_452_n 0.00425741f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_246 N_A_316_47#_c_419_n N_VGND_c_454_n 0.0184819f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_247 N_A_316_47#_c_419_n N_VGND_c_455_n 0.00926951f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_248 N_A_316_47#_c_419_n N_VGND_c_456_n 0.00296958f $X=4.105 $Y=0.74 $X2=0
+ $Y2=0
cc_249 N_A_316_47#_c_431_n N_VGND_c_456_n 0.00447217f $X=4.2 $Y=0.68 $X2=0 $Y2=0
cc_250 N_A_316_47#_M1000_d N_VGND_c_458_n 0.00265018f $X=1.58 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_A_316_47#_M1004_d N_VGND_c_458_n 0.00417027f $X=3.1 $Y=0.235 $X2=0
+ $Y2=0
cc_252 N_A_316_47#_M1009_d N_VGND_c_458_n 0.00674911f $X=4.06 $Y=0.235 $X2=0
+ $Y2=0
cc_253 N_A_316_47#_c_419_n N_VGND_c_458_n 0.032503f $X=4.105 $Y=0.74 $X2=0 $Y2=0
cc_254 N_A_316_47#_c_431_n N_VGND_c_458_n 0.00598996f $X=4.2 $Y=0.68 $X2=0 $Y2=0
