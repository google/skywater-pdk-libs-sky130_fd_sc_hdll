* File: sky130_fd_sc_hdll__xnor2_2.pex.spice
* Created: Wed Sep  2 08:53:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 31 33 34 36 39 40 41 46 51 55
c116 31 0 1.89108e-19 $X=0.925 $Y=1.445
c117 10 0 9.37715e-20 $X=1.005 $Y=0.995
r118 51 52 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=4.395 $Y=1.202
+ $X2=4.42 $Y2=1.202
r119 48 49 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=3.865 $Y=1.202
+ $X2=3.89 $Y2=1.202
r120 46 47 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.005 $Y2=1.202
r121 43 44 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.485 $Y=1.202
+ $X2=0.51 $Y2=1.202
r122 41 55 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=1.145 $Y=1.53
+ $X2=1.15 $Y2=1.53
r123 40 55 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=3.18 $Y=1.53
+ $X2=1.15 $Y2=1.53
r124 39 41 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.01 $Y=1.53
+ $X2=1.145 $Y2=1.53
r125 37 51 36.9788 $w=3.78e-07 $l=2.9e-07 $layer=POLY_cond $X=4.105 $Y=1.202
+ $X2=4.395 $Y2=1.202
r126 37 49 27.4153 $w=3.78e-07 $l=2.15e-07 $layer=POLY_cond $X=4.105 $Y=1.202
+ $X2=3.89 $Y2=1.202
r127 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.16 $X2=4.105 $Y2=1.16
r128 34 36 39.8745 $w=2.08e-07 $l=7.55e-07 $layer=LI1_cond $X=3.35 $Y=1.18
+ $X2=4.105 $Y2=1.18
r129 33 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.265 $Y=1.445
+ $X2=3.18 $Y2=1.53
r130 32 34 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.265 $Y=1.285
+ $X2=3.35 $Y2=1.18
r131 32 33 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.265 $Y=1.285
+ $X2=3.265 $Y2=1.445
r132 31 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.925 $Y=1.445
+ $X2=1.01 $Y2=1.53
r133 30 31 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=0.925 $Y=1.285
+ $X2=0.925 $Y2=1.445
r134 28 46 35.5158 $w=3.8e-07 $l=2.8e-07 $layer=POLY_cond $X=0.7 $Y=1.202
+ $X2=0.98 $Y2=1.202
r135 28 44 24.1 $w=3.8e-07 $l=1.9e-07 $layer=POLY_cond $X=0.7 $Y=1.202 $X2=0.51
+ $Y2=1.202
r136 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.7
+ $Y=1.16 $X2=0.7 $Y2=1.16
r137 25 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=0.84 $Y=1.18
+ $X2=0.925 $Y2=1.285
r138 25 27 7.39394 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=0.84 $Y=1.18
+ $X2=0.7 $Y2=1.18
r139 22 52 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.42 $Y=0.995
+ $X2=4.42 $Y2=1.202
r140 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.42 $Y=0.995
+ $X2=4.42 $Y2=0.56
r141 19 51 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.202
r142 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.395 $Y=1.41
+ $X2=4.395 $Y2=1.985
r143 16 49 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.89 $Y=1.41
+ $X2=3.89 $Y2=1.202
r144 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.89 $Y=1.41
+ $X2=3.89 $Y2=1.985
r145 13 48 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.865 $Y=0.995
+ $X2=3.865 $Y2=1.202
r146 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.865 $Y=0.995
+ $X2=3.865 $Y2=0.56
r147 10 47 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r148 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r149 7 46 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r150 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r151 4 44 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r152 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.985
r153 1 43 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.202
r154 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 28 30 32 40
c93 19 0 1.33039e-19 $X=3.42 $Y=1.41
c94 4 0 1.89108e-19 $X=1.45 $Y=1.41
r95 41 42 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.895 $Y=1.202
+ $X2=1.92 $Y2=1.202
r96 39 41 47.5658 $w=3.8e-07 $l=3.75e-07 $layer=POLY_cond $X=1.52 $Y=1.202
+ $X2=1.895 $Y2=1.202
r97 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.52
+ $Y=1.16 $X2=1.52 $Y2=1.16
r98 37 39 8.87895 $w=3.8e-07 $l=7e-08 $layer=POLY_cond $X=1.45 $Y=1.202 $X2=1.52
+ $Y2=1.202
r99 36 37 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.425 $Y=1.202
+ $X2=1.45 $Y2=1.202
r100 34 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.66
+ $Y=1.16 $X2=2.66 $Y2=1.16
r101 32 42 13.6483 $w=3.8e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=1.92 $Y2=1.202
r102 32 34 111.911 $w=3.3e-07 $l=6.4e-07 $layer=POLY_cond $X=2.02 $Y=1.16
+ $X2=2.66 $Y2=1.16
r103 30 40 0.236129 $w=1.548e-06 $l=3e-08 $layer=LI1_cond $X=2.13 $Y=1.19
+ $X2=2.13 $Y2=1.16
r104 28 29 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.42 $Y=1.202
+ $X2=3.445 $Y2=1.202
r105 27 28 59.6158 $w=3.8e-07 $l=4.7e-07 $layer=POLY_cond $X=2.95 $Y=1.202
+ $X2=3.42 $Y2=1.202
r106 26 27 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.925 $Y=1.202
+ $X2=2.95 $Y2=1.202
r107 25 34 33.2236 $w=3.3e-07 $l=1.9e-07 $layer=POLY_cond $X=2.85 $Y=1.16
+ $X2=2.66 $Y2=1.16
r108 25 26 10.4773 $w=3.8e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.85 $Y=1.16
+ $X2=2.925 $Y2=1.202
r109 22 29 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=1.202
r110 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=0.56
r111 19 28 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.202
r112 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.42 $Y=1.41
+ $X2=3.42 $Y2=1.985
r113 16 27 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.95 $Y2=1.202
r114 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.95 $Y2=1.985
r115 13 26 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.925 $Y=0.995
+ $X2=2.925 $Y2=1.202
r116 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.925 $Y=0.995
+ $X2=2.925 $Y2=0.56
r117 10 42 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.202
r118 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.985
r119 7 41 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=1.202
r120 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.895 $Y=0.995
+ $X2=1.895 $Y2=0.56
r121 4 37 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.202
r122 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.985
r123 1 36 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=1.202
r124 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.425 $Y=0.995
+ $X2=1.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_297# 1 2 3 4 13 15 16 18 19 21 22 24
+ 26 29 31 33 37 41 44 45 46 48 49 51 55 57 59 63
c140 31 0 9.37715e-20 $X=0.745 $Y=0.73
c141 22 0 6.40318e-20 $X=5.88 $Y=0.995
r142 63 64 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.855 $Y=1.202
+ $X2=5.88 $Y2=1.202
r143 60 61 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.36 $Y=1.202
+ $X2=5.385 $Y2=1.202
r144 52 63 34.8816 $w=3.8e-07 $l=2.75e-07 $layer=POLY_cond $X=5.58 $Y=1.202
+ $X2=5.855 $Y2=1.202
r145 52 61 24.7342 $w=3.8e-07 $l=1.95e-07 $layer=POLY_cond $X=5.58 $Y=1.202
+ $X2=5.385 $Y2=1.202
r146 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.58
+ $Y=1.16 $X2=5.58 $Y2=1.16
r147 49 51 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.205 $Y=1.16
+ $X2=5.58 $Y2=1.16
r148 47 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.12 $Y=1.245
+ $X2=5.205 $Y2=1.16
r149 47 48 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.12 $Y=1.245
+ $X2=5.12 $Y2=1.455
r150 45 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.035 $Y=1.54
+ $X2=5.12 $Y2=1.455
r151 45 46 81.877 $w=1.68e-07 $l=1.255e-06 $layer=LI1_cond $X=5.035 $Y=1.54
+ $X2=3.78 $Y2=1.54
r152 43 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.695 $Y=1.625
+ $X2=3.78 $Y2=1.54
r153 43 44 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.695 $Y=1.625
+ $X2=3.695 $Y2=1.785
r154 42 59 6.87424 $w=1.75e-07 $l=1.27475e-07 $layer=LI1_cond $X=2.28 $Y=1.87
+ $X2=2.155 $Y2=1.875
r155 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.61 $Y=1.87
+ $X2=3.695 $Y2=1.785
r156 41 42 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=3.61 $Y=1.87
+ $X2=2.28 $Y2=1.87
r157 38 57 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=1.875
+ $X2=1.215 $Y2=1.875
r158 37 59 6.87424 $w=1.75e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=1.875
+ $X2=2.155 $Y2=1.875
r159 37 38 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=2.03 $Y=1.875
+ $X2=1.34 $Y2=1.875
r160 34 55 2.8704 $w=1.8e-07 $l=1.58e-07 $layer=LI1_cond $X=0.4 $Y=1.875
+ $X2=0.242 $Y2=1.875
r161 33 57 6.72674 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.09 $Y=1.875
+ $X2=1.215 $Y2=1.875
r162 33 34 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=1.09 $Y=1.875
+ $X2=0.4 $Y2=1.875
r163 29 31 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=0.315 $Y=0.77
+ $X2=0.745 $Y2=0.77
r164 26 55 3.61314 $w=2.72e-07 $l=1.08995e-07 $layer=LI1_cond $X=0.2 $Y=1.785
+ $X2=0.242 $Y2=1.875
r165 25 29 6.8319 $w=2.5e-07 $l=1.73205e-07 $layer=LI1_cond $X=0.2 $Y=0.895
+ $X2=0.315 $Y2=0.77
r166 25 26 44.5945 $w=2.28e-07 $l=8.9e-07 $layer=LI1_cond $X=0.2 $Y=0.895
+ $X2=0.2 $Y2=1.785
r167 22 64 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.88 $Y=0.995
+ $X2=5.88 $Y2=1.202
r168 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.88 $Y=0.995
+ $X2=5.88 $Y2=0.56
r169 19 63 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.855 $Y=1.41
+ $X2=5.855 $Y2=1.202
r170 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.855 $Y=1.41
+ $X2=5.855 $Y2=1.985
r171 16 61 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.385 $Y=1.41
+ $X2=5.385 $Y2=1.202
r172 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.385 $Y=1.41
+ $X2=5.385 $Y2=1.985
r173 13 60 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.36 $Y2=1.202
r174 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.36 $Y=0.995
+ $X2=5.36 $Y2=0.56
r175 4 59 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.01
+ $Y=1.485 $X2=2.155 $Y2=1.96
r176 3 57 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.215 $Y2=1.96
r177 2 55 300 $w=1.7e-07 $l=5.40486e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.96
r178 1 31 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=0.56
+ $Y=0.235 $X2=0.745 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%VPWR 1 2 3 4 5 20 22 26 30 34 36 38 41 42
+ 44 45 46 61 66 69 73
c105 44 0 1.96631e-19 $X=5.025 $Y=2.72
r106 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r107 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r108 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r109 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r110 64 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r112 61 72 5.19438 $w=1.7e-07 $l=2.37e-07 $layer=LI1_cond $X=5.965 $Y=2.72
+ $X2=6.202 $Y2=2.72
r113 61 63 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.965 $Y=2.72
+ $X2=5.75 $Y2=2.72
r114 60 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r115 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r116 57 60 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 56 59 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=4.83 $Y2=2.72
r118 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r119 54 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r120 53 54 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r121 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r122 51 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r123 50 53 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r124 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r125 48 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=1.685 $Y2=2.72
r126 48 50 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.81 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 46 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 44 59 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.025 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 44 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.025 $Y=2.72
+ $X2=5.15 $Y2=2.72
r130 43 63 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=5.75 $Y2=2.72
r131 43 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=5.15 $Y2=2.72
r132 41 53 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=2.72 $X2=2.99
+ $Y2=2.72
r133 41 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=3.185 $Y2=2.72
r134 40 56 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=3.45 $Y2=2.72
r135 40 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.31 $Y=2.72
+ $X2=3.185 $Y2=2.72
r136 36 72 2.95882 $w=3.75e-07 $l=1.07121e-07 $layer=LI1_cond $X=6.152 $Y=2.635
+ $X2=6.202 $Y2=2.72
r137 36 38 20.744 $w=3.73e-07 $l=6.75e-07 $layer=LI1_cond $X=6.152 $Y=2.635
+ $X2=6.152 $Y2=1.96
r138 32 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.15 $Y=2.635
+ $X2=5.15 $Y2=2.72
r139 32 34 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.15 $Y=2.635
+ $X2=5.15 $Y2=2.3
r140 28 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=2.635
+ $X2=3.185 $Y2=2.72
r141 28 30 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.185 $Y=2.635
+ $X2=3.185 $Y2=2.3
r142 24 69 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=2.635
+ $X2=1.685 $Y2=2.72
r143 24 26 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.685 $Y=2.635
+ $X2=1.685 $Y2=2.3
r144 23 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.745 $Y2=2.72
r145 22 69 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=1.685 $Y2=2.72
r146 22 23 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.56 $Y=2.72
+ $X2=0.87 $Y2=2.72
r147 18 66 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r148 18 20 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.3
r149 5 38 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.945
+ $Y=1.485 $X2=6.09 $Y2=1.96
r150 4 34 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=5.025
+ $Y=1.485 $X2=5.15 $Y2=2.3
r151 3 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.185 $Y2=2.3
r152 2 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.485 $X2=1.685 $Y2=2.3
r153 1 20 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.745 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%A_514_297# 1 2 3 10 13 17 18 21 24 25
c56 24 0 1.96631e-19 $X=3.77 $Y=2.21
c57 18 0 1.33039e-19 $X=2.895 $Y=2.21
r58 25 34 6.02816 $w=3.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.692 $Y=2.21
+ $X2=3.692 $Y2=2.38
r59 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.77 $Y=2.21
+ $X2=3.77 $Y2=2.21
r60 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.75 $Y=2.21
+ $X2=2.75 $Y2=2.21
r61 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.895 $Y=2.21
+ $X2=2.75 $Y2=2.21
r62 17 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.625 $Y=2.21
+ $X2=3.77 $Y2=2.21
r63 17 18 0.903464 $w=1.4e-07 $l=7.3e-07 $layer=MET1_cond $X=3.625 $Y=2.21
+ $X2=2.895 $Y2=2.21
r64 13 15 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.63 $Y=2.3 $X2=4.63
+ $Y2=2.38
r65 11 34 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=3.855 $Y=2.38
+ $X2=3.692 $Y2=2.38
r66 10 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.505 $Y=2.38
+ $X2=4.63 $Y2=2.38
r67 10 11 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.505 $Y=2.38
+ $X2=3.855 $Y2=2.38
r68 3 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.485
+ $Y=1.485 $X2=4.63 $Y2=2.3
r69 2 25 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.51
+ $Y=1.485 $X2=3.655 $Y2=2.3
r70 1 21 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.57
+ $Y=1.485 $X2=2.715 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%Y 1 2 3 4 13 15 20 21 22 23 32
c55 21 0 6.40318e-20 $X=6.145 $Y=0.475
r56 23 26 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=4.18 $Y=1.88 $X2=4.18
+ $Y2=1.96
r57 22 32 2.64069 $w=2.08e-07 $l=5e-08 $layer=LI1_cond $X=6.145 $Y=1.52
+ $X2=6.195 $Y2=1.52
r58 22 35 27.7273 $w=2.08e-07 $l=5.25e-07 $layer=LI1_cond $X=6.145 $Y=1.52
+ $X2=5.62 $Y2=1.52
r59 21 31 2.51472 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=6.145 $Y=0.475
+ $X2=6.145 $Y2=0.39
r60 21 22 27.7768 $w=3.88e-07 $l=9.4e-07 $layer=LI1_cond $X=6.145 $Y=0.475
+ $X2=6.145 $Y2=1.415
r61 20 29 3.18546 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.62 $Y=1.795
+ $X2=5.62 $Y2=1.96
r62 20 35 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=5.62 $Y=1.795
+ $X2=5.62 $Y2=1.625
r63 15 31 5.76906 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.95 $Y=0.39
+ $X2=6.145 $Y2=0.39
r64 15 17 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=5.95 $Y=0.39 $X2=5.15
+ $Y2=0.39
r65 14 23 1.9771 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=4.285 $Y=1.88
+ $X2=4.18 $Y2=1.88
r66 13 29 3.9577 $w=1.7e-07 $l=1.60078e-07 $layer=LI1_cond $X=5.495 $Y=1.88
+ $X2=5.62 $Y2=1.96
r67 13 14 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=5.495 $Y=1.88
+ $X2=4.285 $Y2=1.88
r68 4 35 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.485 $X2=5.62 $Y2=1.62
r69 4 29 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=5.475
+ $Y=1.485 $X2=5.62 $Y2=1.96
r70 3 26 600 $w=1.7e-07 $l=5.57786e-07 $layer=licon1_PDIFF $count=1 $X=3.98
+ $Y=1.485 $X2=4.16 $Y2=1.96
r71 2 31 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.955
+ $Y=0.235 $X2=6.09 $Y2=0.39
r72 1 17 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.025
+ $Y=0.235 $X2=5.15 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%A_27_47# 1 2 3 10 14 15 16 20
r44 18 20 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.13 $Y=0.725
+ $X2=2.13 $Y2=0.39
r45 17 25 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.38 $Y=0.815
+ $X2=1.255 $Y2=0.815
r46 16 18 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=1.94 $Y=0.815
+ $X2=2.13 $Y2=0.725
r47 16 17 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.94 $Y=0.815
+ $X2=1.38 $Y2=0.815
r48 15 25 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=1.255 $Y=0.725
+ $X2=1.255 $Y2=0.815
r49 14 23 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.255 $Y=0.475
+ $X2=1.255 $Y2=0.365
r50 14 15 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.255 $Y=0.475
+ $X2=1.255 $Y2=0.725
r51 10 23 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.13 $Y=0.365
+ $X2=1.255 $Y2=0.365
r52 10 12 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=1.13 $Y=0.365
+ $X2=0.275 $Y2=0.365
r53 3 20 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.97
+ $Y=0.235 $X2=2.155 $Y2=0.39
r54 2 25 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.215 $Y2=0.73
r55 2 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.215 $Y2=0.39
r56 1 12 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%VGND 1 2 3 4 15 19 23 27 30 31 33 34 36 37
+ 38 40 59 60 63
r90 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r91 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r92 57 60 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r93 56 59 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r94 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r95 54 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r96 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r97 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r98 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r99 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r100 48 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r101 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r102 45 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=0 $X2=1.685
+ $Y2=0
r103 45 47 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=1.77 $Y=0 $X2=2.53
+ $Y2=0
r104 40 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.6 $Y=0 $X2=1.685
+ $Y2=0
r105 40 42 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=1.6 $Y=0 $X2=0.23
+ $Y2=0
r106 38 64 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.61 $Y2=0
r107 38 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r108 36 53 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=4.545 $Y=0
+ $X2=4.37 $Y2=0
r109 36 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.545 $Y=0 $X2=4.63
+ $Y2=0
r110 35 56 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.715 $Y=0
+ $X2=4.83 $Y2=0
r111 35 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.715 $Y=0 $X2=4.63
+ $Y2=0
r112 33 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.45
+ $Y2=0
r113 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0 $X2=3.655
+ $Y2=0
r114 32 53 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.74 $Y=0 $X2=4.37
+ $Y2=0
r115 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.74 $Y=0 $X2=3.655
+ $Y2=0
r116 30 47 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.53
+ $Y2=0
r117 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0 $X2=2.715
+ $Y2=0
r118 29 50 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.8 $Y=0 $X2=3.45
+ $Y2=0
r119 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=0 $X2=2.715
+ $Y2=0
r120 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0
r121 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.63 $Y=0.085
+ $X2=4.63 $Y2=0.39
r122 21 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0
r123 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.655 $Y=0.085
+ $X2=3.655 $Y2=0.39
r124 17 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0
r125 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0.39
r126 13 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0
r127 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.685 $Y=0.085
+ $X2=1.685 $Y2=0.39
r128 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.495
+ $Y=0.235 $X2=4.63 $Y2=0.39
r129 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.235 $X2=3.655 $Y2=0.39
r130 2 19 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=2.57
+ $Y=0.235 $X2=2.715 $Y2=0.39
r131 1 15 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.5
+ $Y=0.235 $X2=1.685 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XNOR2_2%A_600_47# 1 2 3 12 14 15 18 22 24 25
r51 24 25 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.57 $Y=0.775
+ $X2=5.405 $Y2=0.775
r52 21 22 9.6806 $w=1.8e-07 $l=2.08e-07 $layer=LI1_cond $X=4.325 $Y=0.815
+ $X2=4.117 $Y2=0.815
r53 21 25 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=4.325 $Y=0.815
+ $X2=5.405 $Y2=0.815
r54 16 22 1.40968 $w=4.15e-07 $l=9e-08 $layer=LI1_cond $X=4.117 $Y=0.725
+ $X2=4.117 $Y2=0.815
r55 16 18 9.30285 $w=4.13e-07 $l=3.35e-07 $layer=LI1_cond $X=4.117 $Y=0.725
+ $X2=4.117 $Y2=0.39
r56 14 22 9.6806 $w=1.8e-07 $l=2.07e-07 $layer=LI1_cond $X=3.91 $Y=0.815
+ $X2=4.117 $Y2=0.815
r57 14 15 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.91 $Y=0.815
+ $X2=3.35 $Y2=0.815
r58 10 15 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.16 $Y=0.725
+ $X2=3.35 $Y2=0.815
r59 10 12 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.16 $Y=0.725
+ $X2=3.16 $Y2=0.39
r60 3 24 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=5.435
+ $Y=0.235 $X2=5.57 $Y2=0.73
r61 2 18 91 $w=1.7e-07 $l=2.87228e-07 $layer=licon1_NDIFF $count=2 $X=3.94
+ $Y=0.235 $X2=4.16 $Y2=0.39
r62 1 12 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3 $Y=0.235
+ $X2=3.185 $Y2=0.39
.ends

