* File: sky130_fd_sc_hdll__buf_16.pxi.spice
* Created: Wed Sep  2 08:24:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_16%A N_A_M1011_g N_A_c_186_n N_A_M1001_g N_A_M1014_g
+ N_A_c_187_n N_A_M1013_g N_A_M1028_g N_A_c_188_n N_A_M1017_g N_A_M1036_g
+ N_A_c_189_n N_A_M1022_g N_A_M1038_g N_A_c_190_n N_A_M1030_g N_A_c_191_n
+ N_A_M1037_g N_A_M1039_g A A N_A_c_184_n N_A_c_185_n A A
+ PM_SKY130_FD_SC_HDLL__BUF_16%A
x_PM_SKY130_FD_SC_HDLL__BUF_16%A_109_47# N_A_109_47#_M1011_d N_A_109_47#_M1028_d
+ N_A_109_47#_M1038_d N_A_109_47#_M1001_s N_A_109_47#_M1017_s
+ N_A_109_47#_M1030_s N_A_109_47#_M1005_g N_A_109_47#_c_329_n
+ N_A_109_47#_M1000_g N_A_109_47#_M1006_g N_A_109_47#_c_330_n
+ N_A_109_47#_M1002_g N_A_109_47#_M1007_g N_A_109_47#_c_331_n
+ N_A_109_47#_M1003_g N_A_109_47#_M1009_g N_A_109_47#_c_332_n
+ N_A_109_47#_M1004_g N_A_109_47#_M1012_g N_A_109_47#_c_333_n
+ N_A_109_47#_M1008_g N_A_109_47#_M1015_g N_A_109_47#_c_334_n
+ N_A_109_47#_M1010_g N_A_109_47#_M1019_g N_A_109_47#_c_335_n
+ N_A_109_47#_M1016_g N_A_109_47#_M1020_g N_A_109_47#_c_336_n
+ N_A_109_47#_M1018_g N_A_109_47#_M1021_g N_A_109_47#_c_337_n
+ N_A_109_47#_M1026_g N_A_109_47#_M1023_g N_A_109_47#_c_338_n
+ N_A_109_47#_M1027_g N_A_109_47#_M1024_g N_A_109_47#_c_339_n
+ N_A_109_47#_M1031_g N_A_109_47#_M1025_g N_A_109_47#_c_340_n
+ N_A_109_47#_M1032_g N_A_109_47#_M1029_g N_A_109_47#_c_341_n
+ N_A_109_47#_M1033_g N_A_109_47#_M1034_g N_A_109_47#_c_342_n
+ N_A_109_47#_M1035_g N_A_109_47#_M1040_g N_A_109_47#_c_343_n
+ N_A_109_47#_M1042_g N_A_109_47#_c_344_n N_A_109_47#_M1043_g
+ N_A_109_47#_M1041_g N_A_109_47#_c_355_n N_A_109_47#_c_358_n
+ N_A_109_47#_c_318_n N_A_109_47#_c_319_n N_A_109_47#_c_345_n
+ N_A_109_47#_c_346_n N_A_109_47#_c_377_n N_A_109_47#_c_381_n
+ N_A_109_47#_c_320_n N_A_109_47#_c_347_n N_A_109_47#_c_393_n
+ N_A_109_47#_c_395_n N_A_109_47#_c_321_n N_A_109_47#_c_348_n
+ N_A_109_47#_c_322_n N_A_109_47#_c_323_n N_A_109_47#_c_324_n
+ N_A_109_47#_c_325_n N_A_109_47#_c_350_n N_A_109_47#_c_326_n
+ N_A_109_47#_c_351_n N_A_109_47#_c_327_n N_A_109_47#_c_328_n
+ PM_SKY130_FD_SC_HDLL__BUF_16%A_109_47#
x_PM_SKY130_FD_SC_HDLL__BUF_16%VPWR N_VPWR_M1001_d N_VPWR_M1013_d N_VPWR_M1022_d
+ N_VPWR_M1037_d N_VPWR_M1002_d N_VPWR_M1004_d N_VPWR_M1010_d N_VPWR_M1018_d
+ N_VPWR_M1027_d N_VPWR_M1032_d N_VPWR_M1035_d N_VPWR_M1043_d N_VPWR_c_762_n
+ N_VPWR_c_763_n N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n
+ N_VPWR_c_768_n N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n
+ N_VPWR_c_773_n N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n
+ N_VPWR_c_778_n N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n
+ N_VPWR_c_783_n N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n
+ N_VPWR_c_788_n N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n N_VPWR_c_792_n
+ N_VPWR_c_793_n N_VPWR_c_794_n VPWR N_VPWR_c_795_n N_VPWR_c_761_n
+ N_VPWR_c_797_n N_VPWR_c_798_n PM_SKY130_FD_SC_HDLL__BUF_16%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_16%X N_X_M1005_d N_X_M1007_d N_X_M1012_d N_X_M1019_d
+ N_X_M1021_d N_X_M1024_d N_X_M1029_d N_X_M1040_d N_X_M1000_s N_X_M1003_s
+ N_X_M1008_s N_X_M1016_s N_X_M1026_s N_X_M1031_s N_X_M1033_s N_X_M1042_s
+ N_X_c_986_n N_X_c_984_n N_X_c_985_n N_X_c_948_n N_X_c_949_n N_X_c_966_n
+ N_X_c_967_n N_X_c_1013_n N_X_c_1015_n N_X_c_1019_n N_X_c_950_n N_X_c_968_n
+ N_X_c_1031_n N_X_c_1033_n N_X_c_1037_n N_X_c_951_n N_X_c_969_n N_X_c_1049_n
+ N_X_c_1053_n N_X_c_952_n N_X_c_970_n N_X_c_1065_n N_X_c_1069_n N_X_c_953_n
+ N_X_c_971_n N_X_c_1081_n N_X_c_1085_n N_X_c_954_n N_X_c_972_n N_X_c_1097_n
+ N_X_c_1101_n N_X_c_955_n N_X_c_973_n N_X_c_1113_n N_X_c_956_n N_X_c_957_n
+ N_X_c_974_n N_X_c_958_n N_X_c_975_n N_X_c_959_n N_X_c_976_n N_X_c_960_n
+ N_X_c_977_n N_X_c_961_n N_X_c_978_n N_X_c_962_n N_X_c_979_n N_X_c_963_n
+ N_X_c_964_n N_X_c_980_n N_X_c_981_n X X X N_X_c_1178_n
+ PM_SKY130_FD_SC_HDLL__BUF_16%X
x_PM_SKY130_FD_SC_HDLL__BUF_16%VGND N_VGND_M1011_s N_VGND_M1014_s N_VGND_M1036_s
+ N_VGND_M1039_s N_VGND_M1006_s N_VGND_M1009_s N_VGND_M1015_s N_VGND_M1020_s
+ N_VGND_M1023_s N_VGND_M1025_s N_VGND_M1034_s N_VGND_M1041_s N_VGND_c_1318_n
+ N_VGND_c_1319_n N_VGND_c_1320_n N_VGND_c_1321_n N_VGND_c_1322_n
+ N_VGND_c_1323_n N_VGND_c_1324_n N_VGND_c_1325_n N_VGND_c_1326_n
+ N_VGND_c_1327_n N_VGND_c_1328_n N_VGND_c_1329_n N_VGND_c_1330_n
+ N_VGND_c_1331_n N_VGND_c_1332_n N_VGND_c_1333_n N_VGND_c_1334_n
+ N_VGND_c_1335_n N_VGND_c_1336_n N_VGND_c_1337_n N_VGND_c_1338_n
+ N_VGND_c_1339_n N_VGND_c_1340_n N_VGND_c_1341_n N_VGND_c_1342_n
+ N_VGND_c_1343_n N_VGND_c_1344_n N_VGND_c_1345_n N_VGND_c_1346_n
+ N_VGND_c_1347_n N_VGND_c_1348_n N_VGND_c_1349_n N_VGND_c_1350_n VGND
+ N_VGND_c_1351_n N_VGND_c_1352_n N_VGND_c_1353_n N_VGND_c_1354_n
+ PM_SKY130_FD_SC_HDLL__BUF_16%VGND
cc_1 VNB N_A_M1011_g 0.0243087f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_M1014_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.56
cc_3 VNB N_A_M1028_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_4 VNB N_A_M1036_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.56
cc_5 VNB N_A_M1038_g 0.0188753f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_6 VNB N_A_M1039_g 0.0185509f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.56
cc_7 VNB N_A_c_184_n 0.0220589f $X=-0.19 $Y=-0.24 $X2=2.5 $Y2=1.16
cc_8 VNB N_A_c_185_n 0.141956f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.217
cc_9 VNB N_A_109_47#_M1005_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_10 VNB N_A_109_47#_M1006_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_11 VNB N_A_109_47#_M1007_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_12 VNB N_A_109_47#_M1009_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_109_47#_M1012_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.217
cc_14 VNB N_A_109_47#_M1015_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.217
cc_15 VNB N_A_109_47#_M1019_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.217
cc_16 VNB N_A_109_47#_M1020_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=2.075 $Y2=1.175
cc_17 VNB N_A_109_47#_M1021_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_109_47#_M1023_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_109_47#_M1024_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_109_47#_M1025_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_109_47#_M1029_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_109_47#_M1034_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_109_47#_M1040_g 0.0188791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_109_47#_M1041_g 0.0219373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_109_47#_c_318_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_109_47#_c_319_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_109_47#_c_320_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_109_47#_c_321_n 9.58484e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_109_47#_c_322_n 0.00305698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_109_47#_c_323_n 5.27693e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_109_47#_c_324_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_109_47#_c_325_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_109_47#_c_326_n 0.00278347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_109_47#_c_327_n 0.00163661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_109_47#_c_328_n 0.376772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VPWR_c_761_n 0.478484f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_948_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.217
cc_38 VNB N_X_c_949_n 0.00253087f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=1.217
cc_39 VNB N_X_c_950_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=1.62 $Y2=1.175
cc_40 VNB N_X_c_951_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_952_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_953_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_954_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_955_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_956_n 0.00248919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_X_c_957_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_X_c_958_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_X_c_959_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_X_c_960_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_X_c_961_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_X_c_962_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_X_c_963_n 0.00298874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_X_c_964_n 0.0341207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB X 0.0268696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_1318_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.985
cc_56 VNB N_VGND_c_1319_n 0.00713663f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=1.025
cc_57 VNB N_VGND_c_1320_n 0.0200002f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.56
cc_58 VNB N_VGND_c_1321_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_1322_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.217
cc_60 VNB N_VGND_c_1323_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_61 VNB N_VGND_c_1324_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.217
cc_62 VNB N_VGND_c_1325_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.217
cc_63 VNB N_VGND_c_1326_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.217
cc_64 VNB N_VGND_c_1327_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.175
cc_65 VNB N_VGND_c_1328_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.075 $Y2=1.19
cc_66 VNB N_VGND_c_1329_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1330_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1331_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1332_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1333_n 0.0193874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1334_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1335_n 0.0198969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1336_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_VGND_c_1337_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1338_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1339_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1340_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1341_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1342_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1343_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1344_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1345_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1346_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1347_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1348_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1349_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1350_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1351_n 0.02536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1352_n 0.539794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1353_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1354_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VPB N_A_c_186_n 0.0198486f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_93 VPB N_A_c_187_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_94 VPB N_A_c_188_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_95 VPB N_A_c_189_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_96 VPB N_A_c_190_n 0.0158857f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_97 VPB N_A_c_191_n 0.0159692f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_98 VPB N_A_c_185_n 0.0416088f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.217
cc_99 VPB N_A_109_47#_c_329_n 0.0162292f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_100 VPB N_A_109_47#_c_330_n 0.0158858f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=0.56
cc_101 VPB N_A_109_47#_c_331_n 0.0158869f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_102 VPB N_A_109_47#_c_332_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.995 $Y2=1.105
cc_103 VPB N_A_109_47#_c_333_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_104 VPB N_A_109_47#_c_334_n 0.0158869f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=1.217
cc_105 VPB N_A_109_47#_c_335_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.175
cc_106 VPB N_A_109_47#_c_336_n 0.0158869f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.175
cc_107 VPB N_A_109_47#_c_337_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_109_47#_c_338_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_109_47#_c_339_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_A_109_47#_c_340_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_109_47#_c_341_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_A_109_47#_c_342_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_A_109_47#_c_343_n 0.0158865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_A_109_47#_c_344_n 0.0192027f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_A_109_47#_c_345_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_A_109_47#_c_346_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_109_47#_c_347_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_A_109_47#_c_348_n 9.4165e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_109_47#_c_323_n 0.0025308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_109_47#_c_350_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_109_47#_c_351_n 0.00179747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_109_47#_c_328_n 0.102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_VPWR_c_762_n 0.0110239f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_124 VPB N_VPWR_c_763_n 0.00807576f $X=-0.19 $Y=1.305 $X2=2.87 $Y2=1.025
cc_125 VPB N_VPWR_c_764_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.105
cc_126 VPB N_VPWR_c_765_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.217
cc_127 VPB N_VPWR_c_766_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.217
cc_128 VPB N_VPWR_c_767_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_129 VPB N_VPWR_c_768_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_130 VPB N_VPWR_c_769_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.5 $Y2=1.16
cc_131 VPB N_VPWR_c_770_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.175
cc_132 VPB N_VPWR_c_771_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.62 $Y2=1.175
cc_133 VPB N_VPWR_c_772_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.5 $Y2=1.175
cc_134 VPB N_VPWR_c_773_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_VPWR_c_774_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_VPWR_c_775_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_VPWR_c_776_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_VPWR_c_777_n 0.020564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_VPWR_c_778_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_VPWR_c_779_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_780_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_781_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_782_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_783_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_784_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_785_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_786_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_787_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_788_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_789_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_790_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_791_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_792_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_793_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_794_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_795_n 0.025987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_761_n 0.0651591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_797_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_798_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_X_c_966_n 0.00172363f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.217
cc_161 VPB N_X_c_967_n 0.00176159f $X=-0.19 $Y=1.305 $X2=2.5 $Y2=1.217
cc_162 VPB N_X_c_968_n 0.00172363f $X=-0.19 $Y=1.305 $X2=2.075 $Y2=1.19
cc_163 VPB N_X_c_969_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_X_c_970_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_X_c_971_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_X_c_972_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_X_c_973_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_X_c_974_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_X_c_975_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_X_c_976_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_X_c_977_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_X_c_978_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_X_c_979_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_X_c_980_n 0.00231436f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_X_c_981_n 0.0578556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB X 0.00194398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB X 0.0095361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 N_A_M1039_g N_A_109_47#_M1005_g 0.0207158f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A_c_191_n N_A_109_47#_c_329_n 0.0216821f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_M1011_g N_A_109_47#_c_355_n 0.00545788f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A_M1014_g N_A_109_47#_c_355_n 0.00693104f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_182 N_A_M1028_g N_A_109_47#_c_355_n 5.47131e-19 $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_c_186_n N_A_109_47#_c_358_n 0.0128929f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_187_n N_A_109_47#_c_358_n 0.0115459f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_c_188_n N_A_109_47#_c_358_n 7.68612e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_M1014_g N_A_109_47#_c_318_n 0.00879805f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A_M1028_g N_A_109_47#_c_318_n 0.00879805f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A_c_184_n N_A_109_47#_c_318_n 0.03957f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_189 N_A_c_185_n N_A_109_47#_c_318_n 0.0031956f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_190 N_A_M1011_g N_A_109_47#_c_319_n 0.00255105f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_M1014_g N_A_109_47#_c_319_n 0.00113891f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A_c_184_n N_A_109_47#_c_319_n 0.030582f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_c_185_n N_A_109_47#_c_319_n 0.00331919f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_194 N_A_c_187_n N_A_109_47#_c_345_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_188_n N_A_109_47#_c_345_n 0.0101048f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_184_n N_A_109_47#_c_345_n 0.0394547f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_c_185_n N_A_109_47#_c_345_n 0.00720931f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_198 N_A_c_186_n N_A_109_47#_c_346_n 0.00397051f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_187_n N_A_109_47#_c_346_n 0.00107777f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_184_n N_A_109_47#_c_346_n 0.0305808f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_c_185_n N_A_109_47#_c_346_n 0.0074788f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_202 N_A_M1014_g N_A_109_47#_c_377_n 5.25882e-19 $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_M1028_g N_A_109_47#_c_377_n 0.00657592f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_204 N_A_M1036_g N_A_109_47#_c_377_n 0.00693104f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_205 N_A_M1038_g N_A_109_47#_c_377_n 5.47131e-19 $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_c_187_n N_A_109_47#_c_381_n 8.07084e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_c_188_n N_A_109_47#_c_381_n 0.0141618f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_189_n N_A_109_47#_c_381_n 0.0115459f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_c_190_n N_A_109_47#_c_381_n 7.68612e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_M1036_g N_A_109_47#_c_320_n 0.00879805f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A_M1038_g N_A_109_47#_c_320_n 0.00879805f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_212 N_A_c_184_n N_A_109_47#_c_320_n 0.03957f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_c_185_n N_A_109_47#_c_320_n 0.0031956f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_214 N_A_c_189_n N_A_109_47#_c_347_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_190_n N_A_109_47#_c_347_n 0.0101048f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_184_n N_A_109_47#_c_347_n 0.0394547f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_c_185_n N_A_109_47#_c_347_n 0.00720931f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_218 N_A_M1036_g N_A_109_47#_c_393_n 5.25882e-19 $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A_M1038_g N_A_109_47#_c_393_n 0.00657592f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_220 N_A_c_189_n N_A_109_47#_c_395_n 8.07084e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_c_190_n N_A_109_47#_c_395_n 0.0141618f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_191_n N_A_109_47#_c_395_n 0.0115459f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_M1039_g N_A_109_47#_c_321_n 0.0116573f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_c_191_n N_A_109_47#_c_348_n 0.0151183f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_185_n N_A_109_47#_c_348_n 3.58038e-19 $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_226 N_A_M1039_g N_A_109_47#_c_322_n 0.00415408f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_c_191_n N_A_109_47#_c_323_n 8.26658e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_185_n N_A_109_47#_c_323_n 0.00331109f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_229 N_A_M1028_g N_A_109_47#_c_325_n 0.00113891f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_M1036_g N_A_109_47#_c_325_n 0.00113891f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A_c_184_n N_A_109_47#_c_325_n 0.030582f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_c_185_n N_A_109_47#_c_325_n 0.00331919f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_233 N_A_c_188_n N_A_109_47#_c_350_n 0.00260297f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_c_189_n N_A_109_47#_c_350_n 0.00107777f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_184_n N_A_109_47#_c_350_n 0.0305808f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_c_185_n N_A_109_47#_c_350_n 0.0074788f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_237 N_A_M1038_g N_A_109_47#_c_326_n 0.0011682f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A_c_184_n N_A_109_47#_c_326_n 0.0274674f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_c_185_n N_A_109_47#_c_326_n 0.00450461f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_240 N_A_c_190_n N_A_109_47#_c_351_n 0.00259297f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_c_191_n N_A_109_47#_c_351_n 0.00128868f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_c_184_n N_A_109_47#_c_351_n 0.0274092f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_243 N_A_c_185_n N_A_109_47#_c_351_n 0.00735453f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_244 N_A_c_184_n N_A_109_47#_c_327_n 0.0130035f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_c_185_n N_A_109_47#_c_327_n 0.00237077f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_246 N_A_c_185_n N_A_109_47#_c_328_n 0.0207158f $X=2.845 $Y=1.217 $X2=0 $Y2=0
cc_247 N_A_c_186_n N_VPWR_c_763_n 0.0082969f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A_c_184_n N_VPWR_c_763_n 0.0143482f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_249 N_A_c_186_n N_VPWR_c_764_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_c_187_n N_VPWR_c_764_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_c_187_n N_VPWR_c_765_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_188_n N_VPWR_c_765_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_188_n N_VPWR_c_766_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_189_n N_VPWR_c_766_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_189_n N_VPWR_c_767_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_c_190_n N_VPWR_c_767_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_c_191_n N_VPWR_c_768_n 0.0052072f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_190_n N_VPWR_c_777_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_c_191_n N_VPWR_c_777_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_186_n N_VPWR_c_761_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_187_n N_VPWR_c_761_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_188_n N_VPWR_c_761_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_189_n N_VPWR_c_761_n 0.0118438f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_190_n N_VPWR_c_761_n 0.00999457f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_191_n N_VPWR_c_761_n 0.011869f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_M1039_g N_X_c_984_n 4.77587e-19 $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_c_191_n N_X_c_985_n 8.07084e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_M1011_g N_VGND_c_1319_n 0.00482457f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A_c_184_n N_VGND_c_1319_n 0.0143482f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_M1011_g N_VGND_c_1320_n 0.00541562f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A_M1014_g N_VGND_c_1320_n 0.00424619f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_272 N_A_M1014_g N_VGND_c_1321_n 0.00390178f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A_M1028_g N_VGND_c_1321_n 0.00276126f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_M1028_g N_VGND_c_1322_n 0.00424619f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_275 N_A_M1036_g N_VGND_c_1322_n 0.00424619f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A_M1036_g N_VGND_c_1323_n 0.00390178f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A_M1038_g N_VGND_c_1323_n 0.00276126f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A_M1039_g N_VGND_c_1324_n 0.00268723f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_M1038_g N_VGND_c_1333_n 0.00424619f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A_M1039_g N_VGND_c_1333_n 0.00439206f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_M1011_g N_VGND_c_1352_n 0.0105829f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_M1014_g N_VGND_c_1352_n 0.00611295f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_M1028_g N_VGND_c_1352_n 0.00599018f $X=1.41 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_M1036_g N_VGND_c_1352_n 0.00611295f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_M1038_g N_VGND_c_1352_n 0.00610552f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_M1039_g N_VGND_c_1352_n 0.00618081f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_109_47#_c_345_n N_VPWR_M1013_d 0.00199888f $X=1.455 $Y=1.53 $X2=0
+ $Y2=0
cc_288 N_A_109_47#_c_347_n N_VPWR_M1022_d 0.00199888f $X=2.395 $Y=1.53 $X2=0
+ $Y2=0
cc_289 N_A_109_47#_c_348_n N_VPWR_M1037_d 0.00347056f $X=2.99 $Y=1.53 $X2=0
+ $Y2=0
cc_290 N_A_109_47#_c_358_n N_VPWR_c_763_n 0.0634185f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_291 N_A_109_47#_c_346_n N_VPWR_c_763_n 0.013414f $X=0.895 $Y=1.53 $X2=0 $Y2=0
cc_292 N_A_109_47#_c_358_n N_VPWR_c_764_n 0.0223557f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_293 N_A_109_47#_c_358_n N_VPWR_c_765_n 0.0385613f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_294 N_A_109_47#_c_345_n N_VPWR_c_765_n 0.0112848f $X=1.455 $Y=1.53 $X2=0
+ $Y2=0
cc_295 N_A_109_47#_c_381_n N_VPWR_c_765_n 0.0470327f $X=1.67 $Y=1.63 $X2=0 $Y2=0
cc_296 N_A_109_47#_c_381_n N_VPWR_c_766_n 0.0223557f $X=1.67 $Y=1.63 $X2=0 $Y2=0
cc_297 N_A_109_47#_c_381_n N_VPWR_c_767_n 0.0385613f $X=1.67 $Y=1.63 $X2=0 $Y2=0
cc_298 N_A_109_47#_c_347_n N_VPWR_c_767_n 0.0112848f $X=2.395 $Y=1.53 $X2=0
+ $Y2=0
cc_299 N_A_109_47#_c_395_n N_VPWR_c_767_n 0.0470327f $X=2.61 $Y=1.63 $X2=0 $Y2=0
cc_300 N_A_109_47#_c_329_n N_VPWR_c_768_n 0.004751f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_109_47#_c_395_n N_VPWR_c_768_n 0.0385613f $X=2.61 $Y=1.63 $X2=0 $Y2=0
cc_302 N_A_109_47#_c_348_n N_VPWR_c_768_n 0.0124926f $X=2.99 $Y=1.53 $X2=0 $Y2=0
cc_303 N_A_109_47#_c_330_n N_VPWR_c_769_n 0.0052072f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_304 N_A_109_47#_c_331_n N_VPWR_c_769_n 0.004751f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_305 N_A_109_47#_c_332_n N_VPWR_c_770_n 0.0052072f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_306 N_A_109_47#_c_333_n N_VPWR_c_770_n 0.004751f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_109_47#_c_334_n N_VPWR_c_771_n 0.0052072f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_308 N_A_109_47#_c_335_n N_VPWR_c_771_n 0.004751f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_109_47#_c_336_n N_VPWR_c_772_n 0.0052072f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_310 N_A_109_47#_c_337_n N_VPWR_c_772_n 0.004751f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_109_47#_c_338_n N_VPWR_c_773_n 0.0052072f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_312 N_A_109_47#_c_339_n N_VPWR_c_773_n 0.004751f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A_109_47#_c_340_n N_VPWR_c_774_n 0.0052072f $X=8.485 $Y=1.41 $X2=0
+ $Y2=0
cc_314 N_A_109_47#_c_341_n N_VPWR_c_774_n 0.004751f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_109_47#_c_342_n N_VPWR_c_775_n 0.0052072f $X=9.425 $Y=1.41 $X2=0
+ $Y2=0
cc_316 N_A_109_47#_c_343_n N_VPWR_c_775_n 0.004751f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_109_47#_c_344_n N_VPWR_c_776_n 0.00688901f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_109_47#_c_395_n N_VPWR_c_777_n 0.0223557f $X=2.61 $Y=1.63 $X2=0 $Y2=0
cc_319 N_A_109_47#_c_329_n N_VPWR_c_779_n 0.00597712f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_109_47#_c_330_n N_VPWR_c_779_n 0.00673617f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_321 N_A_109_47#_c_331_n N_VPWR_c_781_n 0.00597712f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_322 N_A_109_47#_c_332_n N_VPWR_c_781_n 0.00673617f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_109_47#_c_333_n N_VPWR_c_783_n 0.00597712f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_324 N_A_109_47#_c_334_n N_VPWR_c_783_n 0.00673617f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_325 N_A_109_47#_c_335_n N_VPWR_c_785_n 0.00597712f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_326 N_A_109_47#_c_336_n N_VPWR_c_785_n 0.00673617f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_A_109_47#_c_337_n N_VPWR_c_787_n 0.00597712f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A_109_47#_c_338_n N_VPWR_c_787_n 0.00673617f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_A_109_47#_c_339_n N_VPWR_c_789_n 0.00597712f $X=8.015 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_A_109_47#_c_340_n N_VPWR_c_789_n 0.00673617f $X=8.485 $Y=1.41 $X2=0
+ $Y2=0
cc_331 N_A_109_47#_c_341_n N_VPWR_c_791_n 0.00597712f $X=8.955 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_A_109_47#_c_342_n N_VPWR_c_791_n 0.00673617f $X=9.425 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A_109_47#_c_343_n N_VPWR_c_793_n 0.00597712f $X=9.895 $Y=1.41 $X2=0
+ $Y2=0
cc_334 N_A_109_47#_c_344_n N_VPWR_c_793_n 0.00673617f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_335 N_A_109_47#_M1001_s N_VPWR_c_761_n 0.00231261f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_336 N_A_109_47#_M1017_s N_VPWR_c_761_n 0.00231261f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_337 N_A_109_47#_M1030_s N_VPWR_c_761_n 0.00231261f $X=2.465 $Y=1.485 $X2=0
+ $Y2=0
cc_338 N_A_109_47#_c_329_n N_VPWR_c_761_n 0.0100198f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_339 N_A_109_47#_c_330_n N_VPWR_c_761_n 0.0118438f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_340 N_A_109_47#_c_331_n N_VPWR_c_761_n 0.00999457f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A_109_47#_c_332_n N_VPWR_c_761_n 0.0118438f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_342 N_A_109_47#_c_333_n N_VPWR_c_761_n 0.00999457f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A_109_47#_c_334_n N_VPWR_c_761_n 0.0118438f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_344 N_A_109_47#_c_335_n N_VPWR_c_761_n 0.00999457f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_345 N_A_109_47#_c_336_n N_VPWR_c_761_n 0.0118438f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_346 N_A_109_47#_c_337_n N_VPWR_c_761_n 0.00999457f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_A_109_47#_c_338_n N_VPWR_c_761_n 0.0118438f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_348 N_A_109_47#_c_339_n N_VPWR_c_761_n 0.00999457f $X=8.015 $Y=1.41 $X2=0
+ $Y2=0
cc_349 N_A_109_47#_c_340_n N_VPWR_c_761_n 0.0118438f $X=8.485 $Y=1.41 $X2=0
+ $Y2=0
cc_350 N_A_109_47#_c_341_n N_VPWR_c_761_n 0.00999457f $X=8.955 $Y=1.41 $X2=0
+ $Y2=0
cc_351 N_A_109_47#_c_342_n N_VPWR_c_761_n 0.0118438f $X=9.425 $Y=1.41 $X2=0
+ $Y2=0
cc_352 N_A_109_47#_c_343_n N_VPWR_c_761_n 0.00999457f $X=9.895 $Y=1.41 $X2=0
+ $Y2=0
cc_353 N_A_109_47#_c_344_n N_VPWR_c_761_n 0.0131262f $X=10.365 $Y=1.41 $X2=0
+ $Y2=0
cc_354 N_A_109_47#_c_358_n N_VPWR_c_761_n 0.0140101f $X=0.73 $Y=1.63 $X2=0 $Y2=0
cc_355 N_A_109_47#_c_381_n N_VPWR_c_761_n 0.0140101f $X=1.67 $Y=1.63 $X2=0 $Y2=0
cc_356 N_A_109_47#_c_395_n N_VPWR_c_761_n 0.0140101f $X=2.61 $Y=1.63 $X2=0 $Y2=0
cc_357 N_A_109_47#_M1005_g N_X_c_986_n 0.00229101f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_109_47#_M1006_g N_X_c_986_n 0.00248233f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_109_47#_M1005_g N_X_c_984_n 0.00426764f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_109_47#_M1006_g N_X_c_984_n 0.00445433f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_109_47#_M1007_g N_X_c_984_n 4.84753e-19 $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_109_47#_c_329_n N_X_c_985_n 0.0141618f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_109_47#_c_330_n N_X_c_985_n 0.0115459f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_109_47#_c_331_n N_X_c_985_n 7.68612e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_109_47#_c_395_n N_X_c_985_n 0.00629866f $X=2.61 $Y=1.63 $X2=0 $Y2=0
cc_366 N_A_109_47#_M1006_g N_X_c_948_n 0.00879805f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_367 N_A_109_47#_M1007_g N_X_c_948_n 0.00879805f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_368 N_A_109_47#_c_324_n N_X_c_948_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A_109_47#_c_328_n N_X_c_948_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_370 N_A_109_47#_M1005_g N_X_c_949_n 0.00245067f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_109_47#_M1006_g N_X_c_949_n 0.00115337f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_109_47#_c_321_n N_X_c_949_n 0.00808484f $X=2.99 $Y=0.82 $X2=0 $Y2=0
cc_373 N_A_109_47#_c_324_n N_X_c_949_n 0.0305973f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_109_47#_c_328_n N_X_c_949_n 0.00332f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_375 N_A_109_47#_c_330_n N_X_c_966_n 0.0137916f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_109_47#_c_331_n N_X_c_966_n 0.0101048f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A_109_47#_c_324_n N_X_c_966_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_109_47#_c_328_n N_X_c_966_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_379 N_A_109_47#_c_329_n N_X_c_967_n 0.00386185f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_380 N_A_109_47#_c_330_n N_X_c_967_n 0.00107777f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_381 N_A_109_47#_c_348_n N_X_c_967_n 0.0149281f $X=2.99 $Y=1.53 $X2=0 $Y2=0
cc_382 N_A_109_47#_c_324_n N_X_c_967_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_109_47#_c_328_n N_X_c_967_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_384 N_A_109_47#_M1007_g N_X_c_1013_n 0.00226116f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A_109_47#_M1009_g N_X_c_1013_n 0.00248233f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_386 N_A_109_47#_M1006_g N_X_c_1015_n 4.7681e-19 $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_387 N_A_109_47#_M1007_g N_X_c_1015_n 0.0043216f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_388 N_A_109_47#_M1009_g N_X_c_1015_n 0.00445433f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_389 N_A_109_47#_M1012_g N_X_c_1015_n 4.84753e-19 $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_390 N_A_109_47#_c_330_n N_X_c_1019_n 8.07084e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_391 N_A_109_47#_c_331_n N_X_c_1019_n 0.0141618f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_392 N_A_109_47#_c_332_n N_X_c_1019_n 0.0115459f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A_109_47#_c_333_n N_X_c_1019_n 7.68612e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_394 N_A_109_47#_M1009_g N_X_c_950_n 0.00879805f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_395 N_A_109_47#_M1012_g N_X_c_950_n 0.00879805f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_396 N_A_109_47#_c_324_n N_X_c_950_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_397 N_A_109_47#_c_328_n N_X_c_950_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_398 N_A_109_47#_c_332_n N_X_c_968_n 0.0137916f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_399 N_A_109_47#_c_333_n N_X_c_968_n 0.0101048f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_400 N_A_109_47#_c_324_n N_X_c_968_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_401 N_A_109_47#_c_328_n N_X_c_968_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_402 N_A_109_47#_M1012_g N_X_c_1031_n 0.00226116f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_403 N_A_109_47#_M1015_g N_X_c_1031_n 0.00248233f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_404 N_A_109_47#_M1009_g N_X_c_1033_n 4.7681e-19 $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_405 N_A_109_47#_M1012_g N_X_c_1033_n 0.0043216f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_406 N_A_109_47#_M1015_g N_X_c_1033_n 0.00445433f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_407 N_A_109_47#_M1019_g N_X_c_1033_n 4.84753e-19 $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_408 N_A_109_47#_c_332_n N_X_c_1037_n 8.07084e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_409 N_A_109_47#_c_333_n N_X_c_1037_n 0.0141618f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_410 N_A_109_47#_c_334_n N_X_c_1037_n 0.0115459f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_411 N_A_109_47#_c_335_n N_X_c_1037_n 7.68612e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_412 N_A_109_47#_M1015_g N_X_c_951_n 0.00879805f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_413 N_A_109_47#_M1019_g N_X_c_951_n 0.00879805f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_414 N_A_109_47#_c_324_n N_X_c_951_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_415 N_A_109_47#_c_328_n N_X_c_951_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_416 N_A_109_47#_c_334_n N_X_c_969_n 0.0137916f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_417 N_A_109_47#_c_335_n N_X_c_969_n 0.0101048f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_418 N_A_109_47#_c_324_n N_X_c_969_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_419 N_A_109_47#_c_328_n N_X_c_969_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_420 N_A_109_47#_M1015_g N_X_c_1049_n 5.25882e-19 $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_421 N_A_109_47#_M1019_g N_X_c_1049_n 0.00657592f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_422 N_A_109_47#_M1020_g N_X_c_1049_n 0.00693104f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_423 N_A_109_47#_M1021_g N_X_c_1049_n 5.47131e-19 $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_424 N_A_109_47#_c_334_n N_X_c_1053_n 8.07084e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_425 N_A_109_47#_c_335_n N_X_c_1053_n 0.0141618f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_426 N_A_109_47#_c_336_n N_X_c_1053_n 0.0115459f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_427 N_A_109_47#_c_337_n N_X_c_1053_n 7.68612e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_428 N_A_109_47#_M1020_g N_X_c_952_n 0.00879805f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_429 N_A_109_47#_M1021_g N_X_c_952_n 0.00879805f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_430 N_A_109_47#_c_324_n N_X_c_952_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_431 N_A_109_47#_c_328_n N_X_c_952_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_432 N_A_109_47#_c_336_n N_X_c_970_n 0.0137916f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_433 N_A_109_47#_c_337_n N_X_c_970_n 0.0101048f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_434 N_A_109_47#_c_324_n N_X_c_970_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_435 N_A_109_47#_c_328_n N_X_c_970_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_436 N_A_109_47#_M1020_g N_X_c_1065_n 5.25882e-19 $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_437 N_A_109_47#_M1021_g N_X_c_1065_n 0.00657592f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_438 N_A_109_47#_M1023_g N_X_c_1065_n 0.00693104f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_439 N_A_109_47#_M1024_g N_X_c_1065_n 5.47131e-19 $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_440 N_A_109_47#_c_336_n N_X_c_1069_n 8.07084e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_441 N_A_109_47#_c_337_n N_X_c_1069_n 0.0141618f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_442 N_A_109_47#_c_338_n N_X_c_1069_n 0.0115459f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_443 N_A_109_47#_c_339_n N_X_c_1069_n 7.68612e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_444 N_A_109_47#_M1023_g N_X_c_953_n 0.00879805f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_445 N_A_109_47#_M1024_g N_X_c_953_n 0.00879805f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_446 N_A_109_47#_c_324_n N_X_c_953_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_447 N_A_109_47#_c_328_n N_X_c_953_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_448 N_A_109_47#_c_338_n N_X_c_971_n 0.0137916f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_449 N_A_109_47#_c_339_n N_X_c_971_n 0.0101048f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_450 N_A_109_47#_c_324_n N_X_c_971_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_451 N_A_109_47#_c_328_n N_X_c_971_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_452 N_A_109_47#_M1023_g N_X_c_1081_n 5.25882e-19 $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_453 N_A_109_47#_M1024_g N_X_c_1081_n 0.00657592f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_454 N_A_109_47#_M1025_g N_X_c_1081_n 0.00693104f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_455 N_A_109_47#_M1029_g N_X_c_1081_n 5.47131e-19 $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_456 N_A_109_47#_c_338_n N_X_c_1085_n 8.07084e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_457 N_A_109_47#_c_339_n N_X_c_1085_n 0.0141618f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_458 N_A_109_47#_c_340_n N_X_c_1085_n 0.0115459f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_459 N_A_109_47#_c_341_n N_X_c_1085_n 7.68612e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_109_47#_M1025_g N_X_c_954_n 0.00879805f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_461 N_A_109_47#_M1029_g N_X_c_954_n 0.00879805f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_462 N_A_109_47#_c_324_n N_X_c_954_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_463 N_A_109_47#_c_328_n N_X_c_954_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_464 N_A_109_47#_c_340_n N_X_c_972_n 0.0137916f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_465 N_A_109_47#_c_341_n N_X_c_972_n 0.0101048f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_466 N_A_109_47#_c_324_n N_X_c_972_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_467 N_A_109_47#_c_328_n N_X_c_972_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_468 N_A_109_47#_M1025_g N_X_c_1097_n 5.25882e-19 $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_469 N_A_109_47#_M1029_g N_X_c_1097_n 0.00657592f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_470 N_A_109_47#_M1034_g N_X_c_1097_n 0.00693104f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_471 N_A_109_47#_M1040_g N_X_c_1097_n 5.47131e-19 $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_472 N_A_109_47#_c_340_n N_X_c_1101_n 8.07084e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_473 N_A_109_47#_c_341_n N_X_c_1101_n 0.0141618f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_474 N_A_109_47#_c_342_n N_X_c_1101_n 0.0115459f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_475 N_A_109_47#_c_343_n N_X_c_1101_n 7.68612e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_476 N_A_109_47#_M1034_g N_X_c_955_n 0.00879805f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_477 N_A_109_47#_M1040_g N_X_c_955_n 0.00879805f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_478 N_A_109_47#_c_324_n N_X_c_955_n 0.03957f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_479 N_A_109_47#_c_328_n N_X_c_955_n 0.0031956f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_480 N_A_109_47#_c_342_n N_X_c_973_n 0.0137916f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_481 N_A_109_47#_c_343_n N_X_c_973_n 0.0101048f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_482 N_A_109_47#_c_324_n N_X_c_973_n 0.0394547f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_483 N_A_109_47#_c_328_n N_X_c_973_n 0.00720931f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_484 N_A_109_47#_M1034_g N_X_c_1113_n 5.25882e-19 $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_485 N_A_109_47#_M1040_g N_X_c_1113_n 0.00657592f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_486 N_A_109_47#_M1041_g N_X_c_956_n 0.014164f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_487 N_A_109_47#_M1007_g N_X_c_957_n 0.00115337f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_488 N_A_109_47#_M1009_g N_X_c_957_n 0.00115337f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_489 N_A_109_47#_c_324_n N_X_c_957_n 0.0305905f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_490 N_A_109_47#_c_328_n N_X_c_957_n 0.00331994f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_491 N_A_109_47#_c_331_n N_X_c_974_n 0.00260297f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_492 N_A_109_47#_c_332_n N_X_c_974_n 0.00107777f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A_109_47#_c_324_n N_X_c_974_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_494 N_A_109_47#_c_328_n N_X_c_974_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_495 N_A_109_47#_M1012_g N_X_c_958_n 0.00115337f $X=5.17 $Y=0.56 $X2=0 $Y2=0
cc_496 N_A_109_47#_M1015_g N_X_c_958_n 0.00115337f $X=5.64 $Y=0.56 $X2=0 $Y2=0
cc_497 N_A_109_47#_c_324_n N_X_c_958_n 0.0305905f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_498 N_A_109_47#_c_328_n N_X_c_958_n 0.00331994f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_499 N_A_109_47#_c_333_n N_X_c_975_n 0.00260297f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_500 N_A_109_47#_c_334_n N_X_c_975_n 0.00107777f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_501 N_A_109_47#_c_324_n N_X_c_975_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_502 N_A_109_47#_c_328_n N_X_c_975_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_503 N_A_109_47#_M1019_g N_X_c_959_n 0.00113891f $X=6.11 $Y=0.56 $X2=0 $Y2=0
cc_504 N_A_109_47#_M1020_g N_X_c_959_n 0.00113891f $X=6.58 $Y=0.56 $X2=0 $Y2=0
cc_505 N_A_109_47#_c_324_n N_X_c_959_n 0.030582f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_506 N_A_109_47#_c_328_n N_X_c_959_n 0.00331919f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_507 N_A_109_47#_c_335_n N_X_c_976_n 0.00260297f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_508 N_A_109_47#_c_336_n N_X_c_976_n 0.00107777f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_509 N_A_109_47#_c_324_n N_X_c_976_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_510 N_A_109_47#_c_328_n N_X_c_976_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_511 N_A_109_47#_M1021_g N_X_c_960_n 0.00113891f $X=7.05 $Y=0.56 $X2=0 $Y2=0
cc_512 N_A_109_47#_M1023_g N_X_c_960_n 0.00113891f $X=7.52 $Y=0.56 $X2=0 $Y2=0
cc_513 N_A_109_47#_c_324_n N_X_c_960_n 0.030582f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_514 N_A_109_47#_c_328_n N_X_c_960_n 0.00331919f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_515 N_A_109_47#_c_337_n N_X_c_977_n 0.00260297f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_516 N_A_109_47#_c_338_n N_X_c_977_n 0.00107777f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_517 N_A_109_47#_c_324_n N_X_c_977_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_518 N_A_109_47#_c_328_n N_X_c_977_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_519 N_A_109_47#_M1024_g N_X_c_961_n 0.00113891f $X=7.99 $Y=0.56 $X2=0 $Y2=0
cc_520 N_A_109_47#_M1025_g N_X_c_961_n 0.00113891f $X=8.46 $Y=0.56 $X2=0 $Y2=0
cc_521 N_A_109_47#_c_324_n N_X_c_961_n 0.030582f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_522 N_A_109_47#_c_328_n N_X_c_961_n 0.00331919f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_523 N_A_109_47#_c_339_n N_X_c_978_n 0.00260297f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_524 N_A_109_47#_c_340_n N_X_c_978_n 0.00107777f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_525 N_A_109_47#_c_324_n N_X_c_978_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_526 N_A_109_47#_c_328_n N_X_c_978_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_527 N_A_109_47#_M1029_g N_X_c_962_n 0.00113891f $X=8.93 $Y=0.56 $X2=0 $Y2=0
cc_528 N_A_109_47#_M1034_g N_X_c_962_n 0.00113891f $X=9.4 $Y=0.56 $X2=0 $Y2=0
cc_529 N_A_109_47#_c_324_n N_X_c_962_n 0.030582f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_530 N_A_109_47#_c_328_n N_X_c_962_n 0.00331919f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_531 N_A_109_47#_c_341_n N_X_c_979_n 0.00260297f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_532 N_A_109_47#_c_342_n N_X_c_979_n 0.00107777f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_533 N_A_109_47#_c_324_n N_X_c_979_n 0.0305808f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_534 N_A_109_47#_c_328_n N_X_c_979_n 0.0074788f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_535 N_A_109_47#_M1040_g N_X_c_963_n 0.0011682f $X=9.87 $Y=0.56 $X2=0 $Y2=0
cc_536 N_A_109_47#_c_324_n N_X_c_963_n 0.020973f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_537 N_A_109_47#_c_328_n N_X_c_963_n 0.00478914f $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_538 N_A_109_47#_M1041_g N_X_c_964_n 0.00298298f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_539 N_A_109_47#_c_344_n N_X_c_980_n 0.0175207f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_540 N_A_109_47#_c_328_n N_X_c_980_n 3.58038e-19 $X=10.365 $Y=1.217 $X2=0
+ $Y2=0
cc_541 N_A_109_47#_c_344_n N_X_c_981_n 0.00446503f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_542 N_A_109_47#_c_343_n X 0.00260297f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_543 N_A_109_47#_c_344_n X 0.00128868f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_544 N_A_109_47#_c_324_n X 0.0208858f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_545 N_A_109_47#_c_328_n X 0.00779663f $X=10.365 $Y=1.217 $X2=0 $Y2=0
cc_546 N_A_109_47#_c_344_n X 0.00133975f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_547 N_A_109_47#_M1041_g X 0.018747f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_548 N_A_109_47#_c_324_n X 0.00810115f $X=9.88 $Y=1.16 $X2=0 $Y2=0
cc_549 N_A_109_47#_c_342_n N_X_c_1178_n 8.07084e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_550 N_A_109_47#_c_343_n N_X_c_1178_n 0.0141618f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_551 N_A_109_47#_c_344_n N_X_c_1178_n 0.0124331f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_552 N_A_109_47#_c_318_n N_VGND_M1014_s 0.00251598f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_553 N_A_109_47#_c_320_n N_VGND_M1036_s 0.00251598f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_554 N_A_109_47#_c_321_n N_VGND_M1039_s 0.00193551f $X=2.99 $Y=0.82 $X2=0
+ $Y2=0
cc_555 N_A_109_47#_c_319_n N_VGND_c_1319_n 0.00787895f $X=0.895 $Y=0.82 $X2=0
+ $Y2=0
cc_556 N_A_109_47#_c_355_n N_VGND_c_1320_n 0.0216617f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_557 N_A_109_47#_c_318_n N_VGND_c_1320_n 0.00260082f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_558 N_A_109_47#_c_355_n N_VGND_c_1321_n 0.0186688f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_559 N_A_109_47#_c_318_n N_VGND_c_1321_n 0.0127122f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_560 N_A_109_47#_c_318_n N_VGND_c_1322_n 0.00193763f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_561 N_A_109_47#_c_377_n N_VGND_c_1322_n 0.0216617f $X=1.67 $Y=0.4 $X2=0 $Y2=0
cc_562 N_A_109_47#_c_320_n N_VGND_c_1322_n 0.00260082f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_563 N_A_109_47#_c_377_n N_VGND_c_1323_n 0.0186688f $X=1.67 $Y=0.4 $X2=0 $Y2=0
cc_564 N_A_109_47#_c_320_n N_VGND_c_1323_n 0.0127122f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_565 N_A_109_47#_M1005_g N_VGND_c_1324_n 0.00268723f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_566 N_A_109_47#_c_321_n N_VGND_c_1324_n 0.0135251f $X=2.99 $Y=0.82 $X2=0
+ $Y2=0
cc_567 N_A_109_47#_M1006_g N_VGND_c_1325_n 0.00382673f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_568 N_A_109_47#_M1007_g N_VGND_c_1325_n 0.00276126f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_569 N_A_109_47#_M1009_g N_VGND_c_1326_n 0.00382673f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_570 N_A_109_47#_M1012_g N_VGND_c_1326_n 0.00276126f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_571 N_A_109_47#_M1015_g N_VGND_c_1327_n 0.00382673f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_572 N_A_109_47#_M1019_g N_VGND_c_1327_n 0.00276126f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_573 N_A_109_47#_M1020_g N_VGND_c_1328_n 0.00390178f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_574 N_A_109_47#_M1021_g N_VGND_c_1328_n 0.00276126f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_575 N_A_109_47#_M1023_g N_VGND_c_1329_n 0.00390178f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_576 N_A_109_47#_M1024_g N_VGND_c_1329_n 0.00276126f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_577 N_A_109_47#_M1025_g N_VGND_c_1330_n 0.00390178f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_578 N_A_109_47#_M1029_g N_VGND_c_1330_n 0.00276126f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_579 N_A_109_47#_M1034_g N_VGND_c_1331_n 0.00390178f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_580 N_A_109_47#_M1040_g N_VGND_c_1331_n 0.00276126f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_581 N_A_109_47#_M1041_g N_VGND_c_1332_n 0.00438629f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_582 N_A_109_47#_c_320_n N_VGND_c_1333_n 0.00193763f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_583 N_A_109_47#_c_393_n N_VGND_c_1333_n 0.022456f $X=2.61 $Y=0.4 $X2=0 $Y2=0
cc_584 N_A_109_47#_c_321_n N_VGND_c_1333_n 0.00245178f $X=2.99 $Y=0.82 $X2=0
+ $Y2=0
cc_585 N_A_109_47#_M1005_g N_VGND_c_1335_n 0.00539841f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_586 N_A_109_47#_M1006_g N_VGND_c_1335_n 0.00423108f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_587 N_A_109_47#_M1007_g N_VGND_c_1337_n 0.00423108f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_588 N_A_109_47#_M1009_g N_VGND_c_1337_n 0.00423108f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_589 N_A_109_47#_M1012_g N_VGND_c_1339_n 0.00423108f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_590 N_A_109_47#_M1015_g N_VGND_c_1339_n 0.00423108f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_591 N_A_109_47#_M1019_g N_VGND_c_1341_n 0.00424619f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_592 N_A_109_47#_M1020_g N_VGND_c_1341_n 0.00424619f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_593 N_A_109_47#_M1021_g N_VGND_c_1343_n 0.00424619f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_594 N_A_109_47#_M1023_g N_VGND_c_1343_n 0.00424619f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_595 N_A_109_47#_M1024_g N_VGND_c_1345_n 0.00424619f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_596 N_A_109_47#_M1025_g N_VGND_c_1345_n 0.00424619f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_597 N_A_109_47#_M1029_g N_VGND_c_1347_n 0.00424619f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_598 N_A_109_47#_M1034_g N_VGND_c_1347_n 0.00424619f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_599 N_A_109_47#_M1040_g N_VGND_c_1349_n 0.00424619f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_600 N_A_109_47#_M1041_g N_VGND_c_1349_n 0.00439206f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_601 N_A_109_47#_M1011_d N_VGND_c_1352_n 0.00255524f $X=0.545 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_109_47#_M1028_d N_VGND_c_1352_n 0.00255524f $X=1.485 $Y=0.235 $X2=0
+ $Y2=0
cc_603 N_A_109_47#_M1038_d N_VGND_c_1352_n 0.00304616f $X=2.425 $Y=0.235 $X2=0
+ $Y2=0
cc_604 N_A_109_47#_M1005_g N_VGND_c_1352_n 0.00961873f $X=3.29 $Y=0.56 $X2=0
+ $Y2=0
cc_605 N_A_109_47#_M1006_g N_VGND_c_1352_n 0.00612203f $X=3.76 $Y=0.56 $X2=0
+ $Y2=0
cc_606 N_A_109_47#_M1007_g N_VGND_c_1352_n 0.00599926f $X=4.23 $Y=0.56 $X2=0
+ $Y2=0
cc_607 N_A_109_47#_M1009_g N_VGND_c_1352_n 0.00612203f $X=4.7 $Y=0.56 $X2=0
+ $Y2=0
cc_608 N_A_109_47#_M1012_g N_VGND_c_1352_n 0.00599926f $X=5.17 $Y=0.56 $X2=0
+ $Y2=0
cc_609 N_A_109_47#_M1015_g N_VGND_c_1352_n 0.00612203f $X=5.64 $Y=0.56 $X2=0
+ $Y2=0
cc_610 N_A_109_47#_M1019_g N_VGND_c_1352_n 0.00599018f $X=6.11 $Y=0.56 $X2=0
+ $Y2=0
cc_611 N_A_109_47#_M1020_g N_VGND_c_1352_n 0.00611295f $X=6.58 $Y=0.56 $X2=0
+ $Y2=0
cc_612 N_A_109_47#_M1021_g N_VGND_c_1352_n 0.00599018f $X=7.05 $Y=0.56 $X2=0
+ $Y2=0
cc_613 N_A_109_47#_M1023_g N_VGND_c_1352_n 0.00611295f $X=7.52 $Y=0.56 $X2=0
+ $Y2=0
cc_614 N_A_109_47#_M1024_g N_VGND_c_1352_n 0.00599018f $X=7.99 $Y=0.56 $X2=0
+ $Y2=0
cc_615 N_A_109_47#_M1025_g N_VGND_c_1352_n 0.00611295f $X=8.46 $Y=0.56 $X2=0
+ $Y2=0
cc_616 N_A_109_47#_M1029_g N_VGND_c_1352_n 0.00599018f $X=8.93 $Y=0.56 $X2=0
+ $Y2=0
cc_617 N_A_109_47#_M1034_g N_VGND_c_1352_n 0.00611295f $X=9.4 $Y=0.56 $X2=0
+ $Y2=0
cc_618 N_A_109_47#_M1040_g N_VGND_c_1352_n 0.00610552f $X=9.87 $Y=0.56 $X2=0
+ $Y2=0
cc_619 N_A_109_47#_M1041_g N_VGND_c_1352_n 0.00747968f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_620 N_A_109_47#_c_355_n N_VGND_c_1352_n 0.0140924f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_621 N_A_109_47#_c_318_n N_VGND_c_1352_n 0.00961016f $X=1.455 $Y=0.82 $X2=0
+ $Y2=0
cc_622 N_A_109_47#_c_377_n N_VGND_c_1352_n 0.0140924f $X=1.67 $Y=0.4 $X2=0 $Y2=0
cc_623 N_A_109_47#_c_320_n N_VGND_c_1352_n 0.00961016f $X=2.395 $Y=0.82 $X2=0
+ $Y2=0
cc_624 N_A_109_47#_c_393_n N_VGND_c_1352_n 0.0142976f $X=2.61 $Y=0.4 $X2=0 $Y2=0
cc_625 N_A_109_47#_c_321_n N_VGND_c_1352_n 0.00565014f $X=2.99 $Y=0.82 $X2=0
+ $Y2=0
cc_626 N_VPWR_c_761_n N_X_M1000_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_627 N_VPWR_c_761_n N_X_M1003_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_628 N_VPWR_c_761_n N_X_M1008_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_629 N_VPWR_c_761_n N_X_M1016_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_630 N_VPWR_c_761_n N_X_M1026_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_631 N_VPWR_c_761_n N_X_M1031_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_632 N_VPWR_c_761_n N_X_M1033_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_633 N_VPWR_c_761_n N_X_M1042_s 0.00231261f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_634 N_VPWR_c_768_n N_X_c_985_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_635 N_VPWR_c_769_n N_X_c_985_n 0.0385613f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_636 N_VPWR_c_779_n N_X_c_985_n 0.0223557f $X=3.935 $Y=2.72 $X2=0 $Y2=0
cc_637 N_VPWR_c_761_n N_X_c_985_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_638 N_VPWR_M1002_d N_X_c_966_n 0.00199888f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_639 N_VPWR_c_769_n N_X_c_966_n 0.0112848f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_640 N_VPWR_c_769_n N_X_c_1019_n 0.0470327f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_641 N_VPWR_c_770_n N_X_c_1019_n 0.0385613f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_642 N_VPWR_c_781_n N_X_c_1019_n 0.0223557f $X=4.875 $Y=2.72 $X2=0 $Y2=0
cc_643 N_VPWR_c_761_n N_X_c_1019_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_644 N_VPWR_M1004_d N_X_c_968_n 0.00199888f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_645 N_VPWR_c_770_n N_X_c_968_n 0.0112848f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_646 N_VPWR_c_770_n N_X_c_1037_n 0.0470327f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_647 N_VPWR_c_771_n N_X_c_1037_n 0.0385613f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_648 N_VPWR_c_783_n N_X_c_1037_n 0.0223557f $X=5.815 $Y=2.72 $X2=0 $Y2=0
cc_649 N_VPWR_c_761_n N_X_c_1037_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_650 N_VPWR_M1010_d N_X_c_969_n 0.00199888f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_651 N_VPWR_c_771_n N_X_c_969_n 0.0112848f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_652 N_VPWR_c_771_n N_X_c_1053_n 0.0470327f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_653 N_VPWR_c_772_n N_X_c_1053_n 0.0385613f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_654 N_VPWR_c_785_n N_X_c_1053_n 0.0223557f $X=6.755 $Y=2.72 $X2=0 $Y2=0
cc_655 N_VPWR_c_761_n N_X_c_1053_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_656 N_VPWR_M1018_d N_X_c_970_n 0.00199888f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_657 N_VPWR_c_772_n N_X_c_970_n 0.0112848f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_658 N_VPWR_c_772_n N_X_c_1069_n 0.0470327f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_659 N_VPWR_c_773_n N_X_c_1069_n 0.0385613f $X=7.78 $Y=2 $X2=0 $Y2=0
cc_660 N_VPWR_c_787_n N_X_c_1069_n 0.0223557f $X=7.695 $Y=2.72 $X2=0 $Y2=0
cc_661 N_VPWR_c_761_n N_X_c_1069_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_662 N_VPWR_M1027_d N_X_c_971_n 0.00199888f $X=7.635 $Y=1.485 $X2=0 $Y2=0
cc_663 N_VPWR_c_773_n N_X_c_971_n 0.0112848f $X=7.78 $Y=2 $X2=0 $Y2=0
cc_664 N_VPWR_c_773_n N_X_c_1085_n 0.0470327f $X=7.78 $Y=2 $X2=0 $Y2=0
cc_665 N_VPWR_c_774_n N_X_c_1085_n 0.0385613f $X=8.72 $Y=2 $X2=0 $Y2=0
cc_666 N_VPWR_c_789_n N_X_c_1085_n 0.0223557f $X=8.635 $Y=2.72 $X2=0 $Y2=0
cc_667 N_VPWR_c_761_n N_X_c_1085_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_668 N_VPWR_M1032_d N_X_c_972_n 0.00199888f $X=8.575 $Y=1.485 $X2=0 $Y2=0
cc_669 N_VPWR_c_774_n N_X_c_972_n 0.0112848f $X=8.72 $Y=2 $X2=0 $Y2=0
cc_670 N_VPWR_c_774_n N_X_c_1101_n 0.0470327f $X=8.72 $Y=2 $X2=0 $Y2=0
cc_671 N_VPWR_c_775_n N_X_c_1101_n 0.0385613f $X=9.66 $Y=2 $X2=0 $Y2=0
cc_672 N_VPWR_c_791_n N_X_c_1101_n 0.0223557f $X=9.575 $Y=2.72 $X2=0 $Y2=0
cc_673 N_VPWR_c_761_n N_X_c_1101_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_674 N_VPWR_M1035_d N_X_c_973_n 0.00199888f $X=9.515 $Y=1.485 $X2=0 $Y2=0
cc_675 N_VPWR_c_775_n N_X_c_973_n 0.0112848f $X=9.66 $Y=2 $X2=0 $Y2=0
cc_676 N_VPWR_M1043_d N_X_c_980_n 0.00140398f $X=10.455 $Y=1.485 $X2=0 $Y2=0
cc_677 N_VPWR_c_776_n N_X_c_980_n 0.00796332f $X=10.6 $Y=2 $X2=0 $Y2=0
cc_678 N_VPWR_M1043_d N_X_c_981_n 0.00310471f $X=10.455 $Y=1.485 $X2=0 $Y2=0
cc_679 N_VPWR_c_776_n N_X_c_981_n 0.0431348f $X=10.6 $Y=2 $X2=0 $Y2=0
cc_680 N_VPWR_c_795_n N_X_c_981_n 0.0117265f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_681 N_VPWR_c_761_n N_X_c_981_n 0.00992984f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_682 N_VPWR_c_775_n N_X_c_1178_n 0.0470327f $X=9.66 $Y=2 $X2=0 $Y2=0
cc_683 N_VPWR_c_776_n N_X_c_1178_n 0.0385613f $X=10.6 $Y=2 $X2=0 $Y2=0
cc_684 N_VPWR_c_793_n N_X_c_1178_n 0.0223557f $X=10.515 $Y=2.72 $X2=0 $Y2=0
cc_685 N_VPWR_c_761_n N_X_c_1178_n 0.0140101f $X=11.27 $Y=2.72 $X2=0 $Y2=0
cc_686 N_X_c_948_n N_VGND_M1006_s 0.00251598f $X=4.275 $Y=0.82 $X2=0 $Y2=0
cc_687 N_X_c_950_n N_VGND_M1009_s 0.00251598f $X=5.215 $Y=0.82 $X2=0 $Y2=0
cc_688 N_X_c_951_n N_VGND_M1015_s 0.00251598f $X=6.155 $Y=0.82 $X2=0 $Y2=0
cc_689 N_X_c_952_n N_VGND_M1020_s 0.00251598f $X=7.095 $Y=0.82 $X2=0 $Y2=0
cc_690 N_X_c_953_n N_VGND_M1023_s 0.00251598f $X=8.035 $Y=0.82 $X2=0 $Y2=0
cc_691 N_X_c_954_n N_VGND_M1025_s 0.00251598f $X=8.975 $Y=0.82 $X2=0 $Y2=0
cc_692 N_X_c_955_n N_VGND_M1034_s 0.00251598f $X=9.915 $Y=0.82 $X2=0 $Y2=0
cc_693 N_X_c_956_n N_VGND_M1041_s 0.00116312f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_694 N_X_c_964_n N_VGND_M1041_s 0.00200806f $X=10.885 $Y=0.82 $X2=0 $Y2=0
cc_695 N_X_c_986_n N_VGND_c_1325_n 0.0116752f $X=3.525 $Y=0.45 $X2=0 $Y2=0
cc_696 N_X_c_984_n N_VGND_c_1325_n 0.00700786f $X=3.525 $Y=0.735 $X2=0 $Y2=0
cc_697 N_X_c_948_n N_VGND_c_1325_n 0.0127122f $X=4.275 $Y=0.82 $X2=0 $Y2=0
cc_698 N_X_c_1013_n N_VGND_c_1326_n 0.0116752f $X=4.465 $Y=0.45 $X2=0 $Y2=0
cc_699 N_X_c_1015_n N_VGND_c_1326_n 0.00700786f $X=4.465 $Y=0.735 $X2=0 $Y2=0
cc_700 N_X_c_950_n N_VGND_c_1326_n 0.0127122f $X=5.215 $Y=0.82 $X2=0 $Y2=0
cc_701 N_X_c_1031_n N_VGND_c_1327_n 0.0116752f $X=5.405 $Y=0.45 $X2=0 $Y2=0
cc_702 N_X_c_1033_n N_VGND_c_1327_n 0.00700786f $X=5.405 $Y=0.735 $X2=0 $Y2=0
cc_703 N_X_c_951_n N_VGND_c_1327_n 0.0127122f $X=6.155 $Y=0.82 $X2=0 $Y2=0
cc_704 N_X_c_1049_n N_VGND_c_1328_n 0.0186688f $X=6.37 $Y=0.4 $X2=0 $Y2=0
cc_705 N_X_c_952_n N_VGND_c_1328_n 0.0127122f $X=7.095 $Y=0.82 $X2=0 $Y2=0
cc_706 N_X_c_1065_n N_VGND_c_1329_n 0.0186688f $X=7.31 $Y=0.4 $X2=0 $Y2=0
cc_707 N_X_c_953_n N_VGND_c_1329_n 0.0127122f $X=8.035 $Y=0.82 $X2=0 $Y2=0
cc_708 N_X_c_1081_n N_VGND_c_1330_n 0.0186688f $X=8.25 $Y=0.4 $X2=0 $Y2=0
cc_709 N_X_c_954_n N_VGND_c_1330_n 0.0127122f $X=8.975 $Y=0.82 $X2=0 $Y2=0
cc_710 N_X_c_1097_n N_VGND_c_1331_n 0.0186688f $X=9.19 $Y=0.4 $X2=0 $Y2=0
cc_711 N_X_c_955_n N_VGND_c_1331_n 0.0127122f $X=9.915 $Y=0.82 $X2=0 $Y2=0
cc_712 N_X_c_956_n N_VGND_c_1332_n 0.00883327f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_713 N_X_c_964_n N_VGND_c_1332_n 0.0192925f $X=10.885 $Y=0.82 $X2=0 $Y2=0
cc_714 N_X_c_986_n N_VGND_c_1335_n 0.0223797f $X=3.525 $Y=0.45 $X2=0 $Y2=0
cc_715 N_X_c_948_n N_VGND_c_1335_n 0.00260082f $X=4.275 $Y=0.82 $X2=0 $Y2=0
cc_716 N_X_c_948_n N_VGND_c_1337_n 0.00193763f $X=4.275 $Y=0.82 $X2=0 $Y2=0
cc_717 N_X_c_1013_n N_VGND_c_1337_n 0.0221615f $X=4.465 $Y=0.45 $X2=0 $Y2=0
cc_718 N_X_c_950_n N_VGND_c_1337_n 0.00260082f $X=5.215 $Y=0.82 $X2=0 $Y2=0
cc_719 N_X_c_950_n N_VGND_c_1339_n 0.00193763f $X=5.215 $Y=0.82 $X2=0 $Y2=0
cc_720 N_X_c_1031_n N_VGND_c_1339_n 0.0221615f $X=5.405 $Y=0.45 $X2=0 $Y2=0
cc_721 N_X_c_951_n N_VGND_c_1339_n 0.00260082f $X=6.155 $Y=0.82 $X2=0 $Y2=0
cc_722 N_X_c_951_n N_VGND_c_1341_n 0.00193763f $X=6.155 $Y=0.82 $X2=0 $Y2=0
cc_723 N_X_c_1049_n N_VGND_c_1341_n 0.0216617f $X=6.37 $Y=0.4 $X2=0 $Y2=0
cc_724 N_X_c_952_n N_VGND_c_1341_n 0.00260082f $X=7.095 $Y=0.82 $X2=0 $Y2=0
cc_725 N_X_c_952_n N_VGND_c_1343_n 0.00193763f $X=7.095 $Y=0.82 $X2=0 $Y2=0
cc_726 N_X_c_1065_n N_VGND_c_1343_n 0.0216617f $X=7.31 $Y=0.4 $X2=0 $Y2=0
cc_727 N_X_c_953_n N_VGND_c_1343_n 0.00260082f $X=8.035 $Y=0.82 $X2=0 $Y2=0
cc_728 N_X_c_953_n N_VGND_c_1345_n 0.00193763f $X=8.035 $Y=0.82 $X2=0 $Y2=0
cc_729 N_X_c_1081_n N_VGND_c_1345_n 0.0216617f $X=8.25 $Y=0.4 $X2=0 $Y2=0
cc_730 N_X_c_954_n N_VGND_c_1345_n 0.00260082f $X=8.975 $Y=0.82 $X2=0 $Y2=0
cc_731 N_X_c_954_n N_VGND_c_1347_n 0.00193763f $X=8.975 $Y=0.82 $X2=0 $Y2=0
cc_732 N_X_c_1097_n N_VGND_c_1347_n 0.0216617f $X=9.19 $Y=0.4 $X2=0 $Y2=0
cc_733 N_X_c_955_n N_VGND_c_1347_n 0.00260082f $X=9.915 $Y=0.82 $X2=0 $Y2=0
cc_734 N_X_c_955_n N_VGND_c_1349_n 0.00193763f $X=9.915 $Y=0.82 $X2=0 $Y2=0
cc_735 N_X_c_1113_n N_VGND_c_1349_n 0.022456f $X=10.13 $Y=0.4 $X2=0 $Y2=0
cc_736 N_X_c_956_n N_VGND_c_1349_n 0.00248202f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_737 N_X_c_964_n N_VGND_c_1351_n 0.0143833f $X=10.885 $Y=0.82 $X2=0 $Y2=0
cc_738 N_X_M1005_d N_VGND_c_1352_n 0.00255377f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_739 N_X_M1007_d N_VGND_c_1352_n 0.00255431f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_740 N_X_M1012_d N_VGND_c_1352_n 0.00255431f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_741 N_X_M1019_d N_VGND_c_1352_n 0.00255524f $X=6.185 $Y=0.235 $X2=0 $Y2=0
cc_742 N_X_M1021_d N_VGND_c_1352_n 0.00255524f $X=7.125 $Y=0.235 $X2=0 $Y2=0
cc_743 N_X_M1024_d N_VGND_c_1352_n 0.00255524f $X=8.065 $Y=0.235 $X2=0 $Y2=0
cc_744 N_X_M1029_d N_VGND_c_1352_n 0.00255524f $X=9.005 $Y=0.235 $X2=0 $Y2=0
cc_745 N_X_M1040_d N_VGND_c_1352_n 0.00304616f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_746 N_X_c_986_n N_VGND_c_1352_n 0.0141899f $X=3.525 $Y=0.45 $X2=0 $Y2=0
cc_747 N_X_c_948_n N_VGND_c_1352_n 0.00961016f $X=4.275 $Y=0.82 $X2=0 $Y2=0
cc_748 N_X_c_1013_n N_VGND_c_1352_n 0.0141768f $X=4.465 $Y=0.45 $X2=0 $Y2=0
cc_749 N_X_c_950_n N_VGND_c_1352_n 0.00961016f $X=5.215 $Y=0.82 $X2=0 $Y2=0
cc_750 N_X_c_1031_n N_VGND_c_1352_n 0.0141768f $X=5.405 $Y=0.45 $X2=0 $Y2=0
cc_751 N_X_c_951_n N_VGND_c_1352_n 0.00961016f $X=6.155 $Y=0.82 $X2=0 $Y2=0
cc_752 N_X_c_1049_n N_VGND_c_1352_n 0.0140924f $X=6.37 $Y=0.4 $X2=0 $Y2=0
cc_753 N_X_c_952_n N_VGND_c_1352_n 0.00961016f $X=7.095 $Y=0.82 $X2=0 $Y2=0
cc_754 N_X_c_1065_n N_VGND_c_1352_n 0.0140924f $X=7.31 $Y=0.4 $X2=0 $Y2=0
cc_755 N_X_c_953_n N_VGND_c_1352_n 0.00961016f $X=8.035 $Y=0.82 $X2=0 $Y2=0
cc_756 N_X_c_1081_n N_VGND_c_1352_n 0.0140924f $X=8.25 $Y=0.4 $X2=0 $Y2=0
cc_757 N_X_c_954_n N_VGND_c_1352_n 0.00961016f $X=8.975 $Y=0.82 $X2=0 $Y2=0
cc_758 N_X_c_1097_n N_VGND_c_1352_n 0.0140924f $X=9.19 $Y=0.4 $X2=0 $Y2=0
cc_759 N_X_c_955_n N_VGND_c_1352_n 0.00961016f $X=9.915 $Y=0.82 $X2=0 $Y2=0
cc_760 N_X_c_1113_n N_VGND_c_1352_n 0.0142976f $X=10.13 $Y=0.4 $X2=0 $Y2=0
cc_761 N_X_c_956_n N_VGND_c_1352_n 0.00537127f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_762 N_X_c_964_n N_VGND_c_1352_n 0.0150416f $X=10.885 $Y=0.82 $X2=0 $Y2=0
