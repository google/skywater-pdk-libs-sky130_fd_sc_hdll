* File: sky130_fd_sc_hdll__bufbuf_8.pxi.spice
* Created: Wed Sep  2 08:24:51 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%A N_A_c_129_n N_A_M1010_g N_A_M1018_g A
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%A
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1010_s
+ N_A_27_47#_c_156_n N_A_27_47#_M1021_g N_A_27_47#_c_157_n N_A_27_47#_M1024_g
+ N_A_27_47#_c_158_n N_A_27_47#_c_163_n N_A_27_47#_c_159_n N_A_27_47#_c_160_n
+ N_A_27_47#_c_164_n N_A_27_47#_c_165_n N_A_27_47#_c_161_n
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_224_297# N_A_224_297#_M1024_d
+ N_A_224_297#_M1021_d N_A_224_297#_M1005_g N_A_224_297#_c_228_n
+ N_A_224_297#_M1009_g N_A_224_297#_M1011_g N_A_224_297#_c_229_n
+ N_A_224_297#_M1014_g N_A_224_297#_c_230_n N_A_224_297#_M1017_g
+ N_A_224_297#_M1012_g N_A_224_297#_c_231_n N_A_224_297#_c_222_n
+ N_A_224_297#_c_223_n N_A_224_297#_c_224_n N_A_224_297#_c_232_n
+ N_A_224_297#_c_225_n N_A_224_297#_c_226_n N_A_224_297#_c_227_n
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_224_297#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_338_47# N_A_338_47#_M1005_s
+ N_A_338_47#_M1011_s N_A_338_47#_M1009_s N_A_338_47#_M1014_s
+ N_A_338_47#_M1001_g N_A_338_47#_c_342_n N_A_338_47#_M1000_g
+ N_A_338_47#_M1003_g N_A_338_47#_c_343_n N_A_338_47#_M1002_g
+ N_A_338_47#_M1006_g N_A_338_47#_c_344_n N_A_338_47#_M1004_g
+ N_A_338_47#_M1007_g N_A_338_47#_c_345_n N_A_338_47#_M1008_g
+ N_A_338_47#_M1013_g N_A_338_47#_c_346_n N_A_338_47#_M1016_g
+ N_A_338_47#_M1015_g N_A_338_47#_c_347_n N_A_338_47#_M1019_g
+ N_A_338_47#_M1020_g N_A_338_47#_c_348_n N_A_338_47#_M1022_g
+ N_A_338_47#_c_349_n N_A_338_47#_M1025_g N_A_338_47#_M1023_g
+ N_A_338_47#_c_332_n N_A_338_47#_c_350_n N_A_338_47#_c_333_n
+ N_A_338_47#_c_334_n N_A_338_47#_c_351_n N_A_338_47#_c_352_n
+ N_A_338_47#_c_380_n N_A_338_47#_c_382_n N_A_338_47#_c_335_n
+ N_A_338_47#_c_353_n N_A_338_47#_c_336_n N_A_338_47#_c_337_n
+ N_A_338_47#_c_338_n N_A_338_47#_c_339_n N_A_338_47#_c_355_n
+ N_A_338_47#_c_340_n N_A_338_47#_c_341_n
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%A_338_47#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%VPWR N_VPWR_M1010_d N_VPWR_M1009_d
+ N_VPWR_M1017_d N_VPWR_M1002_d N_VPWR_M1008_d N_VPWR_M1019_d N_VPWR_M1025_d
+ N_VPWR_c_567_n N_VPWR_c_568_n N_VPWR_c_569_n N_VPWR_c_570_n N_VPWR_c_571_n
+ N_VPWR_c_572_n N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n
+ N_VPWR_c_577_n N_VPWR_c_578_n N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n
+ N_VPWR_c_582_n N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n VPWR
+ N_VPWR_c_586_n N_VPWR_c_566_n N_VPWR_c_588_n
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%VPWR
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%X N_X_M1001_s N_X_M1006_s N_X_M1013_s
+ N_X_M1020_s N_X_M1000_s N_X_M1004_s N_X_M1016_s N_X_M1022_s N_X_c_697_n
+ N_X_c_698_n N_X_c_679_n N_X_c_680_n N_X_c_688_n N_X_c_689_n N_X_c_724_n
+ N_X_c_728_n N_X_c_681_n N_X_c_690_n N_X_c_740_n N_X_c_744_n N_X_c_682_n
+ N_X_c_691_n N_X_c_756_n N_X_c_758_n N_X_c_683_n N_X_c_762_n N_X_c_684_n
+ N_X_c_692_n N_X_c_685_n N_X_c_693_n N_X_c_686_n N_X_c_694_n X X
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%X
x_PM_SKY130_FD_SC_HDLL__BUFBUF_8%VGND N_VGND_M1018_d N_VGND_M1005_d
+ N_VGND_M1012_d N_VGND_M1003_d N_VGND_M1007_d N_VGND_M1015_d N_VGND_M1023_d
+ N_VGND_c_850_n N_VGND_c_851_n N_VGND_c_852_n N_VGND_c_853_n N_VGND_c_854_n
+ N_VGND_c_855_n N_VGND_c_856_n N_VGND_c_857_n N_VGND_c_858_n N_VGND_c_859_n
+ N_VGND_c_860_n N_VGND_c_861_n N_VGND_c_862_n N_VGND_c_863_n N_VGND_c_864_n
+ N_VGND_c_865_n N_VGND_c_866_n N_VGND_c_867_n N_VGND_c_868_n VGND
+ N_VGND_c_869_n N_VGND_c_870_n N_VGND_c_871_n VGND
+ PM_SKY130_FD_SC_HDLL__BUFBUF_8%VGND
cc_1 VNB N_A_c_129_n 0.04124f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_M1018_g 0.0367557f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_3 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_27_47#_c_156_n 0.0272708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_c_157_n 0.0204744f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_6 VNB N_A_27_47#_c_158_n 0.0197452f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_159_n 0.00207587f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_160_n 0.00999162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_161_n 0.00963657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_224_297#_M1005_g 0.0221051f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_224_297#_M1011_g 0.0188756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_224_297#_M1012_g 0.0185511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_224_297#_c_222_n 0.00539764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_224_297#_c_223_n 0.0194792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_224_297#_c_224_n 0.00656524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_224_297#_c_225_n 7.03049e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_224_297#_c_226_n 0.00238516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_224_297#_c_227_n 0.0683671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_338_47#_M1001_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_338_47#_M1003_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_338_47#_M1006_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_338_47#_M1007_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_338_47#_M1013_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_338_47#_M1015_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_338_47#_M1020_g 0.0188736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_338_47#_M1023_g 0.0218008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_338_47#_c_332_n 0.00443915f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_338_47#_c_333_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_338_47#_c_334_n 0.00437286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_338_47#_c_335_n 0.00102469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_338_47#_c_336_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_338_47#_c_337_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_338_47#_c_338_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_338_47#_c_339_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_338_47#_c_340_n 0.00153756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_338_47#_c_341_n 0.185241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_566_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_679_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_680_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_681_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_X_c_682_n 0.00327828f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_X_c_683_n 0.0101105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_X_c_684_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_X_c_685_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_X_c_686_n 0.00358644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB X 0.0233377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_850_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_851_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_852_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_853_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_854_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_855_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_856_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_857_n 0.0359836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_858_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_859_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_860_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_861_n 0.0200002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_862_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_863_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_864_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_865_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_866_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_867_n 0.0194238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_868_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_869_n 0.0107554f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_870_n 0.363129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_871_n 0.0220461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VPB N_A_c_129_n 0.0391619f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_70 VPB N_A_27_47#_c_156_n 0.0335377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_163_n 0.0248879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_164_n 9.24119e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_165_n 0.00922579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_161_n 0.00606227f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_224_297#_c_228_n 0.0194229f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_76 VPB N_A_224_297#_c_229_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_224_297#_c_230_n 0.0159693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_224_297#_c_231_n 0.00804088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_224_297#_c_232_n 0.00225685f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_224_297#_c_225_n 0.00522453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_224_297#_c_227_n 0.0202804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_338_47#_c_342_n 0.0162292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_338_47#_c_343_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_338_47#_c_344_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_338_47#_c_345_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_338_47#_c_346_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_338_47#_c_347_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_338_47#_c_348_n 0.0158854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_338_47#_c_349_n 0.0191589f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_338_47#_c_350_n 0.00775188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_338_47#_c_351_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_A_338_47#_c_352_n 0.00452041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_338_47#_c_353_n 0.00100785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_338_47#_c_337_n 0.00252324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_338_47#_c_355_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_338_47#_c_341_n 0.0514147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_567_n 0.0139383f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_568_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_569_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_570_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_571_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_572_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_573_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_574_n 0.0366293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_575_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_576_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_577_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_578_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_579_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_580_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_581_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_582_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_583_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_584_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_585_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_586_n 0.0113717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_566_n 0.0673257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_588_n 0.024218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_X_c_688_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_X_c_689_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_X_c_690_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_X_c_691_n 0.00227769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_X_c_692_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_X_c_693_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_X_c_694_n 0.0022912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB X 0.00778049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB X 0.0131281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 N_A_c_129_n N_A_27_47#_c_156_n 0.037158f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_M1018_g N_A_27_47#_c_157_n 0.0193849f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_130 N_A_M1018_g N_A_27_47#_c_158_n 0.0027061f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_c_129_n N_A_27_47#_c_163_n 0.00873793f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_129_n N_A_27_47#_c_159_n 5.98433e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_M1018_g N_A_27_47#_c_159_n 0.0153935f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_134 A N_A_27_47#_c_159_n 0.001048f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A_c_129_n N_A_27_47#_c_160_n 0.00815792f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_136 A N_A_27_47#_c_160_n 0.0255682f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_137 N_A_c_129_n N_A_27_47#_c_164_n 0.0153477f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 A N_A_27_47#_c_164_n 9.95686e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_139 N_A_c_129_n N_A_27_47#_c_165_n 0.00871413f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 A N_A_27_47#_c_165_n 0.0257053f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A_M1018_g N_A_27_47#_c_161_n 0.0085617f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_142 A N_A_27_47#_c_161_n 0.0134215f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_M1018_g N_A_224_297#_c_224_n 6.82563e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_c_129_n N_A_224_297#_c_232_n 6.91288e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_129_n N_VPWR_c_567_n 0.00385319f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_129_n N_VPWR_c_566_n 0.00569968f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_129_n N_VPWR_c_588_n 0.00504659f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_M1018_g N_VGND_c_850_n 0.0028527f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_M1018_g N_VGND_c_870_n 0.00727708f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_M1018_g N_VGND_c_871_n 0.00439206f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_156_n N_A_224_297#_c_231_n 0.0118703f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_156_n N_A_224_297#_c_222_n 0.0019049f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_157_n N_A_224_297#_c_222_n 0.0027278f $X=1.055 $Y=0.995
+ $X2=0 $Y2=0
cc_154 N_A_27_47#_c_161_n N_A_224_297#_c_222_n 0.0127323f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_27_47#_c_156_n N_A_224_297#_c_224_n 0.0010811f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_157_n N_A_224_297#_c_224_n 0.0118137f $X=1.055 $Y=0.995
+ $X2=0 $Y2=0
cc_157 N_A_27_47#_c_158_n N_A_224_297#_c_224_n 0.00353949f $X=0.26 $Y=0.47 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_161_n N_A_224_297#_c_224_n 0.0127906f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_27_47#_c_156_n N_A_224_297#_c_232_n 0.00680279f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_163_n N_A_224_297#_c_232_n 0.00438999f $X=0.26 $Y=1.63 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_161_n N_A_224_297#_c_232_n 0.0099038f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_156_n N_A_224_297#_c_225_n 0.00514298f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_161_n N_A_224_297#_c_225_n 0.0123099f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_156_n N_A_224_297#_c_226_n 0.00496073f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_A_27_47#_c_161_n N_A_224_297#_c_226_n 0.0173927f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_161_n N_VPWR_M1010_d 0.00427994f $X=1.005 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_27_47#_c_156_n N_VPWR_c_567_n 0.0128344f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_163_n N_VPWR_c_567_n 0.0227518f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_164_n N_VPWR_c_567_n 0.00110254f $X=0.66 $Y=1.53 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_161_n N_VPWR_c_567_n 0.0138849f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_156_n N_VPWR_c_574_n 0.00597712f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_156_n N_VPWR_c_566_n 0.0127841f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_163_n N_VPWR_c_566_n 0.0104244f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_163_n N_VPWR_c_588_n 0.00783104f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_161_n N_VGND_M1018_d 0.00377317f $X=1.005 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_27_47#_c_157_n N_VGND_c_850_n 0.00504453f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_177 N_A_27_47#_c_159_n N_VGND_c_850_n 8.13279e-19 $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_161_n N_VGND_c_850_n 0.0133682f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_157_n N_VGND_c_857_n 0.00466005f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_161_n N_VGND_c_857_n 2.28683e-19 $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1018_s N_VGND_c_870_n 0.00260708f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_157_n N_VGND_c_870_n 0.00947228f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_158_n N_VGND_c_870_n 0.0125844f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_159_n N_VGND_c_870_n 0.00502579f $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_161_n N_VGND_c_870_n 0.00111682f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_158_n N_VGND_c_871_n 0.0211122f $X=0.26 $Y=0.47 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_159_n N_VGND_c_871_n 0.00299761f $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_188 N_A_224_297#_M1012_g N_A_338_47#_M1001_g 0.0207193f $X=3.015 $Y=0.56
+ $X2=0 $Y2=0
cc_189 N_A_224_297#_c_230_n N_A_338_47#_c_342_n 0.0215651f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_224_297#_M1005_g N_A_338_47#_c_332_n 0.00693104f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_191 N_A_224_297#_M1011_g N_A_338_47#_c_332_n 5.47935e-19 $X=2.495 $Y=0.56
+ $X2=0 $Y2=0
cc_192 N_A_224_297#_c_224_n N_A_338_47#_c_332_n 0.0403182f $X=1.265 $Y=0.4 $X2=0
+ $Y2=0
cc_193 N_A_224_297#_c_228_n N_A_338_47#_c_350_n 0.0112091f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_224_297#_c_229_n N_A_338_47#_c_350_n 7.06303e-19 $X=2.52 $Y=1.41
+ $X2=0 $Y2=0
cc_195 N_A_224_297#_c_232_n N_A_338_47#_c_350_n 0.0721381f $X=1.265 $Y=1.63
+ $X2=0 $Y2=0
cc_196 N_A_224_297#_M1005_g N_A_338_47#_c_333_n 0.00879805f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_197 N_A_224_297#_M1011_g N_A_338_47#_c_333_n 0.00879805f $X=2.495 $Y=0.56
+ $X2=0 $Y2=0
cc_198 N_A_224_297#_c_223_n N_A_338_47#_c_333_n 0.03957f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_224_297#_c_227_n N_A_338_47#_c_333_n 0.0031956f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_200 N_A_224_297#_M1005_g N_A_338_47#_c_334_n 0.00126794f $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_201 N_A_224_297#_c_223_n N_A_338_47#_c_334_n 0.0278128f $X=2.625 $Y=1.16
+ $X2=0 $Y2=0
cc_202 N_A_224_297#_c_224_n N_A_338_47#_c_334_n 0.0148339f $X=1.265 $Y=0.4 $X2=0
+ $Y2=0
cc_203 N_A_224_297#_c_228_n N_A_338_47#_c_351_n 0.0137916f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_224_297#_c_229_n N_A_338_47#_c_351_n 0.0101048f $X=2.52 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_224_297#_c_223_n N_A_338_47#_c_351_n 0.0394547f $X=2.625 $Y=1.16
+ $X2=0 $Y2=0
cc_206 N_A_224_297#_c_227_n N_A_338_47#_c_351_n 0.00720931f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_207 N_A_224_297#_c_228_n N_A_338_47#_c_352_n 0.00138874f $X=2.05 $Y=1.41
+ $X2=0 $Y2=0
cc_208 N_A_224_297#_c_223_n N_A_338_47#_c_352_n 0.0279779f $X=2.625 $Y=1.16
+ $X2=0 $Y2=0
cc_209 N_A_224_297#_c_225_n N_A_338_47#_c_352_n 0.0147198f $X=1.265 $Y=1.545
+ $X2=0 $Y2=0
cc_210 N_A_224_297#_c_227_n N_A_338_47#_c_352_n 3.20658e-19 $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_211 N_A_224_297#_M1005_g N_A_338_47#_c_380_n 5.25882e-19 $X=2.025 $Y=0.56
+ $X2=0 $Y2=0
cc_212 N_A_224_297#_M1011_g N_A_338_47#_c_380_n 0.00657592f $X=2.495 $Y=0.56
+ $X2=0 $Y2=0
cc_213 N_A_224_297#_c_228_n N_A_338_47#_c_382_n 7.33057e-19 $X=2.05 $Y=1.41
+ $X2=0 $Y2=0
cc_214 N_A_224_297#_c_229_n N_A_338_47#_c_382_n 0.0137692f $X=2.52 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_224_297#_c_230_n N_A_338_47#_c_382_n 0.0112091f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_224_297#_M1012_g N_A_338_47#_c_335_n 0.0116573f $X=3.015 $Y=0.56
+ $X2=0 $Y2=0
cc_217 N_A_224_297#_c_230_n N_A_338_47#_c_353_n 0.0151183f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_224_297#_c_227_n N_A_338_47#_c_353_n 3.58038e-19 $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_219 N_A_224_297#_M1012_g N_A_338_47#_c_336_n 0.00410511f $X=3.015 $Y=0.56
+ $X2=0 $Y2=0
cc_220 N_A_224_297#_c_230_n N_A_338_47#_c_337_n 8.16926e-19 $X=2.99 $Y=1.41
+ $X2=0 $Y2=0
cc_221 N_A_224_297#_c_227_n N_A_338_47#_c_337_n 0.00327205f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_222 N_A_224_297#_M1011_g N_A_338_47#_c_339_n 0.0011682f $X=2.495 $Y=0.56
+ $X2=0 $Y2=0
cc_223 N_A_224_297#_c_223_n N_A_338_47#_c_339_n 0.0307156f $X=2.625 $Y=1.16
+ $X2=0 $Y2=0
cc_224 N_A_224_297#_c_227_n N_A_338_47#_c_339_n 0.00450461f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_225 N_A_224_297#_c_229_n N_A_338_47#_c_355_n 0.00259297f $X=2.52 $Y=1.41
+ $X2=0 $Y2=0
cc_226 N_A_224_297#_c_230_n N_A_338_47#_c_355_n 0.00107777f $X=2.99 $Y=1.41
+ $X2=0 $Y2=0
cc_227 N_A_224_297#_c_223_n N_A_338_47#_c_355_n 0.0305808f $X=2.625 $Y=1.16
+ $X2=0 $Y2=0
cc_228 N_A_224_297#_c_227_n N_A_338_47#_c_355_n 0.00723098f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_229 N_A_224_297#_c_223_n N_A_338_47#_c_340_n 0.014524f $X=2.625 $Y=1.16 $X2=0
+ $Y2=0
cc_230 N_A_224_297#_c_227_n N_A_338_47#_c_340_n 0.00220849f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_231 N_A_224_297#_c_227_n N_A_338_47#_c_341_n 0.0207193f $X=2.99 $Y=1.217
+ $X2=0 $Y2=0
cc_232 N_A_224_297#_c_231_n N_VPWR_c_567_n 0.039955f $X=1.265 $Y=2.31 $X2=0
+ $Y2=0
cc_233 N_A_224_297#_c_228_n N_VPWR_c_568_n 0.00547044f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_224_297#_c_229_n N_VPWR_c_568_n 0.00497803f $X=2.52 $Y=1.41 $X2=0
+ $Y2=0
cc_235 N_A_224_297#_c_230_n N_VPWR_c_569_n 0.00547044f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_224_297#_c_228_n N_VPWR_c_574_n 0.00673617f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_237 N_A_224_297#_c_231_n N_VPWR_c_574_n 0.0280533f $X=1.265 $Y=2.31 $X2=0
+ $Y2=0
cc_238 N_A_224_297#_c_229_n N_VPWR_c_576_n 0.00597712f $X=2.52 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_224_297#_c_230_n N_VPWR_c_576_n 0.00673617f $X=2.99 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_A_224_297#_M1021_d N_VPWR_c_566_n 0.00217517f $X=1.12 $Y=1.485 $X2=0
+ $Y2=0
cc_241 N_A_224_297#_c_228_n N_VPWR_c_566_n 0.0131262f $X=2.05 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_224_297#_c_229_n N_VPWR_c_566_n 0.00999457f $X=2.52 $Y=1.41 $X2=0
+ $Y2=0
cc_243 N_A_224_297#_c_230_n N_VPWR_c_566_n 0.011869f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_224_297#_c_231_n N_VPWR_c_566_n 0.016095f $X=1.265 $Y=2.31 $X2=0
+ $Y2=0
cc_245 N_A_224_297#_M1012_g N_X_c_697_n 5.33681e-19 $X=3.015 $Y=0.56 $X2=0 $Y2=0
cc_246 N_A_224_297#_c_230_n N_X_c_698_n 7.33057e-19 $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_224_297#_c_224_n N_VGND_c_850_n 0.0179214f $X=1.265 $Y=0.4 $X2=0
+ $Y2=0
cc_248 N_A_224_297#_M1005_g N_VGND_c_851_n 0.00390178f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_249 N_A_224_297#_M1011_g N_VGND_c_851_n 0.00276126f $X=2.495 $Y=0.56 $X2=0
+ $Y2=0
cc_250 N_A_224_297#_M1012_g N_VGND_c_852_n 0.00268723f $X=3.015 $Y=0.56 $X2=0
+ $Y2=0
cc_251 N_A_224_297#_M1005_g N_VGND_c_857_n 0.00424619f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_252 N_A_224_297#_c_224_n N_VGND_c_857_n 0.0269844f $X=1.265 $Y=0.4 $X2=0
+ $Y2=0
cc_253 N_A_224_297#_M1011_g N_VGND_c_859_n 0.00424619f $X=2.495 $Y=0.56 $X2=0
+ $Y2=0
cc_254 N_A_224_297#_M1012_g N_VGND_c_859_n 0.00439206f $X=3.015 $Y=0.56 $X2=0
+ $Y2=0
cc_255 N_A_224_297#_M1024_d N_VGND_c_870_n 0.0020946f $X=1.13 $Y=0.235 $X2=0
+ $Y2=0
cc_256 N_A_224_297#_M1005_g N_VGND_c_870_n 0.00731205f $X=2.025 $Y=0.56 $X2=0
+ $Y2=0
cc_257 N_A_224_297#_M1011_g N_VGND_c_870_n 0.00610552f $X=2.495 $Y=0.56 $X2=0
+ $Y2=0
cc_258 N_A_224_297#_M1012_g N_VGND_c_870_n 0.00618081f $X=3.015 $Y=0.56 $X2=0
+ $Y2=0
cc_259 N_A_224_297#_c_224_n N_VGND_c_870_n 0.0159615f $X=1.265 $Y=0.4 $X2=0
+ $Y2=0
cc_260 N_A_338_47#_c_351_n N_VPWR_M1009_d 0.00178587f $X=2.54 $Y=1.53 $X2=0
+ $Y2=0
cc_261 N_A_338_47#_c_353_n N_VPWR_M1017_d 0.00324655f $X=3.14 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_A_338_47#_c_350_n N_VPWR_c_568_n 0.0411685f $X=1.815 $Y=1.63 $X2=0
+ $Y2=0
cc_263 N_A_338_47#_c_351_n N_VPWR_c_568_n 0.0136682f $X=2.54 $Y=1.53 $X2=0 $Y2=0
cc_264 N_A_338_47#_c_382_n N_VPWR_c_568_n 0.0507655f $X=2.755 $Y=1.63 $X2=0
+ $Y2=0
cc_265 N_A_338_47#_c_342_n N_VPWR_c_569_n 0.00497803f $X=3.46 $Y=1.41 $X2=0
+ $Y2=0
cc_266 N_A_338_47#_c_382_n N_VPWR_c_569_n 0.0416217f $X=2.755 $Y=1.63 $X2=0
+ $Y2=0
cc_267 N_A_338_47#_c_353_n N_VPWR_c_569_n 0.0151472f $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_268 N_A_338_47#_c_343_n N_VPWR_c_570_n 0.0052072f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_338_47#_c_344_n N_VPWR_c_570_n 0.004751f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_338_47#_c_345_n N_VPWR_c_571_n 0.0052072f $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_338_47#_c_346_n N_VPWR_c_571_n 0.004751f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_338_47#_c_347_n N_VPWR_c_572_n 0.0052072f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_338_47#_c_348_n N_VPWR_c_572_n 0.004751f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_338_47#_c_349_n N_VPWR_c_573_n 0.00688901f $X=6.75 $Y=1.41 $X2=0
+ $Y2=0
cc_275 N_A_338_47#_c_350_n N_VPWR_c_574_n 0.0210596f $X=1.815 $Y=1.63 $X2=0
+ $Y2=0
cc_276 N_A_338_47#_c_382_n N_VPWR_c_576_n 0.0223557f $X=2.755 $Y=1.63 $X2=0
+ $Y2=0
cc_277 N_A_338_47#_c_342_n N_VPWR_c_578_n 0.00597712f $X=3.46 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_338_47#_c_343_n N_VPWR_c_578_n 0.00673617f $X=3.93 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_338_47#_c_344_n N_VPWR_c_580_n 0.00597712f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_338_47#_c_345_n N_VPWR_c_580_n 0.00673617f $X=4.87 $Y=1.41 $X2=0
+ $Y2=0
cc_281 N_A_338_47#_c_346_n N_VPWR_c_582_n 0.00597712f $X=5.34 $Y=1.41 $X2=0
+ $Y2=0
cc_282 N_A_338_47#_c_347_n N_VPWR_c_582_n 0.00673617f $X=5.81 $Y=1.41 $X2=0
+ $Y2=0
cc_283 N_A_338_47#_c_348_n N_VPWR_c_584_n 0.00597712f $X=6.28 $Y=1.41 $X2=0
+ $Y2=0
cc_284 N_A_338_47#_c_349_n N_VPWR_c_584_n 0.00673617f $X=6.75 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_338_47#_M1009_s N_VPWR_c_566_n 0.00217517f $X=1.69 $Y=1.485 $X2=0
+ $Y2=0
cc_286 N_A_338_47#_M1014_s N_VPWR_c_566_n 0.00231261f $X=2.61 $Y=1.485 $X2=0
+ $Y2=0
cc_287 N_A_338_47#_c_342_n N_VPWR_c_566_n 0.0100198f $X=3.46 $Y=1.41 $X2=0 $Y2=0
cc_288 N_A_338_47#_c_343_n N_VPWR_c_566_n 0.0118438f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_289 N_A_338_47#_c_344_n N_VPWR_c_566_n 0.00999457f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A_338_47#_c_345_n N_VPWR_c_566_n 0.0118438f $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A_338_47#_c_346_n N_VPWR_c_566_n 0.00999457f $X=5.34 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_338_47#_c_347_n N_VPWR_c_566_n 0.0118438f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_293 N_A_338_47#_c_348_n N_VPWR_c_566_n 0.00999457f $X=6.28 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_338_47#_c_349_n N_VPWR_c_566_n 0.0128459f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A_338_47#_c_350_n N_VPWR_c_566_n 0.0124725f $X=1.815 $Y=1.63 $X2=0
+ $Y2=0
cc_296 N_A_338_47#_c_382_n N_VPWR_c_566_n 0.0140101f $X=2.755 $Y=1.63 $X2=0
+ $Y2=0
cc_297 N_A_338_47#_M1001_g N_X_c_697_n 0.0065059f $X=3.435 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_338_47#_M1003_g N_X_c_697_n 0.00693104f $X=3.905 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A_338_47#_M1006_g N_X_c_697_n 5.47131e-19 $X=4.375 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A_338_47#_c_342_n N_X_c_698_n 0.0137692f $X=3.46 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_338_47#_c_343_n N_X_c_698_n 0.0115459f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_338_47#_c_344_n N_X_c_698_n 7.68612e-19 $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_338_47#_c_382_n N_X_c_698_n 0.00486061f $X=2.755 $Y=1.63 $X2=0 $Y2=0
cc_304 N_A_338_47#_M1003_g N_X_c_679_n 0.00879805f $X=3.905 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A_338_47#_M1006_g N_X_c_679_n 0.00879805f $X=4.375 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_338_47#_c_338_n N_X_c_679_n 0.03957f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A_338_47#_c_341_n N_X_c_679_n 0.0031956f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_308 N_A_338_47#_M1001_g N_X_c_680_n 0.00243606f $X=3.435 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_338_47#_M1003_g N_X_c_680_n 0.00113891f $X=3.905 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A_338_47#_c_335_n N_X_c_680_n 0.00808484f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_311 N_A_338_47#_c_338_n N_X_c_680_n 0.030582f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_338_47#_c_341_n N_X_c_680_n 0.00331919f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_313 N_A_338_47#_c_343_n N_X_c_688_n 0.0137916f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_338_47#_c_344_n N_X_c_688_n 0.0101048f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_338_47#_c_338_n N_X_c_688_n 0.0394547f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_338_47#_c_341_n N_X_c_688_n 0.00720931f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_317 N_A_338_47#_c_342_n N_X_c_689_n 0.00386185f $X=3.46 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_338_47#_c_343_n N_X_c_689_n 0.00107777f $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_338_47#_c_353_n N_X_c_689_n 0.0149281f $X=3.14 $Y=1.53 $X2=0 $Y2=0
cc_320 N_A_338_47#_c_338_n N_X_c_689_n 0.0305808f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_338_47#_c_341_n N_X_c_689_n 0.0074788f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_322 N_A_338_47#_M1003_g N_X_c_724_n 5.25882e-19 $X=3.905 $Y=0.56 $X2=0 $Y2=0
cc_323 N_A_338_47#_M1006_g N_X_c_724_n 0.00657592f $X=4.375 $Y=0.56 $X2=0 $Y2=0
cc_324 N_A_338_47#_M1007_g N_X_c_724_n 0.00693104f $X=4.845 $Y=0.56 $X2=0 $Y2=0
cc_325 N_A_338_47#_M1013_g N_X_c_724_n 5.47131e-19 $X=5.315 $Y=0.56 $X2=0 $Y2=0
cc_326 N_A_338_47#_c_343_n N_X_c_728_n 8.07084e-19 $X=3.93 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_338_47#_c_344_n N_X_c_728_n 0.0141618f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A_338_47#_c_345_n N_X_c_728_n 0.0115459f $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_329 N_A_338_47#_c_346_n N_X_c_728_n 7.68612e-19 $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A_338_47#_M1007_g N_X_c_681_n 0.00879805f $X=4.845 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A_338_47#_M1013_g N_X_c_681_n 0.00879805f $X=5.315 $Y=0.56 $X2=0 $Y2=0
cc_332 N_A_338_47#_c_338_n N_X_c_681_n 0.03957f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_333 N_A_338_47#_c_341_n N_X_c_681_n 0.0031956f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_334 N_A_338_47#_c_345_n N_X_c_690_n 0.0137916f $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A_338_47#_c_346_n N_X_c_690_n 0.0101048f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_338_47#_c_338_n N_X_c_690_n 0.0394547f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_338_47#_c_341_n N_X_c_690_n 0.00720931f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_338 N_A_338_47#_M1007_g N_X_c_740_n 5.25882e-19 $X=4.845 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A_338_47#_M1013_g N_X_c_740_n 0.00657592f $X=5.315 $Y=0.56 $X2=0 $Y2=0
cc_340 N_A_338_47#_M1015_g N_X_c_740_n 0.00693104f $X=5.785 $Y=0.56 $X2=0 $Y2=0
cc_341 N_A_338_47#_M1020_g N_X_c_740_n 5.47131e-19 $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_342 N_A_338_47#_c_345_n N_X_c_744_n 8.07084e-19 $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_338_47#_c_346_n N_X_c_744_n 0.0141618f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_338_47#_c_347_n N_X_c_744_n 0.0115459f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A_338_47#_c_348_n N_X_c_744_n 7.68612e-19 $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A_338_47#_M1015_g N_X_c_682_n 0.00879805f $X=5.785 $Y=0.56 $X2=0 $Y2=0
cc_347 N_A_338_47#_M1020_g N_X_c_682_n 0.0101397f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_338_47#_c_338_n N_X_c_682_n 0.0118227f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_349 N_A_338_47#_c_341_n N_X_c_682_n 0.00378155f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_350 N_A_338_47#_c_347_n N_X_c_691_n 0.0137916f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_338_47#_c_348_n N_X_c_691_n 0.0113484f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_338_47#_c_338_n N_X_c_691_n 0.011672f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_353 N_A_338_47#_c_341_n N_X_c_691_n 0.00832854f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_354 N_A_338_47#_M1015_g N_X_c_756_n 5.25882e-19 $X=5.785 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_338_47#_M1020_g N_X_c_756_n 0.00657592f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_338_47#_c_347_n N_X_c_758_n 8.07084e-19 $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_357 N_A_338_47#_c_348_n N_X_c_758_n 0.0141618f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A_338_47#_c_349_n N_X_c_758_n 0.017566f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_338_47#_M1023_g N_X_c_683_n 0.0137799f $X=6.775 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_338_47#_c_349_n N_X_c_762_n 0.0171489f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_338_47#_c_341_n N_X_c_762_n 3.58038e-19 $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_362 N_A_338_47#_M1006_g N_X_c_684_n 0.00113891f $X=4.375 $Y=0.56 $X2=0 $Y2=0
cc_363 N_A_338_47#_M1007_g N_X_c_684_n 0.00113891f $X=4.845 $Y=0.56 $X2=0 $Y2=0
cc_364 N_A_338_47#_c_338_n N_X_c_684_n 0.030582f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_365 N_A_338_47#_c_341_n N_X_c_684_n 0.00331919f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_366 N_A_338_47#_c_344_n N_X_c_692_n 0.00260297f $X=4.4 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_338_47#_c_345_n N_X_c_692_n 0.00107777f $X=4.87 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_338_47#_c_338_n N_X_c_692_n 0.0305808f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_369 N_A_338_47#_c_341_n N_X_c_692_n 0.0074788f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_370 N_A_338_47#_M1013_g N_X_c_685_n 0.00113891f $X=5.315 $Y=0.56 $X2=0 $Y2=0
cc_371 N_A_338_47#_M1015_g N_X_c_685_n 0.00113891f $X=5.785 $Y=0.56 $X2=0 $Y2=0
cc_372 N_A_338_47#_c_338_n N_X_c_685_n 0.030582f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_373 N_A_338_47#_c_341_n N_X_c_685_n 0.00331919f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_374 N_A_338_47#_c_346_n N_X_c_693_n 0.00260297f $X=5.34 $Y=1.41 $X2=0 $Y2=0
cc_375 N_A_338_47#_c_347_n N_X_c_693_n 0.00107777f $X=5.81 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_338_47#_c_338_n N_X_c_693_n 0.0305808f $X=5.465 $Y=1.16 $X2=0 $Y2=0
cc_377 N_A_338_47#_c_341_n N_X_c_693_n 0.0074788f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_378 N_A_338_47#_M1020_g N_X_c_686_n 0.00147497f $X=6.255 $Y=0.56 $X2=0 $Y2=0
cc_379 N_A_338_47#_c_341_n N_X_c_686_n 0.00558583f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_380 N_A_338_47#_c_348_n N_X_c_694_n 0.00334115f $X=6.28 $Y=1.41 $X2=0 $Y2=0
cc_381 N_A_338_47#_c_349_n N_X_c_694_n 0.00128868f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_382 N_A_338_47#_c_341_n N_X_c_694_n 0.00885963f $X=6.75 $Y=1.217 $X2=0 $Y2=0
cc_383 N_A_338_47#_c_349_n X 0.00154146f $X=6.75 $Y=1.41 $X2=0 $Y2=0
cc_384 N_A_338_47#_M1023_g X 0.0251689f $X=6.775 $Y=0.56 $X2=0 $Y2=0
cc_385 N_A_338_47#_c_333_n N_VGND_M1005_d 0.00251598f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_386 N_A_338_47#_c_335_n N_VGND_M1012_d 0.00193551f $X=3.14 $Y=0.82 $X2=0
+ $Y2=0
cc_387 N_A_338_47#_c_332_n N_VGND_c_851_n 0.0184656f $X=1.815 $Y=0.4 $X2=0 $Y2=0
cc_388 N_A_338_47#_c_333_n N_VGND_c_851_n 0.0127122f $X=2.54 $Y=0.82 $X2=0 $Y2=0
cc_389 N_A_338_47#_M1001_g N_VGND_c_852_n 0.00268723f $X=3.435 $Y=0.56 $X2=0
+ $Y2=0
cc_390 N_A_338_47#_c_335_n N_VGND_c_852_n 0.0135251f $X=3.14 $Y=0.82 $X2=0 $Y2=0
cc_391 N_A_338_47#_M1003_g N_VGND_c_853_n 0.00390178f $X=3.905 $Y=0.56 $X2=0
+ $Y2=0
cc_392 N_A_338_47#_M1006_g N_VGND_c_853_n 0.00276126f $X=4.375 $Y=0.56 $X2=0
+ $Y2=0
cc_393 N_A_338_47#_M1007_g N_VGND_c_854_n 0.00390178f $X=4.845 $Y=0.56 $X2=0
+ $Y2=0
cc_394 N_A_338_47#_M1013_g N_VGND_c_854_n 0.00276126f $X=5.315 $Y=0.56 $X2=0
+ $Y2=0
cc_395 N_A_338_47#_M1015_g N_VGND_c_855_n 0.00390178f $X=5.785 $Y=0.56 $X2=0
+ $Y2=0
cc_396 N_A_338_47#_M1020_g N_VGND_c_855_n 0.00276126f $X=6.255 $Y=0.56 $X2=0
+ $Y2=0
cc_397 N_A_338_47#_M1023_g N_VGND_c_856_n 0.00438629f $X=6.775 $Y=0.56 $X2=0
+ $Y2=0
cc_398 N_A_338_47#_c_332_n N_VGND_c_857_n 0.020318f $X=1.815 $Y=0.4 $X2=0 $Y2=0
cc_399 N_A_338_47#_c_333_n N_VGND_c_857_n 0.00260082f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_400 N_A_338_47#_c_333_n N_VGND_c_859_n 0.00193763f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_401 N_A_338_47#_c_380_n N_VGND_c_859_n 0.022456f $X=2.755 $Y=0.4 $X2=0 $Y2=0
cc_402 N_A_338_47#_c_335_n N_VGND_c_859_n 0.00248202f $X=3.14 $Y=0.82 $X2=0
+ $Y2=0
cc_403 N_A_338_47#_M1001_g N_VGND_c_861_n 0.00541562f $X=3.435 $Y=0.56 $X2=0
+ $Y2=0
cc_404 N_A_338_47#_M1003_g N_VGND_c_861_n 0.00424619f $X=3.905 $Y=0.56 $X2=0
+ $Y2=0
cc_405 N_A_338_47#_M1006_g N_VGND_c_863_n 0.00424619f $X=4.375 $Y=0.56 $X2=0
+ $Y2=0
cc_406 N_A_338_47#_M1007_g N_VGND_c_863_n 0.00424619f $X=4.845 $Y=0.56 $X2=0
+ $Y2=0
cc_407 N_A_338_47#_M1013_g N_VGND_c_865_n 0.00424619f $X=5.315 $Y=0.56 $X2=0
+ $Y2=0
cc_408 N_A_338_47#_M1015_g N_VGND_c_865_n 0.00424619f $X=5.785 $Y=0.56 $X2=0
+ $Y2=0
cc_409 N_A_338_47#_M1020_g N_VGND_c_867_n 0.00424619f $X=6.255 $Y=0.56 $X2=0
+ $Y2=0
cc_410 N_A_338_47#_M1023_g N_VGND_c_867_n 0.00439206f $X=6.775 $Y=0.56 $X2=0
+ $Y2=0
cc_411 N_A_338_47#_M1005_s N_VGND_c_870_n 0.0020946f $X=1.69 $Y=0.235 $X2=0
+ $Y2=0
cc_412 N_A_338_47#_M1011_s N_VGND_c_870_n 0.00304616f $X=2.57 $Y=0.235 $X2=0
+ $Y2=0
cc_413 N_A_338_47#_M1001_g N_VGND_c_870_n 0.00965588f $X=3.435 $Y=0.56 $X2=0
+ $Y2=0
cc_414 N_A_338_47#_M1003_g N_VGND_c_870_n 0.00611295f $X=3.905 $Y=0.56 $X2=0
+ $Y2=0
cc_415 N_A_338_47#_M1006_g N_VGND_c_870_n 0.00599018f $X=4.375 $Y=0.56 $X2=0
+ $Y2=0
cc_416 N_A_338_47#_M1007_g N_VGND_c_870_n 0.00611295f $X=4.845 $Y=0.56 $X2=0
+ $Y2=0
cc_417 N_A_338_47#_M1013_g N_VGND_c_870_n 0.00599018f $X=5.315 $Y=0.56 $X2=0
+ $Y2=0
cc_418 N_A_338_47#_M1015_g N_VGND_c_870_n 0.00611295f $X=5.785 $Y=0.56 $X2=0
+ $Y2=0
cc_419 N_A_338_47#_M1020_g N_VGND_c_870_n 0.00610552f $X=6.255 $Y=0.56 $X2=0
+ $Y2=0
cc_420 N_A_338_47#_M1023_g N_VGND_c_870_n 0.00720128f $X=6.775 $Y=0.56 $X2=0
+ $Y2=0
cc_421 N_A_338_47#_c_332_n N_VGND_c_870_n 0.0123792f $X=1.815 $Y=0.4 $X2=0 $Y2=0
cc_422 N_A_338_47#_c_333_n N_VGND_c_870_n 0.00961016f $X=2.54 $Y=0.82 $X2=0
+ $Y2=0
cc_423 N_A_338_47#_c_380_n N_VGND_c_870_n 0.0142976f $X=2.755 $Y=0.4 $X2=0 $Y2=0
cc_424 N_A_338_47#_c_335_n N_VGND_c_870_n 0.00561929f $X=3.14 $Y=0.82 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_566_n N_X_M1000_s 0.00231261f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_566_n N_X_M1004_s 0.00231261f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_566_n N_X_M1016_s 0.00231261f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_566_n N_X_M1022_s 0.00231261f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_429 N_VPWR_c_569_n N_X_c_698_n 0.0507655f $X=3.225 $Y=2 $X2=0 $Y2=0
cc_430 N_VPWR_c_570_n N_X_c_698_n 0.0385613f $X=4.165 $Y=2 $X2=0 $Y2=0
cc_431 N_VPWR_c_578_n N_X_c_698_n 0.0223557f $X=4.08 $Y=2.72 $X2=0 $Y2=0
cc_432 N_VPWR_c_566_n N_X_c_698_n 0.0140101f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_433 N_VPWR_M1002_d N_X_c_688_n 0.00199888f $X=4.02 $Y=1.485 $X2=0 $Y2=0
cc_434 N_VPWR_c_570_n N_X_c_688_n 0.0112848f $X=4.165 $Y=2 $X2=0 $Y2=0
cc_435 N_VPWR_c_570_n N_X_c_728_n 0.0470327f $X=4.165 $Y=2 $X2=0 $Y2=0
cc_436 N_VPWR_c_571_n N_X_c_728_n 0.0385613f $X=5.105 $Y=2 $X2=0 $Y2=0
cc_437 N_VPWR_c_580_n N_X_c_728_n 0.0223557f $X=5.02 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_c_566_n N_X_c_728_n 0.0140101f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_439 N_VPWR_M1008_d N_X_c_690_n 0.00199888f $X=4.96 $Y=1.485 $X2=0 $Y2=0
cc_440 N_VPWR_c_571_n N_X_c_690_n 0.0112848f $X=5.105 $Y=2 $X2=0 $Y2=0
cc_441 N_VPWR_c_571_n N_X_c_744_n 0.0470327f $X=5.105 $Y=2 $X2=0 $Y2=0
cc_442 N_VPWR_c_572_n N_X_c_744_n 0.0385613f $X=6.045 $Y=2 $X2=0 $Y2=0
cc_443 N_VPWR_c_582_n N_X_c_744_n 0.0223557f $X=5.96 $Y=2.72 $X2=0 $Y2=0
cc_444 N_VPWR_c_566_n N_X_c_744_n 0.0140101f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_M1019_d N_X_c_691_n 0.00199888f $X=5.9 $Y=1.485 $X2=0 $Y2=0
cc_446 N_VPWR_c_572_n N_X_c_691_n 0.0112848f $X=6.045 $Y=2 $X2=0 $Y2=0
cc_447 N_VPWR_c_572_n N_X_c_758_n 0.0470327f $X=6.045 $Y=2 $X2=0 $Y2=0
cc_448 N_VPWR_c_573_n N_X_c_758_n 0.0385613f $X=6.985 $Y=2 $X2=0 $Y2=0
cc_449 N_VPWR_c_584_n N_X_c_758_n 0.0223557f $X=6.9 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_566_n N_X_c_758_n 0.0140101f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_451 N_VPWR_M1025_d X 0.00458027f $X=6.84 $Y=1.485 $X2=0 $Y2=0
cc_452 N_VPWR_c_573_n X 0.0124926f $X=6.985 $Y=2 $X2=0 $Y2=0
cc_453 N_X_c_679_n N_VGND_M1003_d 0.00251598f $X=4.42 $Y=0.82 $X2=0 $Y2=0
cc_454 N_X_c_681_n N_VGND_M1007_d 0.00251598f $X=5.36 $Y=0.82 $X2=0 $Y2=0
cc_455 N_X_c_682_n N_VGND_M1015_d 0.00251598f $X=6.3 $Y=0.82 $X2=0 $Y2=0
cc_456 N_X_c_683_n N_VGND_M1023_d 0.00322964f $X=6.86 $Y=0.82 $X2=0 $Y2=0
cc_457 N_X_c_697_n N_VGND_c_853_n 0.0186688f $X=3.695 $Y=0.4 $X2=0 $Y2=0
cc_458 N_X_c_679_n N_VGND_c_853_n 0.0127122f $X=4.42 $Y=0.82 $X2=0 $Y2=0
cc_459 N_X_c_724_n N_VGND_c_854_n 0.0186688f $X=4.635 $Y=0.4 $X2=0 $Y2=0
cc_460 N_X_c_681_n N_VGND_c_854_n 0.0127122f $X=5.36 $Y=0.82 $X2=0 $Y2=0
cc_461 N_X_c_740_n N_VGND_c_855_n 0.0186688f $X=5.575 $Y=0.4 $X2=0 $Y2=0
cc_462 N_X_c_682_n N_VGND_c_855_n 0.0127122f $X=6.3 $Y=0.82 $X2=0 $Y2=0
cc_463 N_X_c_683_n N_VGND_c_856_n 0.0140453f $X=6.86 $Y=0.82 $X2=0 $Y2=0
cc_464 N_X_c_697_n N_VGND_c_861_n 0.0216617f $X=3.695 $Y=0.4 $X2=0 $Y2=0
cc_465 N_X_c_679_n N_VGND_c_861_n 0.00260082f $X=4.42 $Y=0.82 $X2=0 $Y2=0
cc_466 N_X_c_679_n N_VGND_c_863_n 0.00193763f $X=4.42 $Y=0.82 $X2=0 $Y2=0
cc_467 N_X_c_724_n N_VGND_c_863_n 0.0216617f $X=4.635 $Y=0.4 $X2=0 $Y2=0
cc_468 N_X_c_681_n N_VGND_c_863_n 0.00260082f $X=5.36 $Y=0.82 $X2=0 $Y2=0
cc_469 N_X_c_681_n N_VGND_c_865_n 0.00193763f $X=5.36 $Y=0.82 $X2=0 $Y2=0
cc_470 N_X_c_740_n N_VGND_c_865_n 0.0216617f $X=5.575 $Y=0.4 $X2=0 $Y2=0
cc_471 N_X_c_682_n N_VGND_c_865_n 0.00260082f $X=6.3 $Y=0.82 $X2=0 $Y2=0
cc_472 N_X_c_682_n N_VGND_c_867_n 0.00193763f $X=6.3 $Y=0.82 $X2=0 $Y2=0
cc_473 N_X_c_756_n N_VGND_c_867_n 0.022456f $X=6.515 $Y=0.4 $X2=0 $Y2=0
cc_474 N_X_c_683_n N_VGND_c_867_n 0.00218716f $X=6.86 $Y=0.82 $X2=0 $Y2=0
cc_475 N_X_c_683_n N_VGND_c_869_n 0.00279505f $X=6.86 $Y=0.82 $X2=0 $Y2=0
cc_476 N_X_M1001_s N_VGND_c_870_n 0.00255524f $X=3.51 $Y=0.235 $X2=0 $Y2=0
cc_477 N_X_M1006_s N_VGND_c_870_n 0.00255524f $X=4.45 $Y=0.235 $X2=0 $Y2=0
cc_478 N_X_M1013_s N_VGND_c_870_n 0.00255524f $X=5.39 $Y=0.235 $X2=0 $Y2=0
cc_479 N_X_M1020_s N_VGND_c_870_n 0.00304616f $X=6.33 $Y=0.235 $X2=0 $Y2=0
cc_480 N_X_c_697_n N_VGND_c_870_n 0.0140924f $X=3.695 $Y=0.4 $X2=0 $Y2=0
cc_481 N_X_c_679_n N_VGND_c_870_n 0.00961016f $X=4.42 $Y=0.82 $X2=0 $Y2=0
cc_482 N_X_c_724_n N_VGND_c_870_n 0.0140924f $X=4.635 $Y=0.4 $X2=0 $Y2=0
cc_483 N_X_c_681_n N_VGND_c_870_n 0.00961016f $X=5.36 $Y=0.82 $X2=0 $Y2=0
cc_484 N_X_c_740_n N_VGND_c_870_n 0.0140924f $X=5.575 $Y=0.4 $X2=0 $Y2=0
cc_485 N_X_c_682_n N_VGND_c_870_n 0.00961016f $X=6.3 $Y=0.82 $X2=0 $Y2=0
cc_486 N_X_c_756_n N_VGND_c_870_n 0.0142976f $X=6.515 $Y=0.4 $X2=0 $Y2=0
cc_487 N_X_c_683_n N_VGND_c_870_n 0.0105046f $X=6.86 $Y=0.82 $X2=0 $Y2=0
