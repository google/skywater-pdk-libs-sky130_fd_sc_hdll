* File: sky130_fd_sc_hdll__a32o_1.pex.spice
* Created: Thu Aug 27 18:56:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32O_1%A_93_21# 1 2 7 9 10 12 16 17 18 19 20 22 23
+ 25 29 32 34
c97 16 0 1.17293e-19 $X=0.76 $Y=1.495
r98 32 35 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.707 $Y=1.16
+ $X2=0.707 $Y2=1.325
r99 32 34 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=0.707 $Y=1.16
+ $X2=0.707 $Y2=0.995
r100 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.655
+ $Y=1.16 $X2=0.655 $Y2=1.16
r101 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.24 $Y=1.665
+ $X2=3.24 $Y2=1.96
r102 23 25 93.2941 $w=1.68e-07 $l=1.43e-06 $layer=LI1_cond $X=1.315 $Y=0.4
+ $X2=2.745 $Y2=0.4
r103 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.23 $Y=0.485
+ $X2=1.315 $Y2=0.4
r104 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.23 $Y=0.485
+ $X2=1.23 $Y2=0.655
r105 19 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.155 $Y=1.58
+ $X2=3.24 $Y2=1.665
r106 19 20 150.706 $w=1.68e-07 $l=2.31e-06 $layer=LI1_cond $X=3.155 $Y=1.58
+ $X2=0.845 $Y2=1.58
r107 17 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.145 $Y=0.74
+ $X2=1.23 $Y2=0.655
r108 17 18 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=1.145 $Y=0.74
+ $X2=0.845 $Y2=0.74
r109 16 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=1.495
+ $X2=0.845 $Y2=1.58
r110 16 35 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.76 $Y=1.495
+ $X2=0.76 $Y2=1.325
r111 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=0.825
+ $X2=0.845 $Y2=0.74
r112 13 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.76 $Y=0.825
+ $X2=0.76 $Y2=0.995
r113 10 33 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=0.565 $Y=1.41
+ $X2=0.63 $Y2=1.16
r114 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.565 $Y=1.41
+ $X2=0.565 $Y2=1.985
r115 7 33 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.63 $Y2=1.16
r116 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=0.56
r117 2 29 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=3.09
+ $Y=1.485 $X2=3.24 $Y2=1.96
r118 1 25 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.745 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%A3 1 3 4 6 7 13
r34 7 13 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.205 $Y=1.16 $X2=1.155
+ $Y2=1.16
r35 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r36 4 10 38.5615 $w=3.23e-07 $l=1.71377e-07 $layer=POLY_cond $X=1.305 $Y=0.995
+ $X2=1.292 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.305 $Y=0.995
+ $X2=1.305 $Y2=0.56
r38 1 10 46.6797 $w=3.23e-07 $l=2.70185e-07 $layer=POLY_cond $X=1.25 $Y=1.41
+ $X2=1.292 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.25 $Y=1.41 $X2=1.25
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%A2 1 3 4 6 7 8
c35 1 0 1.44397e-19 $X=1.755 $Y=0.995
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.815
+ $Y=1.16 $X2=1.815 $Y2=1.16
r37 8 13 8.40605 $w=4.23e-07 $l=3.1e-07 $layer=LI1_cond $X=1.737 $Y=0.85
+ $X2=1.737 $Y2=1.16
r38 7 13 0.813489 $w=4.23e-07 $l=3e-08 $layer=LI1_cond $X=1.737 $Y=1.19
+ $X2=1.737 $Y2=1.16
r39 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.78 $Y=1.41
+ $X2=1.84 $Y2=1.16
r40 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.78 $Y=1.41 $X2=1.78
+ $Y2=1.985
r41 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.755 $Y=0.995
+ $X2=1.84 $Y2=1.16
r42 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.755 $Y=0.995
+ $X2=1.755 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%A1 1 3 4 6 7 8 13
c33 13 0 1.44397e-19 $X=2.345 $Y=1.16
r34 13 19 6.8592 $w=4.03e-07 $l=2.05e-07 $layer=LI1_cond $X=2.462 $Y=1.16
+ $X2=2.462 $Y2=0.955
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.345
+ $Y=1.16 $X2=2.345 $Y2=1.16
r36 8 19 4.24584 $w=2.83e-07 $l=1.05e-07 $layer=LI1_cond $X=2.522 $Y=0.85
+ $X2=2.522 $Y2=0.955
r37 7 13 0.853661 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=2.462 $Y=1.19
+ $X2=2.462 $Y2=1.16
r38 4 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.455 $Y=0.995
+ $X2=2.37 $Y2=1.16
r39 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.455 $Y=0.995
+ $X2=2.455 $Y2=0.56
r40 1 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.37 $Y2=1.16
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.41 $X2=2.43
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%B1 1 3 4 6 7 8
r32 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.985
+ $Y=1.16 $X2=2.985 $Y2=1.16
r33 7 8 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=2.985 $Y=0.85
+ $X2=2.985 $Y2=1.16
r34 4 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.01 $Y2=1.16
r35 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.095 $Y=0.995
+ $X2=3.095 $Y2=0.56
r36 1 12 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=3 $Y=1.41
+ $X2=3.01 $Y2=1.16
r37 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3 $Y=1.41 $X2=3
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%B2 1 3 4 6 7 12 13 17
r29 13 17 9.84378 $w=2.38e-07 $l=2.05e-07 $layer=LI1_cond $X=3.91 $Y=1.53
+ $X2=3.91 $Y2=1.325
r30 12 17 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=1.16
+ $X2=3.91 $Y2=1.325
r31 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.515
+ $Y=1.16 $X2=3.515 $Y2=1.16
r32 7 12 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=3.79 $Y=1.16 $X2=3.91
+ $Y2=1.16
r33 7 9 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.79 $Y=1.16
+ $X2=3.515 $Y2=1.16
r34 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.54 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.48 $Y=1.41 $X2=3.48
+ $Y2=1.985
r36 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.54 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%X 1 2 7 8 9 10 11 12 36 42 46
r18 46 47 2.40535 $w=3.33e-07 $l=5e-08 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.56
r19 36 49 2.03372 $w=2.53e-07 $l=4.5e-08 $layer=LI1_cond $X=0.217 $Y=1.87
+ $X2=0.217 $Y2=1.915
r20 12 37 4.40336 $w=3.33e-07 $l=1.28e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.082
r21 11 37 5.05699 $w=3.33e-07 $l=1.47e-07 $layer=LI1_cond $X=0.257 $Y=1.935
+ $X2=0.257 $Y2=2.082
r22 11 49 1.37331 $w=3.33e-07 $l=2e-08 $layer=LI1_cond $X=0.257 $Y=1.935
+ $X2=0.257 $Y2=1.915
r23 11 36 0.903877 $w=2.53e-07 $l=2e-08 $layer=LI1_cond $X=0.217 $Y=1.85
+ $X2=0.217 $Y2=1.87
r24 11 33 8.58683 $w=2.53e-07 $l=1.9e-07 $layer=LI1_cond $X=0.217 $Y=1.85
+ $X2=0.217 $Y2=1.66
r25 10 33 5.8752 $w=2.53e-07 $l=1.3e-07 $layer=LI1_cond $X=0.217 $Y=1.53
+ $X2=0.217 $Y2=1.66
r26 9 10 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=1.19
+ $X2=0.217 $Y2=1.53
r27 8 9 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=1.19
r28 8 25 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.217 $Y=0.85
+ $X2=0.217 $Y2=0.725
r29 7 46 0.619223 $w=3.33e-07 $l=1.8e-08 $layer=LI1_cond $X=0.257 $Y=0.492
+ $X2=0.257 $Y2=0.51
r30 7 42 3.68094 $w=3.33e-07 $l=1.07e-07 $layer=LI1_cond $X=0.257 $Y=0.492
+ $X2=0.257 $Y2=0.385
r31 7 25 6.68869 $w=2.53e-07 $l=1.48e-07 $layer=LI1_cond $X=0.217 $Y=0.577
+ $X2=0.217 $Y2=0.725
r32 7 47 0.768295 $w=2.53e-07 $l=1.7e-08 $layer=LI1_cond $X=0.217 $Y=0.577
+ $X2=0.217 $Y2=0.56
r33 2 11 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
r34 2 33 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r35 1 42 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.385
r36 1 25 182 $w=1.7e-07 $l=5.48954e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%VPWR 1 2 9 13 16 17 18 24 33 34 37
c49 1 0 1.17293e-19 $X=0.655 $Y=1.485
r50 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r52 31 34 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r53 31 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 30 33 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r55 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.105 $Y2=2.72
r57 28 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=2.72
+ $X2=2.53 $Y2=2.72
r58 27 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r60 24 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=2.105 $Y2=2.72
r61 24 26 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=2.72
+ $X2=1.61 $Y2=2.72
r62 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 18 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 16 21 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=0.725 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=2.72
+ $X2=0.89 $Y2=2.72
r67 15 26 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=1.61 $Y2=2.72
r68 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=2.72
+ $X2=0.89 $Y2=2.72
r69 11 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2.72
r70 11 13 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.105 $Y=2.635
+ $X2=2.105 $Y2=2.34
r71 7 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.89 $Y=2.635 $X2=0.89
+ $Y2=2.72
r72 7 9 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.89 $Y=2.635
+ $X2=0.89 $Y2=2
r73 2 13 600 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=1.87
+ $Y=1.485 $X2=2.105 $Y2=2.34
r74 1 9 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=0.655
+ $Y=1.485 $X2=0.89 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%A_268_297# 1 2 3 10 12 14 16 18 19 22
r33 20 22 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=3.765 $Y=2.295
+ $X2=3.765 $Y2=1.96
r34 18 20 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=3.635 $Y=2.38
+ $X2=3.765 $Y2=2.295
r35 18 19 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.635 $Y=2.38
+ $X2=2.875 $Y2=2.38
r36 17 19 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.71 $Y=2.295
+ $X2=2.875 $Y2=2.38
r37 16 27 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=2.045 $X2=2.71
+ $Y2=1.96
r38 16 17 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=2.71 $Y=2.045
+ $X2=2.71 $Y2=2.295
r39 15 25 4.64039 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=1.635 $Y=1.96
+ $X2=1.492 $Y2=1.96
r40 14 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=1.96
+ $X2=2.71 $Y2=1.96
r41 14 15 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.545 $Y=1.96
+ $X2=1.635 $Y2=1.96
r42 10 25 2.75828 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=1.492 $Y=2.045
+ $X2=1.492 $Y2=1.96
r43 10 12 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=1.492 $Y=2.045
+ $X2=1.492 $Y2=2.3
r44 3 22 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=3.57
+ $Y=1.485 $X2=3.72 $Y2=1.96
r45 2 27 300 $w=1.7e-07 $l=6.02557e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=1.485 $X2=2.71 $Y2=2
r46 1 25 600 $w=1.7e-07 $l=5.55653e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.485 $X2=1.515 $Y2=1.96
r47 1 12 600 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=1.34
+ $Y=1.485 $X2=1.515 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_1%VGND 1 2 9 11 13 15 17 22 31 35
r54 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r55 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r57 28 29 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 26 29 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r59 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r60 25 28 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r61 25 26 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 23 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=0.785
+ $Y2=0
r63 23 25 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.975 $Y=0 $X2=1.15
+ $Y2=0
r64 22 34 4.91182 $w=1.7e-07 $l=3.17e-07 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.822
+ $Y2=0
r65 22 28 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.505 $Y=0 $X2=3.45
+ $Y2=0
r66 17 31 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.785
+ $Y2=0
r67 17 19 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.23
+ $Y2=0
r68 15 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 11 34 3.28487 $w=3.8e-07 $l=1.64085e-07 $layer=LI1_cond $X=3.695 $Y=0.085
+ $X2=3.822 $Y2=0
r71 11 13 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.695 $Y=0.085
+ $X2=3.695 $Y2=0.38
r72 7 31 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0
r73 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.785 $Y=0.085
+ $X2=0.785 $Y2=0.4
r74 2 13 91 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=2 $X=3.53
+ $Y=0.235 $X2=3.72 $Y2=0.38
r75 1 9 182 $w=1.7e-07 $l=2.64953e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.81 $Y2=0.4
.ends

