* NGSPICE file created from sky130_fd_sc_hdll__and4b_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4b_4 A_N B C D VGND VNB VPB VPWR X
M1000 a_184_21# a_27_47# a_814_47# VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.47e+11p ps=2.06e+06u
M1001 a_718_47# C a_624_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.08e+11p ps=1.94e+06u
M1002 a_624_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.205e+11p ps=6.17e+06u
M1003 VPWR A_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=1.6157e+12p pd=1.333e+07u as=1.134e+11p ps=1.38e+06u
M1004 a_184_21# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.4e+11p pd=5.28e+06u as=0p ps=0u
M1005 a_814_47# B a_718_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1007 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1009 VPWR C a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR a_27_47# a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1014 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_184_21# D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

