* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nor3b_4 A B C_N VGND VNB VPB VPWR Y
X0 a_605_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_215_297# B a_605_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 Y a_27_47# a_605_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_605_297# B a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_27_47# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND B Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_605_297# a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_27_47# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_215_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_215_297# B a_605_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VPWR A a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_605_297# B a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y a_27_47# a_605_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 Y B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_215_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR A a_215_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Y A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
