# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__isobufsrc_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  18.40000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 0.995000 ;
        RECT 0.085000 0.995000 0.665000 1.325000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.650000 1.075000 17.600000 1.285000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  5.713000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  3.325000 0.255000  3.705000 0.725000 ;
        RECT  3.325000 0.725000 18.305000 0.905000 ;
        RECT  4.265000 0.255000  4.645000 0.725000 ;
        RECT  5.205000 0.255000  5.585000 0.725000 ;
        RECT  6.145000 0.255000  6.525000 0.725000 ;
        RECT  7.085000 0.255000  7.465000 0.725000 ;
        RECT  8.025000 0.255000  8.405000 0.725000 ;
        RECT  8.965000 0.255000  9.345000 0.725000 ;
        RECT  9.905000 0.255000 10.285000 0.725000 ;
        RECT 10.845000 0.255000 11.225000 0.725000 ;
        RECT 10.935000 1.455000 18.305000 1.625000 ;
        RECT 10.935000 1.625000 11.185000 2.125000 ;
        RECT 11.785000 0.255000 12.165000 0.725000 ;
        RECT 11.875000 1.625000 12.125000 2.125000 ;
        RECT 12.725000 0.255000 13.105000 0.725000 ;
        RECT 12.815000 1.625000 13.065000 2.125000 ;
        RECT 13.665000 0.255000 14.045000 0.725000 ;
        RECT 13.755000 1.625000 14.005000 2.125000 ;
        RECT 14.605000 0.255000 14.985000 0.725000 ;
        RECT 14.695000 1.625000 14.945000 2.125000 ;
        RECT 15.545000 0.255000 15.925000 0.725000 ;
        RECT 15.635000 1.625000 15.885000 2.125000 ;
        RECT 16.485000 0.255000 16.865000 0.725000 ;
        RECT 16.575000 1.625000 16.825000 2.125000 ;
        RECT 17.425000 0.255000 17.805000 0.725000 ;
        RECT 17.515000 1.625000 17.765000 2.125000 ;
        RECT 17.770000 0.905000 18.305000 1.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 18.400000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 18.400000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 18.400000 0.085000 ;
      RECT  0.000000  2.635000 18.400000 2.805000 ;
      RECT  0.300000  1.495000  0.515000 2.635000 ;
      RECT  0.485000  0.085000  0.865000 0.825000 ;
      RECT  0.685000  1.495000  1.115000 2.465000 ;
      RECT  0.885000  1.065000  2.385000 1.075000 ;
      RECT  0.885000  1.075000 10.480000 1.285000 ;
      RECT  0.885000  1.285000  1.115000 1.495000 ;
      RECT  1.085000  0.255000  1.345000 1.065000 ;
      RECT  1.335000  1.455000  1.555000 2.635000 ;
      RECT  1.565000  0.085000  1.865000 0.895000 ;
      RECT  1.725000  1.285000  2.155000 2.465000 ;
      RECT  2.085000  0.255000  2.385000 1.065000 ;
      RECT  2.375000  1.455000  2.670000 2.635000 ;
      RECT  2.605000  0.085000  3.155000 0.905000 ;
      RECT  2.875000  1.455000 10.715000 1.665000 ;
      RECT  2.875000  1.665000  3.195000 2.465000 ;
      RECT  3.415000  1.835000  3.665000 2.635000 ;
      RECT  3.885000  1.665000  4.135000 2.465000 ;
      RECT  3.925000  0.085000  4.095000 0.555000 ;
      RECT  4.355000  1.835000  4.605000 2.635000 ;
      RECT  4.825000  1.665000  5.075000 2.465000 ;
      RECT  4.865000  0.085000  5.035000 0.555000 ;
      RECT  5.295000  1.835000  5.545000 2.635000 ;
      RECT  5.765000  1.665000  6.015000 2.465000 ;
      RECT  5.805000  0.085000  5.975000 0.555000 ;
      RECT  6.235000  1.835000  6.485000 2.635000 ;
      RECT  6.705000  1.665000  6.955000 2.465000 ;
      RECT  6.745000  0.085000  6.915000 0.555000 ;
      RECT  7.175000  1.835000  7.425000 2.635000 ;
      RECT  7.645000  1.665000  7.895000 2.465000 ;
      RECT  7.685000  0.085000  7.855000 0.555000 ;
      RECT  8.115000  1.835000  8.365000 2.635000 ;
      RECT  8.585000  1.665000  8.835000 2.465000 ;
      RECT  8.625000  0.085000  8.795000 0.555000 ;
      RECT  9.055000  1.835000  9.305000 2.635000 ;
      RECT  9.525000  1.665000  9.775000 2.465000 ;
      RECT  9.565000  0.085000  9.735000 0.555000 ;
      RECT  9.995000  1.835000 10.245000 2.635000 ;
      RECT 10.465000  1.665000 10.715000 2.295000 ;
      RECT 10.465000  2.295000 18.235000 2.465000 ;
      RECT 10.505000  0.085000 10.675000 0.555000 ;
      RECT 11.405000  1.795000 11.655000 2.295000 ;
      RECT 11.445000  0.085000 11.615000 0.555000 ;
      RECT 12.345000  1.795000 12.595000 2.295000 ;
      RECT 12.385000  0.085000 12.555000 0.555000 ;
      RECT 13.285000  1.795000 13.535000 2.295000 ;
      RECT 13.325000  0.085000 13.495000 0.555000 ;
      RECT 14.225000  1.795000 14.475000 2.295000 ;
      RECT 14.265000  0.085000 14.435000 0.555000 ;
      RECT 15.165000  1.795000 15.415000 2.295000 ;
      RECT 15.205000  0.085000 15.375000 0.555000 ;
      RECT 16.105000  1.795000 16.355000 2.295000 ;
      RECT 16.145000  0.085000 16.315000 0.555000 ;
      RECT 17.045000  1.795000 17.295000 2.295000 ;
      RECT 17.085000  0.085000 17.255000 0.555000 ;
      RECT 17.985000  1.795000 18.235000 2.295000 ;
      RECT 18.025000  0.085000 18.295000 0.555000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_16
END LIBRARY
