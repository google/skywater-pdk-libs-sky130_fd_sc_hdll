* File: sky130_fd_sc_hdll__xor3_4.pex.spice
* Created: Thu Aug 27 19:30:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_80_207# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 34 37 38 39 41 43 45 46 48 50 52 54 55 64
c147 52 0 1.87406e-19 $X=2.132 $Y=1.325
c148 38 0 1.48868e-19 $X=2.575 $Y=1.96
c149 28 0 2.52917e-19 $X=2.005 $Y=1.41
r150 63 64 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.005 $Y2=1.202
r151 62 63 52.1616 $w=3.65e-07 $l=3.95e-07 $layer=POLY_cond $X=1.535 $Y=1.202
+ $X2=1.93 $Y2=1.202
r152 61 62 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.535 $Y2=1.202
r153 60 61 52.1616 $w=3.65e-07 $l=3.95e-07 $layer=POLY_cond $X=1.065 $Y=1.202
+ $X2=1.46 $Y2=1.202
r154 59 60 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.065 $Y2=1.202
r155 58 59 52.1616 $w=3.65e-07 $l=3.95e-07 $layer=POLY_cond $X=0.595 $Y=1.202
+ $X2=0.99 $Y2=1.202
r156 57 58 9.90411 $w=3.65e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.595 $Y2=1.202
r157 54 55 13.3132 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=3.895 $Y=0.355
+ $X2=3.66 $Y2=0.355
r158 50 51 18.4591 $w=2.3e-07 $l=3.48e-07 $layer=LI1_cond $X=2.132 $Y=0.865
+ $X2=2.48 $Y2=0.865
r159 46 48 72.0909 $w=1.68e-07 $l=1.105e-06 $layer=LI1_cond $X=2.795 $Y=2.32
+ $X2=3.9 $Y2=2.32
r160 45 46 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.685 $Y=2.235
+ $X2=2.795 $Y2=2.32
r161 44 45 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=2.685 $Y=2.045
+ $X2=2.685 $Y2=2.235
r162 43 55 71.4385 $w=1.68e-07 $l=1.095e-06 $layer=LI1_cond $X=2.565 $Y=0.34
+ $X2=3.66 $Y2=0.34
r163 41 51 2.50919 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.48 $Y=0.695
+ $X2=2.48 $Y2=0.865
r164 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.48 $Y=0.425
+ $X2=2.565 $Y2=0.34
r165 40 41 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.48 $Y=0.425
+ $X2=2.48 $Y2=0.695
r166 38 44 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.575 $Y=1.96
+ $X2=2.685 $Y2=2.045
r167 38 39 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.575 $Y=1.96
+ $X2=2.245 $Y2=1.96
r168 37 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.16 $Y=1.875
+ $X2=2.245 $Y2=1.96
r169 37 52 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.16 $Y=1.875
+ $X2=2.16 $Y2=1.325
r170 35 64 13.2055 $w=3.65e-07 $l=1e-07 $layer=POLY_cond $X=2.105 $Y=1.202
+ $X2=2.005 $Y2=1.202
r171 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.16 $X2=2.105 $Y2=1.16
r172 32 52 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=2.132 $Y=1.213
+ $X2=2.132 $Y2=1.325
r173 32 34 2.71464 $w=2.23e-07 $l=5.3e-08 $layer=LI1_cond $X=2.132 $Y=1.213
+ $X2=2.132 $Y2=1.16
r174 31 50 0.876693 $w=2.25e-07 $l=2.12e-07 $layer=LI1_cond $X=2.132 $Y=1.077
+ $X2=2.132 $Y2=0.865
r175 31 34 4.25123 $w=2.23e-07 $l=8.3e-08 $layer=LI1_cond $X=2.132 $Y=1.077
+ $X2=2.132 $Y2=1.16
r176 28 64 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.005 $Y=1.41
+ $X2=2.005 $Y2=1.202
r177 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.005 $Y=1.41
+ $X2=2.005 $Y2=1.985
r178 25 63 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r179 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r180 22 62 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.202
r181 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.985
r182 19 61 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r183 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r184 16 60 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.065 $Y=1.41
+ $X2=1.065 $Y2=1.202
r185 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.065 $Y=1.41
+ $X2=1.065 $Y2=1.985
r186 13 59 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r187 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r188 10 58 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.595 $Y=1.41
+ $X2=0.595 $Y2=1.202
r189 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.595 $Y=1.41
+ $X2=0.595 $Y2=1.985
r190 7 57 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r191 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r192 2 48 600 $w=1.7e-07 $l=7.84267e-07 $layer=licon1_PDIFF $count=1 $X=3.71
+ $Y=1.625 $X2=3.9 $Y2=2.32
r193 1 54 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.76
+ $Y=0.245 $X2=3.895 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%C 1 4 5 7 8 10 12 13 15 18 22 26
c63 8 0 1.48868e-19 $X=3.52 $Y=1.16
r64 22 26 4.36531 $w=3.28e-07 $l=1.25e-07 $layer=LI1_cond $X=3.58 $Y=1.16
+ $X2=3.455 $Y2=1.16
r65 18 26 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=3.455 $Y2=1.16
r66 13 15 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=3.685 $Y=0.985
+ $X2=3.685 $Y2=0.565
r67 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.62 $Y=1.55
+ $X2=3.62 $Y2=2.045
r68 8 10 85.013 $w=2.27e-07 $l=4.00849e-07 $layer=POLY_cond $X=3.642 $Y=1.16
+ $X2=3.62 $Y2=1.55
r69 8 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.58 $Y=1.16
+ $X2=3.58 $Y2=1.16
r70 8 13 42.7097 $w=2.27e-07 $l=1.9532e-07 $layer=POLY_cond $X=3.642 $Y=1.16
+ $X2=3.685 $Y2=0.985
r71 8 9 136.392 $w=3.3e-07 $l=7.8e-07 $layer=POLY_cond $X=3.52 $Y=1.16 $X2=2.74
+ $Y2=1.16
r72 5 9 38.8824 $w=2.71e-07 $l=1.96914e-07 $layer=POLY_cond $X=2.665 $Y=0.995
+ $X2=2.595 $Y2=1.16
r73 5 7 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.665 $Y=0.995
+ $X2=2.665 $Y2=0.675
r74 1 9 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.55 $Y=1.41
+ $X2=2.595 $Y2=1.16
r75 1 4 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.55 $Y=1.41 $X2=2.55
+ $Y2=1.805
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_528_297# 1 2 7 9 10 12 13 15 17 20 26
c71 13 0 1.53132e-19 $X=2.875 $Y=1.535
r72 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.16 $X2=4.175 $Y2=1.16
r73 23 26 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=4.07 $Y=1.16
+ $X2=4.175 $Y2=1.16
r74 19 23 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.07 $Y=1.325
+ $X2=4.07 $Y2=1.16
r75 19 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.07 $Y=1.325
+ $X2=4.07 $Y2=1.535
r76 18 22 3.40825 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.96 $Y=1.62
+ $X2=2.765 $Y2=1.62
r77 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.985 $Y=1.62
+ $X2=4.07 $Y2=1.535
r78 17 18 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=3.985 $Y=1.62
+ $X2=2.96 $Y2=1.62
r79 13 22 3.40825 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.875 $Y=1.535
+ $X2=2.765 $Y2=1.62
r80 13 15 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2.875 $Y=1.535
+ $X2=2.875 $Y2=0.76
r81 10 27 38.8824 $w=2.71e-07 $l=2.03101e-07 $layer=POLY_cond $X=4.285 $Y=0.995
+ $X2=4.2 $Y2=1.16
r82 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=4.285 $Y=0.995
+ $X2=4.285 $Y2=0.565
r83 7 27 74.8096 $w=2.71e-07 $l=3.9e-07 $layer=POLY_cond $X=4.2 $Y=1.55 $X2=4.2
+ $Y2=1.16
r84 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=4.2 $Y=1.55 $X2=4.2
+ $Y2=2.045
r85 2 22 600 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.485 $X2=2.825 $Y2=1.62
r86 1 15 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=2.74
+ $Y=0.465 $X2=2.875 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_1109_297# 1 2 7 9 12 14 15 16 18 19 21 22
+ 23 27 35 37 38 39 40 47 49 50 58
c178 14 0 1.24749e-19 $X=8.95 $Y=1.28
r179 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.87
+ $Y=1.11 $X2=8.87 $Y2=1.11
r180 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.8 $Y=0.85 $X2=8.8
+ $Y2=1.11
r181 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.75 $Y=0.85
+ $X2=8.75 $Y2=0.85
r182 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.27 $Y=0.85
+ $X2=7.27 $Y2=0.85
r183 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.79 $Y=0.85
+ $X2=5.79 $Y2=0.85
r184 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.415 $Y=0.85
+ $X2=7.27 $Y2=0.85
r185 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.605 $Y=0.85
+ $X2=8.75 $Y2=0.85
r186 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=8.605 $Y=0.85
+ $X2=7.415 $Y2=0.85
r187 38 42 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.985 $Y=0.85
+ $X2=5.79 $Y2=0.85
r188 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.125 $Y=0.85
+ $X2=7.27 $Y2=0.85
r189 37 38 1.41089 $w=1.4e-07 $l=1.14e-06 $layer=MET1_cond $X=7.125 $Y=0.85
+ $X2=5.985 $Y2=0.85
r190 35 47 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=7.247 $Y=0.995
+ $X2=7.247 $Y2=0.85
r191 31 35 6.36987 $w=2.73e-07 $l=1.52e-07 $layer=LI1_cond $X=7.095 $Y=1.132
+ $X2=7.247 $Y2=1.132
r192 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.095
+ $Y=1.16 $X2=7.095 $Y2=1.16
r193 28 58 28.8111 $w=2.88e-07 $l=7.25e-07 $layer=LI1_cond $X=5.845 $Y=1.445
+ $X2=5.845 $Y2=0.72
r194 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=5.845 $Y=1.58
+ $X2=5.845 $Y2=1.445
r195 25 27 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.69 $Y=1.58
+ $X2=5.845 $Y2=1.58
r196 22 32 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=7.36 $Y=1.16
+ $X2=7.095 $Y2=1.16
r197 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=7.36 $Y=1.16
+ $X2=7.46 $Y2=1.202
r198 19 55 38.5432 $w=3.18e-07 $l=2.03101e-07 $layer=POLY_cond $X=8.98 $Y=0.945
+ $X2=8.895 $Y2=1.11
r199 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.98 $Y=0.945
+ $X2=8.98 $Y2=0.535
r200 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.95 $Y=1.57
+ $X2=8.95 $Y2=2.065
r201 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.95 $Y=1.47 $X2=8.95
+ $Y2=1.57
r202 14 55 32.3713 $w=3.18e-07 $l=1.95576e-07 $layer=POLY_cond $X=8.95 $Y=1.28
+ $X2=8.895 $Y2=1.11
r203 14 15 62.9997 $w=2e-07 $l=1.9e-07 $layer=POLY_cond $X=8.95 $Y=1.28 $X2=8.95
+ $Y2=1.47
r204 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=7.485 $Y=0.995
+ $X2=7.46 $Y2=1.202
r205 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.485 $Y=0.995
+ $X2=7.485 $Y2=0.455
r206 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.202
r207 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.46 $Y=1.41
+ $X2=7.46 $Y2=1.805
r208 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.545
+ $Y=1.485 $X2=5.69 $Y2=1.63
r209 1 58 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.77
+ $Y=0.235 $X2=5.905 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 33
+ 37 38 39 48
r129 37 40 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.365 $Y=1.16
+ $X2=8.365 $Y2=1.325
r130 37 39 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.365 $Y=1.16
+ $X2=8.365 $Y2=0.995
r131 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.34
+ $Y=1.16 $X2=8.34 $Y2=1.16
r132 33 48 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.505 $Y=1.53
+ $X2=8.495 $Y2=1.53
r133 33 48 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=8.365 $Y=1.53
+ $X2=8.495 $Y2=1.53
r134 33 38 12.4376 $w=2.73e-07 $l=2.85e-07 $layer=LI1_cond $X=8.365 $Y=1.445
+ $X2=8.365 $Y2=1.16
r135 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=6.65 $Y=1.16 $X2=6.65
+ $Y2=1.085
r136 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=8.385 $Y=2.415
+ $X2=8.385 $Y2=1.965
r137 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=8.385 $Y=1.57
+ $X2=8.385 $Y2=1.965
r138 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.385 $Y=1.47 $X2=8.385
+ $Y2=1.57
r139 24 40 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.385 $Y=1.47
+ $X2=8.385 $Y2=1.325
r140 22 39 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=8.28 $Y=0.565
+ $X2=8.28 $Y2=0.995
r141 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=8.285 $Y=2.54
+ $X2=8.385 $Y2=2.415
r142 18 19 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=8.285 $Y=2.54
+ $X2=6.75 $Y2=2.54
r143 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=6.675 $Y=0.565
+ $X2=6.675 $Y2=1.085
r144 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=6.65 $Y=2.455
+ $X2=6.75 $Y2=2.54
r145 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=6.65 $Y=2.455
+ $X2=6.65 $Y2=1.905
r146 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=6.65 $Y=1.41 $X2=6.65
+ $Y2=1.16
r147 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=6.65 $Y=1.41
+ $X2=6.65 $Y2=1.905
r148 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=6.55 $Y=1.16 $X2=6.65
+ $Y2=1.16
r149 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=6.55 $Y=1.16 $X2=5.77
+ $Y2=1.16
r150 4 9 21.6409 $w=2.34e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.695 $Y=1.085
+ $X2=5.77 $Y2=1.16
r151 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=5.695 $Y=1.085
+ $X2=5.695 $Y2=0.56
r152 1 4 49.4359 $w=2.34e-07 $l=3.38349e-07 $layer=POLY_cond $X=5.455 $Y=1.322
+ $X2=5.695 $Y2=1.085
r153 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.455 $Y=1.41
+ $X2=5.455 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A 1 3 4 6 7
r37 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.4 $Y=1.16
+ $X2=9.4 $Y2=1.16
r38 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=9.53 $Y=0.995
+ $X2=9.435 $Y2=1.16
r39 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.53 $Y=0.995 $X2=9.53
+ $Y2=0.555
r40 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=9.505 $Y=1.41
+ $X2=9.435 $Y2=1.16
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.505 $Y=1.41
+ $X2=9.505 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_1225_365# 1 2 3 4 13 15 16 18 21 23 27 28
+ 29 30 36 37 40 43 44
c129 30 0 1.07404e-19 $X=9.89 $Y=1.495
c130 29 0 1.15937e-19 $X=9.89 $Y=1.325
r131 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.26 $Y=0.51
+ $X2=9.26 $Y2=0.51
r132 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.3 $Y=0.51 $X2=6.3
+ $Y2=0.51
r133 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.445 $Y=0.51
+ $X2=6.3 $Y2=0.51
r134 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.115 $Y=0.51
+ $X2=9.26 $Y2=0.51
r135 36 37 3.30445 $w=1.4e-07 $l=2.67e-06 $layer=MET1_cond $X=9.115 $Y=0.51
+ $X2=6.445 $Y2=0.51
r136 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.95
+ $Y=1.16 $X2=9.95 $Y2=1.16
r137 32 34 20.4335 $w=2.03e-07 $l=3.4e-07 $layer=LI1_cond $X=9.92 $Y=0.82
+ $X2=9.92 $Y2=1.16
r138 31 44 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=9.29 $Y=0.735
+ $X2=9.29 $Y2=0.51
r139 29 34 10.2745 $w=2.03e-07 $l=1.79374e-07 $layer=LI1_cond $X=9.89 $Y=1.325
+ $X2=9.92 $Y2=1.16
r140 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.89 $Y=1.325
+ $X2=9.89 $Y2=1.495
r141 28 31 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=9.435 $Y=0.82
+ $X2=9.29 $Y2=0.735
r142 27 32 1.77774 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.805 $Y=0.82
+ $X2=9.92 $Y2=0.82
r143 27 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=9.805 $Y=0.82
+ $X2=9.435 $Y2=0.82
r144 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=9.805 $Y=1.6
+ $X2=9.89 $Y2=1.495
r145 23 25 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=9.805 $Y=1.6
+ $X2=9.27 $Y2=1.6
r146 19 40 3.61456 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.25 $Y=0.595
+ $X2=6.25 $Y2=0.43
r147 19 21 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=6.25 $Y=0.595
+ $X2=6.25 $Y2=1.94
r148 16 35 38.578 $w=2.95e-07 $l=1.94808e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=9.975 $Y2=1.16
r149 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=10.04 $Y=0.995
+ $X2=10.04 $Y2=0.555
r150 13 35 48.1208 $w=2.95e-07 $l=2.69258e-07 $layer=POLY_cond $X=10.015 $Y=1.41
+ $X2=9.975 $Y2=1.16
r151 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.015 $Y=1.41
+ $X2=10.015 $Y2=1.985
r152 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=9.04
+ $Y=1.645 $X2=9.27 $Y2=1.62
r153 3 21 600 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_PDIFF $count=1 $X=6.125
+ $Y=1.825 $X2=6.25 $Y2=1.94
r154 2 44 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.235 $X2=9.27 $Y2=0.625
r155 1 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=6.29
+ $Y=0.245 $X2=6.415 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%VPWR 1 2 3 4 5 18 20 24 28 32 36 38 39 41
+ 42 44 45 46 55 70 71 74 77 80 83
c124 5 0 1.07404e-19 $X=9.595 $Y=1.485
r125 80 83 0.000284542 $w=4.8e-07 $l=1e-09 $layer=MET1_cond $X=0.229 $Y=2.72
+ $X2=0.23 $Y2=2.72
r126 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r127 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r128 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r129 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r130 67 68 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r131 65 68 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=9.43 $Y2=2.72
r132 65 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 64 67 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=2.72
+ $X2=9.43 $Y2=2.72
r134 64 65 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r135 62 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.22 $Y2=2.72
r136 62 64 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=5.385 $Y=2.72
+ $X2=5.75 $Y2=2.72
r137 61 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r138 60 61 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r139 58 61 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r140 57 60 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=4.83 $Y2=2.72
r141 57 58 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r142 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.055 $Y=2.72
+ $X2=5.22 $Y2=2.72
r143 55 60 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.055 $Y=2.72
+ $X2=4.83 $Y2=2.72
r144 54 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r145 54 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r146 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r147 51 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=2.72
+ $X2=1.3 $Y2=2.72
r148 51 53 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.465 $Y=2.72
+ $X2=2.07 $Y2=2.72
r149 49 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r150 46 75 0.23617 $w=4.8e-07 $l=8.3e-07 $layer=MET1_cond $X=0.32 $Y=2.72
+ $X2=1.15 $Y2=2.72
r151 46 83 0.0256088 $w=4.8e-07 $l=9e-08 $layer=MET1_cond $X=0.32 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 44 67 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.615 $Y=2.72
+ $X2=9.43 $Y2=2.72
r153 44 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.615 $Y=2.72
+ $X2=9.78 $Y2=2.72
r154 43 70 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.945 $Y=2.72
+ $X2=10.35 $Y2=2.72
r155 43 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.945 $Y=2.72
+ $X2=9.78 $Y2=2.72
r156 41 53 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.07 $Y2=2.72
r157 41 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.075 $Y=2.72
+ $X2=2.24 $Y2=2.72
r158 40 57 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.405 $Y=2.72
+ $X2=2.53 $Y2=2.72
r159 40 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.405 $Y=2.72
+ $X2=2.24 $Y2=2.72
r160 38 49 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.23 $Y2=2.72
r161 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.275 $Y=2.72
+ $X2=0.36 $Y2=2.72
r162 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.78 $Y=2.635
+ $X2=9.78 $Y2=2.72
r163 34 36 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.78 $Y=2.635
+ $X2=9.78 $Y2=2.36
r164 30 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.22 $Y=2.635
+ $X2=5.22 $Y2=2.72
r165 30 32 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.22 $Y=2.635
+ $X2=5.22 $Y2=2.32
r166 26 42 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=2.635
+ $X2=2.24 $Y2=2.72
r167 26 28 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.24 $Y=2.635
+ $X2=2.24 $Y2=2.3
r168 22 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=2.635 $X2=1.3
+ $Y2=2.72
r169 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.3 $Y=2.635
+ $X2=1.3 $Y2=2.3
r170 21 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.36 $Y2=2.72
r171 20 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=2.72
+ $X2=1.3 $Y2=2.72
r172 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.135 $Y=2.72
+ $X2=0.445 $Y2=2.72
r173 16 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.36 $Y=2.635
+ $X2=0.36 $Y2=2.72
r174 16 18 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.36 $Y=2.635
+ $X2=0.36 $Y2=2.3
r175 5 36 600 $w=1.7e-07 $l=9.63068e-07 $layer=licon1_PDIFF $count=1 $X=9.595
+ $Y=1.485 $X2=9.78 $Y2=2.36
r176 4 32 600 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=5.095
+ $Y=1.485 $X2=5.22 $Y2=2.32
r177 3 28 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.095
+ $Y=1.485 $X2=2.24 $Y2=2.3
r178 2 24 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.155
+ $Y=1.485 $X2=1.3 $Y2=2.3
r179 1 18 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.235
+ $Y=1.485 $X2=0.36 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%X 1 2 3 4 15 19 21 22 24 27 31 33 34 39 44
c64 24 0 9.97846e-20 $X=1.387 $Y=1.44
r65 42 44 7.77471 $w=6.01e-07 $l=3.83e-07 $layer=LI1_cond $X=1.387 $Y=1.742
+ $X2=1.77 $Y2=1.742
r66 37 39 4.36439 $w=6.01e-07 $l=2.15e-07 $layer=LI1_cond $X=0.83 $Y=1.742
+ $X2=1.045 $Y2=1.742
r67 34 42 4.91248 $w=6.01e-07 $l=2.42e-07 $layer=LI1_cond $X=1.145 $Y=1.742
+ $X2=1.387 $Y2=1.742
r68 34 39 2.02995 $w=6.01e-07 $l=1e-07 $layer=LI1_cond $X=1.145 $Y=1.742
+ $X2=1.045 $Y2=1.742
r69 29 44 8.32752 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=1.77 $Y=2.045
+ $X2=1.77 $Y2=1.742
r70 29 31 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.77 $Y=2.045
+ $X2=1.77 $Y2=2.3
r71 25 33 5.12578 $w=2.67e-07 $l=2.47346e-07 $layer=LI1_cond $X=1.67 $Y=0.66
+ $X2=1.48 $Y2=0.792
r72 25 27 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.67 $Y=0.66 $X2=1.67
+ $Y2=0.56
r73 24 42 3.66491 $w=3.65e-07 $l=3.02e-07 $layer=LI1_cond $X=1.387 $Y=1.44
+ $X2=1.387 $Y2=1.742
r74 23 33 5.12578 $w=2.67e-07 $l=1.73372e-07 $layer=LI1_cond $X=1.387 $Y=0.925
+ $X2=1.48 $Y2=0.792
r75 23 24 16.2605 $w=3.63e-07 $l=5.15e-07 $layer=LI1_cond $X=1.387 $Y=0.925
+ $X2=1.387 $Y2=1.44
r76 21 33 1.3764 $w=2.65e-07 $l=2.75e-07 $layer=LI1_cond $X=1.205 $Y=0.792
+ $X2=1.48 $Y2=0.792
r77 21 22 16.9605 $w=2.63e-07 $l=3.9e-07 $layer=LI1_cond $X=1.205 $Y=0.792
+ $X2=0.815 $Y2=0.792
r78 17 37 8.32752 $w=1.7e-07 $l=3.03e-07 $layer=LI1_cond $X=0.83 $Y=2.045
+ $X2=0.83 $Y2=1.742
r79 17 19 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.83 $Y=2.045
+ $X2=0.83 $Y2=2.3
r80 13 22 7.24806 $w=2.65e-07 $l=1.69245e-07 $layer=LI1_cond $X=0.73 $Y=0.66
+ $X2=0.815 $Y2=0.792
r81 13 15 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=0.73 $Y=0.66 $X2=0.73
+ $Y2=0.56
r82 4 44 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.625
+ $Y=1.485 $X2=1.77 $Y2=1.62
r83 4 31 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.485 $X2=1.77 $Y2=2.3
r84 3 37 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.685
+ $Y=1.485 $X2=0.83 $Y2=1.62
r85 3 19 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.685
+ $Y=1.485 $X2=0.83 $Y2=2.3
r86 2 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.56
r87 1 15 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_652_325# 1 2 3 4 13 18 21 23 25 27 30 32
+ 33 35 37 38 39 45 49
c147 35 0 1.24749e-19 $X=8.55 $Y=0.38
r148 48 49 11.956 $w=2.5e-07 $l=2.45e-07 $layer=LI1_cond $X=4.46 $Y=1.535
+ $X2=4.705 $Y2=1.535
r149 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.27 $Y=1.53
+ $X2=7.27 $Y2=1.53
r150 42 49 5.612 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=4.82 $Y=1.535
+ $X2=4.705 $Y2=1.535
r151 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.82 $Y=1.53
+ $X2=4.82 $Y2=1.53
r152 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.965 $Y=1.53
+ $X2=4.82 $Y2=1.53
r153 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.125 $Y=1.53
+ $X2=7.27 $Y2=1.53
r154 38 39 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=7.125 $Y=1.53
+ $X2=4.965 $Y2=1.53
r155 33 37 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=8.465 $Y=0.36
+ $X2=8.255 $Y2=0.36
r156 33 35 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=8.465 $Y=0.36
+ $X2=8.55 $Y2=0.36
r157 32 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.745 $Y=0.34
+ $X2=8.255 $Y2=0.34
r158 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.66 $Y=0.425
+ $X2=7.745 $Y2=0.34
r159 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=7.66 $Y=0.425
+ $X2=7.66 $Y2=1.445
r160 28 46 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=7.33 $Y=1.53
+ $X2=7.122 $Y2=1.53
r161 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.575 $Y=1.53
+ $X2=7.66 $Y2=1.445
r162 27 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=7.575 $Y=1.53
+ $X2=7.33 $Y2=1.53
r163 23 46 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.122 $Y=1.615
+ $X2=7.122 $Y2=1.53
r164 23 25 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=7.122 $Y=1.615
+ $X2=7.122 $Y2=1.62
r165 19 49 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.705 $Y=1.375
+ $X2=4.705 $Y2=1.535
r166 19 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.705 $Y=1.375
+ $X2=4.705 $Y2=0.76
r167 17 48 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.46 $Y=1.695
+ $X2=4.46 $Y2=1.535
r168 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.46 $Y=1.695
+ $X2=4.46 $Y2=1.895
r169 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.375 $Y=1.98
+ $X2=4.46 $Y2=1.895
r170 13 15 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=4.375 $Y=1.98
+ $X2=3.385 $Y2=1.98
r171 4 25 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=6.74
+ $Y=1.485 $X2=7.09 $Y2=1.62
r172 3 15 600 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_PDIFF $count=1 $X=3.26
+ $Y=1.625 $X2=3.385 $Y2=1.98
r173 2 35 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=8.355
+ $Y=0.245 $X2=8.55 $Y2=0.38
r174 1 21 182 $w=1.7e-07 $l=6.65507e-07 $layer=licon1_NDIFF $count=1 $X=4.36
+ $Y=0.245 $X2=4.705 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_658_49# 1 2 3 4 13 18 19 20 22 23 24 26
+ 28 29 32 33 34 36 39 43 48 50 52 53 55
r185 53 54 16.6089 $w=2.02e-07 $l=2.75e-07 $layer=LI1_cond $X=6.61 $Y=0.772
+ $X2=6.885 $Y2=0.772
r186 50 51 8.30177 $w=1.69e-07 $l=1.15e-07 $layer=LI1_cond $X=5.045 $Y=1.12
+ $X2=5.16 $Y2=1.12
r187 46 48 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.685 $Y=2.32
+ $X2=4.8 $Y2=2.32
r188 41 54 1.74864 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.885 $Y=0.655
+ $X2=6.885 $Y2=0.772
r189 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.885 $Y=0.655
+ $X2=6.885 $Y2=0.545
r190 37 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.695 $Y=2.36
+ $X2=6.61 $Y2=2.36
r191 37 39 131.134 $w=1.68e-07 $l=2.01e-06 $layer=LI1_cond $X=6.695 $Y=2.36
+ $X2=8.705 $Y2=2.36
r192 36 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=2.275
+ $X2=6.61 $Y2=2.36
r193 35 53 1.74864 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=6.61 $Y=0.89
+ $X2=6.61 $Y2=0.772
r194 35 36 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=6.61 $Y=0.89
+ $X2=6.61 $Y2=2.275
r195 33 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.525 $Y=2.36
+ $X2=6.61 $Y2=2.36
r196 33 34 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.525 $Y=2.36
+ $X2=5.99 $Y2=2.36
r197 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.905 $Y=2.275
+ $X2=5.99 $Y2=2.36
r198 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.905 $Y=2.065
+ $X2=5.905 $Y2=2.275
r199 30 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.245 $Y=1.98
+ $X2=5.16 $Y2=1.98
r200 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.82 $Y=1.98
+ $X2=5.905 $Y2=2.065
r201 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.82 $Y=1.98
+ $X2=5.245 $Y2=1.98
r202 28 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=1.895
+ $X2=5.16 $Y2=1.98
r203 27 51 0.680474 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=1.205
+ $X2=5.16 $Y2=1.12
r204 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.16 $Y=1.205
+ $X2=5.16 $Y2=1.895
r205 26 50 0.680474 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=1.035
+ $X2=5.045 $Y2=1.12
r206 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.045 $Y=0.425
+ $X2=5.045 $Y2=1.035
r207 23 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.075 $Y=1.98
+ $X2=5.16 $Y2=1.98
r208 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=5.075 $Y=1.98
+ $X2=4.885 $Y2=1.98
r209 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.8 $Y=2.235
+ $X2=4.8 $Y2=2.32
r210 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.8 $Y=2.065
+ $X2=4.885 $Y2=1.98
r211 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.8 $Y=2.065
+ $X2=4.8 $Y2=2.235
r212 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.96 $Y=0.34
+ $X2=5.045 $Y2=0.425
r213 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.96 $Y=0.34
+ $X2=4.45 $Y2=0.34
r214 17 20 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.34 $Y=0.425
+ $X2=4.45 $Y2=0.34
r215 17 18 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=4.34 $Y=0.425
+ $X2=4.34 $Y2=0.655
r216 13 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=4.23 $Y=0.74
+ $X2=4.34 $Y2=0.655
r217 13 15 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=4.23 $Y=0.74
+ $X2=3.425 $Y2=0.74
r218 4 39 600 $w=1.7e-07 $l=8.21995e-07 $layer=licon1_PDIFF $count=1 $X=8.475
+ $Y=1.645 $X2=8.705 $Y2=2.36
r219 3 46 600 $w=1.7e-07 $l=8.70373e-07 $layer=licon1_PDIFF $count=1 $X=4.29
+ $Y=1.625 $X2=4.685 $Y2=2.32
r220 2 43 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=6.75
+ $Y=0.245 $X2=6.885 $Y2=0.545
r221 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.29
+ $Y=0.245 $X2=3.425 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%A_1510_297# 1 2 3 4 15 18 23 26 29 31 36
r64 34 36 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=10.25 $Y=0.42
+ $X2=10.34 $Y2=0.42
r65 28 29 18.846 $w=2.28e-07 $l=3.6e-07 $layer=LI1_cond $X=10.25 $Y=1.99
+ $X2=9.89 $Y2=1.99
r66 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=10.34 $Y=1.875
+ $X2=10.34 $Y2=1.99
r67 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.34 $Y=0.585
+ $X2=10.34 $Y2=0.42
r68 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=10.34 $Y=0.585
+ $X2=10.34 $Y2=1.875
r69 21 31 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=10.295 $Y=1.99
+ $X2=10.34 $Y2=1.99
r70 21 28 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=10.295 $Y=1.99
+ $X2=10.25 $Y2=1.99
r71 21 23 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=10.295 $Y=2.105
+ $X2=10.295 $Y2=2.3
r72 20 29 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=8.15 $Y=2.02
+ $X2=9.89 $Y2=2.02
r73 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=8.085 $Y=2.02
+ $X2=8.15 $Y2=2.02
r74 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8 $Y=1.935
+ $X2=8.085 $Y2=2.02
r75 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=8 $Y=1.935 $X2=8
+ $Y2=0.76
r76 4 28 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=10.105
+ $Y=1.485 $X2=10.25 $Y2=1.96
r77 4 23 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.105
+ $Y=1.485 $X2=10.25 $Y2=2.3
r78 3 20 600 $w=1.7e-07 $l=8.25227e-07 $layer=licon1_PDIFF $count=1 $X=7.55
+ $Y=1.485 $X2=8.15 $Y2=2.02
r79 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=10.115
+ $Y=0.235 $X2=10.25 $Y2=0.42
r80 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=7.56
+ $Y=0.245 $X2=8 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_4%VGND 1 2 3 4 5 16 18 20 24 28 32 35 36 38
+ 39 40 42 61 62 69 75 78
r131 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r132 70 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r133 69 72 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.175 $Y=0
+ $X2=1.175 $Y2=0.38
r134 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r135 65 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r136 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r137 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r138 58 59 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r139 56 59 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r140 55 58 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=9.43
+ $Y2=0
r141 55 56 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r142 53 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r143 52 53 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r144 50 53 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=5.29 $Y2=0
r145 50 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r146 49 52 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=5.29
+ $Y2=0
r147 49 50 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r148 47 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0 $X2=2.14
+ $Y2=0
r149 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.53 $Y2=0
r150 46 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r151 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r152 43 65 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r153 43 45 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.69
+ $Y2=0
r154 42 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=1.175
+ $Y2=0
r155 42 45 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.985 $Y=0 $X2=0.69
+ $Y2=0
r156 40 46 0.10528 $w=4.8e-07 $l=3.7e-07 $layer=MET1_cond $X=0.32 $Y=0 $X2=0.69
+ $Y2=0
r157 40 78 0.0284542 $w=4.8e-07 $l=1e-07 $layer=MET1_cond $X=0.32 $Y=0 $X2=0.22
+ $Y2=0
r158 38 58 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=9.695 $Y=0
+ $X2=9.43 $Y2=0
r159 38 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.695 $Y=0 $X2=9.78
+ $Y2=0
r160 37 61 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=9.865 $Y=0
+ $X2=10.35 $Y2=0
r161 37 39 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.865 $Y=0 $X2=9.78
+ $Y2=0
r162 35 52 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.29
+ $Y2=0
r163 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.3 $Y=0 $X2=5.385
+ $Y2=0
r164 34 55 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.75
+ $Y2=0
r165 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=0 $X2=5.385
+ $Y2=0
r166 30 39 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.78 $Y=0.085
+ $X2=9.78 $Y2=0
r167 30 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.78 $Y=0.085
+ $X2=9.78 $Y2=0.4
r168 26 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.385 $Y=0.085
+ $X2=5.385 $Y2=0
r169 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.385 $Y=0.085
+ $X2=5.385 $Y2=0.38
r170 22 75 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r171 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.36
r172 21 69 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.365 $Y=0 $X2=1.175
+ $Y2=0
r173 20 75 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r174 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=1.365
+ $Y2=0
r175 16 65 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r176 16 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r177 5 32 182 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_NDIFF $count=1 $X=9.605
+ $Y=0.235 $X2=9.78 $Y2=0.4
r178 4 28 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=5.26
+ $Y=0.235 $X2=5.385 $Y2=0.38
r179 3 24 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.36
r180 2 72 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r181 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

