* File: sky130_fd_sc_hdll__a211oi_4.pxi.spice
* Created: Thu Aug 27 18:51:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211OI_4%A2 N_A2_c_109_n N_A2_M16_noxref_g N_A2_M1003_g
+ N_A2_c_110_n N_A2_M17_noxref_g N_A2_M1011_g N_A2_c_111_n N_A2_M18_noxref_g
+ N_A2_M1020_g N_A2_c_103_n N_A2_M23_noxref_g N_A2_c_104_n N_A2_M1031_g
+ N_A2_c_113_n N_A2_c_105_n A2 N_A2_c_107_n N_A2_c_108_n
+ PM_SKY130_FD_SC_HDLL__A211OI_4%A2
x_PM_SKY130_FD_SC_HDLL__A211OI_4%A1 N_A1_M1012_g N_A1_c_225_n N_A1_M19_noxref_g
+ N_A1_M1025_g N_A1_c_226_n N_A1_M20_noxref_g N_A1_M1028_g N_A1_c_227_n
+ N_A1_M21_noxref_g N_A1_c_228_n N_A1_M22_noxref_g N_A1_M1030_g A1 N_A1_c_223_n
+ N_A1_c_224_n A1 PM_SKY130_FD_SC_HDLL__A211OI_4%A1
x_PM_SKY130_FD_SC_HDLL__A211OI_4%B1 N_B1_c_290_n N_B1_M1005_g N_B1_c_298_n
+ N_B1_M24_noxref_g N_B1_c_299_n N_B1_M25_noxref_g N_B1_c_291_n N_B1_M1008_g
+ N_B1_c_300_n N_B1_M26_noxref_g N_B1_c_292_n N_B1_M1021_g N_B1_c_293_n
+ N_B1_M31_noxref_g N_B1_c_294_n N_B1_M1024_g N_B1_c_325_p N_B1_c_295_n
+ N_B1_c_303_n N_B1_c_311_n N_B1_c_304_n N_B1_c_305_n B1 N_B1_c_296_n
+ N_B1_c_297_n PM_SKY130_FD_SC_HDLL__A211OI_4%B1
x_PM_SKY130_FD_SC_HDLL__A211OI_4%C1 N_C1_c_432_n N_C1_M27_noxref_g N_C1_c_426_n
+ N_C1_M1001_g N_C1_c_433_n N_C1_M28_noxref_g N_C1_c_427_n N_C1_M1004_g
+ N_C1_c_434_n N_C1_M29_noxref_g N_C1_c_428_n N_C1_M1013_g N_C1_c_435_n
+ N_C1_M30_noxref_g N_C1_c_429_n N_C1_M1022_g N_C1_c_430_n N_C1_c_436_n C1
+ N_C1_c_431_n PM_SKY130_FD_SC_HDLL__A211OI_4%C1
x_PM_SKY130_FD_SC_HDLL__A211OI_4%noxref_7 N_noxref_7_M16_noxref_s
+ N_noxref_7_M17_noxref_d N_noxref_7_M19_noxref_d N_noxref_7_M21_noxref_d
+ N_noxref_7_M23_noxref_d N_noxref_7_M25_noxref_d N_noxref_7_M31_noxref_d
+ N_noxref_7_c_514_n N_noxref_7_c_515_n N_noxref_7_c_524_n N_noxref_7_c_561_p
+ N_noxref_7_c_528_n N_noxref_7_c_564_p N_noxref_7_c_530_n N_noxref_7_c_567_p
+ N_noxref_7_c_531_n N_noxref_7_c_533_n N_noxref_7_c_570_p N_noxref_7_c_516_n
+ N_noxref_7_c_534_n N_noxref_7_c_536_n N_noxref_7_c_537_n
+ PM_SKY130_FD_SC_HDLL__A211OI_4%noxref_7
x_PM_SKY130_FD_SC_HDLL__A211OI_4%VPWR N_VPWR_M16_noxref_d N_VPWR_M18_noxref_d
+ N_VPWR_M20_noxref_d N_VPWR_M22_noxref_d VPWR N_VPWR_c_616_n N_VPWR_c_617_n
+ N_VPWR_c_618_n N_VPWR_c_619_n N_VPWR_c_620_n N_VPWR_c_615_n N_VPWR_c_622_n
+ N_VPWR_c_623_n N_VPWR_c_624_n N_VPWR_c_625_n
+ PM_SKY130_FD_SC_HDLL__A211OI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__A211OI_4%noxref_9 N_noxref_9_M24_noxref_d
+ N_noxref_9_M28_noxref_d N_noxref_9_c_736_n N_noxref_9_c_732_n
+ N_noxref_9_c_733_n PM_SKY130_FD_SC_HDLL__A211OI_4%noxref_9
x_PM_SKY130_FD_SC_HDLL__A211OI_4%Y N_Y_M1012_s N_Y_M1028_s N_Y_M1005_s
+ N_Y_M1021_s N_Y_M1004_s N_Y_M1022_s N_Y_M27_noxref_d N_Y_M29_noxref_d
+ N_Y_c_786_n N_Y_c_787_n N_Y_c_801_n N_Y_c_882_p N_Y_c_834_n N_Y_c_807_n
+ N_Y_c_884_p N_Y_c_812_n N_Y_c_782_n N_Y_c_789_n N_Y_c_791_n N_Y_c_823_n
+ N_Y_c_852_n N_Y_c_876_p Y N_Y_c_783_n PM_SKY130_FD_SC_HDLL__A211OI_4%Y
x_PM_SKY130_FD_SC_HDLL__A211OI_4%VGND N_VGND_M1003_d N_VGND_M1011_d
+ N_VGND_M1031_d N_VGND_M1008_d N_VGND_M1001_d N_VGND_M1013_d N_VGND_M1024_d
+ N_VGND_c_924_n N_VGND_c_925_n N_VGND_c_926_n N_VGND_c_927_n N_VGND_c_928_n
+ N_VGND_c_929_n N_VGND_c_930_n N_VGND_c_931_n N_VGND_c_932_n N_VGND_c_933_n
+ N_VGND_c_934_n N_VGND_c_935_n N_VGND_c_936_n N_VGND_c_937_n N_VGND_c_938_n
+ VGND N_VGND_c_939_n N_VGND_c_940_n N_VGND_c_941_n N_VGND_c_942_n
+ N_VGND_c_943_n PM_SKY130_FD_SC_HDLL__A211OI_4%VGND
x_PM_SKY130_FD_SC_HDLL__A211OI_4%A_119_47# N_A_119_47#_M1003_s
+ N_A_119_47#_M1020_s N_A_119_47#_M1025_d N_A_119_47#_M1030_d
+ N_A_119_47#_c_1052_n N_A_119_47#_c_1058_n N_A_119_47#_c_1059_n
+ N_A_119_47#_c_1063_n N_A_119_47#_c_1061_n
+ PM_SKY130_FD_SC_HDLL__A211OI_4%A_119_47#
cc_1 VNB N_A2_M1003_g 0.0249276f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_A2_M1011_g 0.0181696f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_A2_M1020_g 0.0183466f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_A2_c_103_n 0.0214479f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_5 VNB N_A2_c_104_n 0.01695f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_6 VNB N_A2_c_105_n 0.00425679f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.16
cc_7 VNB A2 0.0157817f $X=-0.19 $Y=-0.24 $X2=1.07 $Y2=1.445
cc_8 VNB N_A2_c_107_n 0.0721733f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.217
cc_9 VNB N_A2_c_108_n 0.0021746f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.33
cc_10 VNB N_A1_M1012_g 0.0183466f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_11 VNB N_A1_M1025_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_12 VNB N_A1_M1028_g 0.0190961f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_13 VNB N_A1_M1030_g 0.0192359f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_14 VNB N_A1_c_223_n 0.00179333f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.16
cc_15 VNB N_A1_c_224_n 0.0875027f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.217
cc_16 VNB N_B1_c_290_n 0.0177008f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_B1_c_291_n 0.0178287f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_18 VNB N_B1_c_292_n 0.0173251f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_19 VNB N_B1_c_293_n 0.0254146f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_20 VNB N_B1_c_294_n 0.0189775f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_21 VNB N_B1_c_295_n 0.00372159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B1_c_296_n 0.0583184f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_B1_c_297_n 0.0017689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C1_c_426_n 0.0170033f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.025
cc_25 VNB N_C1_c_427_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_26 VNB N_C1_c_428_n 0.0167427f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_27 VNB N_C1_c_429_n 0.0172739f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_28 VNB N_C1_c_430_n 0.00215472f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_29 VNB N_C1_c_431_n 0.0767995f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.217
cc_30 VNB N_VPWR_c_615_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.16
cc_31 VNB N_Y_c_782_n 0.0111406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_783_n 0.0243148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_924_n 0.0109754f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_34 VNB N_VGND_c_925_n 0.0186333f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_35 VNB N_VGND_c_926_n 0.00224819f $X=-0.19 $Y=-0.24 $X2=3.595 $Y2=1.535
cc_36 VNB N_VGND_c_927_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.16
cc_37 VNB N_VGND_c_928_n 0.00224653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_929_n 0.00213178f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=1.217
cc_39 VNB N_VGND_c_930_n 0.00209192f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.217
cc_40 VNB N_VGND_c_931_n 0.0608139f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=1.16
cc_41 VNB N_VGND_c_932_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.217
cc_42 VNB N_VGND_c_933_n 0.0177818f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.16
cc_43 VNB N_VGND_c_934_n 0.00510002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_935_n 0.0149619f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_936_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.33
cc_46 VNB N_VGND_c_937_n 0.0146899f $X=-0.19 $Y=-0.24 $X2=1.32 $Y2=1.33
cc_47 VNB N_VGND_c_938_n 0.00507043f $X=-0.19 $Y=-0.24 $X2=1.24 $Y2=1.33
cc_48 VNB N_VGND_c_939_n 0.0163029f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_940_n 0.0146683f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_941_n 0.00399928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_942_n 0.0264203f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_943_n 0.391849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_A2_c_109_n 0.0188351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_A2_c_110_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_55 VPB N_A2_c_111_n 0.0151596f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_56 VPB N_A2_c_103_n 0.0245018f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_57 VPB N_A2_c_113_n 0.0134802f $X=-0.19 $Y=1.305 $X2=3.595 $Y2=1.535
cc_58 VPB N_A2_c_105_n 0.00230756f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.16
cc_59 VPB A2 0.0141397f $X=-0.19 $Y=1.305 $X2=1.07 $Y2=1.445
cc_60 VPB N_A2_c_107_n 0.0181642f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.217
cc_61 VPB N_A2_c_108_n 0.00172565f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.33
cc_62 VPB N_A1_c_225_n 0.0157656f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_63 VPB N_A1_c_226_n 0.0154404f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_64 VPB N_A1_c_227_n 0.0157014f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_65 VPB N_A1_c_228_n 0.0154834f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_66 VPB N_A1_c_224_n 0.0255351f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_67 VPB N_B1_c_298_n 0.0156532f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.025
cc_68 VPB N_B1_c_299_n 0.0155301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B1_c_300_n 0.0162101f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_70 VPB N_B1_c_293_n 0.0305154f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_71 VPB N_B1_c_295_n 5.09812e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_B1_c_303_n 0.00279869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B1_c_304_n 0.0016588f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.217
cc_74 VPB N_B1_c_305_n 0.00256406f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.16
cc_75 VPB N_B1_c_296_n 0.0352752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_B1_c_297_n 0.00265635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_C1_c_432_n 0.0163182f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_78 VPB N_C1_c_433_n 0.0160541f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_C1_c_434_n 0.0162115f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_80 VPB N_C1_c_435_n 0.01663f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_81 VPB N_C1_c_436_n 0.00228439f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.535
cc_82 VPB N_C1_c_431_n 0.0491383f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_83 VPB N_noxref_7_c_514_n 0.0125686f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_84 VPB N_noxref_7_c_515_n 0.0144536f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.985
cc_85 VPB N_noxref_7_c_516_n 0.00955326f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.33
cc_86 VPB N_VPWR_c_616_n 0.0143912f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_87 VPB N_VPWR_c_617_n 0.0123455f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_88 VPB N_VPWR_c_618_n 0.0123059f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.995
cc_89 VPB N_VPWR_c_619_n 0.0123059f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.445
cc_90 VPB N_VPWR_c_620_n 0.104974f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.217
cc_91 VPB N_VPWR_c_615_n 0.0470746f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=1.16
cc_92 VPB N_VPWR_c_622_n 0.00547281f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.217
cc_93 VPB N_VPWR_c_623_n 0.00537738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_624_n 0.00537738f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.33
cc_95 VPB N_VPWR_c_625_n 0.00547137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_noxref_9_c_732_n 0.00541979f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_97 VPB N_noxref_9_c_733_n 0.00218946f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_98 VPB Y 0.0275049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_Y_c_783_n 0.00967841f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 N_A2_M1020_g N_A1_M1012_g 0.0232139f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_101 N_A2_c_111_n N_A1_c_225_n 0.039255f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A2_c_113_n N_A1_c_225_n 0.0122923f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_103 N_A2_c_108_n N_A1_c_225_n 8.51953e-19 $X=1.535 $Y=1.33 $X2=0 $Y2=0
cc_104 N_A2_c_113_n N_A1_c_226_n 0.012338f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_105 N_A2_c_113_n N_A1_c_227_n 0.012338f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_106 N_A2_c_103_n N_A1_c_228_n 0.0392284f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A2_c_113_n N_A1_c_228_n 0.0136085f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_108 N_A2_c_105_n N_A1_c_228_n 8.11693e-19 $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A2_c_103_n N_A1_M1030_g 0.0219233f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A2_c_104_n N_A1_M1030_g 0.0240028f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A2_c_103_n N_A1_c_223_n 2.41204e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A2_c_113_n N_A1_c_223_n 0.108205f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_113 N_A2_c_105_n N_A1_c_223_n 0.0135224f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A2_c_107_n N_A1_c_223_n 3.004e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_115 N_A2_c_108_n N_A1_c_223_n 0.0138716f $X=1.535 $Y=1.33 $X2=0 $Y2=0
cc_116 N_A2_c_103_n N_A1_c_224_n 0.00370403f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_113_n N_A1_c_224_n 0.0220802f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_118 N_A2_c_105_n N_A1_c_224_n 0.00513015f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A2_c_107_n N_A1_c_224_n 0.0232139f $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_120 N_A2_c_108_n N_A1_c_224_n 0.00119682f $X=1.535 $Y=1.33 $X2=0 $Y2=0
cc_121 N_A2_c_104_n N_B1_c_290_n 0.0281372f $X=3.81 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_122 N_A2_c_103_n N_B1_c_298_n 0.0225535f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_113_n N_B1_c_298_n 9.48119e-19 $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_124 N_A2_c_113_n N_B1_c_311_n 0.00166216f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_125 N_A2_c_103_n N_B1_c_296_n 0.0260682f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_105_n N_B1_c_296_n 0.00124065f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_127 N_A2_c_103_n N_B1_c_297_n 0.00162342f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_113_n N_B1_c_297_n 0.0083273f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_129 N_A2_c_105_n N_B1_c_297_n 0.0363011f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_130 A2 N_noxref_7_M16_noxref_s 0.00295363f $X=1.07 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_131 A2 N_noxref_7_M17_noxref_d 0.0013695f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_132 N_A2_c_108_n N_noxref_7_M17_noxref_d 4.96997e-19 $X=1.535 $Y=1.33 $X2=0
+ $Y2=0
cc_133 N_A2_c_113_n N_noxref_7_M19_noxref_d 0.00181032f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_134 N_A2_c_113_n N_noxref_7_M21_noxref_d 0.00181032f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_135 N_A2_c_113_n N_noxref_7_M23_noxref_d 0.00153522f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_136 A2 N_noxref_7_c_514_n 0.0218555f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_137 N_A2_c_109_n N_noxref_7_c_524_n 0.0143534f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A2_c_110_n N_noxref_7_c_524_n 0.0148071f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 A2 N_noxref_7_c_524_n 0.0428155f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_140 N_A2_c_107_n N_noxref_7_c_524_n 8.48578e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_141 N_A2_c_111_n N_noxref_7_c_528_n 0.0148013f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A2_c_108_n N_noxref_7_c_528_n 0.0405214f $X=1.535 $Y=1.33 $X2=0 $Y2=0
cc_143 N_A2_c_113_n N_noxref_7_c_530_n 0.0392728f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_144 N_A2_c_103_n N_noxref_7_c_531_n 0.0153796f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_113_n N_noxref_7_c_531_n 0.040879f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_146 N_A2_c_113_n N_noxref_7_c_533_n 0.00356588f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_147 A2 N_noxref_7_c_534_n 0.0150366f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_148 N_A2_c_107_n N_noxref_7_c_534_n 6.76214e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_149 N_A2_c_113_n N_noxref_7_c_536_n 0.0138678f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_150 N_A2_c_113_n N_noxref_7_c_537_n 0.0138678f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_151 A2 N_VPWR_M16_noxref_d 0.00194857f $X=1.07 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_152 N_A2_c_113_n N_VPWR_M18_noxref_d 0.00187879f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_153 N_A2_c_113_n N_VPWR_M20_noxref_d 0.00187879f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_154 N_A2_c_113_n N_VPWR_M22_noxref_d 0.001873f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_155 N_A2_c_109_n N_VPWR_c_616_n 0.00311736f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A2_c_110_n N_VPWR_c_617_n 0.00453434f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A2_c_111_n N_VPWR_c_617_n 0.00309549f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_103_n N_VPWR_c_620_n 0.00450253f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A2_c_109_n N_VPWR_c_615_n 0.0046225f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A2_c_110_n N_VPWR_c_615_n 0.00513756f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A2_c_111_n N_VPWR_c_615_n 0.00367588f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_103_n N_VPWR_c_615_n 0.00511159f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_109_n N_VPWR_c_622_n 0.0110296f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_110_n N_VPWR_c_622_n 0.0067928f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A2_c_111_n N_VPWR_c_622_n 4.88209e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_110_n N_VPWR_c_623_n 5.3082e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_111_n N_VPWR_c_623_n 0.00911887f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_103_n N_VPWR_c_625_n 0.00756943f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A2_c_113_n N_Y_c_786_n 0.00748359f $X=3.595 $Y=1.535 $X2=0 $Y2=0
cc_170 N_A2_c_103_n N_Y_c_787_n 0.00127448f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A2_c_104_n N_Y_c_787_n 0.0121896f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A2_c_103_n N_Y_c_789_n 0.00262806f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A2_c_105_n N_Y_c_789_n 0.0251565f $X=3.76 $Y=1.16 $X2=0 $Y2=0
cc_174 N_A2_c_104_n N_Y_c_791_n 9.00022e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A2_M1003_g N_VGND_c_925_n 0.00335108f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_176 A2 N_VGND_c_925_n 0.0130826f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_177 N_A2_c_107_n N_VGND_c_925_n 3.33405e-19 $X=1.435 $Y=1.217 $X2=0 $Y2=0
cc_178 N_A2_M1003_g N_VGND_c_926_n 0.00138649f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_179 N_A2_M1011_g N_VGND_c_926_n 0.0117833f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_180 N_A2_M1020_g N_VGND_c_926_n 0.00377152f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_181 N_A2_c_104_n N_VGND_c_927_n 0.00268723f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_M1020_g N_VGND_c_931_n 0.00393157f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A2_c_104_n N_VGND_c_931_n 0.00433717f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A2_M1003_g N_VGND_c_939_n 0.00585385f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A2_M1011_g N_VGND_c_939_n 0.00245007f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A2_M1003_g N_VGND_c_943_n 0.0117437f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_187 N_A2_M1011_g N_VGND_c_943_n 0.00323974f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_188 N_A2_M1020_g N_VGND_c_943_n 0.00568988f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_189 N_A2_c_104_n N_VGND_c_943_n 0.00598582f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_M1011_g N_A_119_47#_c_1052_n 0.00951185f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A2_M1020_g N_A_119_47#_c_1052_n 0.00982742f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_192 N_A2_c_113_n N_A_119_47#_c_1052_n 0.0063014f $X=3.595 $Y=1.535 $X2=0
+ $Y2=0
cc_193 A2 N_A_119_47#_c_1052_n 0.0418614f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_194 N_A2_c_107_n N_A_119_47#_c_1052_n 0.00304778f $X=1.435 $Y=1.217 $X2=0
+ $Y2=0
cc_195 N_A2_c_108_n N_A_119_47#_c_1052_n 0.00661089f $X=1.535 $Y=1.33 $X2=0
+ $Y2=0
cc_196 N_A2_M1020_g N_A_119_47#_c_1058_n 0.00415162f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_197 N_A2_M1011_g N_A_119_47#_c_1059_n 5.18971e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_198 N_A2_M1020_g N_A_119_47#_c_1059_n 0.00535368f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_199 A2 N_A_119_47#_c_1061_n 0.0155201f $X=1.07 $Y=1.445 $X2=0 $Y2=0
cc_200 N_A2_c_107_n N_A_119_47#_c_1061_n 0.00308075f $X=1.435 $Y=1.217 $X2=0
+ $Y2=0
cc_201 N_A1_c_225_n N_noxref_7_c_528_n 0.0152244f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A1_c_226_n N_noxref_7_c_530_n 0.0148803f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A1_c_227_n N_noxref_7_c_530_n 0.0153033f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A1_c_228_n N_noxref_7_c_531_n 0.0148013f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_225_n N_VPWR_c_618_n 0.00450253f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A1_c_226_n N_VPWR_c_618_n 0.00309549f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A1_c_227_n N_VPWR_c_619_n 0.00450253f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A1_c_228_n N_VPWR_c_619_n 0.00309549f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A1_c_225_n N_VPWR_c_615_n 0.00508637f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A1_c_226_n N_VPWR_c_615_n 0.00367588f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A1_c_227_n N_VPWR_c_615_n 0.00508637f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A1_c_228_n N_VPWR_c_615_n 0.00367588f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A1_c_225_n N_VPWR_c_623_n 0.00652571f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A1_c_226_n N_VPWR_c_623_n 4.81844e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A1_c_225_n N_VPWR_c_624_n 5.3082e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A1_c_226_n N_VPWR_c_624_n 0.00915194f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A1_c_227_n N_VPWR_c_624_n 0.00655878f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A1_c_228_n N_VPWR_c_624_n 4.81844e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A1_c_227_n N_VPWR_c_625_n 5.3082e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A1_c_228_n N_VPWR_c_625_n 0.00911887f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A1_M1012_g N_Y_c_786_n 0.00275966f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A1_M1025_g N_Y_c_786_n 0.00922564f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A1_M1028_g N_Y_c_786_n 0.00922564f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A1_M1030_g N_Y_c_786_n 0.0105489f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A1_c_223_n N_Y_c_786_n 0.086599f $X=3.14 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A1_c_224_n N_Y_c_786_n 0.0102592f $X=3.315 $Y=1.217 $X2=0 $Y2=0
cc_227 N_A1_M1012_g N_VGND_c_931_n 0.00357877f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A1_M1025_g N_VGND_c_931_n 0.00357877f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A1_M1028_g N_VGND_c_931_n 0.00357877f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A1_M1030_g N_VGND_c_931_n 0.00357877f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_231 N_A1_M1012_g N_VGND_c_943_n 0.00538422f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_232 N_A1_M1025_g N_VGND_c_943_n 0.00548399f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A1_M1028_g N_VGND_c_943_n 0.00560377f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A1_M1030_g N_VGND_c_943_n 0.00562222f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_235 N_A1_M1012_g N_A_119_47#_c_1063_n 0.0115833f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_236 N_A1_M1025_g N_A_119_47#_c_1063_n 0.0101441f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A1_M1028_g N_A_119_47#_c_1063_n 0.0105263f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_238 N_A1_M1030_g N_A_119_47#_c_1063_n 0.0105263f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_239 N_A1_c_223_n N_A_119_47#_c_1063_n 0.00337712f $X=3.14 $Y=1.16 $X2=0 $Y2=0
cc_240 N_B1_c_300_n N_C1_c_432_n 0.046689f $X=5.195 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_241 N_B1_c_292_n N_C1_c_426_n 0.0103831f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B1_c_303_n N_C1_c_434_n 0.00367117f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_243 N_B1_c_293_n N_C1_c_435_n 0.0456716f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_244 N_B1_c_303_n N_C1_c_435_n 0.0110937f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_245 N_B1_c_304_n N_C1_c_435_n 0.00156497f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_246 N_B1_c_305_n N_C1_c_435_n 0.00165848f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_247 N_B1_c_294_n N_C1_c_429_n 0.0212301f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_c_325_p N_C1_c_430_n 0.0161108f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_249 N_B1_c_303_n N_C1_c_430_n 0.0136562f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_250 N_B1_c_296_n N_C1_c_430_n 0.00185061f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_251 N_B1_c_295_n N_C1_c_436_n 0.0183176f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B1_c_303_n N_C1_c_436_n 0.0139703f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_253 N_B1_c_304_n N_C1_c_436_n 0.00253014f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_254 N_B1_c_305_n N_C1_c_436_n 0.0119466f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_255 N_B1_c_293_n N_C1_c_431_n 0.0242647f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B1_c_325_p N_C1_c_431_n 2.52572e-19 $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_257 N_B1_c_295_n N_C1_c_431_n 0.00396132f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_258 N_B1_c_303_n N_C1_c_431_n 0.00322928f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_259 N_B1_c_305_n N_C1_c_431_n 7.84743e-19 $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_260 N_B1_c_296_n N_C1_c_431_n 0.0273394f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_261 N_B1_c_303_n N_noxref_7_M25_noxref_d 0.00116348f $X=7.28 $Y=1.53 $X2=0
+ $Y2=0
cc_262 N_B1_c_297_n N_noxref_7_M25_noxref_d 0.00163863f $X=4.96 $Y=1.325 $X2=0
+ $Y2=0
cc_263 N_B1_c_298_n N_noxref_7_c_516_n 0.01165f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B1_c_299_n N_noxref_7_c_516_n 0.0100267f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B1_c_300_n N_noxref_7_c_516_n 0.0102134f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B1_c_293_n N_noxref_7_c_516_n 0.0102822f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B1_c_311_n N_noxref_7_c_516_n 0.00114739f $X=4.515 $Y=1.53 $X2=0 $Y2=0
cc_268 N_B1_c_297_n N_noxref_7_c_516_n 0.0020586f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_269 N_B1_c_298_n N_VPWR_c_620_n 0.00429453f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B1_c_299_n N_VPWR_c_620_n 0.00429453f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B1_c_300_n N_VPWR_c_620_n 0.00429453f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B1_c_293_n N_VPWR_c_620_n 0.00429453f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B1_c_298_n N_VPWR_c_615_n 0.00609021f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B1_c_299_n N_VPWR_c_615_n 0.00606499f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B1_c_300_n N_VPWR_c_615_n 0.00615459f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B1_c_293_n N_VPWR_c_615_n 0.00718326f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B1_c_298_n N_VPWR_c_625_n 0.00100567f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B1_c_311_n N_noxref_9_M24_noxref_d 0.0018074f $X=4.515 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_279 N_B1_c_297_n N_noxref_9_M24_noxref_d 0.00123452f $X=4.96 $Y=1.325
+ $X2=-0.19 $Y2=-0.24
cc_280 N_B1_c_298_n N_noxref_9_c_736_n 0.00638325f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_281 N_B1_c_299_n N_noxref_9_c_736_n 0.0138426f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B1_c_300_n N_noxref_9_c_736_n 0.00620876f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B1_c_325_p N_noxref_9_c_736_n 0.0019017f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B1_c_303_n N_noxref_9_c_736_n 0.00842081f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_285 N_B1_c_311_n N_noxref_9_c_736_n 0.00660439f $X=4.515 $Y=1.53 $X2=0 $Y2=0
cc_286 N_B1_c_296_n N_noxref_9_c_736_n 0.00378307f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_287 N_B1_c_297_n N_noxref_9_c_736_n 0.0372219f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_288 N_B1_c_300_n N_noxref_9_c_732_n 2.71904e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_289 N_B1_c_303_n N_noxref_9_c_732_n 0.0549799f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_290 N_B1_c_299_n N_noxref_9_c_733_n 0.00144139f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B1_c_300_n N_noxref_9_c_733_n 0.0228638f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B1_c_325_p N_noxref_9_c_733_n 0.0124633f $X=5.09 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B1_c_303_n N_noxref_9_c_733_n 0.0270528f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_294 N_B1_c_311_n N_noxref_9_c_733_n 0.0010382f $X=4.515 $Y=1.53 $X2=0 $Y2=0
cc_295 N_B1_c_296_n N_noxref_9_c_733_n 0.00288506f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_296 N_B1_c_297_n N_noxref_9_c_733_n 0.0119831f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_297 N_B1_c_303_n N_Y_M29_noxref_d 8.82306e-19 $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_298 N_B1_c_290_n N_Y_c_787_n 0.00889752f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_299 N_B1_c_297_n N_Y_c_787_n 0.00932849f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_300 N_B1_c_290_n N_Y_c_801_n 2.03469e-19 $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_301 N_B1_c_291_n N_Y_c_801_n 0.0143323f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_302 N_B1_c_292_n N_Y_c_801_n 0.0127823f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_303 N_B1_c_303_n N_Y_c_801_n 0.00200247f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_304 N_B1_c_296_n N_Y_c_801_n 0.00381167f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_305 N_B1_c_297_n N_Y_c_801_n 0.0424934f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_306 N_B1_c_293_n N_Y_c_807_n 0.0108914f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_307 N_B1_c_295_n N_Y_c_807_n 0.00345904f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_308 N_B1_c_303_n N_Y_c_807_n 0.0206449f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_309 N_B1_c_304_n N_Y_c_807_n 0.0043469f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_310 N_B1_c_305_n N_Y_c_807_n 0.0122579f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_311 N_B1_c_303_n N_Y_c_812_n 0.00105829f $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_312 N_B1_c_293_n N_Y_c_782_n 0.00262257f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_313 N_B1_c_294_n N_Y_c_782_n 0.012219f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B1_c_295_n N_Y_c_782_n 0.0299036f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_315 N_B1_c_304_n N_Y_c_782_n 6.72968e-19 $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_316 N_B1_c_290_n N_Y_c_791_n 0.016256f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B1_c_291_n N_Y_c_791_n 0.00715102f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B1_c_303_n N_Y_c_791_n 4.8542e-19 $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_319 N_B1_c_311_n N_Y_c_791_n 9.38335e-19 $X=4.515 $Y=1.53 $X2=0 $Y2=0
cc_320 N_B1_c_296_n N_Y_c_791_n 0.00610569f $X=5.195 $Y=1.202 $X2=0 $Y2=0
cc_321 N_B1_c_297_n N_Y_c_791_n 0.0280361f $X=4.96 $Y=1.325 $X2=0 $Y2=0
cc_322 N_B1_c_303_n N_Y_c_823_n 9.96425e-19 $X=7.28 $Y=1.53 $X2=0 $Y2=0
cc_323 N_B1_c_293_n Y 0.0245765f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_324 N_B1_c_295_n Y 0.00426192f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_325 N_B1_c_304_n Y 0.00513795f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_326 N_B1_c_305_n Y 0.0106725f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_327 N_B1_c_293_n N_Y_c_783_n 0.0119812f $X=7.665 $Y=1.41 $X2=0 $Y2=0
cc_328 N_B1_c_294_n N_Y_c_783_n 0.00607288f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_329 N_B1_c_295_n N_Y_c_783_n 0.0260895f $X=7.6 $Y=1.16 $X2=0 $Y2=0
cc_330 N_B1_c_304_n N_Y_c_783_n 0.00228238f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_331 N_B1_c_305_n N_Y_c_783_n 0.00618043f $X=7.425 $Y=1.53 $X2=0 $Y2=0
cc_332 N_B1_c_303_n noxref_12 2.99984e-19 $X=7.28 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_333 N_B1_c_304_n noxref_12 0.00247248f $X=7.425 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_334 N_B1_c_305_n noxref_12 0.00501617f $X=7.425 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_335 N_B1_c_290_n N_VGND_c_927_n 0.00268723f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B1_c_290_n N_VGND_c_928_n 0.00104422f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_337 N_B1_c_291_n N_VGND_c_928_n 0.00767007f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_338 N_B1_c_292_n N_VGND_c_928_n 0.00168617f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B1_c_292_n N_VGND_c_929_n 5.21577e-19 $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B1_c_290_n N_VGND_c_933_n 0.00420025f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B1_c_291_n N_VGND_c_933_n 0.00351072f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B1_c_292_n N_VGND_c_935_n 0.00422112f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_343 N_B1_c_294_n N_VGND_c_940_n 0.00224438f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_344 N_B1_c_294_n N_VGND_c_942_n 0.011654f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_345 N_B1_c_290_n N_VGND_c_943_n 0.00611438f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_346 N_B1_c_291_n N_VGND_c_943_n 0.00448048f $X=4.815 $Y=0.995 $X2=0 $Y2=0
cc_347 N_B1_c_292_n N_VGND_c_943_n 0.00586577f $X=5.295 $Y=0.995 $X2=0 $Y2=0
cc_348 N_B1_c_294_n N_VGND_c_943_n 0.00302906f $X=7.66 $Y=0.995 $X2=0 $Y2=0
cc_349 N_C1_c_432_n N_noxref_7_c_516_n 0.0143764f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_350 N_C1_c_433_n N_noxref_7_c_516_n 0.0128283f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_351 N_C1_c_434_n N_noxref_7_c_516_n 0.0129691f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_352 N_C1_c_435_n N_noxref_7_c_516_n 0.0131148f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_353 N_C1_c_432_n N_VPWR_c_620_n 0.00429453f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_354 N_C1_c_433_n N_VPWR_c_620_n 0.00429453f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_355 N_C1_c_434_n N_VPWR_c_620_n 0.00429453f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_356 N_C1_c_435_n N_VPWR_c_620_n 0.00429453f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_357 N_C1_c_432_n N_VPWR_c_615_n 0.00623092f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_358 N_C1_c_433_n N_VPWR_c_615_n 0.00615861f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_359 N_C1_c_434_n N_VPWR_c_615_n 0.00620984f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_360 N_C1_c_435_n N_VPWR_c_615_n 0.00630544f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_361 N_C1_c_432_n N_noxref_9_c_732_n 0.0158668f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_362 N_C1_c_433_n N_noxref_9_c_732_n 0.0127349f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_363 N_C1_c_434_n N_noxref_9_c_732_n 0.00457561f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_364 N_C1_c_430_n N_noxref_9_c_732_n 0.0717187f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_365 N_C1_c_436_n N_noxref_9_c_732_n 0.0143237f $X=6.885 $Y=1.16 $X2=0 $Y2=0
cc_366 N_C1_c_431_n N_noxref_9_c_732_n 0.0164942f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_367 N_C1_c_432_n N_noxref_9_c_733_n 0.00636651f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_368 N_C1_c_436_n N_Y_M29_noxref_d 0.00528592f $X=6.885 $Y=1.16 $X2=0 $Y2=0
cc_369 N_C1_c_426_n N_Y_c_834_n 0.0116741f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_370 N_C1_c_427_n N_Y_c_834_n 0.0119432f $X=6.24 $Y=0.995 $X2=0 $Y2=0
cc_371 N_C1_c_430_n N_Y_c_834_n 0.0466473f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_372 N_C1_c_431_n N_Y_c_834_n 0.00591975f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_373 N_C1_c_432_n N_Y_c_807_n 0.00518552f $X=5.695 $Y=1.41 $X2=0 $Y2=0
cc_374 N_C1_c_433_n N_Y_c_807_n 0.0112999f $X=6.175 $Y=1.41 $X2=0 $Y2=0
cc_375 N_C1_c_434_n N_Y_c_807_n 0.0128645f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_376 N_C1_c_435_n N_Y_c_807_n 0.012216f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_377 N_C1_c_430_n N_Y_c_807_n 0.00197922f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_378 N_C1_c_436_n N_Y_c_807_n 0.0136151f $X=6.885 $Y=1.16 $X2=0 $Y2=0
cc_379 N_C1_c_431_n N_Y_c_807_n 0.00203065f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_380 N_C1_c_428_n N_Y_c_812_n 0.0117921f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_381 N_C1_c_430_n N_Y_c_812_n 0.0171332f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_382 N_C1_c_436_n N_Y_c_812_n 0.0167606f $X=6.885 $Y=1.16 $X2=0 $Y2=0
cc_383 N_C1_c_431_n N_Y_c_812_n 0.00355113f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_384 N_C1_c_429_n N_Y_c_782_n 0.0157488f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_385 N_C1_c_430_n N_Y_c_823_n 0.00362434f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_386 N_C1_c_431_n N_Y_c_823_n 3.65018e-19 $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_387 N_C1_c_430_n N_Y_c_852_n 0.0129498f $X=6.83 $Y=1.155 $X2=0 $Y2=0
cc_388 N_C1_c_431_n N_Y_c_852_n 0.00316255f $X=7.155 $Y=1.202 $X2=0 $Y2=0
cc_389 N_C1_c_435_n Y 0.00113842f $X=7.155 $Y=1.41 $X2=0 $Y2=0
cc_390 N_C1_c_426_n N_VGND_c_929_n 0.00690582f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_391 N_C1_c_427_n N_VGND_c_929_n 0.00167984f $X=6.24 $Y=0.995 $X2=0 $Y2=0
cc_392 N_C1_c_427_n N_VGND_c_930_n 5.21725e-19 $X=6.24 $Y=0.995 $X2=0 $Y2=0
cc_393 N_C1_c_428_n N_VGND_c_930_n 0.00686982f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_394 N_C1_c_429_n N_VGND_c_930_n 0.00163785f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_395 N_C1_c_426_n N_VGND_c_935_n 0.00338189f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_396 N_C1_c_427_n N_VGND_c_937_n 0.0042361f $X=6.24 $Y=0.995 $X2=0 $Y2=0
cc_397 N_C1_c_428_n N_VGND_c_937_n 0.00337001f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_398 N_C1_c_429_n N_VGND_c_940_n 0.00422112f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_399 N_C1_c_429_n N_VGND_c_942_n 0.00117123f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_400 N_C1_c_426_n N_VGND_c_943_n 0.00408147f $X=5.77 $Y=0.995 $X2=0 $Y2=0
cc_401 N_C1_c_427_n N_VGND_c_943_n 0.00582317f $X=6.24 $Y=0.995 $X2=0 $Y2=0
cc_402 N_C1_c_428_n N_VGND_c_943_n 0.00403265f $X=6.71 $Y=0.995 $X2=0 $Y2=0
cc_403 N_C1_c_429_n N_VGND_c_943_n 0.00588951f $X=7.18 $Y=0.995 $X2=0 $Y2=0
cc_404 N_noxref_7_c_524_n N_VPWR_M16_noxref_d 0.00352421f $X=1.115 $Y=1.94
+ $X2=-0.19 $Y2=1.305
cc_405 N_noxref_7_c_528_n N_VPWR_M18_noxref_d 0.00373688f $X=2.055 $Y=1.95 $X2=0
+ $Y2=0
cc_406 N_noxref_7_c_530_n N_VPWR_M20_noxref_d 0.00352431f $X=2.995 $Y=1.95 $X2=0
+ $Y2=0
cc_407 N_noxref_7_c_531_n N_VPWR_M22_noxref_d 0.00371889f $X=3.935 $Y=1.95 $X2=0
+ $Y2=0
cc_408 N_noxref_7_c_515_n N_VPWR_c_616_n 0.017474f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_409 N_noxref_7_c_524_n N_VPWR_c_616_n 0.0024418f $X=1.115 $Y=1.94 $X2=0 $Y2=0
cc_410 N_noxref_7_c_524_n N_VPWR_c_617_n 0.0032881f $X=1.115 $Y=1.94 $X2=0 $Y2=0
cc_411 N_noxref_7_c_561_p N_VPWR_c_617_n 0.011801f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_412 N_noxref_7_c_528_n N_VPWR_c_617_n 0.00257067f $X=2.055 $Y=1.95 $X2=0
+ $Y2=0
cc_413 N_noxref_7_c_528_n N_VPWR_c_618_n 0.00346124f $X=2.055 $Y=1.95 $X2=0
+ $Y2=0
cc_414 N_noxref_7_c_564_p N_VPWR_c_618_n 0.011801f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_415 N_noxref_7_c_530_n N_VPWR_c_618_n 0.00257067f $X=2.995 $Y=1.95 $X2=0
+ $Y2=0
cc_416 N_noxref_7_c_530_n N_VPWR_c_619_n 0.00346124f $X=2.995 $Y=1.95 $X2=0
+ $Y2=0
cc_417 N_noxref_7_c_567_p N_VPWR_c_619_n 0.011801f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_418 N_noxref_7_c_531_n N_VPWR_c_619_n 0.00257067f $X=3.935 $Y=1.95 $X2=0
+ $Y2=0
cc_419 N_noxref_7_c_531_n N_VPWR_c_620_n 0.00346124f $X=3.935 $Y=1.95 $X2=0
+ $Y2=0
cc_420 N_noxref_7_c_570_p N_VPWR_c_620_n 0.0119415f $X=4.02 $Y=2.255 $X2=0 $Y2=0
cc_421 N_noxref_7_c_516_n N_VPWR_c_620_n 0.225533f $X=7.9 $Y=2.34 $X2=0 $Y2=0
cc_422 N_noxref_7_M16_noxref_s N_VPWR_c_615_n 0.00238238f $X=0.135 $Y=1.485
+ $X2=0 $Y2=0
cc_423 N_noxref_7_M17_noxref_d N_VPWR_c_615_n 0.00271014f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_424 N_noxref_7_M19_noxref_d N_VPWR_c_615_n 0.00269325f $X=1.995 $Y=1.485
+ $X2=0 $Y2=0
cc_425 N_noxref_7_M21_noxref_d N_VPWR_c_615_n 0.00269325f $X=2.935 $Y=1.485
+ $X2=0 $Y2=0
cc_426 N_noxref_7_M23_noxref_d N_VPWR_c_615_n 0.00251101f $X=3.875 $Y=1.485
+ $X2=0 $Y2=0
cc_427 N_noxref_7_M25_noxref_d N_VPWR_c_615_n 0.00231289f $X=4.815 $Y=1.485
+ $X2=0 $Y2=0
cc_428 N_noxref_7_M31_noxref_d N_VPWR_c_615_n 0.00217543f $X=7.755 $Y=1.485
+ $X2=0 $Y2=0
cc_429 N_noxref_7_c_515_n N_VPWR_c_615_n 0.00954719f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_430 N_noxref_7_c_524_n N_VPWR_c_615_n 0.0115793f $X=1.115 $Y=1.94 $X2=0 $Y2=0
cc_431 N_noxref_7_c_561_p N_VPWR_c_615_n 0.00646745f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_432 N_noxref_7_c_528_n N_VPWR_c_615_n 0.0118582f $X=2.055 $Y=1.95 $X2=0 $Y2=0
cc_433 N_noxref_7_c_564_p N_VPWR_c_615_n 0.00646745f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_434 N_noxref_7_c_530_n N_VPWR_c_615_n 0.0118582f $X=2.995 $Y=1.95 $X2=0 $Y2=0
cc_435 N_noxref_7_c_567_p N_VPWR_c_615_n 0.00646745f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_436 N_noxref_7_c_531_n N_VPWR_c_615_n 0.0118582f $X=3.935 $Y=1.95 $X2=0 $Y2=0
cc_437 N_noxref_7_c_570_p N_VPWR_c_615_n 0.00654444f $X=4.02 $Y=2.255 $X2=0
+ $Y2=0
cc_438 N_noxref_7_c_516_n N_VPWR_c_615_n 0.141495f $X=7.9 $Y=2.34 $X2=0 $Y2=0
cc_439 N_noxref_7_c_515_n N_VPWR_c_622_n 0.016131f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_440 N_noxref_7_c_524_n N_VPWR_c_622_n 0.0203416f $X=1.115 $Y=1.94 $X2=0 $Y2=0
cc_441 N_noxref_7_c_561_p N_VPWR_c_622_n 0.0128538f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_442 N_noxref_7_c_561_p N_VPWR_c_623_n 0.0141845f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_443 N_noxref_7_c_528_n N_VPWR_c_623_n 0.0203018f $X=2.055 $Y=1.95 $X2=0 $Y2=0
cc_444 N_noxref_7_c_564_p N_VPWR_c_623_n 0.0116296f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_445 N_noxref_7_c_564_p N_VPWR_c_624_n 0.0141845f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_446 N_noxref_7_c_530_n N_VPWR_c_624_n 0.0203018f $X=2.995 $Y=1.95 $X2=0 $Y2=0
cc_447 N_noxref_7_c_567_p N_VPWR_c_624_n 0.0116296f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_448 N_noxref_7_c_567_p N_VPWR_c_625_n 0.0141845f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_449 N_noxref_7_c_531_n N_VPWR_c_625_n 0.0203018f $X=3.935 $Y=1.95 $X2=0 $Y2=0
cc_450 N_noxref_7_c_570_p N_VPWR_c_625_n 0.0129886f $X=4.02 $Y=2.255 $X2=0 $Y2=0
cc_451 N_noxref_7_c_516_n N_noxref_9_M24_noxref_d 0.00353637f $X=7.9 $Y=2.34
+ $X2=-0.19 $Y2=1.305
cc_452 N_noxref_7_c_516_n N_noxref_9_M28_noxref_d 0.00375335f $X=7.9 $Y=2.34
+ $X2=0 $Y2=0
cc_453 N_noxref_7_M25_noxref_d N_noxref_9_c_736_n 0.00375343f $X=4.815 $Y=1.485
+ $X2=0 $Y2=0
cc_454 N_noxref_7_c_533_n N_noxref_9_c_736_n 0.0252594f $X=4.02 $Y=2.105 $X2=0
+ $Y2=0
cc_455 N_noxref_7_c_516_n N_noxref_9_c_736_n 0.044002f $X=7.9 $Y=2.34 $X2=0
+ $Y2=0
cc_456 N_noxref_7_c_516_n N_noxref_9_c_732_n 0.00581426f $X=7.9 $Y=2.34 $X2=0
+ $Y2=0
cc_457 N_noxref_7_c_516_n N_noxref_9_c_733_n 0.0202793f $X=7.9 $Y=2.34 $X2=0
+ $Y2=0
cc_458 N_noxref_7_c_516_n noxref_10 0.00489103f $X=7.9 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_459 N_noxref_7_c_516_n N_Y_M27_noxref_d 0.00375335f $X=7.9 $Y=2.34 $X2=0
+ $Y2=0
cc_460 N_noxref_7_c_516_n N_Y_M29_noxref_d 0.00415694f $X=7.9 $Y=2.34 $X2=0
+ $Y2=0
cc_461 N_noxref_7_c_516_n N_Y_c_807_n 0.103509f $X=7.9 $Y=2.34 $X2=0 $Y2=0
cc_462 N_noxref_7_M31_noxref_d Y 0.00705879f $X=7.755 $Y=1.485 $X2=0 $Y2=0
cc_463 N_noxref_7_c_516_n Y 0.0254904f $X=7.9 $Y=2.34 $X2=0 $Y2=0
cc_464 N_noxref_7_c_516_n noxref_12 0.0043297f $X=7.9 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_465 N_VPWR_c_615_n N_noxref_9_M24_noxref_d 0.00232895f $X=8.05 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_466 N_VPWR_c_615_n N_noxref_9_M28_noxref_d 0.00240926f $X=8.05 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_615_n noxref_10 0.00256987f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_468 N_VPWR_c_615_n N_Y_M27_noxref_d 0.00240926f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_469 N_VPWR_c_615_n N_Y_M29_noxref_d 0.00256987f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_470 N_VPWR_c_620_n Y 0.00180709f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_c_615_n Y 0.00362255f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_472 N_VPWR_c_615_n noxref_12 0.00265018f $X=8.05 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_473 N_noxref_9_c_732_n noxref_10 0.00193908f $X=6.415 $Y=1.61 $X2=-0.19
+ $Y2=1.305
cc_474 N_noxref_9_c_733_n noxref_10 0.00578553f $X=5.295 $Y=1.57 $X2=-0.19
+ $Y2=1.305
cc_475 N_noxref_9_c_732_n N_Y_M27_noxref_d 0.00200574f $X=6.415 $Y=1.61 $X2=0
+ $Y2=0
cc_476 N_noxref_9_c_733_n N_Y_c_801_n 0.00283531f $X=5.295 $Y=1.57 $X2=0 $Y2=0
cc_477 N_noxref_9_M28_noxref_d N_Y_c_807_n 0.00359876f $X=6.265 $Y=1.485 $X2=0
+ $Y2=0
cc_478 N_noxref_9_c_732_n N_Y_c_807_n 0.0452041f $X=6.415 $Y=1.61 $X2=0 $Y2=0
cc_479 N_noxref_9_c_733_n N_Y_c_807_n 0.012939f $X=5.295 $Y=1.57 $X2=0 $Y2=0
cc_480 N_noxref_9_c_732_n N_Y_c_823_n 0.00246739f $X=6.415 $Y=1.61 $X2=0 $Y2=0
cc_481 N_noxref_9_c_733_n N_Y_c_823_n 0.00100183f $X=5.295 $Y=1.57 $X2=0 $Y2=0
cc_482 N_Y_c_807_n noxref_12 0.00453035f $X=7.68 $Y=1.975 $X2=-0.19 $Y2=-0.24
cc_483 N_Y_c_787_n N_VGND_M1031_d 0.00665097f $X=4.275 $Y=0.78 $X2=0 $Y2=0
cc_484 N_Y_c_801_n N_VGND_M1008_d 0.00415578f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_485 N_Y_c_834_n N_VGND_M1001_d 0.00402934f $X=6.365 $Y=0.745 $X2=0 $Y2=0
cc_486 N_Y_c_812_n N_VGND_M1013_d 0.00169165f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_487 N_Y_c_876_p N_VGND_M1013_d 0.00226647f $X=7.055 $Y=0.74 $X2=0 $Y2=0
cc_488 N_Y_c_782_n N_VGND_M1024_d 0.00594168f $X=7.905 $Y=0.72 $X2=0 $Y2=0
cc_489 N_Y_c_783_n N_VGND_M1024_d 0.00107792f $X=7.92 $Y=1.495 $X2=0 $Y2=0
cc_490 N_Y_c_787_n N_VGND_c_927_n 0.012114f $X=4.275 $Y=0.78 $X2=0 $Y2=0
cc_491 N_Y_c_801_n N_VGND_c_928_n 0.0184994f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_492 N_Y_c_791_n N_VGND_c_928_n 0.0122063f $X=4.51 $Y=0.42 $X2=0 $Y2=0
cc_493 N_Y_c_882_p N_VGND_c_929_n 0.0115031f $X=5.51 $Y=0.42 $X2=0 $Y2=0
cc_494 N_Y_c_834_n N_VGND_c_929_n 0.0171863f $X=6.365 $Y=0.745 $X2=0 $Y2=0
cc_495 N_Y_c_884_p N_VGND_c_930_n 0.0115031f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_496 N_Y_c_812_n N_VGND_c_930_n 0.0180515f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_497 N_Y_c_787_n N_VGND_c_931_n 0.00272119f $X=4.275 $Y=0.78 $X2=0 $Y2=0
cc_498 N_Y_c_787_n N_VGND_c_933_n 0.00212504f $X=4.275 $Y=0.78 $X2=0 $Y2=0
cc_499 N_Y_c_801_n N_VGND_c_933_n 0.00348728f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_500 N_Y_c_791_n N_VGND_c_933_n 0.0236575f $X=4.51 $Y=0.42 $X2=0 $Y2=0
cc_501 N_Y_c_801_n N_VGND_c_935_n 0.00344289f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_502 N_Y_c_882_p N_VGND_c_935_n 0.011686f $X=5.51 $Y=0.42 $X2=0 $Y2=0
cc_503 N_Y_c_834_n N_VGND_c_935_n 0.00338855f $X=6.365 $Y=0.745 $X2=0 $Y2=0
cc_504 N_Y_c_834_n N_VGND_c_937_n 0.00325342f $X=6.365 $Y=0.745 $X2=0 $Y2=0
cc_505 N_Y_c_884_p N_VGND_c_937_n 0.0115146f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_506 N_Y_c_812_n N_VGND_c_937_n 0.00347761f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_507 N_Y_c_782_n N_VGND_c_940_n 0.00935325f $X=7.905 $Y=0.72 $X2=0 $Y2=0
cc_508 N_Y_c_782_n N_VGND_c_942_n 0.0295198f $X=7.905 $Y=0.72 $X2=0 $Y2=0
cc_509 N_Y_M1012_s N_VGND_c_943_n 0.00256987f $X=1.955 $Y=0.235 $X2=0 $Y2=0
cc_510 N_Y_M1028_s N_VGND_c_943_n 0.00297142f $X=2.895 $Y=0.235 $X2=0 $Y2=0
cc_511 N_Y_M1005_s N_VGND_c_943_n 0.00381696f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_512 N_Y_M1021_s N_VGND_c_943_n 0.00310609f $X=5.37 $Y=0.235 $X2=0 $Y2=0
cc_513 N_Y_M1004_s N_VGND_c_943_n 0.00304199f $X=6.315 $Y=0.235 $X2=0 $Y2=0
cc_514 N_Y_M1022_s N_VGND_c_943_n 0.00378113f $X=7.255 $Y=0.235 $X2=0 $Y2=0
cc_515 N_Y_c_787_n N_VGND_c_943_n 0.00981342f $X=4.275 $Y=0.78 $X2=0 $Y2=0
cc_516 N_Y_c_801_n N_VGND_c_943_n 0.0132461f $X=5.425 $Y=0.74 $X2=0 $Y2=0
cc_517 N_Y_c_882_p N_VGND_c_943_n 0.0064465f $X=5.51 $Y=0.42 $X2=0 $Y2=0
cc_518 N_Y_c_834_n N_VGND_c_943_n 0.0128042f $X=6.365 $Y=0.745 $X2=0 $Y2=0
cc_519 N_Y_c_884_p N_VGND_c_943_n 0.00645162f $X=6.45 $Y=0.42 $X2=0 $Y2=0
cc_520 N_Y_c_812_n N_VGND_c_943_n 0.00734441f $X=6.93 $Y=0.74 $X2=0 $Y2=0
cc_521 N_Y_c_782_n N_VGND_c_943_n 0.0203112f $X=7.905 $Y=0.72 $X2=0 $Y2=0
cc_522 N_Y_c_791_n N_VGND_c_943_n 0.0139995f $X=4.51 $Y=0.42 $X2=0 $Y2=0
cc_523 N_Y_c_786_n N_A_119_47#_M1025_d 0.00401123f $X=3.585 $Y=0.77 $X2=0 $Y2=0
cc_524 N_Y_c_786_n N_A_119_47#_M1030_d 0.00335846f $X=3.585 $Y=0.77 $X2=0 $Y2=0
cc_525 N_Y_c_789_n N_A_119_47#_M1030_d 0.00190753f $X=3.68 $Y=0.77 $X2=0 $Y2=0
cc_526 N_Y_M1012_s N_A_119_47#_c_1063_n 0.00401967f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_527 N_Y_M1028_s N_A_119_47#_c_1063_n 0.00511433f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_528 N_Y_c_786_n N_A_119_47#_c_1063_n 0.0950953f $X=3.585 $Y=0.77 $X2=0 $Y2=0
cc_529 N_VGND_c_943_n N_A_119_47#_M1003_s 0.00417445f $X=8.05 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_530 N_VGND_c_943_n N_A_119_47#_M1020_s 0.00215206f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_943_n N_A_119_47#_M1025_d 0.00255381f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_943_n N_A_119_47#_M1030_d 0.00263978f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_M1011_d N_A_119_47#_c_1052_n 0.00434543f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_VGND_c_926_n N_A_119_47#_c_1052_n 0.0171911f $X=1.2 $Y=0.36 $X2=0 $Y2=0
cc_535 N_VGND_c_931_n N_A_119_47#_c_1052_n 0.00212526f $X=3.935 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_939_n N_A_119_47#_c_1052_n 0.00218565f $X=1 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_943_n N_A_119_47#_c_1052_n 0.00968351f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_538 N_VGND_c_926_n N_A_119_47#_c_1058_n 0.0203829f $X=1.2 $Y=0.36 $X2=0 $Y2=0
cc_539 N_VGND_c_931_n N_A_119_47#_c_1058_n 0.0185333f $X=3.935 $Y=0 $X2=0 $Y2=0
cc_540 N_VGND_c_943_n N_A_119_47#_c_1058_n 0.0110827f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_541 N_VGND_c_926_n N_A_119_47#_c_1059_n 0.00148728f $X=1.2 $Y=0.36 $X2=0
+ $Y2=0
cc_542 N_VGND_c_931_n N_A_119_47#_c_1063_n 0.111767f $X=3.935 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_943_n N_A_119_47#_c_1063_n 0.0705956f $X=8.05 $Y=0 $X2=0 $Y2=0
cc_544 N_VGND_c_939_n N_A_119_47#_c_1061_n 0.00451429f $X=1 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_943_n N_A_119_47#_c_1061_n 0.00655826f $X=8.05 $Y=0 $X2=0 $Y2=0
