* File: sky130_fd_sc_hdll__nor4_8.pex.spice
* Created: Thu Aug 27 19:17:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 70 71
r145 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r146 69 71 17.0272 $w=3.68e-07 $l=1.3e-07 $layer=POLY_cond $X=3.63 $Y=1.202
+ $X2=3.76 $Y2=1.202
r147 69 70 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r148 67 69 37.9837 $w=3.68e-07 $l=2.9e-07 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.63 $Y2=1.202
r149 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.34 $Y2=1.202
r150 65 66 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.315 $Y2=1.202
r151 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r152 63 64 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=2.4 $Y=1.202
+ $X2=2.82 $Y2=1.202
r153 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r154 61 62 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=2.375 $Y2=1.202
r155 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r156 59 60 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.88 $Y2=1.202
r157 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r158 57 58 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.435 $Y2=1.202
r159 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r160 54 56 48.462 $w=3.68e-07 $l=3.7e-07 $layer=POLY_cond $X=0.57 $Y=1.202
+ $X2=0.94 $Y2=1.202
r161 54 55 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=0.57
+ $Y=1.16 $X2=0.57 $Y2=1.16
r162 52 54 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.57 $Y2=1.202
r163 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r164 49 70 82.3896 $w=2.08e-07 $l=1.56e-06 $layer=LI1_cond $X=2.07 $Y=1.18
+ $X2=3.63 $Y2=1.18
r165 49 55 79.2208 $w=2.08e-07 $l=1.5e-06 $layer=LI1_cond $X=2.07 $Y=1.18
+ $X2=0.57 $Y2=1.18
r166 46 72 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r167 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r168 43 71 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r169 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.56
r170 40 67 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r171 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r172 37 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r173 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r174 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r175 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r176 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r177 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r178 28 63 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=1.202
r179 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=0.56
r180 25 62 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r181 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r182 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r183 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r184 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r185 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.56
r186 16 59 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r187 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r188 13 58 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r189 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r190 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r191 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r192 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r193 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r194 4 52 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r195 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r196 1 51 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r197 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 70 71
r146 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.52 $Y=1.202
+ $X2=7.545 $Y2=1.202
r147 69 71 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=7.47 $Y=1.202
+ $X2=7.52 $Y2=1.202
r148 69 70 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=7.47
+ $Y=1.16 $X2=7.47 $Y2=1.16
r149 67 69 48.462 $w=3.68e-07 $l=3.7e-07 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.47 $Y2=1.202
r150 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.075 $Y=1.202
+ $X2=7.1 $Y2=1.202
r151 65 66 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=6.605 $Y=1.202
+ $X2=7.075 $Y2=1.202
r152 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.202
+ $X2=6.605 $Y2=1.202
r153 63 64 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.58 $Y2=1.202
r154 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.135 $Y=1.202
+ $X2=6.16 $Y2=1.202
r155 61 62 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=6.135 $Y2=1.202
r156 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.202
+ $X2=5.665 $Y2=1.202
r157 59 60 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.64 $Y2=1.202
r158 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.22 $Y2=1.202
r159 57 58 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=5.195 $Y2=1.202
r160 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.202
+ $X2=4.725 $Y2=1.202
r161 54 56 37.9837 $w=3.68e-07 $l=2.9e-07 $layer=POLY_cond $X=4.41 $Y=1.202
+ $X2=4.7 $Y2=1.202
r162 54 55 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=4.41
+ $Y=1.16 $X2=4.41 $Y2=1.16
r163 52 54 17.0272 $w=3.68e-07 $l=1.3e-07 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.41 $Y2=1.202
r164 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.28 $Y2=1.202
r165 49 70 90.8398 $w=2.08e-07 $l=1.72e-06 $layer=LI1_cond $X=5.75 $Y=1.18
+ $X2=7.47 $Y2=1.18
r166 49 55 70.7706 $w=2.08e-07 $l=1.34e-06 $layer=LI1_cond $X=5.75 $Y=1.18
+ $X2=4.41 $Y2=1.18
r167 46 72 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.202
r168 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r169 43 71 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.52 $Y=0.995
+ $X2=7.52 $Y2=1.202
r170 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.52 $Y=0.995
+ $X2=7.52 $Y2=0.56
r171 40 67 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r172 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r173 37 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.202
r174 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r175 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.202
r176 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r177 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=1.202
r178 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=0.56
r179 28 63 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r180 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r181 25 62 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.202
r182 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r183 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r184 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r185 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.64 $Y=0.995
+ $X2=5.64 $Y2=1.202
r186 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.64 $Y=0.995
+ $X2=5.64 $Y2=0.56
r187 16 59 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r188 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r189 13 58 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r190 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r191 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r192 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r193 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=1.202
r194 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.7 $Y=0.995 $X2=4.7
+ $Y2=0.56
r195 4 52 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r196 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r197 1 51 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r198 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%C 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 70 71
r149 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=11.8 $Y=1.202
+ $X2=11.825 $Y2=1.202
r150 69 71 17.0272 $w=3.68e-07 $l=1.3e-07 $layer=POLY_cond $X=11.67 $Y=1.202
+ $X2=11.8 $Y2=1.202
r151 69 70 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=11.67
+ $Y=1.16 $X2=11.67 $Y2=1.16
r152 67 69 37.9837 $w=3.68e-07 $l=2.9e-07 $layer=POLY_cond $X=11.38 $Y=1.202
+ $X2=11.67 $Y2=1.202
r153 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=11.355 $Y=1.202
+ $X2=11.38 $Y2=1.202
r154 65 66 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=10.885 $Y=1.202
+ $X2=11.355 $Y2=1.202
r155 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=10.86 $Y=1.202
+ $X2=10.885 $Y2=1.202
r156 63 64 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=10.44 $Y=1.202
+ $X2=10.86 $Y2=1.202
r157 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=10.415 $Y=1.202
+ $X2=10.44 $Y2=1.202
r158 61 62 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=9.945 $Y=1.202
+ $X2=10.415 $Y2=1.202
r159 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=9.92 $Y=1.202
+ $X2=9.945 $Y2=1.202
r160 59 60 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=9.5 $Y=1.202
+ $X2=9.92 $Y2=1.202
r161 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=9.475 $Y=1.202
+ $X2=9.5 $Y2=1.202
r162 57 58 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=9.005 $Y=1.202
+ $X2=9.475 $Y2=1.202
r163 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.98 $Y=1.202
+ $X2=9.005 $Y2=1.202
r164 54 56 48.462 $w=3.68e-07 $l=3.7e-07 $layer=POLY_cond $X=8.61 $Y=1.202
+ $X2=8.98 $Y2=1.202
r165 54 55 29.056 $w=1.7e-07 $l=8.5e-07 $layer=licon1_POLY $count=5 $X=8.61
+ $Y=1.16 $X2=8.61 $Y2=1.16
r166 52 54 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=8.56 $Y=1.202
+ $X2=8.61 $Y2=1.202
r167 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.535 $Y=1.202
+ $X2=8.56 $Y2=1.202
r168 49 70 69.7143 $w=2.08e-07 $l=1.32e-06 $layer=LI1_cond $X=10.35 $Y=1.18
+ $X2=11.67 $Y2=1.18
r169 49 55 91.8961 $w=2.08e-07 $l=1.74e-06 $layer=LI1_cond $X=10.35 $Y=1.18
+ $X2=8.61 $Y2=1.18
r170 46 72 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.825 $Y=1.41
+ $X2=11.825 $Y2=1.202
r171 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.825 $Y=1.41
+ $X2=11.825 $Y2=1.985
r172 43 71 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.8 $Y=0.995
+ $X2=11.8 $Y2=1.202
r173 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.8 $Y=0.995
+ $X2=11.8 $Y2=0.56
r174 40 67 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.38 $Y=0.995
+ $X2=11.38 $Y2=1.202
r175 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.38 $Y=0.995
+ $X2=11.38 $Y2=0.56
r176 37 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.355 $Y=1.41
+ $X2=11.355 $Y2=1.202
r177 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.355 $Y=1.41
+ $X2=11.355 $Y2=1.985
r178 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.885 $Y=1.41
+ $X2=10.885 $Y2=1.202
r179 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.885 $Y=1.41
+ $X2=10.885 $Y2=1.985
r180 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.86 $Y=0.995
+ $X2=10.86 $Y2=1.202
r181 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.86 $Y=0.995
+ $X2=10.86 $Y2=0.56
r182 28 63 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.44 $Y=0.995
+ $X2=10.44 $Y2=1.202
r183 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.44 $Y=0.995
+ $X2=10.44 $Y2=0.56
r184 25 62 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.415 $Y=1.41
+ $X2=10.415 $Y2=1.202
r185 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.415 $Y=1.41
+ $X2=10.415 $Y2=1.985
r186 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.202
r187 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.945 $Y=1.41
+ $X2=9.945 $Y2=1.985
r188 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.92 $Y=0.995
+ $X2=9.92 $Y2=1.202
r189 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.92 $Y=0.995
+ $X2=9.92 $Y2=0.56
r190 16 59 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=1.202
r191 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=0.56
r192 13 58 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.202
r193 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.475 $Y=1.41
+ $X2=9.475 $Y2=1.985
r194 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.202
r195 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.005 $Y=1.41
+ $X2=9.005 $Y2=1.985
r196 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.98 $Y=0.995
+ $X2=8.98 $Y2=1.202
r197 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.98 $Y=0.995
+ $X2=8.98 $Y2=0.56
r198 4 52 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=1.202
r199 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=0.56
r200 1 51 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.202
r201 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.535 $Y=1.41
+ $X2=8.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%D 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 70 71
r140 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=15.56 $Y=1.202
+ $X2=15.585 $Y2=1.202
r141 69 71 48.462 $w=3.68e-07 $l=3.7e-07 $layer=POLY_cond $X=15.19 $Y=1.202
+ $X2=15.56 $Y2=1.202
r142 69 70 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=15.19
+ $Y=1.16 $X2=15.19 $Y2=1.16
r143 67 69 6.54891 $w=3.68e-07 $l=5e-08 $layer=POLY_cond $X=15.14 $Y=1.202
+ $X2=15.19 $Y2=1.202
r144 66 67 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=15.115 $Y=1.202
+ $X2=15.14 $Y2=1.202
r145 65 66 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=14.645 $Y=1.202
+ $X2=15.115 $Y2=1.202
r146 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=14.62 $Y=1.202
+ $X2=14.645 $Y2=1.202
r147 63 64 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=14.2 $Y=1.202
+ $X2=14.62 $Y2=1.202
r148 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=14.175 $Y=1.202
+ $X2=14.2 $Y2=1.202
r149 61 62 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=13.705 $Y=1.202
+ $X2=14.175 $Y2=1.202
r150 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=13.68 $Y=1.202
+ $X2=13.705 $Y2=1.202
r151 59 60 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=13.26 $Y=1.202
+ $X2=13.68 $Y2=1.202
r152 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=13.235 $Y=1.202
+ $X2=13.26 $Y2=1.202
r153 56 58 11.1332 $w=3.68e-07 $l=8.5e-08 $layer=POLY_cond $X=13.15 $Y=1.202
+ $X2=13.235 $Y2=1.202
r154 56 57 41.5086 $w=1.7e-07 $l=5.95e-07 $layer=licon1_POLY $count=3 $X=13.15
+ $Y=1.16 $X2=13.15 $Y2=1.16
r155 54 56 50.4266 $w=3.68e-07 $l=3.85e-07 $layer=POLY_cond $X=12.765 $Y=1.202
+ $X2=13.15 $Y2=1.202
r156 53 54 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=12.74 $Y=1.202
+ $X2=12.765 $Y2=1.202
r157 52 53 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=12.32 $Y=1.202
+ $X2=12.74 $Y2=1.202
r158 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=12.295 $Y=1.202
+ $X2=12.32 $Y2=1.202
r159 49 70 36.9697 $w=2.08e-07 $l=7e-07 $layer=LI1_cond $X=14.49 $Y=1.18
+ $X2=15.19 $Y2=1.18
r160 49 57 70.7706 $w=2.08e-07 $l=1.34e-06 $layer=LI1_cond $X=14.49 $Y=1.18
+ $X2=13.15 $Y2=1.18
r161 46 72 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.585 $Y=1.41
+ $X2=15.585 $Y2=1.202
r162 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.585 $Y=1.41
+ $X2=15.585 $Y2=1.985
r163 43 71 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.56 $Y=0.995
+ $X2=15.56 $Y2=1.202
r164 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.56 $Y=0.995
+ $X2=15.56 $Y2=0.56
r165 40 67 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.14 $Y=0.995
+ $X2=15.14 $Y2=1.202
r166 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.14 $Y=0.995
+ $X2=15.14 $Y2=0.56
r167 37 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.115 $Y=1.41
+ $X2=15.115 $Y2=1.202
r168 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.115 $Y=1.41
+ $X2=15.115 $Y2=1.985
r169 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.645 $Y=1.41
+ $X2=14.645 $Y2=1.202
r170 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.645 $Y=1.41
+ $X2=14.645 $Y2=1.985
r171 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.62 $Y=0.995
+ $X2=14.62 $Y2=1.202
r172 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.62 $Y=0.995
+ $X2=14.62 $Y2=0.56
r173 28 63 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.2 $Y=0.995
+ $X2=14.2 $Y2=1.202
r174 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.2 $Y=0.995
+ $X2=14.2 $Y2=0.56
r175 25 62 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.175 $Y=1.41
+ $X2=14.175 $Y2=1.202
r176 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.175 $Y=1.41
+ $X2=14.175 $Y2=1.985
r177 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.705 $Y=1.41
+ $X2=13.705 $Y2=1.202
r178 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.705 $Y=1.41
+ $X2=13.705 $Y2=1.985
r179 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.68 $Y=0.995
+ $X2=13.68 $Y2=1.202
r180 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.68 $Y=0.995
+ $X2=13.68 $Y2=0.56
r181 16 59 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.26 $Y=0.995
+ $X2=13.26 $Y2=1.202
r182 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.26 $Y=0.995
+ $X2=13.26 $Y2=0.56
r183 13 58 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.235 $Y=1.41
+ $X2=13.235 $Y2=1.202
r184 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.235 $Y=1.41
+ $X2=13.235 $Y2=1.985
r185 10 54 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.765 $Y=1.41
+ $X2=12.765 $Y2=1.202
r186 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.765 $Y=1.41
+ $X2=12.765 $Y2=1.985
r187 7 53 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.74 $Y=0.995
+ $X2=12.74 $Y2=1.202
r188 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.74 $Y=0.995
+ $X2=12.74 $Y2=0.56
r189 4 52 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.32 $Y=0.995
+ $X2=12.32 $Y2=1.202
r190 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.32 $Y=0.995
+ $X2=12.32 $Y2=0.56
r191 1 51 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.295 $Y=1.41
+ $X2=12.295 $Y2=1.202
r192 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.295 $Y=1.41
+ $X2=12.295 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%A_27_297# 1 2 3 4 5 6 7 8 9 30 34 35 38 40
+ 44 46 50 52 54 55 56 60 62 66 68 72 74 78 81 83 85 90 91 92
r118 76 78 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=7.8 $Y=2.295
+ $X2=7.8 $Y2=1.96
r119 75 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.965 $Y=2.38
+ $X2=6.84 $Y2=2.38
r120 74 76 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=7.655 $Y=2.38
+ $X2=7.8 $Y2=2.295
r121 74 75 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.655 $Y=2.38
+ $X2=6.965 $Y2=2.38
r122 70 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.295
+ $X2=6.84 $Y2=2.38
r123 70 72 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.84 $Y=2.295
+ $X2=6.84 $Y2=1.96
r124 69 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.025 $Y=2.38
+ $X2=5.9 $Y2=2.38
r125 68 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.715 $Y=2.38
+ $X2=6.84 $Y2=2.38
r126 68 69 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.715 $Y=2.38
+ $X2=6.025 $Y2=2.38
r127 64 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.295
+ $X2=5.9 $Y2=2.38
r128 64 66 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.9 $Y=2.295
+ $X2=5.9 $Y2=1.96
r129 63 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.085 $Y=2.38
+ $X2=4.96 $Y2=2.38
r130 62 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.9 $Y2=2.38
r131 62 63 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.775 $Y=2.38
+ $X2=5.085 $Y2=2.38
r132 58 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.295
+ $X2=4.96 $Y2=2.38
r133 58 60 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.96 $Y=2.295
+ $X2=4.96 $Y2=1.96
r134 57 89 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.145 $Y=2.38
+ $X2=4.02 $Y2=2.38
r135 56 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.835 $Y=2.38
+ $X2=4.96 $Y2=2.38
r136 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.835 $Y=2.38
+ $X2=4.145 $Y2=2.38
r137 55 89 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.295
+ $X2=4.02 $Y2=2.38
r138 54 87 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=1.625
+ $X2=4.02 $Y2=1.54
r139 54 55 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=4.02 $Y=1.625
+ $X2=4.02 $Y2=2.295
r140 53 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.205 $Y=1.54
+ $X2=3.08 $Y2=1.54
r141 52 87 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.895 $Y=1.54
+ $X2=4.02 $Y2=1.54
r142 52 53 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.895 $Y=1.54
+ $X2=3.205 $Y2=1.54
r143 48 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.625
+ $X2=3.08 $Y2=1.54
r144 48 50 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.08 $Y=1.625
+ $X2=3.08 $Y2=2.3
r145 47 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=1.54
+ $X2=2.14 $Y2=1.54
r146 46 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.955 $Y=1.54
+ $X2=3.08 $Y2=1.54
r147 46 47 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.955 $Y=1.54
+ $X2=2.265 $Y2=1.54
r148 42 83 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=1.54
r149 42 44 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.14 $Y=1.625
+ $X2=2.14 $Y2=2.3
r150 41 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.54
+ $X2=1.2 $Y2=1.54
r151 40 83 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=1.54
+ $X2=2.14 $Y2=1.54
r152 40 41 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.015 $Y=1.54
+ $X2=1.325 $Y2=1.54
r153 36 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.625
+ $X2=1.2 $Y2=1.54
r154 36 38 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.2 $Y=1.625
+ $X2=1.2 $Y2=2.3
r155 34 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=1.2 $Y2=1.54
r156 34 35 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=1.075 $Y=1.54
+ $X2=0.425 $Y2=1.54
r157 30 32 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r158 28 35 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.425 $Y2=1.54
r159 28 30 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.63
r160 9 78 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=1.96
r161 8 72 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=1.96
r162 7 66 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.96
r163 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.96
r164 5 89 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.3
r165 5 87 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.62
r166 4 85 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.62
r167 4 50 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.3
r168 3 83 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.62
r169 3 44 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.3
r170 2 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.62
r171 2 38 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.3
r172 1 32 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r173 1 30 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%VPWR 1 2 3 4 15 17 21 23 27 29 33 35 37 47
+ 48 51 54 57 60 65
r183 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r184 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r185 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r186 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r187 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r188 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r189 52 65 0.125198 $w=4.8e-07 $l=4.4e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.25 $Y2=2.72
r190 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r191 47 48 0.688889 $w=1.7e-07 $l=2.295e-06 $layer=mcon $count=13 $X=15.87
+ $Y=2.72 $X2=15.87 $Y2=2.72
r192 45 48 3.40312 $w=4.8e-07 $l=1.196e-05 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=15.87 $Y2=2.72
r193 45 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r194 44 47 780.278 $w=1.68e-07 $l=1.196e-05 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=15.87 $Y2=2.72
r195 44 45 0.688889 $w=1.7e-07 $l=2.295e-06 $layer=mcon $count=13 $X=3.91
+ $Y=2.72 $X2=3.91 $Y2=2.72
r196 42 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.55 $Y2=2.72
r197 42 44 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=3.675 $Y=2.72
+ $X2=3.91 $Y2=2.72
r198 37 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.73 $Y2=2.72
r199 37 39 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r200 35 65 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.25 $Y2=2.72
r201 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r202 31 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r203 31 33 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=1.96
r204 30 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=2.61 $Y2=2.72
r205 29 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=3.55 $Y2=2.72
r206 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.425 $Y=2.72
+ $X2=2.735 $Y2=2.72
r207 25 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.72
r208 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=1.96
r209 24 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.795 $Y=2.72
+ $X2=1.67 $Y2=2.72
r210 23 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.61 $Y2=2.72
r211 23 24 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=1.795 $Y2=2.72
r212 19 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r213 19 21 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=1.96
r214 18 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.73 $Y2=2.72
r215 17 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=1.67 $Y2=2.72
r216 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.72
+ $X2=0.855 $Y2=2.72
r217 13 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r218 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=1.96
r219 4 33 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.96
r220 3 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r221 2 21 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r222 1 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%A_869_297# 1 2 3 4 5 6 7 8 27 31 35 39 43
+ 47 51 56 58 60 62 64 66 68 70
r120 52 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.775 $Y=1.54
+ $X2=10.65 $Y2=1.54
r121 51 70 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.465 $Y=1.54
+ $X2=11.59 $Y2=1.54
r122 51 52 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.465 $Y=1.54
+ $X2=10.775 $Y2=1.54
r123 48 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.835 $Y=1.54
+ $X2=9.71 $Y2=1.54
r124 47 68 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.525 $Y=1.54
+ $X2=10.65 $Y2=1.54
r125 47 48 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.525 $Y=1.54
+ $X2=9.835 $Y2=1.54
r126 44 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.895 $Y=1.54
+ $X2=8.77 $Y2=1.54
r127 43 66 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.585 $Y=1.54
+ $X2=9.71 $Y2=1.54
r128 43 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.585 $Y=1.54
+ $X2=8.895 $Y2=1.54
r129 40 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.435 $Y=1.54
+ $X2=7.31 $Y2=1.54
r130 39 64 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.645 $Y=1.54
+ $X2=8.77 $Y2=1.54
r131 39 40 78.9412 $w=1.68e-07 $l=1.21e-06 $layer=LI1_cond $X=8.645 $Y=1.54
+ $X2=7.435 $Y2=1.54
r132 36 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.495 $Y=1.54
+ $X2=6.37 $Y2=1.54
r133 35 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.185 $Y=1.54
+ $X2=7.31 $Y2=1.54
r134 35 36 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.185 $Y=1.54
+ $X2=6.495 $Y2=1.54
r135 32 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.555 $Y=1.54
+ $X2=5.43 $Y2=1.54
r136 31 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.245 $Y=1.54
+ $X2=6.37 $Y2=1.54
r137 31 32 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.245 $Y=1.54
+ $X2=5.555 $Y2=1.54
r138 28 56 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.615 $Y=1.54
+ $X2=4.49 $Y2=1.54
r139 27 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.305 $Y=1.54
+ $X2=5.43 $Y2=1.54
r140 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.305 $Y=1.54
+ $X2=4.615 $Y2=1.54
r141 8 70 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=11.445
+ $Y=1.485 $X2=11.59 $Y2=1.62
r142 7 68 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=10.505
+ $Y=1.485 $X2=10.65 $Y2=1.62
r143 6 66 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=9.565
+ $Y=1.485 $X2=9.71 $Y2=1.62
r144 5 64 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.625
+ $Y=1.485 $X2=8.77 $Y2=1.62
r145 4 62 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.62
r146 3 60 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.62
r147 2 58 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.62
r148 1 56 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%A_1635_297# 1 2 3 4 5 6 7 8 9 30 32 33 36
+ 38 42 44 48 50 54 56 60 62 66 68 72 74 76 78 80 81 82 84 85 86 87
r120 76 89 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.845 $Y=2.295
+ $X2=15.845 $Y2=2.38
r121 76 78 25.5458 $w=2.98e-07 $l=6.65e-07 $layer=LI1_cond $X=15.845 $Y=2.295
+ $X2=15.845 $Y2=1.63
r122 75 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.005 $Y=2.38
+ $X2=14.88 $Y2=2.38
r123 74 89 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=15.695 $Y=2.38
+ $X2=15.845 $Y2=2.38
r124 74 75 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.695 $Y=2.38
+ $X2=15.005 $Y2=2.38
r125 70 87 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=14.88 $Y=2.295
+ $X2=14.88 $Y2=2.38
r126 70 72 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=14.88 $Y=2.295
+ $X2=14.88 $Y2=1.96
r127 69 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.065 $Y=2.38
+ $X2=13.94 $Y2=2.38
r128 68 87 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.755 $Y=2.38
+ $X2=14.88 $Y2=2.38
r129 68 69 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.755 $Y=2.38
+ $X2=14.065 $Y2=2.38
r130 64 86 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13.94 $Y=2.295
+ $X2=13.94 $Y2=2.38
r131 64 66 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=13.94 $Y=2.295
+ $X2=13.94 $Y2=1.96
r132 63 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.125 $Y=2.38
+ $X2=13 $Y2=2.38
r133 62 86 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.815 $Y=2.38
+ $X2=13.94 $Y2=2.38
r134 62 63 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=13.815 $Y=2.38
+ $X2=13.125 $Y2=2.38
r135 58 85 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=13 $Y=2.295
+ $X2=13 $Y2=2.38
r136 58 60 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=13 $Y=2.295 $X2=13
+ $Y2=1.96
r137 57 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.185 $Y=2.38
+ $X2=12.06 $Y2=2.38
r138 56 85 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=12.875 $Y=2.38
+ $X2=13 $Y2=2.38
r139 56 57 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=12.875 $Y=2.38
+ $X2=12.185 $Y2=2.38
r140 52 84 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=12.06 $Y=2.295
+ $X2=12.06 $Y2=2.38
r141 52 54 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=12.06 $Y=2.295
+ $X2=12.06 $Y2=1.62
r142 51 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.245 $Y=2.38
+ $X2=11.12 $Y2=2.38
r143 50 84 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.935 $Y=2.38
+ $X2=12.06 $Y2=2.38
r144 50 51 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=11.935 $Y=2.38
+ $X2=11.245 $Y2=2.38
r145 46 82 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.12 $Y=2.295
+ $X2=11.12 $Y2=2.38
r146 46 48 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=11.12 $Y=2.295
+ $X2=11.12 $Y2=1.96
r147 45 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.305 $Y=2.38
+ $X2=10.18 $Y2=2.38
r148 44 82 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.995 $Y=2.38
+ $X2=11.12 $Y2=2.38
r149 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.995 $Y=2.38
+ $X2=10.305 $Y2=2.38
r150 40 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=2.295
+ $X2=10.18 $Y2=2.38
r151 40 42 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=10.18 $Y=2.295
+ $X2=10.18 $Y2=1.96
r152 39 80 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.365 $Y=2.38
+ $X2=9.22 $Y2=2.38
r153 38 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.055 $Y=2.38
+ $X2=10.18 $Y2=2.38
r154 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.055 $Y=2.38
+ $X2=9.365 $Y2=2.38
r155 34 80 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=2.295
+ $X2=9.22 $Y2=2.38
r156 34 36 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=9.22 $Y=2.295
+ $X2=9.22 $Y2=1.96
r157 32 80 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=9.075 $Y=2.38
+ $X2=9.22 $Y2=2.38
r158 32 33 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=9.075 $Y=2.38
+ $X2=8.425 $Y2=2.38
r159 28 33 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.28 $Y=2.295
+ $X2=8.425 $Y2=2.38
r160 28 30 13.3127 $w=2.88e-07 $l=3.35e-07 $layer=LI1_cond $X=8.28 $Y=2.295
+ $X2=8.28 $Y2=1.96
r161 9 89 400 $w=1.7e-07 $l=8.99166e-07 $layer=licon1_PDIFF $count=1 $X=15.675
+ $Y=1.485 $X2=15.83 $Y2=2.31
r162 9 78 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=15.675
+ $Y=1.485 $X2=15.83 $Y2=1.63
r163 8 72 300 $w=1.7e-07 $l=5.47037e-07 $layer=licon1_PDIFF $count=2 $X=14.735
+ $Y=1.485 $X2=14.89 $Y2=1.96
r164 7 66 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=13.795
+ $Y=1.485 $X2=13.94 $Y2=1.96
r165 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=12.855
+ $Y=1.485 $X2=13 $Y2=1.96
r166 5 84 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=11.915
+ $Y=1.485 $X2=12.06 $Y2=2.3
r167 5 54 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=11.915
+ $Y=1.485 $X2=12.06 $Y2=1.62
r168 4 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.975
+ $Y=1.485 $X2=11.12 $Y2=1.96
r169 3 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.035
+ $Y=1.485 $X2=10.18 $Y2=1.96
r170 2 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.095
+ $Y=1.485 $X2=9.24 $Y2=1.96
r171 1 30 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=8.175
+ $Y=1.485 $X2=8.3 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17
+ 18 19 20 63 65 66 69 71 75 77 81 83 87 89 93 95 99 101 105 107 111 113 117 119
+ 123 125 129 131 135 139 141 145 149 151 155 159 161 165 169 170 171 172 173
+ 174 175 176 177 178 179 181 184 185 187 188 190 192 193
c408 184 0 1.85425e-19 $X=12.53 $Y=1.62
r409 182 193 7.44872 $w=4.08e-07 $l=2.65e-07 $layer=LI1_cond $X=12.61 $Y=1.455
+ $X2=12.61 $Y2=1.19
r410 182 184 2.88756 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.61 $Y=1.455
+ $X2=12.61 $Y2=1.54
r411 180 193 8.01088 $w=4.08e-07 $l=2.85e-07 $layer=LI1_cond $X=12.61 $Y=0.905
+ $X2=12.61 $Y2=1.19
r412 180 181 1.17876 $w=4.1e-07 $l=9.94987e-08 $layer=LI1_cond $X=12.61 $Y=0.905
+ $X2=12.59 $Y2=0.815
r413 163 165 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.35 $Y=0.725
+ $X2=15.35 $Y2=0.39
r414 162 188 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.575 $Y=0.815
+ $X2=14.41 $Y2=0.815
r415 161 163 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=15.185
+ $Y=0.815 $X2=15.35 $Y2=0.725
r416 161 162 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=15.185 $Y=0.815
+ $X2=14.575 $Y2=0.815
r417 160 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.535 $Y=1.54
+ $X2=14.41 $Y2=1.54
r418 159 192 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.225 $Y=1.54
+ $X2=15.35 $Y2=1.54
r419 159 160 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=15.225 $Y=1.54
+ $X2=14.535 $Y2=1.54
r420 153 188 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.41 $Y=0.725
+ $X2=14.41 $Y2=0.815
r421 153 155 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.41 $Y=0.725
+ $X2=14.41 $Y2=0.39
r422 152 185 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.635 $Y=0.815
+ $X2=13.47 $Y2=0.815
r423 151 188 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.245 $Y=0.815
+ $X2=14.41 $Y2=0.815
r424 151 152 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=14.245 $Y=0.815
+ $X2=13.635 $Y2=0.815
r425 150 187 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.595 $Y=1.54
+ $X2=13.47 $Y2=1.54
r426 149 190 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=14.285 $Y=1.54
+ $X2=14.41 $Y2=1.54
r427 149 150 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=14.285 $Y=1.54
+ $X2=13.595 $Y2=1.54
r428 143 185 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=13.47 $Y=0.725
+ $X2=13.47 $Y2=0.815
r429 143 145 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.47 $Y=0.725
+ $X2=13.47 $Y2=0.39
r430 142 184 3.80956 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=12.815 $Y=1.54
+ $X2=12.61 $Y2=1.54
r431 141 187 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=13.345 $Y=1.54
+ $X2=13.47 $Y2=1.54
r432 141 142 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.345 $Y=1.54
+ $X2=12.815 $Y2=1.54
r433 140 181 5.47904 $w=1.8e-07 $l=2.25e-07 $layer=LI1_cond $X=12.815 $Y=0.815
+ $X2=12.59 $Y2=0.815
r434 139 185 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.305 $Y=0.815
+ $X2=13.47 $Y2=0.815
r435 139 140 30.1919 $w=1.78e-07 $l=4.9e-07 $layer=LI1_cond $X=13.305 $Y=0.815
+ $X2=12.815 $Y2=0.815
r436 133 181 1.17876 $w=3.3e-07 $l=1.16189e-07 $layer=LI1_cond $X=12.53 $Y=0.725
+ $X2=12.59 $Y2=0.815
r437 133 135 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.53 $Y=0.725
+ $X2=12.53 $Y2=0.39
r438 132 179 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.755 $Y=0.815
+ $X2=11.59 $Y2=0.815
r439 131 181 5.47904 $w=1.8e-07 $l=2.25e-07 $layer=LI1_cond $X=12.365 $Y=0.815
+ $X2=12.59 $Y2=0.815
r440 131 132 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=12.365 $Y=0.815
+ $X2=11.755 $Y2=0.815
r441 127 179 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=11.59 $Y=0.725
+ $X2=11.59 $Y2=0.815
r442 127 129 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=11.59 $Y=0.725
+ $X2=11.59 $Y2=0.39
r443 126 178 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.815 $Y=0.815
+ $X2=10.65 $Y2=0.815
r444 125 179 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.425 $Y=0.815
+ $X2=11.59 $Y2=0.815
r445 125 126 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=11.425 $Y=0.815
+ $X2=10.815 $Y2=0.815
r446 121 178 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=10.65 $Y=0.725
+ $X2=10.65 $Y2=0.815
r447 121 123 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.65 $Y=0.725
+ $X2=10.65 $Y2=0.39
r448 120 177 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.875 $Y=0.815
+ $X2=9.71 $Y2=0.815
r449 119 178 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=10.485 $Y=0.815
+ $X2=10.65 $Y2=0.815
r450 119 120 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=10.485 $Y=0.815
+ $X2=9.875 $Y2=0.815
r451 115 177 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=9.71 $Y=0.725
+ $X2=9.71 $Y2=0.815
r452 115 117 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.71 $Y=0.725
+ $X2=9.71 $Y2=0.39
r453 114 176 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.935 $Y=0.815
+ $X2=8.77 $Y2=0.815
r454 113 177 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=9.545 $Y=0.815
+ $X2=9.71 $Y2=0.815
r455 113 114 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=9.545 $Y=0.815
+ $X2=8.935 $Y2=0.815
r456 109 176 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=8.77 $Y=0.725
+ $X2=8.77 $Y2=0.815
r457 109 111 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=8.77 $Y=0.725
+ $X2=8.77 $Y2=0.39
r458 108 175 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=0.815
+ $X2=7.31 $Y2=0.815
r459 107 176 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=8.605 $Y=0.815
+ $X2=8.77 $Y2=0.815
r460 107 108 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=8.605 $Y=0.815
+ $X2=7.475 $Y2=0.815
r461 103 175 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=7.31 $Y=0.725
+ $X2=7.31 $Y2=0.815
r462 103 105 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.31 $Y=0.725
+ $X2=7.31 $Y2=0.39
r463 102 174 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.535 $Y=0.815
+ $X2=6.37 $Y2=0.815
r464 101 175 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=0.815
+ $X2=7.31 $Y2=0.815
r465 101 102 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=7.145 $Y=0.815
+ $X2=6.535 $Y2=0.815
r466 97 174 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.37 $Y=0.725
+ $X2=6.37 $Y2=0.815
r467 97 99 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.37 $Y=0.725
+ $X2=6.37 $Y2=0.39
r468 96 173 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=0.815
+ $X2=5.43 $Y2=0.815
r469 95 174 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.205 $Y=0.815
+ $X2=6.37 $Y2=0.815
r470 95 96 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=6.205 $Y=0.815
+ $X2=5.595 $Y2=0.815
r471 91 173 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=5.43 $Y=0.725
+ $X2=5.43 $Y2=0.815
r472 91 93 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.43 $Y=0.725
+ $X2=5.43 $Y2=0.39
r473 90 172 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=0.815
+ $X2=4.49 $Y2=0.815
r474 89 173 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=0.815
+ $X2=5.43 $Y2=0.815
r475 89 90 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=5.265 $Y=0.815
+ $X2=4.655 $Y2=0.815
r476 85 172 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=4.49 $Y=0.725
+ $X2=4.49 $Y2=0.815
r477 85 87 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.49 $Y=0.725
+ $X2=4.49 $Y2=0.39
r478 84 171 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=0.815
+ $X2=3.55 $Y2=0.815
r479 83 172 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=0.815
+ $X2=4.49 $Y2=0.815
r480 83 84 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=4.325 $Y=0.815
+ $X2=3.715 $Y2=0.815
r481 79 171 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.55 $Y=0.725
+ $X2=3.55 $Y2=0.815
r482 79 81 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.55 $Y=0.725
+ $X2=3.55 $Y2=0.39
r483 78 170 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=0.815
+ $X2=2.61 $Y2=0.815
r484 77 171 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=3.55 $Y2=0.815
r485 77 78 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=0.815
+ $X2=2.775 $Y2=0.815
r486 73 170 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.61 $Y=0.725
+ $X2=2.61 $Y2=0.815
r487 73 75 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.61 $Y=0.725
+ $X2=2.61 $Y2=0.39
r488 72 169 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=0.815
+ $X2=1.67 $Y2=0.815
r489 71 170 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=0.815
+ $X2=2.61 $Y2=0.815
r490 71 72 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=0.815
+ $X2=1.835 $Y2=0.815
r491 67 169 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=1.67 $Y=0.725
+ $X2=1.67 $Y2=0.815
r492 67 69 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=0.725
+ $X2=1.67 $Y2=0.39
r493 65 169 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=1.67 $Y2=0.815
r494 65 66 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=0.815
+ $X2=0.895 $Y2=0.815
r495 61 66 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.895 $Y2=0.815
r496 61 63 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=0.725
+ $X2=0.73 $Y2=0.39
r497 20 192 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=15.205
+ $Y=1.485 $X2=15.35 $Y2=1.62
r498 19 190 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=14.265
+ $Y=1.485 $X2=14.41 $Y2=1.62
r499 18 187 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=13.325
+ $Y=1.485 $X2=13.47 $Y2=1.62
r500 17 184 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=12.385
+ $Y=1.485 $X2=12.53 $Y2=1.62
r501 16 165 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=15.215
+ $Y=0.235 $X2=15.35 $Y2=0.39
r502 15 155 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=14.275
+ $Y=0.235 $X2=14.41 $Y2=0.39
r503 14 145 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=13.335
+ $Y=0.235 $X2=13.47 $Y2=0.39
r504 13 135 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=12.395
+ $Y=0.235 $X2=12.53 $Y2=0.39
r505 12 129 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=11.455
+ $Y=0.235 $X2=11.59 $Y2=0.39
r506 11 123 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.515
+ $Y=0.235 $X2=10.65 $Y2=0.39
r507 10 117 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=9.575
+ $Y=0.235 $X2=9.71 $Y2=0.39
r508 9 111 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.635
+ $Y=0.235 $X2=8.77 $Y2=0.39
r509 8 105 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=7.175
+ $Y=0.235 $X2=7.31 $Y2=0.39
r510 7 99 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.235
+ $Y=0.235 $X2=6.37 $Y2=0.39
r511 6 93 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.235 $X2=5.43 $Y2=0.39
r512 5 87 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.235 $X2=4.49 $Y2=0.39
r513 4 81 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.39
r514 3 75 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.39
r515 2 69 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.39
r516 1 63 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4_8%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 52 54 58 60 64 66 70 72 76 78 82 86 90 94 98 102 106 110 114 118 120 122
+ 125 126 128 129 131 132 134 135 137 138 140 141 143 144 146 147 149 150 151
+ 153 191 199 202 205 208 211 216 219 222
r274 221 222 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r275 218 219 9.8562 $w=6.38e-07 $l=1.35e-07 $layer=LI1_cond $X=8.3 $Y=0.235
+ $X2=8.435 $Y2=0.235
r276 214 218 4.67218 $w=6.38e-07 $l=2.5e-07 $layer=LI1_cond $X=8.05 $Y=0.235
+ $X2=8.3 $Y2=0.235
r277 214 216 14.9022 $w=6.38e-07 $l=4.05e-07 $layer=LI1_cond $X=8.05 $Y=0.235
+ $X2=7.645 $Y2=0.235
r278 214 215 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r279 211 212 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r280 209 212 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r281 208 209 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r282 206 209 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r283 205 206 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r284 203 206 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r285 202 203 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r286 200 203 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r287 199 200 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r288 194 222 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=15.87 $Y2=0
r289 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r290 191 221 4.24382 $w=1.7e-07 $l=2.07e-07 $layer=LI1_cond $X=15.685 $Y=0
+ $X2=15.892 $Y2=0
r291 191 193 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=15.685 $Y=0
+ $X2=15.41 $Y2=0
r292 190 194 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=15.41 $Y2=0
r293 189 190 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r294 187 190 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.49 $Y2=0
r295 186 187 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r296 184 187 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r297 183 184 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r298 181 184 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.65 $Y2=0
r299 180 181 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r300 178 181 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r301 177 178 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r302 175 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r303 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r304 172 175 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.89 $Y2=0
r305 172 215 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=8.05 $Y2=0
r306 171 219 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=8.435 $Y2=0
r307 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r308 168 215 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r309 167 216 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=7.645 $Y2=0
r310 167 168 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r311 164 168 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r312 163 164 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r313 161 164 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r314 161 212 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=4.83 $Y2=0
r315 160 161 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r316 158 211 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=4.96 $Y2=0
r317 158 160 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.095 $Y=0
+ $X2=5.75 $Y2=0
r318 157 200 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.15 $Y2=0
r319 156 157 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r320 154 196 4.06843 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.197 $Y2=0
r321 154 156 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0
+ $X2=0.69 $Y2=0
r322 153 199 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=1.2 $Y2=0
r323 153 156 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=0
+ $X2=0.69 $Y2=0
r324 151 157 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r325 151 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r326 149 189 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=14.745 $Y=0
+ $X2=14.49 $Y2=0
r327 149 150 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.745 $Y=0
+ $X2=14.88 $Y2=0
r328 148 193 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=15.015 $Y=0
+ $X2=15.41 $Y2=0
r329 148 150 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.015 $Y=0
+ $X2=14.88 $Y2=0
r330 146 186 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=13.57 $Y2=0
r331 146 147 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.805 $Y=0
+ $X2=13.94 $Y2=0
r332 145 189 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=14.075 $Y=0
+ $X2=14.49 $Y2=0
r333 145 147 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.075 $Y=0
+ $X2=13.94 $Y2=0
r334 143 183 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=12.865 $Y=0
+ $X2=12.65 $Y2=0
r335 143 144 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.865 $Y=0
+ $X2=13 $Y2=0
r336 142 186 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=13.135 $Y=0
+ $X2=13.57 $Y2=0
r337 142 144 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.135 $Y=0
+ $X2=13 $Y2=0
r338 140 180 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=11.73 $Y2=0
r339 140 141 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.925 $Y=0
+ $X2=12.06 $Y2=0
r340 139 183 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=12.195 $Y=0
+ $X2=12.65 $Y2=0
r341 139 141 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.195 $Y=0
+ $X2=12.06 $Y2=0
r342 137 177 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=10.81 $Y2=0
r343 137 138 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.985 $Y=0
+ $X2=11.12 $Y2=0
r344 136 180 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=11.255 $Y=0
+ $X2=11.73 $Y2=0
r345 136 138 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.255 $Y=0
+ $X2=11.12 $Y2=0
r346 134 174 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=9.89 $Y2=0
r347 134 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.045 $Y=0
+ $X2=10.18 $Y2=0
r348 133 177 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.81 $Y2=0
r349 133 135 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.315 $Y=0
+ $X2=10.18 $Y2=0
r350 131 171 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=9.105 $Y=0
+ $X2=8.97 $Y2=0
r351 131 132 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.105 $Y=0
+ $X2=9.24 $Y2=0
r352 130 174 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=9.375 $Y=0
+ $X2=9.89 $Y2=0
r353 130 132 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.375 $Y=0
+ $X2=9.24 $Y2=0
r354 128 163 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.67 $Y2=0
r355 128 129 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=0
+ $X2=6.84 $Y2=0
r356 127 167 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=7.59 $Y2=0
r357 127 129 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.975 $Y=0
+ $X2=6.84 $Y2=0
r358 125 160 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.765 $Y=0
+ $X2=5.75 $Y2=0
r359 125 126 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.765 $Y=0
+ $X2=5.9 $Y2=0
r360 124 163 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.035 $Y=0
+ $X2=6.67 $Y2=0
r361 124 126 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.035 $Y=0
+ $X2=5.9 $Y2=0
r362 120 221 3.11623 $w=2.8e-07 $l=1.13666e-07 $layer=LI1_cond $X=15.825
+ $Y=0.085 $X2=15.892 $Y2=0
r363 120 122 12.5534 $w=2.78e-07 $l=3.05e-07 $layer=LI1_cond $X=15.825 $Y=0.085
+ $X2=15.825 $Y2=0.39
r364 116 150 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.88 $Y=0.085
+ $X2=14.88 $Y2=0
r365 116 118 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=14.88 $Y=0.085
+ $X2=14.88 $Y2=0.39
r366 112 147 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.94 $Y=0.085
+ $X2=13.94 $Y2=0
r367 112 114 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13.94 $Y=0.085
+ $X2=13.94 $Y2=0.39
r368 108 144 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13 $Y=0.085
+ $X2=13 $Y2=0
r369 108 110 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=13 $Y=0.085
+ $X2=13 $Y2=0.39
r370 104 141 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.06 $Y=0.085
+ $X2=12.06 $Y2=0
r371 104 106 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=12.06 $Y=0.085
+ $X2=12.06 $Y2=0.39
r372 100 138 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.12 $Y=0.085
+ $X2=11.12 $Y2=0
r373 100 102 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=11.12 $Y=0.085
+ $X2=11.12 $Y2=0.39
r374 96 135 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0
r375 96 98 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.18 $Y=0.085
+ $X2=10.18 $Y2=0.39
r376 92 132 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0
r377 92 94 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.24 $Y=0.085
+ $X2=9.24 $Y2=0.39
r378 88 129 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r379 88 90 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.39
r380 84 126 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0
r381 84 86 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0.39
r382 80 211 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r383 80 82 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.39
r384 79 208 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=0
+ $X2=4.02 $Y2=0
r385 78 211 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.96 $Y2=0
r386 78 79 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.825 $Y=0
+ $X2=4.155 $Y2=0
r387 74 208 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r388 74 76 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.39
r389 73 205 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=0
+ $X2=3.08 $Y2=0
r390 72 208 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=4.02 $Y2=0
r391 72 73 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=0
+ $X2=3.215 $Y2=0
r392 68 205 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r393 68 70 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.39
r394 67 202 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=0
+ $X2=2.14 $Y2=0
r395 66 205 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=3.08 $Y2=0
r396 66 67 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=0
+ $X2=2.275 $Y2=0
r397 62 202 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r398 62 64 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.39
r399 61 199 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.2
+ $Y2=0
r400 60 202 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=2.14 $Y2=0
r401 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0
+ $X2=1.335 $Y2=0
r402 56 199 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r403 56 58 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.39
r404 52 196 3.14379 $w=2.6e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.197 $Y2=0
r405 52 54 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=0.085
+ $X2=0.265 $Y2=0.39
r406 17 122 91 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=2 $X=15.635
+ $Y=0.235 $X2=15.83 $Y2=0.39
r407 16 118 182 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=1 $X=14.695
+ $Y=0.235 $X2=14.89 $Y2=0.39
r408 15 114 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=13.755
+ $Y=0.235 $X2=13.94 $Y2=0.39
r409 14 110 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=12.815
+ $Y=0.235 $X2=13 $Y2=0.39
r410 13 106 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=11.875
+ $Y=0.235 $X2=12.06 $Y2=0.39
r411 12 102 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=10.935
+ $Y=0.235 $X2=11.12 $Y2=0.39
r412 11 98 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.995
+ $Y=0.235 $X2=10.18 $Y2=0.39
r413 10 94 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.055
+ $Y=0.235 $X2=9.24 $Y2=0.39
r414 9 218 91 $w=1.7e-07 $l=7.78653e-07 $layer=licon1_NDIFF $count=2 $X=7.595
+ $Y=0.235 $X2=8.3 $Y2=0.39
r415 8 90 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.39
r416 7 86 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.39
r417 6 82 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.39
r418 5 76 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.39
r419 4 70 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.39
r420 3 64 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.39
r421 2 58 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.39
r422 1 54 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

