* File: sky130_fd_sc_hdll__muxb16to1_1.spice
* Created: Thu Aug 27 19:11:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb16to1_1.pex.spice"
.subckt sky130_fd_sc_hdll__muxb16to1_1  VNB VPB D[0] D[8] S[0] S[8] S[1] S[9]
+ D[1] D[9] D[2] D[10] S[2] S[10] S[3] S[11] D[3] D[11] D[4] D[12] S[4] S[12]
+ S[5] S[13] D[5] D[13] D[6] D[14] S[6] S[14] S[7] S[15] D[7] D[15] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[15]	D[15]
* D[7]	D[7]
* S[15]	S[15]
* S[7]	S[7]
* S[14]	S[14]
* S[6]	S[6]
* D[14]	D[14]
* D[6]	D[6]
* D[13]	D[13]
* D[5]	D[5]
* S[13]	S[13]
* S[5]	S[5]
* S[12]	S[12]
* S[4]	S[4]
* D[12]	D[12]
* D[4]	D[4]
* D[11]	D[11]
* D[3]	D[3]
* S[11]	S[11]
* S[3]	S[3]
* S[10]	S[10]
* S[2]	S[2]
* D[10]	D[10]
* D[2]	D[2]
* D[9]	D[9]
* D[1]	D[1]
* S[9]	S[9]
* S[1]	S[1]
* S[8]	S[8]
* S[0]	S[0]
* D[8]	D[8]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1086 A_109_47# N_D[0]_M1086_g N_VGND_M1086_s VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.169 PD=1.08333 PS=1.82 NRD=21.636 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1025 A_109_911# N_D[8]_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.169 PD=1.08333 PS=1.82 NRD=21.636 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1092 N_Z_M1092_d N_S[0]_M1092_g A_109_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75000.7
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1056 N_Z_M1056_d N_S[8]_M1056_g A_109_911# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75000.7
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1058 N_VGND_M1058_d N_S[0]_M1058_g N_A_184_265#_M1058_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1067 N_VGND_M1067_d N_S[8]_M1067_g N_A_184_793#_M1067_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1055 N_A_533_47#_M1055_d N_S[1]_M1055_g N_VGND_M1058_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1031 N_A_533_937#_M1031_d N_S[9]_M1031_g N_VGND_M1067_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1023 A_746_47# N_S[1]_M1023_g N_Z_M1023_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1047 A_746_937# N_S[9]_M1047_g N_Z_M1047_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1062 N_VGND_M1062_d N_D[1]_M1062_g A_746_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1057 N_VGND_M1057_d N_D[9]_M1057_g A_746_937# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1002 A_937_47# N_D[2]_M1002_g N_VGND_M1062_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1011 A_937_911# N_D[10]_M1011_g N_VGND_M1057_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1018 N_Z_M1018_d N_S[2]_M1018_g A_937_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1065 N_Z_M1065_d N_S[10]_M1065_g A_937_911# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1088 N_VGND_M1088_d N_S[2]_M1088_g N_A_1012_265#_M1088_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1082 N_VGND_M1082_d N_S[10]_M1082_g N_A_1012_793#_M1082_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1052 N_A_1361_47#_M1052_d N_S[3]_M1052_g N_VGND_M1088_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1061 N_A_1361_937#_M1061_d N_S[11]_M1061_g N_VGND_M1082_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1015 A_1574_47# N_S[3]_M1015_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1068 A_1574_937# N_S[11]_M1068_g N_Z_M1068_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1081 N_VGND_M1081_d N_D[3]_M1081_g A_1574_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1043 N_VGND_M1043_d N_D[11]_M1043_g A_1574_937# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1001 A_1765_47# N_D[4]_M1001_g N_VGND_M1081_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1037 A_1765_911# N_D[12]_M1037_g N_VGND_M1043_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1030 N_Z_M1030_d N_S[4]_M1030_g A_1765_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1069 N_Z_M1069_d N_S[12]_M1069_g A_1765_911# VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667
+ SA=75001.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1094 N_VGND_M1094_d N_S[4]_M1094_g N_A_1840_265#_M1094_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1024 N_VGND_M1024_d N_S[12]_M1024_g N_A_1840_793#_M1024_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1078 N_A_2189_47#_M1078_d N_S[5]_M1078_g N_VGND_M1094_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1070 N_A_2189_937#_M1070_d N_S[13]_M1070_g N_VGND_M1024_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1020 A_2402_47# N_S[5]_M1020_g N_Z_M1020_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1016 A_2402_937# N_S[13]_M1016_g N_Z_M1016_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1087 N_VGND_M1087_d N_D[5]_M1087_g A_2402_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1091 N_VGND_M1091_d N_D[13]_M1091_g A_2402_937# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.111944 PD=0.98 PS=1.08333 NRD=4.608 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75001 A=0.0975 P=1.6 MULT=1
MM1003 A_2593_47# N_D[6]_M1003_g N_VGND_M1087_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1083 A_2593_911# N_D[14]_M1083_g N_VGND_M1091_d VNB NSHORT L=0.15 W=0.65
+ AD=0.111944 AS=0.10725 PD=1.08333 PS=0.98 NRD=21.636 NRS=4.608 M=1 R=4.33333
+ SA=75001 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1063 N_Z_M1063_d N_S[6]_M1063_g A_2593_47# VNB NSHORT L=0.15 W=0.52 AD=0.1352
+ AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1084 N_Z_M1084_d N_S[14]_M1084_g A_2593_911# VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0895556 PD=1.56 PS=0.866667 NRD=0 NRS=27.048 M=1 R=3.46667
+ SA=75001.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1007 N_VGND_M1007_d N_S[6]_M1007_g N_A_2668_265#_M1007_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1026 N_VGND_M1026_d N_S[14]_M1026_g N_A_2668_793#_M1026_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1118 AS=0.1482 PD=0.95 PS=1.61 NRD=17.304 NRS=4.608 M=1 R=3.46667
+ SA=75000.2 SB=75000.8 A=0.078 P=1.34 MULT=1
MM1095 N_A_3017_47#_M1095_d N_S[7]_M1095_g N_VGND_M1007_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1073 N_A_3017_937#_M1073_d N_S[15]_M1073_g N_VGND_M1026_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1482 AS=0.1118 PD=1.61 PS=0.95 NRD=4.608 NRS=17.304 M=1 R=3.46667
+ SA=75000.8 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1060 A_3230_47# N_S[7]_M1060_g N_Z_M1060_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.7 A=0.078 P=1.34 MULT=1
MM1054 A_3230_937# N_S[15]_M1054_g N_Z_M1054_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0895556 AS=0.1352 PD=0.866667 PS=1.56 NRD=27.048 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.7 A=0.078 P=1.34 MULT=1
MM1089 N_VGND_M1089_d N_D[7]_M1089_g A_3230_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.111944 PD=1.82 PS=1.08333 NRD=0 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1034_d N_D[15]_M1034_g A_3230_937# VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.111944 PD=1.82 PS=1.08333 NRD=0 NRS=21.636 M=1 R=4.33333
+ SA=75000.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1027 A_117_297# N_D[0]_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.27 PD=1.47802 PS=2.54 NRD=24.8417 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1032 A_117_591# N_D[8]_M1032_g N_VPWR_M1032_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.27 PD=1.47802 PS=2.54 NRD=24.8417 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1036 N_Z_M1036_d N_A_184_265#_M1036_g A_117_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90000.7 SB=90000.2 A=0.1476 P=2 MULT=1
MM1090 N_Z_M1090_d N_A_184_793#_M1090_g A_117_591# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90000.7 SB=90000.2 A=0.1476 P=2 MULT=1
MM1045 N_VPWR_M1045_d N_S[0]_M1045_g N_A_184_265#_M1045_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1048 N_VPWR_M1048_d N_S[8]_M1048_g N_A_184_793#_M1048_s VPB PHIGHVT L=0.18 W=1
+ AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1039 N_A_533_47#_M1039_d N_S[1]_M1039_g N_VPWR_M1045_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1042 N_A_533_937#_M1042_d N_S[9]_M1042_g N_VPWR_M1048_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1017 A_734_333# N_A_533_47#_M1017_g N_Z_M1017_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1071 A_734_591# N_A_533_937#_M1071_g N_Z_M1071_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1075 N_VPWR_M1075_d N_D[1]_M1075_g A_734_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1076 N_VPWR_M1076_d N_D[9]_M1076_g A_734_591# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1040 A_945_297# N_D[2]_M1040_g N_VPWR_M1075_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1044 A_945_591# N_D[10]_M1044_g N_VPWR_M1076_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1041 N_Z_M1041_d N_A_1012_265#_M1041_g A_945_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1000 N_Z_M1000_d N_A_1012_793#_M1000_g A_945_591# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1050 N_VPWR_M1050_d N_S[2]_M1050_g N_A_1012_265#_M1050_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1053 N_VPWR_M1053_d N_S[10]_M1053_g N_A_1012_793#_M1053_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1009 N_A_1361_47#_M1009_d N_S[3]_M1009_g N_VPWR_M1050_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1012 N_A_1361_937#_M1012_d N_S[11]_M1012_g N_VPWR_M1053_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1022 A_1562_333# N_A_1361_47#_M1022_g N_Z_M1022_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1074 A_1562_591# N_A_1361_937#_M1074_g N_Z_M1074_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1028 N_VPWR_M1028_d N_D[3]_M1028_g A_1562_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1033 N_VPWR_M1033_d N_D[11]_M1033_g A_1562_591# VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 A_1773_297# N_D[4]_M1005_g N_VPWR_M1028_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 A_1773_591# N_D[12]_M1006_g N_VPWR_M1033_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1014 N_Z_M1014_d N_A_1840_265#_M1014_g A_1773_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1064 N_Z_M1064_d N_A_1840_793#_M1064_g A_1773_591# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1080 N_VPWR_M1080_d N_S[4]_M1080_g N_A_1840_265#_M1080_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1085 N_VPWR_M1085_d N_S[12]_M1085_g N_A_1840_793#_M1085_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1046 N_A_2189_47#_M1046_d N_S[5]_M1046_g N_VPWR_M1080_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1049 N_A_2189_937#_M1049_d N_S[13]_M1049_g N_VPWR_M1085_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1059 A_2390_333# N_A_2189_47#_M1059_g N_Z_M1059_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1008 A_2390_591# N_A_2189_937#_M1008_g N_Z_M1008_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.8 A=0.1476 P=2 MULT=1
MM1077 N_VPWR_M1077_d N_D[5]_M1077_g A_2390_333# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1079 N_VPWR_M1079_d N_D[13]_M1079_g A_2390_591# VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.181154 PD=1.35 PS=1.47802 NRD=6.8753 NRS=24.8417 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1029 A_2601_297# N_D[6]_M1029_g N_VPWR_M1077_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1035 A_2601_591# N_D[14]_M1035_g N_VPWR_M1079_d VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.175 PD=1.47802 PS=1.35 NRD=24.8417 NRS=6.8753 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1051 N_Z_M1051_d N_A_2668_265#_M1051_g A_2601_297# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1004 N_Z_M1004_d N_A_2668_793#_M1004_g A_2601_591# VPB PHIGHVT L=0.18 W=0.82
+ AD=0.2214 AS=0.148546 PD=2.18 PS=1.21198 NRD=1.182 NRS=30.2986 M=1 R=4.55556
+ SA=90001.8 SB=90000.2 A=0.1476 P=2 MULT=1
MM1066 N_VPWR_M1066_d N_S[6]_M1066_g N_A_2668_265#_M1066_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1072 N_VPWR_M1072_d N_S[14]_M1072_g N_A_2668_793#_M1072_s VPB PHIGHVT L=0.18
+ W=1 AD=0.2 AS=0.27 PD=1.4 PS=2.54 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1019 N_A_3017_47#_M1019_d N_S[7]_M1019_g N_VPWR_M1066_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90000.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1021 N_A_3017_937#_M1021_d N_S[15]_M1021_g N_VPWR_M1072_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.2 PD=2.54 PS=1.4 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1093 A_3218_333# N_A_3017_47#_M1093_g N_Z_M1093_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.7 A=0.1476 P=2 MULT=1
MM1038 A_3218_591# N_A_3017_937#_M1038_g N_Z_M1038_s VPB PHIGHVT L=0.18 W=0.82
+ AD=0.148546 AS=0.2214 PD=1.21198 PS=2.18 NRD=30.2986 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.7 A=0.1476 P=2 MULT=1
MM1010 N_VPWR_M1010_d N_D[7]_M1010_g A_3218_333# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.181154 PD=2.54 PS=1.47802 NRD=0.9653 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_D[15]_M1013_g A_3218_591# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.181154 PD=2.54 PS=1.47802 NRD=0.9653 NRS=24.8417 M=1 R=5.55556 SA=90000.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX96_noxref VNB VPB NWDIODE A=49.242 P=40.46
*
.include "sky130_fd_sc_hdll__muxb16to1_1.pxi.spice"
*
.ends
*
*
