* File: sky130_fd_sc_hdll__xnor3_1.spice
* Created: Wed Sep  2 08:53:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xnor3_1.pex.spice"
.subckt sky130_fd_sc_hdll__xnor3_1  VNB VPB C B A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1012 N_VGND_M1012_d N_A_83_21#_M1012_g N_X_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.153388 AS=0.182 PD=1.29393 PS=1.86 NRD=4.608 NRS=2.76 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1020 N_A_226_93#_M1020_d N_C_M1020_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1995 AS=0.0991121 PD=1.79 PS=0.836075 NRD=54.276 NRS=51.708 M=1 R=2.8
+ SA=75000.8 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1002 N_A_83_21#_M1002_d N_C_M1002_g N_A_375_49#_M1002_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1088 AS=0.2048 PD=0.98 PS=1.92 NRD=0.936 NRS=8.436 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1013 N_A_351_325#_M1013_d N_A_226_93#_M1013_g N_A_83_21#_M1002_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.224 AS=0.1088 PD=1.98 PS=0.98 NRD=12.18 NRS=10.308 M=1
+ R=4.26667 SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1008 N_A_783_297#_M1008_d N_B_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.16515 AS=0.2535 PD=1.82 PS=2.08 NRD=0 NRS=17.532 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_351_325#_M1006_d N_B_M1006_g N_A_901_297#_M1006_s VNB NSHORT L=0.15
+ W=0.64 AD=0.232513 AS=0.19475 PD=1.56377 PS=1.9 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75000.2 SB=75002.7 A=0.096 P=1.58 MULT=1
MM1016 N_A_1184_297#_M1016_d N_A_783_297#_M1016_g N_A_351_325#_M1006_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.152666 AS=0.152587 PD=1.0183 PS=1.02623 NRD=88.14
+ NRS=108.564 M=1 R=2.8 SA=75001 SB=75003 A=0.063 P=1.14 MULT=1
MM1019 N_A_375_49#_M1019_d N_B_M1019_g N_A_1184_297#_M1016_d VNB NSHORT L=0.15
+ W=0.64 AD=0.175819 AS=0.232634 PD=1.23355 PS=1.5517 NRD=10.308 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1001 N_A_901_297#_M1001_d N_A_783_297#_M1001_g N_A_375_49#_M1019_d VNB NSHORT
+ L=0.15 W=0.6 AD=0.123387 AS=0.164831 PD=1.01129 PS=1.15645 NRD=15.996
+ NRS=41.988 M=1 R=4 SA=75002.1 SB=75001.6 A=0.09 P=1.5 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_901_297#_M1001_d VNB NSHORT L=0.15 W=0.64
+ AD=0.2032 AS=0.131613 PD=1.275 PS=1.07871 NRD=31.872 NRS=8.436 M=1 R=4.26667
+ SA=75002.5 SB=75001 A=0.096 P=1.58 MULT=1
MM1003 N_A_1184_297#_M1003_d N_A_901_297#_M1003_g N_VGND_M1009_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.1824 AS=0.2032 PD=1.85 PS=1.275 NRD=0 NRS=34.68 M=1
+ R=4.26667 SA=75003.3 SB=75000.2 A=0.096 P=1.58 MULT=1
MM1000 N_VPWR_M1000_d N_A_83_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.216098 AS=0.29 PD=1.68902 PS=2.58 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1017 N_A_226_93#_M1017_d N_C_M1017_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1856 AS=0.138302 PD=1.86 PS=1.08098 NRD=1.5366 NRS=49.5849 M=1 R=3.55556
+ SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1015 N_A_83_21#_M1015_d N_C_M1015_g N_A_351_325#_M1015_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.16135 AS=0.2814 PD=1.335 PS=2.35 NRD=1.1623 NRS=1.1623 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1021 N_A_375_49#_M1021_d N_A_226_93#_M1021_g N_A_83_21#_M1015_d VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.33075 AS=0.16135 PD=2.47 PS=1.335 NRD=25.7873 NRS=17.5724
+ M=1 R=4.66667 SA=90000.7 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1004 N_A_783_297#_M1004_d N_B_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.32 AS=0.26655 PD=2.64 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1010 N_A_375_49#_M1010_d N_B_M1010_g N_A_901_297#_M1010_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.284351 AS=0.3612 PD=1.66297 PS=2.54 NRD=48.068 NRS=38.6908 M=1
+ R=4.66667 SA=90000.3 SB=90002.5 A=0.1512 P=2.04 MULT=1
MM1018 N_A_1184_297#_M1018_d N_A_783_297#_M1018_g N_A_375_49#_M1010_d VPB
+ PHIGHVT L=0.18 W=0.64 AD=0.2524 AS=0.216649 PD=1.545 PS=1.26703 NRD=141.584
+ NRS=43.0839 M=1 R=3.55556 SA=90001.1 SB=90002.4 A=0.1152 P=1.64 MULT=1
MM1011 N_A_351_325#_M1011_d N_B_M1011_g N_A_1184_297#_M1018_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.132497 AS=0.2524 PD=1.05946 PS=1.545 NRD=46.7875 NRS=0 M=1
+ R=3.55556 SA=90001.6 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1005 N_A_901_297#_M1005_d N_A_783_297#_M1005_g N_A_351_325#_M1011_d VPB
+ PHIGHVT L=0.18 W=0.84 AD=0.164987 AS=0.173903 PD=1.25543 PS=1.39054
+ NRD=33.1551 NRS=0 M=1 R=4.66667 SA=90001.7 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_901_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.3025 AS=0.196413 PD=1.605 PS=1.49457 NRD=33.4703 NRS=0.9653 M=1 R=5.55556
+ SA=90002 SB=90001 A=0.18 P=2.36 MULT=1
MM1007 N_A_1184_297#_M1007_d N_A_901_297#_M1007_g N_VPWR_M1014_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.295 AS=0.3025 PD=2.59 PS=1.605 NRD=1.9503 NRS=30.535 M=1
+ R=5.55556 SA=90002.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX22_noxref VNB VPB NWDIODE A=15.3759 P=22.37
pX23_noxref noxref_16 B B PROBETYPE=1
c_151 VPB 0 4.99043e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__xnor3_1.pxi.spice"
*
.ends
*
*
