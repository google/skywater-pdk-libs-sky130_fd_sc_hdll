* File: sky130_fd_sc_hdll__o221a_4.pxi.spice
* Created: Thu Aug 27 19:20:31 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221A_4%C1 N_C1_c_115_n N_C1_M1001_g N_C1_c_111_n
+ N_C1_M1002_g N_C1_c_116_n N_C1_M1009_g N_C1_c_112_n N_C1_M1019_g C1
+ N_C1_c_114_n C1 PM_SKY130_FD_SC_HDLL__O221A_4%C1
x_PM_SKY130_FD_SC_HDLL__O221A_4%B1 N_B1_c_151_n N_B1_M1006_g N_B1_c_152_n
+ N_B1_M1014_g N_B1_c_153_n N_B1_M1022_g N_B1_c_154_n N_B1_M1027_g N_B1_c_159_n
+ N_B1_c_155_n B1 B1 N_B1_c_156_n PM_SKY130_FD_SC_HDLL__O221A_4%B1
x_PM_SKY130_FD_SC_HDLL__O221A_4%B2 N_B2_c_226_n N_B2_M1015_g N_B2_c_230_n
+ N_B2_M1011_g N_B2_c_231_n N_B2_M1016_g N_B2_c_227_n N_B2_M1024_g B2
+ N_B2_c_229_n B2 PM_SKY130_FD_SC_HDLL__O221A_4%B2
x_PM_SKY130_FD_SC_HDLL__O221A_4%A1 N_A1_c_268_n N_A1_M1005_g N_A1_c_269_n
+ N_A1_M1000_g N_A1_c_270_n N_A1_M1026_g N_A1_c_271_n N_A1_M1010_g N_A1_c_277_n
+ N_A1_c_272_n N_A1_c_273_n A1 A1 PM_SKY130_FD_SC_HDLL__O221A_4%A1
x_PM_SKY130_FD_SC_HDLL__O221A_4%A2 N_A2_c_345_n N_A2_M1018_g N_A2_c_349_n
+ N_A2_M1013_g N_A2_c_350_n N_A2_M1020_g N_A2_c_346_n N_A2_M1025_g A2
+ N_A2_c_347_n N_A2_c_348_n A2 PM_SKY130_FD_SC_HDLL__O221A_4%A2
x_PM_SKY130_FD_SC_HDLL__O221A_4%A_117_297# N_A_117_297#_M1002_s
+ N_A_117_297#_M1001_s N_A_117_297#_M1011_s N_A_117_297#_M1013_s
+ N_A_117_297#_c_395_n N_A_117_297#_M1003_g N_A_117_297#_c_401_n
+ N_A_117_297#_M1004_g N_A_117_297#_c_396_n N_A_117_297#_M1007_g
+ N_A_117_297#_c_402_n N_A_117_297#_M1012_g N_A_117_297#_c_397_n
+ N_A_117_297#_M1008_g N_A_117_297#_c_403_n N_A_117_297#_M1017_g
+ N_A_117_297#_c_404_n N_A_117_297#_M1023_g N_A_117_297#_c_398_n
+ N_A_117_297#_M1021_g N_A_117_297#_c_399_n N_A_117_297#_c_451_p
+ N_A_117_297#_c_414_n N_A_117_297#_c_434_n N_A_117_297#_c_406_n
+ N_A_117_297#_c_439_n N_A_117_297#_c_491_p N_A_117_297#_c_415_n
+ N_A_117_297#_c_416_n N_A_117_297#_c_400_n
+ PM_SKY130_FD_SC_HDLL__O221A_4%A_117_297#
x_PM_SKY130_FD_SC_HDLL__O221A_4%VPWR N_VPWR_M1001_d N_VPWR_M1009_d
+ N_VPWR_M1022_d N_VPWR_M1026_d N_VPWR_M1012_s N_VPWR_M1023_s N_VPWR_c_547_n
+ N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n
+ N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n
+ N_VPWR_c_558_n N_VPWR_c_559_n VPWR N_VPWR_c_560_n N_VPWR_c_546_n
+ N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n
+ PM_SKY130_FD_SC_HDLL__O221A_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O221A_4%A_305_297# N_A_305_297#_M1006_s
+ N_A_305_297#_M1016_d N_A_305_297#_c_660_n N_A_305_297#_c_666_n
+ N_A_305_297#_c_667_n PM_SKY130_FD_SC_HDLL__O221A_4%A_305_297#
x_PM_SKY130_FD_SC_HDLL__O221A_4%A_785_297# N_A_785_297#_M1005_s
+ N_A_785_297#_M1020_d N_A_785_297#_c_678_n N_A_785_297#_c_684_n
+ N_A_785_297#_c_685_n PM_SKY130_FD_SC_HDLL__O221A_4%A_785_297#
x_PM_SKY130_FD_SC_HDLL__O221A_4%X N_X_M1003_d N_X_M1008_d N_X_M1004_d
+ N_X_M1017_d N_X_c_705_n N_X_c_748_n N_X_c_708_n N_X_c_711_n N_X_c_694_n
+ N_X_c_695_n N_X_c_724_n N_X_c_699_n N_X_c_700_n N_X_c_732_n N_X_c_756_n
+ N_X_c_701_n N_X_c_696_n N_X_c_697_n N_X_c_702_n X
+ PM_SKY130_FD_SC_HDLL__O221A_4%X
x_PM_SKY130_FD_SC_HDLL__O221A_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1019_d
+ N_A_27_47#_M1015_s N_A_27_47#_M1027_d N_A_27_47#_c_780_n N_A_27_47#_c_781_n
+ N_A_27_47#_c_787_n N_A_27_47#_c_782_n N_A_27_47#_c_783_n N_A_27_47#_c_815_p
+ PM_SKY130_FD_SC_HDLL__O221A_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O221A_4%A_307_47# N_A_307_47#_M1014_s
+ N_A_307_47#_M1024_d N_A_307_47#_M1000_d N_A_307_47#_M1025_d
+ N_A_307_47#_c_824_n N_A_307_47#_c_847_n N_A_307_47#_c_825_n
+ N_A_307_47#_c_853_n N_A_307_47#_c_826_n
+ PM_SKY130_FD_SC_HDLL__O221A_4%A_307_47#
x_PM_SKY130_FD_SC_HDLL__O221A_4%VGND N_VGND_M1000_s N_VGND_M1018_s
+ N_VGND_M1010_s N_VGND_M1007_s N_VGND_M1021_s N_VGND_c_885_n N_VGND_c_886_n
+ N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n N_VGND_c_890_n N_VGND_c_891_n
+ N_VGND_c_892_n N_VGND_c_893_n N_VGND_c_894_n N_VGND_c_895_n N_VGND_c_896_n
+ N_VGND_c_897_n VGND N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n
+ N_VGND_c_901_n PM_SKY130_FD_SC_HDLL__O221A_4%VGND
cc_1 VNB N_C1_c_111_n 0.0221633f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_C1_c_112_n 0.0171139f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB C1 0.00832616f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_C1_c_114_n 0.0596535f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_5 VNB N_B1_c_151_n 0.0227132f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_6 VNB N_B1_c_152_n 0.0168034f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_7 VNB N_B1_c_153_n 0.02582f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_8 VNB N_B1_c_154_n 0.022163f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_9 VNB N_B1_c_155_n 0.00407735f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_10 VNB N_B1_c_156_n 0.0053542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B2_c_226_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_B2_c_227_n 0.0173947f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_13 VNB B2 0.00159679f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_14 VNB N_B2_c_229_n 0.0357741f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_15 VNB N_A1_c_268_n 0.0270649f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB N_A1_c_269_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_17 VNB N_A1_c_270_n 0.0241005f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_18 VNB N_A1_c_271_n 0.0169343f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_19 VNB N_A1_c_272_n 0.00735792f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_20 VNB N_A1_c_273_n 2.8054e-19 $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_21 VNB A1 0.00624415f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.175
cc_22 VNB N_A2_c_345_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_23 VNB N_A2_c_346_n 0.0173889f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_24 VNB N_A2_c_347_n 0.00269793f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_25 VNB N_A2_c_348_n 0.036456f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_26 VNB N_A_117_297#_c_395_n 0.0166243f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_27 VNB N_A_117_297#_c_396_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_28 VNB N_A_117_297#_c_397_n 0.0172f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_29 VNB N_A_117_297#_c_398_n 0.02013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_117_297#_c_399_n 0.00199769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_117_297#_c_400_n 0.0771388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_546_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_694_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_34 VNB N_X_c_695_n 0.00252077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_696_n 0.0135579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_697_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB X 0.0232342f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_27_47#_c_780_n 0.00972331f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_39 VNB N_A_27_47#_c_781_n 0.0176817f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.202
cc_40 VNB N_A_27_47#_c_782_n 0.0018401f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_41 VNB N_A_27_47#_c_783_n 0.00294344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_307_47#_c_824_n 0.0295035f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_43 VNB N_A_307_47#_c_825_n 0.00603871f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_44 VNB N_A_307_47#_c_826_n 0.00290513f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_885_n 0.00814995f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_46 VNB N_VGND_c_886_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.175
cc_47 VNB N_VGND_c_887_n 0.00668757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_888_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_889_n 0.0179581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_890_n 0.0176387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_891_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_892_n 0.0201004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_893_n 0.00326658f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_894_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_895_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_896_n 0.0193072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_897_n 0.0048778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_898_n 0.0800581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_899_n 0.0107189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_900_n 0.376114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_901_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VPB N_C1_c_115_n 0.0202694f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_63 VPB N_C1_c_116_n 0.0160914f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_64 VPB N_C1_c_114_n 0.0323232f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_65 VPB N_B1_c_151_n 0.0247986f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_66 VPB N_B1_c_153_n 0.0300116f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_67 VPB N_B1_c_159_n 0.00578212f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_68 VPB N_B1_c_155_n 0.00336065f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_69 VPB N_B1_c_156_n 0.00208789f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B2_c_230_n 0.0159735f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_71 VPB N_B2_c_231_n 0.0159779f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_72 VPB N_B2_c_229_n 0.0192969f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_73 VPB N_A1_c_268_n 0.0303637f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_74 VPB N_A1_c_270_n 0.0259281f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_75 VPB N_A1_c_277_n 0.00670376f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_76 VPB N_A1_c_272_n 0.00397875f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_77 VPB N_A1_c_273_n 0.00134618f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_78 VPB N_A2_c_349_n 0.0159801f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_79 VPB N_A2_c_350_n 0.0159745f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_80 VPB N_A2_c_348_n 0.0193456f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_81 VPB N_A_117_297#_c_401_n 0.015823f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_82 VPB N_A_117_297#_c_402_n 0.0162131f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.175
cc_83 VPB N_A_117_297#_c_403_n 0.0158542f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_117_297#_c_404_n 0.019194f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_117_297#_c_399_n 0.00143102f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_117_297#_c_406_n 0.00516793f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_117_297#_c_400_n 0.0470159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_547_n 0.0116091f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_89 VPB N_VPWR_c_548_n 0.00824019f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.202
cc_90 VPB N_VPWR_c_549_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_91 VPB N_VPWR_c_550_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_551_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_552_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_553_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_554_n 0.0403375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_555_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_556_n 0.0199367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_557_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_558_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_559_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_560_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_546_n 0.0552276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_562_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_563_n 0.0403375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_564_n 0.0226624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_X_c_699_n 4.86412e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_X_c_700_n 0.00138651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_X_c_701_n 0.00202786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_X_c_702_n 0.00150464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB X 0.0258474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 N_C1_c_116_n N_B1_c_151_n 0.0361755f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_112 N_C1_c_114_n N_B1_c_151_n 0.0262361f $X=0.965 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_113 N_C1_c_112_n N_B1_c_152_n 0.00979464f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_114 N_C1_c_116_n N_B1_c_156_n 0.00132328f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_115 N_C1_c_114_n N_B1_c_156_n 0.00314703f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_116 N_C1_c_115_n N_A_117_297#_c_399_n 0.00149306f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_C1_c_111_n N_A_117_297#_c_399_n 0.00289179f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_C1_c_116_n N_A_117_297#_c_399_n 0.00597741f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_C1_c_112_n N_A_117_297#_c_399_n 0.00269744f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_120 C1 N_A_117_297#_c_399_n 0.0144753f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_121 N_C1_c_114_n N_A_117_297#_c_399_n 0.0355952f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_122 N_C1_c_116_n N_A_117_297#_c_414_n 0.0150566f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_123 N_C1_c_111_n N_A_117_297#_c_415_n 0.00775566f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_C1_c_116_n N_A_117_297#_c_416_n 7.63508e-19 $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_125 N_C1_c_115_n N_VPWR_c_548_n 0.00562819f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_126 C1 N_VPWR_c_548_n 0.0193718f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_127 N_C1_c_114_n N_VPWR_c_548_n 0.00610779f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_128 N_C1_c_115_n N_VPWR_c_549_n 0.00702461f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C1_c_116_n N_VPWR_c_549_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_130 N_C1_c_116_n N_VPWR_c_550_n 0.00294959f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C1_c_115_n N_VPWR_c_546_n 0.0132955f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C1_c_116_n N_VPWR_c_546_n 0.00698456f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_133 N_C1_c_111_n N_A_27_47#_c_781_n 0.00440997f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_134 C1 N_A_27_47#_c_781_n 0.0198144f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_135 N_C1_c_114_n N_A_27_47#_c_781_n 0.00595621f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_136 N_C1_c_111_n N_A_27_47#_c_787_n 0.0115292f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C1_c_112_n N_A_27_47#_c_787_n 0.0140389f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_138 C1 N_A_27_47#_c_787_n 0.0017805f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_139 N_C1_c_114_n N_A_27_47#_c_787_n 0.00215693f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_140 N_C1_c_111_n N_VGND_c_898_n 0.00357877f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_141 N_C1_c_112_n N_VGND_c_898_n 0.00357877f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_142 N_C1_c_111_n N_VGND_c_900_n 0.00635588f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_143 N_C1_c_112_n N_VGND_c_900_n 0.00550244f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B1_c_152_n N_B2_c_226_n 0.0267679f $X=1.46 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_145 N_B1_c_151_n N_B2_c_230_n 0.0385271f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B1_c_159_n N_B2_c_230_n 0.013461f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_147 N_B1_c_156_n N_B2_c_230_n 0.00105708f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_148 N_B1_c_153_n N_B2_c_231_n 0.0385408f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B1_c_159_n N_B2_c_231_n 0.0113203f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_150 N_B1_c_155_n N_B2_c_231_n 9.98177e-19 $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_151 N_B1_c_154_n N_B2_c_227_n 0.0223535f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B1_c_153_n B2 6.6954e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B1_c_159_n B2 0.0386816f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_154 N_B1_c_155_n B2 0.0173853f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_155 N_B1_c_156_n B2 0.0142733f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_156 N_B1_c_151_n N_B2_c_229_n 0.0262094f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_157 N_B1_c_153_n N_B2_c_229_n 0.0251351f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B1_c_159_n N_B2_c_229_n 0.00803891f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_159 N_B1_c_155_n N_B2_c_229_n 0.00388221f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_160 N_B1_c_156_n N_B2_c_229_n 0.00594076f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_161 N_B1_c_153_n N_A1_c_268_n 0.00583907f $X=2.845 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_162 N_B1_c_155_n N_A1_c_268_n 9.05184e-19 $X=2.83 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_163 N_B1_c_153_n N_A1_c_272_n 0.00290896f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_164 N_B1_c_155_n N_A1_c_272_n 0.0351503f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_165 N_B1_c_159_n N_A_117_297#_M1011_s 0.00187547f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_166 N_B1_c_151_n N_A_117_297#_c_399_n 0.00154949f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_B1_c_156_n N_A_117_297#_c_399_n 0.0372081f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_168 N_B1_c_151_n N_A_117_297#_c_414_n 0.0136317f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B1_c_153_n N_A_117_297#_c_414_n 0.015667f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B1_c_155_n N_A_117_297#_c_414_n 0.0201576f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_171 N_B1_c_156_n N_A_117_297#_c_414_n 0.0886333f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_172 N_B1_c_156_n N_VPWR_M1009_d 0.00219254f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_173 N_B1_c_155_n N_VPWR_M1022_d 0.00229269f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_174 N_B1_c_151_n N_VPWR_c_550_n 0.0030665f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B1_c_151_n N_VPWR_c_546_n 0.00695991f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B1_c_153_n N_VPWR_c_546_n 0.00826476f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B1_c_151_n N_VPWR_c_563_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B1_c_153_n N_VPWR_c_563_n 0.00702461f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B1_c_153_n N_VPWR_c_564_n 0.00505472f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_159_n N_A_305_297#_M1006_s 2.87715e-19 $X=2.665 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_181 N_B1_c_156_n N_A_305_297#_M1006_s 0.00163414f $X=1.73 $Y=1.345 $X2=-0.19
+ $Y2=-0.24
cc_182 N_B1_c_159_n N_A_305_297#_M1016_d 0.00182938f $X=2.665 $Y=1.53 $X2=0
+ $Y2=0
cc_183 N_B1_c_155_n N_A_305_297#_M1016_d 6.67308e-19 $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_184 N_B1_c_151_n N_A_27_47#_c_782_n 2.30339e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B1_c_152_n N_A_27_47#_c_782_n 0.00393466f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B1_c_156_n N_A_27_47#_c_782_n 0.0153113f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_187 N_B1_c_151_n N_A_27_47#_c_783_n 0.00167844f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B1_c_152_n N_A_27_47#_c_783_n 0.0098207f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_189 N_B1_c_154_n N_A_27_47#_c_783_n 0.00923997f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_190 N_B1_c_156_n N_A_27_47#_c_783_n 0.00389822f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_191 N_B1_c_151_n N_A_307_47#_c_824_n 0.00149476f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B1_c_152_n N_A_307_47#_c_824_n 0.00599667f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_193 N_B1_c_153_n N_A_307_47#_c_824_n 0.0044163f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B1_c_154_n N_A_307_47#_c_824_n 0.0142117f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_195 N_B1_c_159_n N_A_307_47#_c_824_n 0.0125151f $X=2.665 $Y=1.53 $X2=0 $Y2=0
cc_196 N_B1_c_155_n N_A_307_47#_c_824_n 0.0302712f $X=2.83 $Y=1.16 $X2=0 $Y2=0
cc_197 N_B1_c_156_n N_A_307_47#_c_824_n 0.0224424f $X=1.73 $Y=1.345 $X2=0 $Y2=0
cc_198 N_B1_c_154_n N_VGND_c_885_n 0.00236436f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_199 N_B1_c_152_n N_VGND_c_898_n 0.00357877f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_200 N_B1_c_154_n N_VGND_c_898_n 0.00357877f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_152_n N_VGND_c_900_n 0.00539883f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_202 N_B1_c_154_n N_VGND_c_900_n 0.00670225f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_203 N_B2_c_230_n N_A_117_297#_c_414_n 0.0108425f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B2_c_231_n N_A_117_297#_c_414_n 0.0108425f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B2_c_230_n N_VPWR_c_546_n 0.00609021f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B2_c_231_n N_VPWR_c_546_n 0.00609021f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B2_c_230_n N_VPWR_c_563_n 0.00429453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B2_c_231_n N_VPWR_c_563_n 0.00429453f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B2_c_230_n N_A_305_297#_c_660_n 0.0099733f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B2_c_231_n N_A_305_297#_c_660_n 0.0099733f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B2_c_226_n N_A_27_47#_c_783_n 0.00881459f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B2_c_227_n N_A_27_47#_c_783_n 0.00923997f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B2_c_226_n N_A_307_47#_c_824_n 0.0135773f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B2_c_227_n N_A_307_47#_c_824_n 0.0118409f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_215 B2 N_A_307_47#_c_824_n 0.0402792f $X=2.19 $Y=1.105 $X2=0 $Y2=0
cc_216 N_B2_c_229_n N_A_307_47#_c_824_n 0.0047334f $X=2.375 $Y=1.202 $X2=0 $Y2=0
cc_217 N_B2_c_226_n N_VGND_c_898_n 0.00357877f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B2_c_227_n N_VGND_c_898_n 0.00357877f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B2_c_226_n N_VGND_c_900_n 0.00549573f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B2_c_227_n N_VGND_c_900_n 0.00561849f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A1_c_269_n N_A2_c_345_n 0.0165763f $X=3.86 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_222 N_A1_c_268_n N_A2_c_349_n 0.0385591f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A1_c_277_n N_A2_c_349_n 0.0115164f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_224 N_A1_c_272_n N_A2_c_349_n 9.9831e-19 $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A1_c_270_n N_A2_c_350_n 0.0379119f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A1_c_277_n N_A2_c_350_n 0.0131991f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_227 N_A1_c_273_n N_A2_c_350_n 8.25237e-19 $X=5.1 $Y=1.445 $X2=0 $Y2=0
cc_228 N_A1_c_271_n N_A2_c_346_n 0.0103136f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A1_c_268_n N_A2_c_347_n 7.32803e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A1_c_277_n N_A2_c_347_n 0.0449721f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_231 N_A1_c_272_n N_A2_c_347_n 0.0182967f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_232 A1 N_A2_c_347_n 0.0142244f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_233 N_A1_c_268_n N_A2_c_348_n 0.0165763f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A1_c_270_n N_A2_c_348_n 0.0262494f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A1_c_277_n N_A2_c_348_n 0.0080388f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_236 N_A1_c_272_n N_A2_c_348_n 0.00403136f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A1_c_273_n N_A2_c_348_n 0.00328579f $X=5.1 $Y=1.445 $X2=0 $Y2=0
cc_238 A1 N_A2_c_348_n 0.00171552f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A1_c_277_n N_A_117_297#_M1013_s 0.00187547f $X=4.975 $Y=1.53 $X2=0
+ $Y2=0
cc_240 N_A1_c_271_n N_A_117_297#_c_395_n 0.012217f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A1_c_270_n N_A_117_297#_c_401_n 0.0352481f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A1_c_268_n N_A_117_297#_c_414_n 0.0157639f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A1_c_270_n N_A_117_297#_c_414_n 0.0156384f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A1_c_277_n N_A_117_297#_c_414_n 0.0687248f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_245 N_A1_c_272_n N_A_117_297#_c_414_n 0.0439529f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_246 A1 N_A_117_297#_c_414_n 0.00663869f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A1_c_270_n N_A_117_297#_c_434_n 0.00367495f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A1_c_270_n N_A_117_297#_c_406_n 0.00188746f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A1_c_277_n N_A_117_297#_c_406_n 0.0106198f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_250 N_A1_c_273_n N_A_117_297#_c_406_n 0.00512702f $X=5.1 $Y=1.445 $X2=0 $Y2=0
cc_251 A1 N_A_117_297#_c_406_n 0.00457456f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_252 A1 N_A_117_297#_c_439_n 0.0173838f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A1_c_270_n N_A_117_297#_c_400_n 0.0265394f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A1_c_273_n N_A_117_297#_c_400_n 4.17602e-19 $X=5.1 $Y=1.445 $X2=0 $Y2=0
cc_255 A1 N_A_117_297#_c_400_n 0.0015569f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_256 N_A1_c_272_n N_VPWR_M1022_d 0.00731812f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A1_c_270_n N_VPWR_c_551_n 0.00300743f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A1_c_268_n N_VPWR_c_554_n 0.00702461f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A1_c_270_n N_VPWR_c_554_n 0.00702461f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A1_c_268_n N_VPWR_c_546_n 0.00823967f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A1_c_270_n N_VPWR_c_546_n 0.006985f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A1_c_268_n N_VPWR_c_564_n 0.00514457f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A1_c_277_n N_A_785_297#_M1005_s 0.00187547f $X=4.975 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_264 N_A1_c_277_n N_A_785_297#_M1020_d 0.00190905f $X=4.975 $Y=1.53 $X2=0
+ $Y2=0
cc_265 N_A1_c_268_n N_A_307_47#_c_824_n 0.00466528f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A1_c_269_n N_A_307_47#_c_824_n 0.0155787f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A1_c_277_n N_A_307_47#_c_824_n 0.00102987f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_268 N_A1_c_272_n N_A_307_47#_c_824_n 0.0532824f $X=3.74 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A1_c_270_n N_A_307_47#_c_825_n 0.00239967f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A1_c_271_n N_A_307_47#_c_825_n 2.01812e-19 $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A1_c_277_n N_A_307_47#_c_825_n 0.00717418f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_272 A1 N_A_307_47#_c_825_n 0.0179599f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_273 N_A1_c_277_n N_A_307_47#_c_826_n 0.00527349f $X=4.975 $Y=1.53 $X2=0 $Y2=0
cc_274 N_A1_c_269_n N_VGND_c_885_n 0.00482545f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A1_c_270_n N_VGND_c_887_n 2.31083e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A1_c_271_n N_VGND_c_887_n 0.00283672f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_277 A1 N_VGND_c_887_n 0.0118366f $X=5.21 $Y=1.105 $X2=0 $Y2=0
cc_278 N_A1_c_269_n N_VGND_c_890_n 0.00426565f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A1_c_271_n N_VGND_c_892_n 0.00585385f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A1_c_269_n N_VGND_c_900_n 0.00697014f $X=3.86 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A1_c_271_n N_VGND_c_900_n 0.0107097f $X=5.27 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A2_c_349_n N_A_117_297#_c_414_n 0.0108425f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_283 N_A2_c_350_n N_A_117_297#_c_414_n 0.0108425f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_284 N_A2_c_349_n N_VPWR_c_554_n 0.00429453f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_285 N_A2_c_350_n N_VPWR_c_554_n 0.00429453f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A2_c_349_n N_VPWR_c_546_n 0.00609021f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A2_c_350_n N_VPWR_c_546_n 0.00609021f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_288 N_A2_c_349_n N_A_785_297#_c_678_n 0.0099733f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_289 N_A2_c_350_n N_A_785_297#_c_678_n 0.0099733f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A2_c_345_n N_A_307_47#_c_847_n 0.00543771f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A2_c_346_n N_A_307_47#_c_847_n 2.9078e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A2_c_345_n N_A_307_47#_c_825_n 0.00929182f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A2_c_346_n N_A_307_47#_c_825_n 0.0106577f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A2_c_347_n N_A_307_47#_c_825_n 0.0372111f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A2_c_348_n N_A_307_47#_c_825_n 0.00468948f $X=4.775 $Y=1.202 $X2=0
+ $Y2=0
cc_296 N_A2_c_345_n N_A_307_47#_c_853_n 5.69179e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A2_c_346_n N_A_307_47#_c_853_n 0.00856992f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A2_c_345_n N_A_307_47#_c_826_n 0.00262985f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A2_c_346_n N_A_307_47#_c_826_n 2.4448e-19 $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A2_c_347_n N_A_307_47#_c_826_n 0.00911001f $X=4.54 $Y=1.16 $X2=0 $Y2=0
cc_301 N_A2_c_345_n N_VGND_c_886_n 0.00385467f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A2_c_346_n N_VGND_c_886_n 0.00365402f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A2_c_345_n N_VGND_c_890_n 0.00423334f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A2_c_346_n N_VGND_c_892_n 0.00396605f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A2_c_345_n N_VGND_c_900_n 0.00610858f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A2_c_346_n N_VGND_c_900_n 0.00594864f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_117_297#_c_414_n N_VPWR_M1009_d 0.00369247f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_308 N_A_117_297#_c_414_n N_VPWR_M1022_d 0.0259264f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_309 N_A_117_297#_c_414_n N_VPWR_M1026_d 0.00328773f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_310 N_A_117_297#_c_434_n N_VPWR_M1026_d 0.00219605f $X=5.56 $Y=1.785 $X2=0
+ $Y2=0
cc_311 N_A_117_297#_c_406_n N_VPWR_M1026_d 0.00155253f $X=5.815 $Y=1.445 $X2=0
+ $Y2=0
cc_312 N_A_117_297#_c_399_n N_VPWR_c_548_n 0.00194745f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_313 N_A_117_297#_c_451_p N_VPWR_c_549_n 0.0149311f $X=0.73 $Y=1.96 $X2=0
+ $Y2=0
cc_314 N_A_117_297#_c_414_n N_VPWR_c_550_n 0.0139109f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_315 N_A_117_297#_c_401_n N_VPWR_c_551_n 0.00300743f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_316 N_A_117_297#_c_414_n N_VPWR_c_551_n 0.0142681f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_317 N_A_117_297#_c_402_n N_VPWR_c_552_n 0.00300743f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_318 N_A_117_297#_c_403_n N_VPWR_c_552_n 0.00300743f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_117_297#_c_404_n N_VPWR_c_553_n 0.00479105f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_117_297#_c_401_n N_VPWR_c_556_n 0.00702461f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_321 N_A_117_297#_c_402_n N_VPWR_c_556_n 0.00702461f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_322 N_A_117_297#_c_403_n N_VPWR_c_558_n 0.00702461f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_323 N_A_117_297#_c_404_n N_VPWR_c_558_n 0.00702461f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_324 N_A_117_297#_M1001_s N_VPWR_c_546_n 0.00339604f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_325 N_A_117_297#_M1011_s N_VPWR_c_546_n 0.00232895f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_326 N_A_117_297#_M1013_s N_VPWR_c_546_n 0.00232895f $X=4.395 $Y=1.485 $X2=0
+ $Y2=0
cc_327 N_A_117_297#_c_401_n N_VPWR_c_546_n 0.0118497f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_328 N_A_117_297#_c_402_n N_VPWR_c_546_n 0.00693457f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_329 N_A_117_297#_c_403_n N_VPWR_c_546_n 0.0124092f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_330 N_A_117_297#_c_404_n N_VPWR_c_546_n 0.0134606f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_331 N_A_117_297#_c_451_p N_VPWR_c_546_n 0.00955092f $X=0.73 $Y=1.96 $X2=0
+ $Y2=0
cc_332 N_A_117_297#_c_414_n N_VPWR_c_546_n 0.043839f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_333 N_A_117_297#_c_416_n N_VPWR_c_546_n 0.00100653f $X=0.755 $Y=1.87 $X2=0
+ $Y2=0
cc_334 N_A_117_297#_c_414_n N_VPWR_c_564_n 0.0547305f $X=5.475 $Y=1.87 $X2=0
+ $Y2=0
cc_335 N_A_117_297#_c_414_n N_A_305_297#_M1006_s 0.00369247f $X=5.475 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_336 N_A_117_297#_c_414_n N_A_305_297#_M1016_d 0.00365569f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_337 N_A_117_297#_M1011_s N_A_305_297#_c_660_n 0.00424775f $X=1.995 $Y=1.485
+ $X2=0 $Y2=0
cc_338 N_A_117_297#_c_414_n N_A_305_297#_c_660_n 0.0188794f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_339 N_A_117_297#_c_414_n N_A_305_297#_c_666_n 0.0131392f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_340 N_A_117_297#_c_414_n N_A_305_297#_c_667_n 0.0130645f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_341 N_A_117_297#_c_414_n N_A_785_297#_M1005_s 0.00370949f $X=5.475 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_342 N_A_117_297#_c_414_n N_A_785_297#_M1020_d 0.00368934f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_343 N_A_117_297#_M1013_s N_A_785_297#_c_678_n 0.00424775f $X=4.395 $Y=1.485
+ $X2=0 $Y2=0
cc_344 N_A_117_297#_c_414_n N_A_785_297#_c_678_n 0.0188794f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_345 N_A_117_297#_c_414_n N_A_785_297#_c_684_n 0.0131392f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_346 N_A_117_297#_c_414_n N_A_785_297#_c_685_n 0.0131392f $X=5.475 $Y=1.87
+ $X2=0 $Y2=0
cc_347 N_A_117_297#_c_406_n N_X_M1004_d 0.00223383f $X=5.815 $Y=1.445 $X2=0
+ $Y2=0
cc_348 N_A_117_297#_c_395_n N_X_c_705_n 0.00513121f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_349 N_A_117_297#_c_396_n N_X_c_705_n 0.00686626f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_350 N_A_117_297#_c_397_n N_X_c_705_n 5.45498e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_351 N_A_117_297#_c_402_n N_X_c_708_n 0.0127987f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_117_297#_c_403_n N_X_c_708_n 0.00168782f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A_117_297#_c_491_p N_X_c_708_n 0.00608731f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_354 N_A_117_297#_c_414_n N_X_c_711_n 0.0120976f $X=5.475 $Y=1.87 $X2=0 $Y2=0
cc_355 N_A_117_297#_c_406_n N_X_c_711_n 0.00488151f $X=5.815 $Y=1.445 $X2=0
+ $Y2=0
cc_356 N_A_117_297#_c_491_p N_X_c_711_n 0.00435403f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_357 N_A_117_297#_c_400_n N_X_c_711_n 0.00302225f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_358 N_A_117_297#_c_396_n N_X_c_694_n 0.00901745f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_359 N_A_117_297#_c_397_n N_X_c_694_n 0.00901745f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_360 N_A_117_297#_c_491_p N_X_c_694_n 0.0397461f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A_117_297#_c_400_n N_X_c_694_n 0.00345541f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_362 N_A_117_297#_c_395_n N_X_c_695_n 0.002559f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A_117_297#_c_396_n N_X_c_695_n 0.00116636f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_117_297#_c_439_n N_X_c_695_n 0.0160387f $X=5.925 $Y=1.175 $X2=0 $Y2=0
cc_365 N_A_117_297#_c_491_p N_X_c_695_n 0.0152659f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_366 N_A_117_297#_c_400_n N_X_c_695_n 0.00358172f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_367 N_A_117_297#_c_403_n N_X_c_724_n 0.00143499f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_117_297#_c_403_n N_X_c_699_n 0.0152802f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_369 N_A_117_297#_c_491_p N_X_c_699_n 0.0184316f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_370 N_A_117_297#_c_400_n N_X_c_699_n 0.00242942f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_371 N_A_117_297#_c_402_n N_X_c_700_n 0.00111277f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_372 N_A_117_297#_c_406_n N_X_c_700_n 0.00476901f $X=5.815 $Y=1.445 $X2=0
+ $Y2=0
cc_373 N_A_117_297#_c_491_p N_X_c_700_n 0.0135262f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_374 N_A_117_297#_c_400_n N_X_c_700_n 0.00430965f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_375 N_A_117_297#_c_396_n N_X_c_732_n 5.24597e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_376 N_A_117_297#_c_397_n N_X_c_732_n 0.00651696f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A_117_297#_c_404_n N_X_c_701_n 0.0192758f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_378 N_A_117_297#_c_491_p N_X_c_701_n 0.00278263f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_379 N_A_117_297#_c_400_n N_X_c_701_n 9.44081e-19 $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_380 N_A_117_297#_c_398_n N_X_c_696_n 0.0139504f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A_117_297#_c_397_n N_X_c_697_n 0.00119564f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A_117_297#_c_491_p N_X_c_697_n 0.0307352f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_383 N_A_117_297#_c_400_n N_X_c_697_n 0.00486271f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_384 N_A_117_297#_c_491_p N_X_c_702_n 0.020385f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_385 N_A_117_297#_c_400_n N_X_c_702_n 0.00643699f $X=7.125 $Y=1.202 $X2=0
+ $Y2=0
cc_386 N_A_117_297#_c_404_n X 0.00132098f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_387 N_A_117_297#_c_398_n X 0.0187563f $X=7.15 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A_117_297#_c_491_p X 0.0106198f $X=6.89 $Y=1.16 $X2=0 $Y2=0
cc_389 N_A_117_297#_c_399_n N_A_27_47#_c_781_n 0.00110546f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_390 N_A_117_297#_c_415_n N_A_27_47#_c_781_n 0.0169491f $X=0.73 $Y=0.73 $X2=0
+ $Y2=0
cc_391 N_A_117_297#_M1002_s N_A_27_47#_c_787_n 0.00399909f $X=0.595 $Y=0.235
+ $X2=0 $Y2=0
cc_392 N_A_117_297#_c_415_n N_A_27_47#_c_787_n 0.0214489f $X=0.73 $Y=0.73 $X2=0
+ $Y2=0
cc_393 N_A_117_297#_c_399_n N_A_27_47#_c_782_n 0.00123997f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_394 N_A_117_297#_c_395_n N_VGND_c_887_n 0.00282267f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_395 N_A_117_297#_c_406_n N_VGND_c_887_n 0.00109643f $X=5.815 $Y=1.445 $X2=0
+ $Y2=0
cc_396 N_A_117_297#_c_396_n N_VGND_c_888_n 0.00379224f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_397 N_A_117_297#_c_397_n N_VGND_c_888_n 0.00276126f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_398 N_A_117_297#_c_398_n N_VGND_c_889_n 0.00450113f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_399 N_A_117_297#_c_395_n N_VGND_c_894_n 0.00541359f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_400 N_A_117_297#_c_396_n N_VGND_c_894_n 0.00423334f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_401 N_A_117_297#_c_397_n N_VGND_c_896_n 0.00423334f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_402 N_A_117_297#_c_398_n N_VGND_c_896_n 0.00439206f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_403 N_A_117_297#_M1002_s N_VGND_c_900_n 0.00256987f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_404 N_A_117_297#_c_395_n N_VGND_c_900_n 0.00965571f $X=5.69 $Y=0.995 $X2=0
+ $Y2=0
cc_405 N_A_117_297#_c_396_n N_VGND_c_900_n 0.006093f $X=6.16 $Y=0.995 $X2=0
+ $Y2=0
cc_406 N_A_117_297#_c_397_n N_VGND_c_900_n 0.00608558f $X=6.63 $Y=0.995 $X2=0
+ $Y2=0
cc_407 N_A_117_297#_c_398_n N_VGND_c_900_n 0.00725214f $X=7.15 $Y=0.995 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_546_n N_A_305_297#_M1006_s 0.00247166f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_409 N_VPWR_c_546_n N_A_305_297#_M1016_d 0.0023603f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_546_n N_A_305_297#_c_660_n 0.0239224f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_563_n N_A_305_297#_c_660_n 0.0386815f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_546_n N_A_305_297#_c_666_n 0.00938745f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_563_n N_A_305_297#_c_666_n 0.014332f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_546_n N_A_305_297#_c_667_n 0.00938288f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_563_n N_A_305_297#_c_667_n 0.0143006f $X=2.965 $Y=2.465 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_546_n N_A_785_297#_M1005_s 0.00241598f $X=7.59 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_417 N_VPWR_c_546_n N_A_785_297#_M1020_d 0.00241598f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_554_n N_A_785_297#_c_678_n 0.0386815f $X=5.355 $Y=2.72 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_546_n N_A_785_297#_c_678_n 0.0239224f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_554_n N_A_785_297#_c_684_n 0.014332f $X=5.355 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_546_n N_A_785_297#_c_684_n 0.00938745f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_554_n N_A_785_297#_c_685_n 0.014332f $X=5.355 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_546_n N_A_785_297#_c_685_n 0.00938745f $X=7.59 $Y=2.72 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_546_n N_X_M1004_d 0.00449333f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_425 N_VPWR_c_546_n N_X_M1017_d 0.00370124f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_426 N_VPWR_c_556_n N_X_c_748_n 0.0133725f $X=6.295 $Y=2.72 $X2=0 $Y2=0
cc_427 N_VPWR_c_546_n N_X_c_748_n 0.00801045f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_M1012_s N_X_c_708_n 0.00360212f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_429 N_VPWR_c_552_n N_X_c_708_n 0.0143751f $X=6.42 $Y=2.3 $X2=0 $Y2=0
cc_430 N_VPWR_c_546_n N_X_c_708_n 0.0074233f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_431 N_VPWR_M1012_s N_X_c_724_n 0.00138147f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_432 N_VPWR_c_552_n N_X_c_699_n 2.71364e-19 $X=6.42 $Y=2.3 $X2=0 $Y2=0
cc_433 N_VPWR_M1012_s N_X_c_700_n 3.54961e-19 $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_434 N_VPWR_c_558_n N_X_c_756_n 0.0149311f $X=7.235 $Y=2.72 $X2=0 $Y2=0
cc_435 N_VPWR_c_546_n N_X_c_756_n 0.00955092f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_436 N_VPWR_M1023_s N_X_c_701_n 0.00100172f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_437 N_VPWR_c_553_n N_X_c_701_n 0.00721472f $X=7.36 $Y=1.96 $X2=0 $Y2=0
cc_438 N_VPWR_M1023_s X 0.00199676f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_439 N_VPWR_c_553_n X 0.0102775f $X=7.36 $Y=1.96 $X2=0 $Y2=0
cc_440 N_X_c_694_n N_VGND_M1007_s 0.00251047f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_441 N_X_c_696_n N_VGND_M1021_s 0.00281303f $X=7.365 $Y=0.82 $X2=0 $Y2=0
cc_442 N_X_c_695_n N_VGND_c_887_n 0.00830019f $X=6.115 $Y=0.815 $X2=0 $Y2=0
cc_443 N_X_c_705_n N_VGND_c_888_n 0.0183628f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_444 N_X_c_694_n N_VGND_c_888_n 0.0127273f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_445 N_X_c_696_n N_VGND_c_889_n 0.0208473f $X=7.365 $Y=0.82 $X2=0 $Y2=0
cc_446 N_X_c_705_n N_VGND_c_894_n 0.0223596f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_447 N_X_c_694_n N_VGND_c_894_n 0.00266636f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_448 N_X_c_694_n N_VGND_c_896_n 0.00198695f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_449 N_X_c_732_n N_VGND_c_896_n 0.0231806f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_450 N_X_c_696_n N_VGND_c_896_n 0.00248202f $X=7.365 $Y=0.82 $X2=0 $Y2=0
cc_451 N_X_c_696_n N_VGND_c_899_n 0.00300062f $X=7.365 $Y=0.82 $X2=0 $Y2=0
cc_452 N_X_M1003_d N_VGND_c_900_n 0.0025535f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_453 N_X_M1008_d N_VGND_c_900_n 0.00304426f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_454 N_X_c_705_n N_VGND_c_900_n 0.0141302f $X=5.95 $Y=0.39 $X2=0 $Y2=0
cc_455 N_X_c_694_n N_VGND_c_900_n 0.00972452f $X=6.675 $Y=0.815 $X2=0 $Y2=0
cc_456 N_X_c_732_n N_VGND_c_900_n 0.0143352f $X=6.89 $Y=0.39 $X2=0 $Y2=0
cc_457 N_X_c_696_n N_VGND_c_900_n 0.0110296f $X=7.365 $Y=0.82 $X2=0 $Y2=0
cc_458 N_A_27_47#_c_783_n N_A_307_47#_M1014_s 0.00312026f $X=3.08 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_459 N_A_27_47#_c_783_n N_A_307_47#_M1024_d 0.00411406f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_460 N_A_27_47#_M1015_s N_A_307_47#_c_824_n 0.00279596f $X=1.955 $Y=0.235
+ $X2=0 $Y2=0
cc_461 N_A_27_47#_M1027_d N_A_307_47#_c_824_n 0.0031705f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_462 N_A_27_47#_c_782_n N_A_307_47#_c_824_n 0.0203033f $X=1.2 $Y=0.73 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_783_n N_A_307_47#_c_824_n 0.0991323f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_464 N_A_27_47#_c_783_n N_VGND_c_885_n 0.0177537f $X=3.08 $Y=0.38 $X2=0 $Y2=0
cc_465 N_A_27_47#_c_780_n N_VGND_c_898_n 0.0182708f $X=0.215 $Y=0.475 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_c_787_n N_VGND_c_898_n 0.0425444f $X=1.115 $Y=0.365 $X2=0
+ $Y2=0
cc_467 N_A_27_47#_c_783_n N_VGND_c_898_n 0.112499f $X=3.08 $Y=0.38 $X2=0 $Y2=0
cc_468 N_A_27_47#_c_815_p N_VGND_c_898_n 0.011673f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_469 N_A_27_47#_M1002_d N_VGND_c_900_n 0.00250318f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_M1019_d N_VGND_c_900_n 0.00255365f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_471 N_A_27_47#_M1015_s N_VGND_c_900_n 0.00295535f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_472 N_A_27_47#_M1027_d N_VGND_c_900_n 0.00209344f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_473 N_A_27_47#_c_780_n N_VGND_c_900_n 0.00999725f $X=0.215 $Y=0.475 $X2=0
+ $Y2=0
cc_474 N_A_27_47#_c_787_n N_VGND_c_900_n 0.0273233f $X=1.115 $Y=0.365 $X2=0
+ $Y2=0
cc_475 N_A_27_47#_c_783_n N_VGND_c_900_n 0.070764f $X=3.08 $Y=0.38 $X2=0 $Y2=0
cc_476 N_A_27_47#_c_815_p N_VGND_c_900_n 0.00653933f $X=1.2 $Y=0.39 $X2=0 $Y2=0
cc_477 N_A_307_47#_c_824_n N_VGND_M1000_s 0.00440719f $X=3.985 $Y=0.775
+ $X2=-0.19 $Y2=-0.24
cc_478 N_A_307_47#_c_825_n N_VGND_M1018_s 0.00348805f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_479 N_A_307_47#_c_824_n N_VGND_c_885_n 0.0219584f $X=3.985 $Y=0.775 $X2=0
+ $Y2=0
cc_480 N_A_307_47#_c_847_n N_VGND_c_886_n 0.0177813f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_481 N_A_307_47#_c_825_n N_VGND_c_886_n 0.0131987f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_482 N_A_307_47#_c_853_n N_VGND_c_886_n 0.0223967f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_483 N_A_307_47#_c_825_n N_VGND_c_887_n 0.00133683f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_484 N_A_307_47#_c_824_n N_VGND_c_890_n 0.00311455f $X=3.985 $Y=0.775 $X2=0
+ $Y2=0
cc_485 N_A_307_47#_c_847_n N_VGND_c_890_n 0.0151073f $X=4.07 $Y=0.42 $X2=0 $Y2=0
cc_486 N_A_307_47#_c_825_n N_VGND_c_890_n 0.00266636f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_487 N_A_307_47#_c_825_n N_VGND_c_892_n 0.00199443f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_488 N_A_307_47#_c_853_n N_VGND_c_892_n 0.023074f $X=5.01 $Y=0.39 $X2=0 $Y2=0
cc_489 N_A_307_47#_c_824_n N_VGND_c_898_n 0.00331169f $X=3.985 $Y=0.775 $X2=0
+ $Y2=0
cc_490 N_A_307_47#_M1014_s N_VGND_c_900_n 0.00216833f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_491 N_A_307_47#_M1024_d N_VGND_c_900_n 0.00256987f $X=2.475 $Y=0.235 $X2=0
+ $Y2=0
cc_492 N_A_307_47#_M1000_d N_VGND_c_900_n 0.00232983f $X=3.935 $Y=0.235 $X2=0
+ $Y2=0
cc_493 N_A_307_47#_M1025_d N_VGND_c_900_n 0.00324782f $X=4.875 $Y=0.235 $X2=0
+ $Y2=0
cc_494 N_A_307_47#_c_824_n N_VGND_c_900_n 0.0156742f $X=3.985 $Y=0.775 $X2=0
+ $Y2=0
cc_495 N_A_307_47#_c_847_n N_VGND_c_900_n 0.00933462f $X=4.07 $Y=0.42 $X2=0
+ $Y2=0
cc_496 N_A_307_47#_c_825_n N_VGND_c_900_n 0.0100158f $X=4.795 $Y=0.815 $X2=0
+ $Y2=0
cc_497 N_A_307_47#_c_853_n N_VGND_c_900_n 0.0141066f $X=5.01 $Y=0.39 $X2=0 $Y2=0
