* NGSPICE file created from sky130_fd_sc_hdll__nor2b_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nor2b_1 A B_N VGND VNB VPB VPWR Y
M1000 a_253_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.3e+11p pd=2.46e+06u as=3.666e+11p ps=3e+06u
M1001 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1002 VGND a_27_47# Y VNB nshort w=650000u l=150000u
+  ad=4.912e+11p pd=4.26e+06u as=1.755e+11p ps=1.84e+06u
M1003 Y A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_47# a_253_297# VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1005 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends

