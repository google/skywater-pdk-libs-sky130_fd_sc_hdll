* File: sky130_fd_sc_hdll__o22a_1.pxi.spice
* Created: Wed Sep  2 08:45:14 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22A_1%A_83_21# N_A_83_21#_M1008_d N_A_83_21#_M1003_d
+ N_A_83_21#_c_49_n N_A_83_21#_M1006_g N_A_83_21#_c_50_n N_A_83_21#_M1001_g
+ N_A_83_21#_c_51_n N_A_83_21#_c_52_n N_A_83_21#_c_59_p N_A_83_21#_c_84_p
+ N_A_83_21#_c_71_p N_A_83_21#_c_60_p N_A_83_21#_c_53_n N_A_83_21#_c_54_n
+ PM_SKY130_FD_SC_HDLL__O22A_1%A_83_21#
x_PM_SKY130_FD_SC_HDLL__O22A_1%B1 N_B1_c_115_n N_B1_M1005_g N_B1_c_116_n
+ N_B1_M1008_g B1 B1 PM_SKY130_FD_SC_HDLL__O22A_1%B1
x_PM_SKY130_FD_SC_HDLL__O22A_1%B2 N_B2_c_144_n N_B2_M1009_g N_B2_c_145_n
+ N_B2_M1003_g B2 PM_SKY130_FD_SC_HDLL__O22A_1%B2
x_PM_SKY130_FD_SC_HDLL__O22A_1%A2 N_A2_c_177_n N_A2_M1000_g N_A2_c_178_n
+ N_A2_M1007_g N_A2_c_179_n A2 PM_SKY130_FD_SC_HDLL__O22A_1%A2
x_PM_SKY130_FD_SC_HDLL__O22A_1%A1 N_A1_c_216_n N_A1_M1004_g N_A1_c_217_n
+ N_A1_M1002_g A1 A1 PM_SKY130_FD_SC_HDLL__O22A_1%A1
x_PM_SKY130_FD_SC_HDLL__O22A_1%X N_X_M1006_s N_X_M1001_s X N_X_c_238_n
+ PM_SKY130_FD_SC_HDLL__O22A_1%X
x_PM_SKY130_FD_SC_HDLL__O22A_1%VPWR N_VPWR_M1001_d N_VPWR_M1002_d N_VPWR_c_253_n
+ N_VPWR_c_254_n N_VPWR_c_255_n VPWR N_VPWR_c_256_n N_VPWR_c_257_n
+ N_VPWR_c_258_n N_VPWR_c_252_n PM_SKY130_FD_SC_HDLL__O22A_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O22A_1%VGND N_VGND_M1006_d N_VGND_M1000_d N_VGND_c_298_n
+ N_VGND_c_299_n N_VGND_c_300_n N_VGND_c_301_n VGND N_VGND_c_302_n
+ N_VGND_c_303_n N_VGND_c_304_n PM_SKY130_FD_SC_HDLL__O22A_1%VGND
x_PM_SKY130_FD_SC_HDLL__O22A_1%A_219_47# N_A_219_47#_M1008_s N_A_219_47#_M1009_d
+ N_A_219_47#_M1004_d N_A_219_47#_c_348_n N_A_219_47#_c_363_n
+ N_A_219_47#_c_355_n N_A_219_47#_c_349_n N_A_219_47#_c_350_n
+ PM_SKY130_FD_SC_HDLL__O22A_1%A_219_47#
cc_1 VNB N_A_83_21#_c_49_n 0.0230702f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_83_21#_c_50_n 0.0298615f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_3 VNB N_A_83_21#_c_51_n 0.00401692f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_4 VNB N_A_83_21#_c_52_n 6.40298e-19 $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=0.805
cc_5 VNB N_A_83_21#_c_53_n 0.00347005f $X=-0.19 $Y=-0.24 $X2=1.64 $Y2=0.73
cc_6 VNB N_A_83_21#_c_54_n 0.00967959f $X=-0.19 $Y=-0.24 $X2=1.44 $Y2=0.77
cc_7 VNB N_B1_c_115_n 0.0228999f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.235
cc_8 VNB N_B1_c_116_n 0.0200261f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB B1 0.00498786f $X=-0.19 $Y=-0.24 $X2=0.697 $Y2=1.16
cc_10 VNB N_B2_c_144_n 0.0178342f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.235
cc_11 VNB N_B2_c_145_n 0.0223375f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB B2 0.00457865f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_13 VNB N_A2_c_177_n 0.0184455f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.235
cc_14 VNB N_A2_c_178_n 0.0205627f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A2_c_179_n 0.00361766f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_16 VNB N_A1_c_216_n 0.0227688f $X=-0.19 $Y=-0.24 $X2=1.505 $Y2=0.235
cc_17 VNB N_A1_c_217_n 0.0281186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB A1 0.0127686f $X=-0.19 $Y=-0.24 $X2=0.697 $Y2=1.16
cc_19 VNB N_X_c_238_n 0.04234f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_20 VNB N_VPWR_c_252_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_298_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_22 VNB N_VGND_c_299_n 0.00468873f $X=-0.19 $Y=-0.24 $X2=0.697 $Y2=1.16
cc_23 VNB N_VGND_c_300_n 0.0449254f $X=-0.19 $Y=-0.24 $X2=1.44 $Y2=0.805
cc_24 VNB N_VGND_c_301_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.86 $Y2=0.805
cc_25 VNB N_VGND_c_302_n 0.0261505f $X=-0.19 $Y=-0.24 $X2=2.04 $Y2=1.6
cc_26 VNB N_VGND_c_303_n 0.212905f $X=-0.19 $Y=-0.24 $X2=2.11 $Y2=1.62
cc_27 VNB N_VGND_c_304_n 0.0225479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_219_47#_c_348_n 0.00250617f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_29 VNB N_A_219_47#_c_349_n 0.00799997f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_30 VNB N_A_219_47#_c_350_n 0.0168702f $X=-0.19 $Y=-0.24 $X2=1.805 $Y2=1.6
cc_31 VPB N_A_83_21#_c_50_n 0.0330877f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_32 VPB N_A_83_21#_c_51_n 0.00225933f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_33 VPB N_B1_c_115_n 0.0278592f $X=-0.19 $Y=1.305 $X2=1.505 $Y2=0.235
cc_34 VPB B1 0.00210698f $X=-0.19 $Y=1.305 $X2=0.697 $Y2=1.16
cc_35 VPB N_B2_c_145_n 0.0261379f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB B2 0.00167528f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.995
cc_37 VPB N_A2_c_178_n 0.0259053f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A2_c_179_n 0.00138015f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_39 VPB A2 0.00151654f $X=-0.19 $Y=1.305 $X2=0.697 $Y2=0.895
cc_40 VPB N_A1_c_217_n 0.0321024f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_X_c_238_n 0.0473448f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_42 VPB N_VPWR_c_253_n 0.0050754f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_43 VPB N_VPWR_c_254_n 0.0159551f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_44 VPB N_VPWR_c_255_n 0.0642572f $X=-0.19 $Y=1.305 $X2=0.697 $Y2=0.895
cc_45 VPB N_VPWR_c_256_n 0.0187803f $X=-0.19 $Y=1.305 $X2=0.86 $Y2=0.805
cc_46 VPB N_VPWR_c_257_n 0.0431545f $X=-0.19 $Y=1.305 $X2=2.11 $Y2=2.3
cc_47 VPB N_VPWR_c_258_n 0.0131648f $X=-0.19 $Y=1.305 $X2=2.04 $Y2=1.6
cc_48 VPB N_VPWR_c_252_n 0.0452896f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 N_A_83_21#_c_50_n N_B1_c_115_n 0.0134394f $X=0.515 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_50 N_A_83_21#_c_51_n N_B1_c_115_n 0.00567225f $X=0.62 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_51 N_A_83_21#_c_59_p N_B1_c_115_n 0.021092f $X=1.805 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_52 N_A_83_21#_c_60_p N_B1_c_115_n 0.00316705f $X=2.11 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_53 N_A_83_21#_c_54_n N_B1_c_115_n 0.00312484f $X=1.44 $Y=0.77 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_83_21#_c_51_n N_B1_c_116_n 0.00260652f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A_83_21#_c_53_n N_B1_c_116_n 0.00623759f $X=1.64 $Y=0.73 $X2=0 $Y2=0
cc_56 N_A_83_21#_c_54_n N_B1_c_116_n 0.00825457f $X=1.44 $Y=0.77 $X2=0 $Y2=0
cc_57 N_A_83_21#_c_50_n B1 8.56035e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_83_21#_c_51_n B1 0.0186525f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_83_21#_c_59_p B1 0.0312297f $X=1.805 $Y=1.6 $X2=0 $Y2=0
cc_60 N_A_83_21#_c_54_n B1 0.0336453f $X=1.44 $Y=0.77 $X2=0 $Y2=0
cc_61 N_A_83_21#_c_53_n N_B2_c_144_n 0.00439747f $X=1.64 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A_83_21#_c_59_p N_B2_c_145_n 0.00400212f $X=1.805 $Y=1.6 $X2=0 $Y2=0
cc_63 N_A_83_21#_c_71_p N_B2_c_145_n 0.00693649f $X=2.04 $Y=1.705 $X2=0 $Y2=0
cc_64 N_A_83_21#_c_60_p N_B2_c_145_n 0.0215465f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_65 N_A_83_21#_c_59_p B2 0.00354041f $X=1.805 $Y=1.6 $X2=0 $Y2=0
cc_66 N_A_83_21#_c_71_p B2 0.0257479f $X=2.04 $Y=1.705 $X2=0 $Y2=0
cc_67 N_A_83_21#_c_53_n B2 0.00551193f $X=1.64 $Y=0.73 $X2=0 $Y2=0
cc_68 N_A_83_21#_c_71_p N_A2_c_178_n 0.00190779f $X=2.04 $Y=1.705 $X2=0 $Y2=0
cc_69 N_A_83_21#_c_60_p N_A2_c_178_n 0.0078776f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_70 N_A_83_21#_c_71_p A2 0.0168645f $X=2.04 $Y=1.705 $X2=0 $Y2=0
cc_71 N_A_83_21#_c_60_p A2 0.0542317f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_72 N_A_83_21#_c_49_n N_X_c_238_n 0.0156626f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_83_21#_c_50_n N_X_c_238_n 0.00858854f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_83_21#_c_51_n N_X_c_238_n 0.0466468f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_83_21#_c_52_n N_X_c_238_n 0.00794913f $X=0.86 $Y=0.805 $X2=0 $Y2=0
cc_76 N_A_83_21#_c_84_p N_X_c_238_n 0.0170997f $X=0.86 $Y=1.6 $X2=0 $Y2=0
cc_77 N_A_83_21#_c_59_p N_VPWR_M1001_d 0.0131637f $X=1.805 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_83_21#_c_84_p N_VPWR_M1001_d 0.00296326f $X=0.86 $Y=1.6 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_83_21#_c_50_n N_VPWR_c_253_n 0.00447425f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_83_21#_c_59_p N_VPWR_c_253_n 0.0361694f $X=1.805 $Y=1.6 $X2=0 $Y2=0
cc_81 N_A_83_21#_c_84_p N_VPWR_c_253_n 0.0178069f $X=0.86 $Y=1.6 $X2=0 $Y2=0
cc_82 N_A_83_21#_c_60_p N_VPWR_c_253_n 0.0220646f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_83 N_A_83_21#_c_50_n N_VPWR_c_256_n 0.00700684f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_83_21#_c_60_p N_VPWR_c_257_n 0.0305511f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_85 N_A_83_21#_M1003_d N_VPWR_c_252_n 0.00679892f $X=1.965 $Y=1.485 $X2=0
+ $Y2=0
cc_86 N_A_83_21#_c_50_n N_VPWR_c_252_n 0.0140041f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_83_21#_c_60_p N_VPWR_c_252_n 0.0172239f $X=2.11 $Y=2.3 $X2=0 $Y2=0
cc_88 N_A_83_21#_c_59_p A_299_297# 0.010182f $X=1.805 $Y=1.6 $X2=-0.19 $Y2=-0.24
cc_89 N_A_83_21#_c_52_n N_VGND_M1006_d 0.00298767f $X=0.86 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_83_21#_c_49_n N_VGND_c_298_n 0.00438629f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_83_21#_c_50_n N_VGND_c_298_n 5.78894e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_83_21#_c_52_n N_VGND_c_298_n 0.0139733f $X=0.86 $Y=0.805 $X2=0 $Y2=0
cc_93 N_A_83_21#_c_52_n N_VGND_c_300_n 0.00125429f $X=0.86 $Y=0.805 $X2=0 $Y2=0
cc_94 N_A_83_21#_c_54_n N_VGND_c_300_n 0.00303519f $X=1.44 $Y=0.77 $X2=0 $Y2=0
cc_95 N_A_83_21#_M1008_d N_VGND_c_303_n 0.00219239f $X=1.505 $Y=0.235 $X2=0
+ $Y2=0
cc_96 N_A_83_21#_c_49_n N_VGND_c_303_n 0.0120328f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_83_21#_c_52_n N_VGND_c_303_n 0.00498677f $X=0.86 $Y=0.805 $X2=0 $Y2=0
cc_98 N_A_83_21#_c_54_n N_VGND_c_303_n 0.00607201f $X=1.44 $Y=0.77 $X2=0 $Y2=0
cc_99 N_A_83_21#_c_49_n N_VGND_c_304_n 0.00555578f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_83_21#_c_52_n N_VGND_c_304_n 8.42882e-19 $X=0.86 $Y=0.805 $X2=0 $Y2=0
cc_101 N_A_83_21#_c_54_n N_A_219_47#_M1008_s 0.0031941f $X=1.44 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_102 N_A_83_21#_M1008_d N_A_219_47#_c_348_n 0.00326408f $X=1.505 $Y=0.235
+ $X2=0 $Y2=0
cc_103 N_A_83_21#_c_53_n N_A_219_47#_c_348_n 0.0173867f $X=1.64 $Y=0.73 $X2=0
+ $Y2=0
cc_104 N_A_83_21#_c_54_n N_A_219_47#_c_348_n 0.0167975f $X=1.44 $Y=0.77 $X2=0
+ $Y2=0
cc_105 N_A_83_21#_c_71_p N_A_219_47#_c_355_n 0.00397424f $X=2.04 $Y=1.705 $X2=0
+ $Y2=0
cc_106 N_A_83_21#_c_53_n N_A_219_47#_c_355_n 0.0133845f $X=1.64 $Y=0.73 $X2=0
+ $Y2=0
cc_107 N_B1_c_116_n N_B2_c_144_n 0.0240908f $X=1.43 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_108 N_B1_c_115_n N_B2_c_145_n 0.0751566f $X=1.405 $Y=1.41 $X2=0 $Y2=0
cc_109 B1 N_B2_c_145_n 8.53413e-19 $X=1.415 $Y=1.19 $X2=0 $Y2=0
cc_110 N_B1_c_115_n B2 8.67257e-19 $X=1.405 $Y=1.41 $X2=0 $Y2=0
cc_111 B1 B2 0.0197812f $X=1.415 $Y=1.19 $X2=0 $Y2=0
cc_112 N_B1_c_115_n N_VPWR_c_253_n 0.0183304f $X=1.405 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_115_n N_VPWR_c_257_n 0.00525069f $X=1.405 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B1_c_115_n N_VPWR_c_252_n 0.00896952f $X=1.405 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B1_c_116_n N_VGND_c_298_n 0.00241512f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_116 N_B1_c_116_n N_VGND_c_300_n 0.00366111f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B1_c_116_n N_VGND_c_303_n 0.0065944f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B1_c_116_n N_A_219_47#_c_348_n 0.00833791f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_119 N_B2_c_144_n N_A2_c_177_n 0.0145313f $X=1.85 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_120 N_B2_c_145_n N_A2_c_178_n 0.03339f $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_121 B2 N_A2_c_178_n 8.83711e-19 $X=1.85 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B2_c_145_n N_A2_c_179_n 7.01707e-19 $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_123 B2 N_A2_c_179_n 0.0203031f $X=1.85 $Y=1.105 $X2=0 $Y2=0
cc_124 N_B2_c_145_n A2 8.46959e-19 $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B2_c_145_n N_VPWR_c_253_n 0.0028413f $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B2_c_145_n N_VPWR_c_257_n 0.00461082f $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_127 N_B2_c_145_n N_VPWR_c_252_n 0.00715067f $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B2_c_144_n N_VGND_c_300_n 0.00366111f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B2_c_144_n N_VGND_c_303_n 0.0057112f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_130 N_B2_c_144_n N_A_219_47#_c_348_n 0.0126817f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B2_c_145_n N_A_219_47#_c_348_n 0.00202776f $X=1.875 $Y=1.41 $X2=0 $Y2=0
cc_132 B2 N_A_219_47#_c_348_n 0.00598879f $X=1.85 $Y=1.105 $X2=0 $Y2=0
cc_133 N_B2_c_144_n N_A_219_47#_c_355_n 0.006589f $X=1.85 $Y=0.995 $X2=0 $Y2=0
cc_134 B2 N_A_219_47#_c_355_n 0.00647116f $X=1.85 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A2_c_177_n N_A1_c_216_n 0.0219414f $X=2.44 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_136 N_A2_c_178_n N_A1_c_217_n 0.0721688f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A2_c_179_n N_A1_c_217_n 0.0036294f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_138 A2 N_A1_c_217_n 0.0081133f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_139 N_A2_c_178_n A1 6.47926e-19 $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A2_c_179_n A1 0.0170239f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A2_c_178_n N_VPWR_c_255_n 0.00228399f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_142 A2 N_VPWR_c_255_n 0.0458233f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_143 N_A2_c_178_n N_VPWR_c_257_n 0.00545889f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_144 A2 N_VPWR_c_257_n 0.00944848f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_145 N_A2_c_178_n N_VPWR_c_252_n 0.00909663f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_146 A2 N_VPWR_c_252_n 0.00762415f $X=2.445 $Y=1.785 $X2=0 $Y2=0
cc_147 A2 A_511_297# 0.0107086f $X=2.445 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_148 N_A2_c_177_n N_VGND_c_299_n 0.00428153f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_177_n N_VGND_c_300_n 0.00420155f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_177_n N_VGND_c_303_n 0.00634859f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A2_c_177_n N_A_219_47#_c_363_n 0.00245595f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A2_c_177_n N_A_219_47#_c_355_n 0.00467302f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A2_c_179_n N_A_219_47#_c_355_n 0.00293259f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_154 N_A2_c_177_n N_A_219_47#_c_349_n 0.00885861f $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A2_c_178_n N_A_219_47#_c_349_n 0.00289163f $X=2.465 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A2_c_179_n N_A_219_47#_c_349_n 0.0157304f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A2_c_177_n N_A_219_47#_c_350_n 5.10857e-19 $X=2.44 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A1_c_217_n N_VPWR_c_255_n 0.0278025f $X=2.945 $Y=1.41 $X2=0 $Y2=0
cc_159 A1 N_VPWR_c_255_n 0.0257682f $X=3.085 $Y=1.19 $X2=0 $Y2=0
cc_160 N_A1_c_217_n N_VPWR_c_257_n 0.00505556f $X=2.945 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A1_c_217_n N_VPWR_c_252_n 0.00868699f $X=2.945 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A1_c_216_n N_VGND_c_299_n 0.00277568f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_216_n N_VGND_c_302_n 0.00421028f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A1_c_216_n N_VGND_c_303_n 0.00696607f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A1_c_216_n N_A_219_47#_c_355_n 4.66393e-19 $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_216_n N_A_219_47#_c_349_n 0.00977838f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_217_n N_A_219_47#_c_349_n 0.00345407f $X=2.945 $Y=1.41 $X2=0 $Y2=0
cc_168 A1 N_A_219_47#_c_349_n 0.0288039f $X=3.085 $Y=1.19 $X2=0 $Y2=0
cc_169 N_A1_c_216_n N_A_219_47#_c_350_n 0.00601017f $X=2.92 $Y=0.995 $X2=0 $Y2=0
cc_170 N_X_c_238_n N_VPWR_c_253_n 0.0394127f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_171 N_X_c_238_n N_VPWR_c_256_n 0.0196165f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_172 N_X_M1001_s N_VPWR_c_252_n 0.00442207f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_173 N_X_c_238_n N_VPWR_c_252_n 0.0107063f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_174 N_X_M1006_s N_VGND_c_303_n 0.00414151f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_175 N_X_c_238_n N_VGND_c_303_n 0.0100809f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_176 N_X_c_238_n N_VGND_c_304_n 0.01133f $X=0.26 $Y=0.595 $X2=0 $Y2=0
cc_177 N_VPWR_c_252_n A_299_297# 0.0123962f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_178 N_VPWR_c_252_n A_511_297# 0.00905777f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_179 N_VPWR_c_255_n N_A_219_47#_c_349_n 0.00174633f $X=3.18 $Y=1.66 $X2=0
+ $Y2=0
cc_180 N_VGND_c_303_n N_A_219_47#_M1008_s 0.00211652f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_181 N_VGND_c_303_n N_A_219_47#_M1009_d 0.0035771f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_182 N_VGND_c_303_n N_A_219_47#_M1004_d 0.00251629f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_183 N_VGND_c_298_n N_A_219_47#_c_348_n 0.0106215f $X=0.7 $Y=0.38 $X2=0 $Y2=0
cc_184 N_VGND_c_300_n N_A_219_47#_c_348_n 0.0456961f $X=2.625 $Y=0 $X2=0 $Y2=0
cc_185 N_VGND_c_303_n N_A_219_47#_c_348_n 0.0352856f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_186 N_VGND_c_299_n N_A_219_47#_c_363_n 0.0111926f $X=2.71 $Y=0.36 $X2=0 $Y2=0
cc_187 N_VGND_c_300_n N_A_219_47#_c_363_n 0.0166263f $X=2.625 $Y=0 $X2=0 $Y2=0
cc_188 N_VGND_c_303_n N_A_219_47#_c_363_n 0.0121819f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_189 N_VGND_c_299_n N_A_219_47#_c_355_n 0.00289632f $X=2.71 $Y=0.36 $X2=0
+ $Y2=0
cc_190 N_VGND_M1000_d N_A_219_47#_c_349_n 0.00829366f $X=2.515 $Y=0.235 $X2=0
+ $Y2=0
cc_191 N_VGND_c_299_n N_A_219_47#_c_349_n 0.0125799f $X=2.71 $Y=0.36 $X2=0 $Y2=0
cc_192 N_VGND_c_300_n N_A_219_47#_c_349_n 0.0029937f $X=2.625 $Y=0 $X2=0 $Y2=0
cc_193 N_VGND_c_302_n N_A_219_47#_c_349_n 0.00211912f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_194 N_VGND_c_303_n N_A_219_47#_c_349_n 0.0102404f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_195 N_VGND_c_302_n N_A_219_47#_c_350_n 0.021576f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_196 N_VGND_c_303_n N_A_219_47#_c_350_n 0.0144931f $X=3.45 $Y=0 $X2=0 $Y2=0
