* File: sky130_fd_sc_hdll__einvn_8.pex.spice
* Created: Wed Sep  2 08:31:26 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%TE_B 1 3 4 6 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 27 29 31 32 34 36 37 39 41 42 44 46 47 50 51 52 53 54 55 56
c137 55 0 7.37965e-20 $X=3.84 $Y=1.395
c138 54 0 7.37964e-20 $X=3.37 $Y=1.395
c139 53 0 7.37965e-20 $X=2.9 $Y=1.395
c140 52 0 7.37964e-20 $X=2.43 $Y=1.395
c141 51 0 7.37965e-20 $X=1.96 $Y=1.395
c142 50 0 7.37964e-20 $X=1.49 $Y=1.395
c143 42 0 2.16486e-19 $X=4.22 $Y=1.395
c144 37 0 1.65302e-19 $X=3.75 $Y=1.395
c145 32 0 1.64536e-19 $X=3.28 $Y=1.395
c146 27 0 1.65302e-19 $X=2.81 $Y=1.395
c147 22 0 1.64536e-19 $X=2.34 $Y=1.395
c148 17 0 1.78583e-19 $X=1.87 $Y=1.395
c149 1 0 1.15275e-19 $X=0.495 $Y=1.41
r150 61 62 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r151 59 61 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.495 $Y2=1.202
r152 56 59 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r153 47 49 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=1.02 $Y=1.25
+ $X2=1.02 $Y2=1.395
r154 44 46 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=4.31 $Y=1.47
+ $X2=4.31 $Y2=2.015
r155 43 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.93 $Y=1.395
+ $X2=3.84 $Y2=1.395
r156 42 44 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.22 $Y=1.395
+ $X2=4.31 $Y2=1.47
r157 42 43 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.22 $Y=1.395
+ $X2=3.93 $Y2=1.395
r158 39 55 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.84 $Y=1.47
+ $X2=3.84 $Y2=1.395
r159 39 41 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.84 $Y=1.47
+ $X2=3.84 $Y2=2.015
r160 38 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.46 $Y=1.395
+ $X2=3.37 $Y2=1.395
r161 37 55 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.75 $Y=1.395
+ $X2=3.84 $Y2=1.395
r162 37 38 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.75 $Y=1.395
+ $X2=3.46 $Y2=1.395
r163 34 54 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.37 $Y=1.47
+ $X2=3.37 $Y2=1.395
r164 34 36 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.37 $Y=1.47
+ $X2=3.37 $Y2=2.015
r165 33 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.99 $Y=1.395 $X2=2.9
+ $Y2=1.395
r166 32 54 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.28 $Y=1.395
+ $X2=3.37 $Y2=1.395
r167 32 33 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.28 $Y=1.395
+ $X2=2.99 $Y2=1.395
r168 29 53 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.9 $Y=1.47 $X2=2.9
+ $Y2=1.395
r169 29 31 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.9 $Y=1.47
+ $X2=2.9 $Y2=2.015
r170 28 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.52 $Y=1.395
+ $X2=2.43 $Y2=1.395
r171 27 53 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.81 $Y=1.395 $X2=2.9
+ $Y2=1.395
r172 27 28 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.81 $Y=1.395
+ $X2=2.52 $Y2=1.395
r173 24 52 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.43 $Y=1.47
+ $X2=2.43 $Y2=1.395
r174 24 26 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.43 $Y=1.47
+ $X2=2.43 $Y2=2.015
r175 23 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.05 $Y=1.395
+ $X2=1.96 $Y2=1.395
r176 22 52 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.34 $Y=1.395
+ $X2=2.43 $Y2=1.395
r177 22 23 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.34 $Y=1.395
+ $X2=2.05 $Y2=1.395
r178 19 51 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=1.47
+ $X2=1.96 $Y2=1.395
r179 19 21 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.96 $Y=1.47
+ $X2=1.96 $Y2=2.015
r180 18 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.58 $Y=1.395
+ $X2=1.49 $Y2=1.395
r181 17 51 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.87 $Y=1.395
+ $X2=1.96 $Y2=1.395
r182 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=1.395
+ $X2=1.58 $Y2=1.395
r183 14 50 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.49 $Y=1.47
+ $X2=1.49 $Y2=1.395
r184 14 16 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.49 $Y=1.47
+ $X2=1.49 $Y2=2.015
r185 13 49 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.12 $Y=1.395
+ $X2=1.02 $Y2=1.395
r186 12 50 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.4 $Y=1.395 $X2=1.49
+ $Y2=1.395
r187 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.4 $Y=1.395
+ $X2=1.12 $Y2=1.395
r188 9 49 25.676 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.47 $X2=1.02
+ $Y2=1.395
r189 9 11 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.02 $Y=1.47
+ $X2=1.02 $Y2=2.015
r190 8 62 27.0958 $w=3.65e-07 $l=9.60469e-08 $layer=POLY_cond $X=0.595 $Y=1.25
+ $X2=0.52 $Y2=1.202
r191 7 47 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.92 $Y=1.25 $X2=1.02
+ $Y2=1.25
r192 7 8 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.92 $Y=1.25
+ $X2=0.595 $Y2=1.25
r193 4 62 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r194 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r195 1 61 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r196 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 27 29 30 32 34 35 37 39 42 44 45 46 47 48 49 50 51 54 56 60 65
c157 49 0 1.07001e-19 $X=3.91 $Y=1.035
c158 47 0 1.07001e-19 $X=2.97 $Y=1.035
c159 45 0 1.07001e-19 $X=2.03 $Y=1.035
c160 42 0 7.54923e-20 $X=4.865 $Y=0.96
c161 35 0 3.79794e-19 $X=4.305 $Y=1.035
c162 30 0 1.17964e-19 $X=3.835 $Y=1.035
c163 25 0 3.79794e-19 $X=3.365 $Y=1.035
c164 20 0 1.17964e-19 $X=2.895 $Y=1.035
c165 15 0 3.79794e-19 $X=2.425 $Y=1.035
c166 10 0 1.17964e-19 $X=1.955 $Y=1.035
r167 61 65 41.9243 $w=3.65e-07 $l=1.35e-07 $layer=POLY_cond $X=4.755 $Y=1.142
+ $X2=4.62 $Y2=1.142
r168 60 61 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.16 $X2=4.755 $Y2=1.16
r169 58 63 3.43149 $w=3.3e-07 $l=3.8e-07 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=0.515 $Y2=1.16
r170 58 60 134.801 $w=3.28e-07 $l=3.86e-06 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=4.755 $Y2=1.16
r171 54 63 14.9901 $w=5.23e-07 $l=6.36801e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.515 $Y2=1.16
r172 54 56 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.815
r173 51 63 14.9901 $w=5.23e-07 $l=6.36801e-07 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.515 $Y2=1.16
r174 51 53 4.5451 $w=2.55e-07 $l=9.5e-08 $layer=LI1_cond $X=0.217 $Y=0.655
+ $X2=0.217 $Y2=0.56
r175 42 61 17.3903 $w=3.65e-07 $l=1.1e-07 $layer=POLY_cond $X=4.865 $Y=1.142
+ $X2=4.755 $Y2=1.142
r176 42 44 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.865 $Y=0.96
+ $X2=4.865 $Y2=0.56
r177 41 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.455 $Y=1.035
+ $X2=4.38 $Y2=1.035
r178 41 65 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=1.035
+ $X2=4.62 $Y2=1.035
r179 37 50 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.38 $Y=0.96
+ $X2=4.38 $Y2=1.035
r180 37 39 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=4.38 $Y=0.96 $X2=4.38
+ $Y2=0.56
r181 36 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.985 $Y=1.035
+ $X2=3.91 $Y2=1.035
r182 35 50 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.305 $Y=1.035
+ $X2=4.38 $Y2=1.035
r183 35 36 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.305 $Y=1.035
+ $X2=3.985 $Y2=1.035
r184 32 49 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.91 $Y=0.96
+ $X2=3.91 $Y2=1.035
r185 32 34 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.91 $Y=0.96 $X2=3.91
+ $Y2=0.56
r186 31 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.515 $Y=1.035
+ $X2=3.44 $Y2=1.035
r187 30 49 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.835 $Y=1.035
+ $X2=3.91 $Y2=1.035
r188 30 31 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.835 $Y=1.035
+ $X2=3.515 $Y2=1.035
r189 27 48 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.44 $Y=0.96
+ $X2=3.44 $Y2=1.035
r190 27 29 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=3.44 $Y=0.96 $X2=3.44
+ $Y2=0.56
r191 26 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.045 $Y=1.035
+ $X2=2.97 $Y2=1.035
r192 25 48 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.365 $Y=1.035
+ $X2=3.44 $Y2=1.035
r193 25 26 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=3.365 $Y=1.035
+ $X2=3.045 $Y2=1.035
r194 22 47 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.97 $Y=0.96
+ $X2=2.97 $Y2=1.035
r195 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.97 $Y=0.96 $X2=2.97
+ $Y2=0.56
r196 21 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.575 $Y=1.035
+ $X2=2.5 $Y2=1.035
r197 20 47 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=2.97 $Y2=1.035
r198 20 21 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.895 $Y=1.035
+ $X2=2.575 $Y2=1.035
r199 17 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.5 $Y=0.96 $X2=2.5
+ $Y2=1.035
r200 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.5 $Y=0.96 $X2=2.5
+ $Y2=0.56
r201 16 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.105 $Y=1.035
+ $X2=2.03 $Y2=1.035
r202 15 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.425 $Y=1.035
+ $X2=2.5 $Y2=1.035
r203 15 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=1.035
+ $X2=2.105 $Y2=1.035
r204 12 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.03 $Y=0.96
+ $X2=2.03 $Y2=1.035
r205 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.03 $Y=0.96 $X2=2.03
+ $Y2=0.56
r206 10 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=1.035
+ $X2=2.03 $Y2=1.035
r207 10 11 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=1.955 $Y=1.035
+ $X2=1.585 $Y2=1.035
r208 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.51 $Y=0.96
+ $X2=1.585 $Y2=1.035
r209 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.51 $Y=0.96 $X2=1.51
+ $Y2=0.56
r210 2 56 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
r211 1 53 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 50 51 52 53 54 55 56 85
+ 88 93 96 99 102 105 108 111
r135 85 86 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.64 $Y=1.202
+ $X2=8.665 $Y2=1.202
r136 83 85 20.3016 $w=3.68e-07 $l=1.55e-07 $layer=POLY_cond $X=8.485 $Y=1.202
+ $X2=8.64 $Y2=1.202
r137 81 83 41.2582 $w=3.68e-07 $l=3.15e-07 $layer=POLY_cond $X=8.17 $Y=1.202
+ $X2=8.485 $Y2=1.202
r138 80 81 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.145 $Y=1.202
+ $X2=8.17 $Y2=1.202
r139 79 80 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=7.7 $Y=1.202
+ $X2=8.145 $Y2=1.202
r140 78 79 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.675 $Y=1.202
+ $X2=7.7 $Y2=1.202
r141 77 78 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=7.23 $Y=1.202
+ $X2=7.675 $Y2=1.202
r142 76 77 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.205 $Y=1.202
+ $X2=7.23 $Y2=1.202
r143 75 76 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=6.76 $Y=1.202
+ $X2=7.205 $Y2=1.202
r144 74 75 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.735 $Y=1.202
+ $X2=6.76 $Y2=1.202
r145 73 74 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=6.29 $Y=1.202
+ $X2=6.735 $Y2=1.202
r146 72 73 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.265 $Y=1.202
+ $X2=6.29 $Y2=1.202
r147 71 72 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=5.82 $Y=1.202
+ $X2=6.265 $Y2=1.202
r148 70 71 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.795 $Y=1.202
+ $X2=5.82 $Y2=1.202
r149 68 70 49.7717 $w=3.68e-07 $l=3.8e-07 $layer=POLY_cond $X=5.415 $Y=1.202
+ $X2=5.795 $Y2=1.202
r150 66 68 8.51359 $w=3.68e-07 $l=6.5e-08 $layer=POLY_cond $X=5.35 $Y=1.202
+ $X2=5.415 $Y2=1.202
r151 65 66 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.325 $Y=1.202
+ $X2=5.35 $Y2=1.202
r152 56 111 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=8.485 $Y=1.14
+ $X2=8.525 $Y2=1.14
r153 56 108 16.6906 $w=2.88e-07 $l=4.2e-07 $layer=LI1_cond $X=8.485 $Y=1.14
+ $X2=8.065 $Y2=1.14
r154 56 83 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=8.485
+ $Y=1.16 $X2=8.485 $Y2=1.16
r155 55 108 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=8.05 $Y=1.14
+ $X2=8.065 $Y2=1.14
r156 55 105 18.0814 $w=2.88e-07 $l=4.55e-07 $layer=LI1_cond $X=8.05 $Y=1.14
+ $X2=7.595 $Y2=1.14
r157 54 105 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=7.58 $Y=1.14
+ $X2=7.595 $Y2=1.14
r158 54 102 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=7.58 $Y=1.14
+ $X2=7.135 $Y2=1.14
r159 53 102 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=7.115 $Y=1.14
+ $X2=7.135 $Y2=1.14
r160 53 99 17.4853 $w=2.88e-07 $l=4.4e-07 $layer=LI1_cond $X=7.115 $Y=1.14
+ $X2=6.675 $Y2=1.14
r161 52 99 0.397394 $w=2.88e-07 $l=1e-08 $layer=LI1_cond $X=6.665 $Y=1.14
+ $X2=6.675 $Y2=1.14
r162 52 96 17.8827 $w=2.88e-07 $l=4.5e-07 $layer=LI1_cond $X=6.665 $Y=1.14
+ $X2=6.215 $Y2=1.14
r163 51 96 0.596091 $w=2.88e-07 $l=1.5e-08 $layer=LI1_cond $X=6.2 $Y=1.14
+ $X2=6.215 $Y2=1.14
r164 51 93 17.684 $w=2.88e-07 $l=4.45e-07 $layer=LI1_cond $X=6.2 $Y=1.14
+ $X2=5.755 $Y2=1.14
r165 50 93 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=5.75 $Y=1.14
+ $X2=5.755 $Y2=1.14
r166 49 50 16.4919 $w=2.88e-07 $l=4.15e-07 $layer=LI1_cond $X=5.335 $Y=1.14
+ $X2=5.75 $Y2=1.14
r167 49 88 1.58958 $w=2.88e-07 $l=4e-08 $layer=LI1_cond $X=5.335 $Y=1.14
+ $X2=5.295 $Y2=1.14
r168 49 68 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=5.415
+ $Y=1.16 $X2=5.415 $Y2=1.16
r169 46 86 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.665 $Y=0.995
+ $X2=8.665 $Y2=1.202
r170 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.665 $Y=0.995
+ $X2=8.665 $Y2=0.56
r171 43 85 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.64 $Y=1.41
+ $X2=8.64 $Y2=1.202
r172 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.64 $Y=1.41
+ $X2=8.64 $Y2=1.985
r173 40 81 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.17 $Y=1.41
+ $X2=8.17 $Y2=1.202
r174 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.17 $Y=1.41
+ $X2=8.17 $Y2=1.985
r175 37 80 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.145 $Y=0.995
+ $X2=8.145 $Y2=1.202
r176 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.145 $Y=0.995
+ $X2=8.145 $Y2=0.56
r177 34 79 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.7 $Y=1.41 $X2=7.7
+ $Y2=1.202
r178 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.7 $Y=1.41
+ $X2=7.7 $Y2=1.985
r179 31 78 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.675 $Y=0.995
+ $X2=7.675 $Y2=1.202
r180 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.675 $Y=0.995
+ $X2=7.675 $Y2=0.56
r181 28 77 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.23 $Y=1.41
+ $X2=7.23 $Y2=1.202
r182 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.23 $Y=1.41
+ $X2=7.23 $Y2=1.985
r183 25 76 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.205 $Y=0.995
+ $X2=7.205 $Y2=1.202
r184 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.205 $Y=0.995
+ $X2=7.205 $Y2=0.56
r185 22 75 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.76 $Y=1.41
+ $X2=6.76 $Y2=1.202
r186 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.76 $Y=1.41
+ $X2=6.76 $Y2=1.985
r187 19 74 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.735 $Y=0.995
+ $X2=6.735 $Y2=1.202
r188 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.735 $Y=0.995
+ $X2=6.735 $Y2=0.56
r189 16 73 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.202
r190 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.985
r191 13 72 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.265 $Y=0.995
+ $X2=6.265 $Y2=1.202
r192 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.265 $Y=0.995
+ $X2=6.265 $Y2=0.56
r193 10 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.202
r194 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.985
r195 7 70 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=1.202
r196 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.795 $Y=0.995
+ $X2=5.795 $Y2=0.56
r197 4 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.202
r198 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.985
r199 1 65 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.325 $Y=0.995
+ $X2=5.325 $Y2=1.202
r200 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.325 $Y=0.995
+ $X2=5.325 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%VPWR 1 2 3 4 5 18 22 24 28 30 34 36 40 42
+ 44 49 59 60 63 66 69 72 75
r130 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r132 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r134 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r135 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 59 60 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r139 57 60 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=8.97 $Y2=2.72
r140 57 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 56 59 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=8.97 $Y2=2.72
r142 56 57 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r143 54 75 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.73 $Y=2.72 $X2=4.53
+ $Y2=2.72
r144 54 56 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.73 $Y=2.72 $X2=4.83
+ $Y2=2.72
r145 53 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r146 53 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r147 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r148 50 63 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r149 50 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r150 49 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=2.72 $X2=1.7
+ $Y2=2.72
r151 49 52 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r152 44 63 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r153 44 46 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r154 42 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r155 42 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r156 38 75 1.46811 $w=4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.53 $Y=2.635 $X2=4.53
+ $Y2=2.72
r157 38 40 18.295 $w=3.98e-07 $l=6.35e-07 $layer=LI1_cond $X=4.53 $Y=2.635
+ $X2=4.53 $Y2=2
r158 37 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.77 $Y=2.72
+ $X2=3.58 $Y2=2.72
r159 36 75 9.81116 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=4.33 $Y=2.72 $X2=4.53
+ $Y2=2.72
r160 36 37 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.33 $Y=2.72
+ $X2=3.77 $Y2=2.72
r161 32 72 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.58 $Y=2.635
+ $X2=3.58 $Y2=2.72
r162 32 34 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=3.58 $Y=2.635
+ $X2=3.58 $Y2=2.02
r163 31 69 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=2.64 $Y2=2.72
r164 30 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=3.58 $Y2=2.72
r165 30 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=2.83 $Y2=2.72
r166 26 69 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=2.635
+ $X2=2.64 $Y2=2.72
r167 26 28 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=2.64 $Y=2.635
+ $X2=2.64 $Y2=2.02
r168 25 66 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=2.72 $X2=1.7
+ $Y2=2.72
r169 24 69 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=2.64 $Y2=2.72
r170 24 25 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=1.89 $Y2=2.72
r171 20 66 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.635 $X2=1.7
+ $Y2=2.72
r172 20 22 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=1.7 $Y=2.635
+ $X2=1.7 $Y2=2.02
r173 16 63 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r174 16 18 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.02
r175 5 40 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=1.545 $X2=4.545 $Y2=2
r176 4 34 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.46
+ $Y=1.545 $X2=3.605 $Y2=2.02
r177 3 28 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=1.545 $X2=2.665 $Y2=2.02
r178 2 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.545 $X2=1.725 $Y2=2.02
r179 1 18 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%A_222_309# 1 2 3 4 5 6 7 8 9 30 32 33 36
+ 38 42 44 48 50 55 56 57 60 62 66 68 72 74 78 80 81 82 83 84 85
c149 82 0 1.83107e-19 $X=4.075 $Y=1.58
c150 81 0 1.83107e-19 $X=3.135 $Y=1.58
c151 80 0 1.83107e-19 $X=2.195 $Y=1.58
c152 44 0 2.24965e-19 $X=3.99 $Y=1.58
c153 38 0 2.24965e-19 $X=3.05 $Y=1.58
c154 33 0 1.15275e-19 $X=1.34 $Y=1.58
c155 32 0 2.24965e-19 $X=2.11 $Y=1.58
r156 76 78 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.942 $Y=2.295
+ $X2=8.942 $Y2=1.96
r157 75 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.02 $Y=2.38
+ $X2=7.935 $Y2=2.38
r158 74 76 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=8.79 $Y=2.38
+ $X2=8.942 $Y2=2.295
r159 74 75 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.79 $Y=2.38
+ $X2=8.02 $Y2=2.38
r160 70 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=7.935 $Y2=2.38
r161 70 72 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=7.935 $Y=2.295
+ $X2=7.935 $Y2=1.96
r162 69 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.08 $Y=2.38
+ $X2=6.995 $Y2=2.38
r163 68 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.85 $Y=2.38
+ $X2=7.935 $Y2=2.38
r164 68 69 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=7.85 $Y=2.38
+ $X2=7.08 $Y2=2.38
r165 64 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.995 $Y=2.295
+ $X2=6.995 $Y2=2.38
r166 64 66 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.995 $Y=2.295
+ $X2=6.995 $Y2=1.96
r167 63 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.14 $Y=2.38
+ $X2=6.055 $Y2=2.38
r168 62 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=2.38
+ $X2=6.995 $Y2=2.38
r169 62 63 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=6.91 $Y=2.38
+ $X2=6.14 $Y2=2.38
r170 58 83 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.295
+ $X2=6.055 $Y2=2.38
r171 58 60 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.055 $Y=2.295
+ $X2=6.055 $Y2=1.96
r172 56 83 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.97 $Y=2.38
+ $X2=6.055 $Y2=2.38
r173 56 57 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.97 $Y=2.38
+ $X2=5.2 $Y2=2.38
r174 53 57 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.075 $Y=2.295
+ $X2=5.2 $Y2=2.38
r175 53 55 22.1269 $w=2.48e-07 $l=4.8e-07 $layer=LI1_cond $X=5.075 $Y=2.295
+ $X2=5.075 $Y2=1.815
r176 52 55 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.075 $Y=1.665
+ $X2=5.075 $Y2=1.815
r177 51 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.16 $Y=1.58
+ $X2=4.075 $Y2=1.58
r178 50 52 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.95 $Y=1.58
+ $X2=5.075 $Y2=1.665
r179 50 51 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.95 $Y=1.58
+ $X2=4.16 $Y2=1.58
r180 46 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=1.665
+ $X2=4.075 $Y2=1.58
r181 46 48 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=4.075 $Y=1.665
+ $X2=4.075 $Y2=1.815
r182 45 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=1.58
+ $X2=3.135 $Y2=1.58
r183 44 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.58
+ $X2=4.075 $Y2=1.58
r184 44 45 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.99 $Y=1.58
+ $X2=3.22 $Y2=1.58
r185 40 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.135 $Y=1.665
+ $X2=3.135 $Y2=1.58
r186 40 42 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.135 $Y=1.665
+ $X2=3.135 $Y2=1.815
r187 39 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=1.58
+ $X2=2.195 $Y2=1.58
r188 38 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.05 $Y=1.58
+ $X2=3.135 $Y2=1.58
r189 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.05 $Y=1.58
+ $X2=2.28 $Y2=1.58
r190 34 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.58
r191 34 36 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.815
r192 32 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=1.58
+ $X2=2.195 $Y2=1.58
r193 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.11 $Y=1.58
+ $X2=1.34 $Y2=1.58
r194 28 33 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=1.202 $Y=1.665
+ $X2=1.34 $Y2=1.58
r195 28 30 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=1.202 $Y=1.665
+ $X2=1.202 $Y2=1.815
r196 9 78 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.73
+ $Y=1.485 $X2=8.875 $Y2=1.96
r197 8 72 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.79
+ $Y=1.485 $X2=7.935 $Y2=1.96
r198 7 66 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.85
+ $Y=1.485 $X2=6.995 $Y2=1.96
r199 6 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.485 $X2=6.055 $Y2=1.96
r200 5 55 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=4.99
+ $Y=1.485 $X2=5.115 $Y2=1.815
r201 4 48 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.93
+ $Y=1.545 $X2=4.075 $Y2=1.815
r202 3 42 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.99
+ $Y=1.545 $X2=3.135 $Y2=1.815
r203 2 36 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.545 $X2=2.195 $Y2=1.815
r204 1 30 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.545 $X2=1.255 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%Z 1 2 3 4 5 6 7 8 27 29 30 33 35 37 39 41
+ 43 45 47 48 49 50 58 63 67 69
c122 49 0 7.54923e-20 $X=8.87 $Y=0.765
r123 80 82 50.8559 $w=2.03e-07 $l=9.4e-07 $layer=LI1_cond $X=7.465 $Y=0.722
+ $X2=8.405 $Y2=0.722
r124 78 80 50.8559 $w=2.03e-07 $l=9.4e-07 $layer=LI1_cond $X=6.525 $Y=0.722
+ $X2=7.465 $Y2=0.722
r125 75 78 50.8559 $w=2.03e-07 $l=9.4e-07 $layer=LI1_cond $X=5.585 $Y=0.722
+ $X2=6.525 $Y2=0.722
r126 67 69 1.28049 $w=2.23e-07 $l=2.5e-08 $layer=LI1_cond $X=8.982 $Y=0.825
+ $X2=8.982 $Y2=0.85
r127 49 67 3.27477 $w=2.25e-07 $l=1.03e-07 $layer=LI1_cond $X=8.982 $Y=0.722
+ $X2=8.982 $Y2=0.825
r128 49 82 20.843 $w=2.63e-07 $l=4.65e-07 $layer=LI1_cond $X=8.87 $Y=0.722
+ $X2=8.405 $Y2=0.722
r129 49 50 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=8.982 $Y=0.88
+ $X2=8.982 $Y2=1.19
r130 49 69 1.53659 $w=2.23e-07 $l=3e-08 $layer=LI1_cond $X=8.982 $Y=0.88
+ $X2=8.982 $Y2=0.85
r131 48 63 5.15567 $w=3.78e-07 $l=1.7e-07 $layer=LI1_cond $X=8.38 $Y=1.87
+ $X2=8.38 $Y2=1.7
r132 47 58 5.15567 $w=3.78e-07 $l=1.7e-07 $layer=LI1_cond $X=7.44 $Y=1.87
+ $X2=7.44 $Y2=1.7
r133 46 50 13.5732 $w=2.23e-07 $l=2.65e-07 $layer=LI1_cond $X=8.982 $Y=1.455
+ $X2=8.982 $Y2=1.19
r134 44 63 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=8.38 $Y=1.625
+ $X2=8.38 $Y2=1.7
r135 44 45 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.38 $Y=1.625
+ $X2=8.38 $Y2=1.54
r136 42 58 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=7.44 $Y=1.625
+ $X2=7.44 $Y2=1.7
r137 42 43 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.44 $Y=1.625
+ $X2=7.44 $Y2=1.54
r138 40 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.57 $Y=1.54
+ $X2=8.38 $Y2=1.54
r139 39 46 6.9898 $w=1.7e-07 $l=1.4854e-07 $layer=LI1_cond $X=8.87 $Y=1.54
+ $X2=8.982 $Y2=1.455
r140 39 40 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.87 $Y=1.54 $X2=8.57
+ $Y2=1.54
r141 38 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.63 $Y=1.54
+ $X2=7.44 $Y2=1.54
r142 37 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.19 $Y=1.54
+ $X2=8.38 $Y2=1.54
r143 37 38 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.19 $Y=1.54
+ $X2=7.63 $Y2=1.54
r144 36 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.69 $Y=1.54 $X2=6.5
+ $Y2=1.54
r145 35 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.25 $Y=1.54
+ $X2=7.44 $Y2=1.54
r146 35 36 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.25 $Y=1.54
+ $X2=6.69 $Y2=1.54
r147 31 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.5 $Y=1.625 $X2=6.5
+ $Y2=1.54
r148 31 33 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=6.5 $Y=1.625
+ $X2=6.5 $Y2=1.7
r149 29 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.31 $Y=1.54 $X2=6.5
+ $Y2=1.54
r150 29 30 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.31 $Y=1.54
+ $X2=5.75 $Y2=1.54
r151 25 30 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=5.56 $Y=1.625
+ $X2=5.75 $Y2=1.54
r152 25 27 2.27456 $w=3.78e-07 $l=7.5e-08 $layer=LI1_cond $X=5.56 $Y=1.625
+ $X2=5.56 $Y2=1.7
r153 8 63 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=8.26
+ $Y=1.485 $X2=8.405 $Y2=1.7
r154 7 58 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=7.32
+ $Y=1.485 $X2=7.465 $Y2=1.7
r155 6 33 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=6.38
+ $Y=1.485 $X2=6.525 $Y2=1.7
r156 5 27 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.485 $X2=5.585 $Y2=1.7
r157 4 82 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=8.22
+ $Y=0.235 $X2=8.405 $Y2=0.74
r158 3 80 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=7.28
+ $Y=0.235 $X2=7.465 $Y2=0.74
r159 2 78 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=6.34
+ $Y=0.235 $X2=6.525 $Y2=0.74
r160 1 75 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=5.4
+ $Y=0.235 $X2=5.585 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%VGND 1 2 3 4 5 18 20 24 28 32 36 39 40 42
+ 43 45 46 47 49 68 69 72 75
r122 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r123 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r124 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r125 68 69 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r126 66 69 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=8.97
+ $Y2=0
r127 65 68 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=8.97
+ $Y2=0
r128 65 66 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r129 63 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r130 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r131 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r132 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r133 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r134 57 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r135 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r136 54 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.77
+ $Y2=0
r137 54 56 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.935 $Y=0
+ $X2=2.53 $Y2=0
r138 49 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r139 49 51 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r140 47 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r141 47 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r142 45 62 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.37
+ $Y2=0
r143 45 46 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.595
+ $Y2=0
r144 44 65 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.83
+ $Y2=0
r145 44 46 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.765 $Y=0 $X2=4.595
+ $Y2=0
r146 42 59 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.45
+ $Y2=0
r147 42 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.65
+ $Y2=0
r148 41 62 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.815 $Y=0
+ $X2=4.37 $Y2=0
r149 41 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=0 $X2=3.65
+ $Y2=0
r150 39 56 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r151 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.71
+ $Y2=0
r152 38 59 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.875 $Y=0
+ $X2=3.45 $Y2=0
r153 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.71
+ $Y2=0
r154 34 46 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=0.085
+ $X2=4.595 $Y2=0
r155 34 36 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=4.595 $Y=0.085
+ $X2=4.595 $Y2=0.36
r156 30 43 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.65 $Y=0.085
+ $X2=3.65 $Y2=0
r157 30 32 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.65 $Y=0.085
+ $X2=3.65 $Y2=0.36
r158 26 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0
r159 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0.36
r160 22 75 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0
r161 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0.36
r162 21 72 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r163 20 75 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.77
+ $Y2=0
r164 20 21 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.895 $Y2=0
r165 16 72 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r166 16 18 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.38
r167 5 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.235 $X2=4.59 $Y2=0.36
r168 4 32 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.36
r169 3 28 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.235 $X2=2.71 $Y2=0.36
r170 2 24 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.77 $Y2=0.36
r171 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_8%A_235_47# 1 2 3 4 5 6 7 8 9 28 31 32 33 36
+ 38 41 43 46 52 60 62 63 64
c102 64 0 9.85391e-20 $X=4.12 $Y=0.74
c103 63 0 9.85391e-20 $X=3.18 $Y=0.74
c104 62 0 9.85391e-20 $X=2.24 $Y=0.74
c105 46 0 3.14634e-19 $X=4.985 $Y=0.74
c106 41 0 5.75579e-19 $X=4.035 $Y=0.74
c107 36 0 5.75579e-19 $X=3.095 $Y=0.74
c108 31 0 3.26175e-19 $X=2.155 $Y=0.74
r109 58 60 53.4639 $w=1.93e-07 $l=9.4e-07 $layer=LI1_cond $X=7.935 $Y=0.352
+ $X2=8.875 $Y2=0.352
r110 56 58 53.4639 $w=1.93e-07 $l=9.4e-07 $layer=LI1_cond $X=6.995 $Y=0.352
+ $X2=7.935 $Y2=0.352
r111 54 56 53.4639 $w=1.93e-07 $l=9.4e-07 $layer=LI1_cond $X=6.055 $Y=0.352
+ $X2=6.995 $Y2=0.352
r112 52 54 48.6294 $w=1.93e-07 $l=8.55e-07 $layer=LI1_cond $X=5.2 $Y=0.352
+ $X2=6.055 $Y2=0.352
r113 49 51 5.09219 $w=2.13e-07 $l=9.5e-08 $layer=LI1_cond $X=5.092 $Y=0.655
+ $X2=5.092 $Y2=0.56
r114 48 52 6.83761 $w=1.95e-07 $l=1.49158e-07 $layer=LI1_cond $X=5.092 $Y=0.45
+ $X2=5.2 $Y2=0.352
r115 48 51 5.89622 $w=2.13e-07 $l=1.1e-07 $layer=LI1_cond $X=5.092 $Y=0.45
+ $X2=5.092 $Y2=0.56
r116 47 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0.74
+ $X2=4.12 $Y2=0.74
r117 46 49 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=4.985 $Y=0.74
+ $X2=5.092 $Y2=0.655
r118 46 47 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=4.985 $Y=0.74
+ $X2=4.205 $Y2=0.74
r119 43 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0.655
+ $X2=4.12 $Y2=0.74
r120 43 45 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.12 $Y=0.655
+ $X2=4.12 $Y2=0.56
r121 42 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.265 $Y=0.74
+ $X2=3.18 $Y2=0.74
r122 41 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.74
+ $X2=4.12 $Y2=0.74
r123 41 42 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.035 $Y=0.74
+ $X2=3.265 $Y2=0.74
r124 38 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=0.655
+ $X2=3.18 $Y2=0.74
r125 38 40 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.18 $Y=0.655
+ $X2=3.18 $Y2=0.56
r126 37 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=0.74
+ $X2=2.24 $Y2=0.74
r127 36 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=0.74
+ $X2=3.18 $Y2=0.74
r128 36 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.095 $Y=0.74
+ $X2=2.325 $Y2=0.74
r129 33 62 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.655
+ $X2=2.24 $Y2=0.74
r130 33 35 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.24 $Y=0.655
+ $X2=2.24 $Y2=0.56
r131 31 62 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.74
+ $X2=2.24 $Y2=0.74
r132 31 32 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.155 $Y=0.74
+ $X2=1.385 $Y2=0.74
r133 28 32 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.225 $Y=0.655
+ $X2=1.385 $Y2=0.74
r134 28 30 3.62188 $w=3.2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.225 $Y=0.655
+ $X2=1.225 $Y2=0.56
r135 9 60 182 $w=1.7e-07 $l=1.89143e-07 $layer=licon1_NDIFF $count=1 $X=8.74
+ $Y=0.235 $X2=8.875 $Y2=0.365
r136 8 58 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=7.75
+ $Y=0.235 $X2=7.935 $Y2=0.365
r137 7 56 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=6.81
+ $Y=0.235 $X2=6.995 $Y2=0.365
r138 6 54 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=5.87
+ $Y=0.235 $X2=6.055 $Y2=0.365
r139 5 51 182 $w=1.7e-07 $l=3.92906e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.235 $X2=5.09 $Y2=0.56
r140 4 45 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.12 $Y2=0.56
r141 3 40 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=3.045
+ $Y=0.235 $X2=3.18 $Y2=0.56
r142 2 35 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.105
+ $Y=0.235 $X2=2.24 $Y2=0.56
r143 1 30 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.56
.ends

