* File: sky130_fd_sc_hdll__nand3_4.pxi.spice
* Created: Thu Aug 27 19:13:51 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3_4%C N_C_c_101_n N_C_M1001_g N_C_M1002_g
+ N_C_c_102_n N_C_M1010_g N_C_M1017_g N_C_c_103_n N_C_M1015_g N_C_M1018_g
+ N_C_c_104_n N_C_M1021_g N_C_M1023_g C C C C N_C_c_99_n N_C_c_100_n C C
+ PM_SKY130_FD_SC_HDLL__NAND3_4%C
x_PM_SKY130_FD_SC_HDLL__NAND3_4%B N_B_M1009_g N_B_c_183_n N_B_M1000_g
+ N_B_M1013_g N_B_c_184_n N_B_M1005_g N_B_M1019_g N_B_c_185_n N_B_M1008_g
+ N_B_c_186_n N_B_M1012_g N_B_M1020_g B B B B N_B_c_181_n B B B B
+ PM_SKY130_FD_SC_HDLL__NAND3_4%B
x_PM_SKY130_FD_SC_HDLL__NAND3_4%A N_A_c_269_n N_A_M1003_g N_A_M1004_g
+ N_A_c_270_n N_A_M1007_g N_A_M1006_g N_A_c_271_n N_A_M1014_g N_A_M1011_g
+ N_A_c_272_n N_A_M1022_g N_A_M1016_g A A A A N_A_c_266_n N_A_c_267_n A A A
+ PM_SKY130_FD_SC_HDLL__NAND3_4%A
x_PM_SKY130_FD_SC_HDLL__NAND3_4%VPWR N_VPWR_M1001_d N_VPWR_M1010_d
+ N_VPWR_M1021_d N_VPWR_M1005_d N_VPWR_M1012_d N_VPWR_M1003_s N_VPWR_M1007_s
+ N_VPWR_M1022_s N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n N_VPWR_c_349_n
+ N_VPWR_c_350_n N_VPWR_c_351_n N_VPWR_c_352_n N_VPWR_c_353_n N_VPWR_c_354_n
+ N_VPWR_c_355_n N_VPWR_c_356_n VPWR N_VPWR_c_357_n N_VPWR_c_358_n
+ N_VPWR_c_340_n N_VPWR_c_360_n N_VPWR_c_361_n N_VPWR_c_362_n
+ PM_SKY130_FD_SC_HDLL__NAND3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3_4%Y N_Y_M1004_s N_Y_M1011_s N_Y_M1001_s
+ N_Y_M1015_s N_Y_M1000_s N_Y_M1008_s N_Y_M1003_d N_Y_M1014_d N_Y_c_450_n
+ N_Y_c_468_n N_Y_c_451_n N_Y_c_475_n N_Y_c_452_n N_Y_c_481_n N_Y_c_453_n
+ N_Y_c_497_n N_Y_c_454_n N_Y_c_447_n N_Y_c_521_n N_Y_c_455_n N_Y_c_528_n
+ N_Y_c_456_n N_Y_c_457_n N_Y_c_458_n N_Y_c_459_n N_Y_c_460_n N_Y_c_461_n Y Y Y
+ N_Y_c_449_n PM_SKY130_FD_SC_HDLL__NAND3_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND3_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1017_d
+ N_A_27_47#_M1023_d N_A_27_47#_M1013_d N_A_27_47#_M1020_d N_A_27_47#_c_604_n
+ N_A_27_47#_c_605_n N_A_27_47#_c_606_n N_A_27_47#_c_620_n N_A_27_47#_c_607_n
+ N_A_27_47#_c_608_n N_A_27_47#_c_609_n N_A_27_47#_c_610_n N_A_27_47#_c_611_n
+ N_A_27_47#_c_612_n N_A_27_47#_c_613_n PM_SKY130_FD_SC_HDLL__NAND3_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND3_4%VGND N_VGND_M1002_s N_VGND_M1018_s
+ N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n VGND N_VGND_c_687_n
+ N_VGND_c_688_n N_VGND_c_689_n N_VGND_c_690_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND3_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND3_4%A_485_47# N_A_485_47#_M1009_s
+ N_A_485_47#_M1019_s N_A_485_47#_M1004_d N_A_485_47#_M1006_d
+ N_A_485_47#_M1016_d N_A_485_47#_c_755_n
+ PM_SKY130_FD_SC_HDLL__NAND3_4%A_485_47#
cc_1 VNB N_C_M1002_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_C_M1017_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_C_M1018_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_C_M1023_g 0.018112f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_5 VNB C 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.105
cc_6 VNB N_C_c_99_n 0.0322984f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_7 VNB N_C_c_100_n 0.0848306f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.217
cc_8 VNB N_B_M1009_g 0.018112f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_9 VNB N_B_M1013_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_10 VNB N_B_M1019_g 0.0188863f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_11 VNB N_B_M1020_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_12 VNB N_B_c_181_n 0.0890066f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_13 VNB B 0.00579823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_M1004_g 0.0244807f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_A_M1006_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_16 VNB N_A_M1011_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_17 VNB N_A_M1016_g 0.0216212f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_18 VNB N_A_c_266_n 0.032981f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.16
cc_19 VNB N_A_c_267_n 0.0877027f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.217
cc_20 VNB A 0.00733316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_340_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_Y_c_447_n 0.0107685f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_23 VNB Y 0.0210462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_449_n 0.0152082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_604_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.025
cc_26 VNB N_A_27_47#_c_605_n 0.00258986f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_27 VNB N_A_27_47#_c_606_n 0.00942711f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_607_n 0.00233388f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.105
cc_29 VNB N_A_27_47#_c_608_n 0.00268189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_609_n 0.00410109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_610_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_32 VNB N_A_27_47#_c_611_n 0.00249456f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_33 VNB N_A_27_47#_c_612_n 0.00750224f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.217
cc_34 VNB N_A_27_47#_c_613_n 0.00277241f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.217
cc_35 VNB N_VGND_c_684_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.025
cc_36 VNB N_VGND_c_685_n 0.019303f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_37 VNB N_VGND_c_686_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_38 VNB N_VGND_c_687_n 0.121918f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_39 VNB N_VGND_c_688_n 0.338984f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_40 VNB N_VGND_c_689_n 0.0219658f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=1.105
cc_41 VNB N_VGND_c_690_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_485_47#_c_755_n 0.0196317f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_43 VPB N_C_c_101_n 0.0198486f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_44 VPB N_C_c_102_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_45 VPB N_C_c_103_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_46 VPB N_C_c_104_n 0.0160015f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_47 VPB N_C_c_100_n 0.028998f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_48 VPB N_B_c_183_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_49 VPB N_B_c_184_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_50 VPB N_B_c_185_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_51 VPB N_B_c_186_n 0.0201049f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_52 VPB N_B_c_181_n 0.0287283f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_53 VPB N_A_c_269_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_54 VPB N_A_c_270_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_55 VPB N_A_c_271_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_56 VPB N_A_c_272_n 0.0192567f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_57 VPB N_A_c_267_n 0.0292992f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_58 VPB N_VPWR_c_341_n 0.00994749f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.025
cc_59 VPB N_VPWR_c_342_n 0.0464745f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_60 VPB N_VPWR_c_343_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.075 $Y2=1.105
cc_61 VPB N_VPWR_c_344_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_345_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.16
cc_63 VPB N_VPWR_c_346_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_347_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.217
cc_65 VPB N_VPWR_c_348_n 0.0164978f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_66 VPB N_VPWR_c_349_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_350_n 0.0302042f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_68 VPB N_VPWR_c_351_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.175
cc_69 VPB N_VPWR_c_352_n 0.00324069f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.19
cc_70 VPB N_VPWR_c_353_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_354_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_355_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_356_n 0.00507132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_357_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_358_n 0.0116899f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_340_n 0.0518269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_360_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_361_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_362_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_Y_c_450_n 0.00176159f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.025
cc_81 VPB N_Y_c_451_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_82 VPB N_Y_c_452_n 0.00423523f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_Y_c_453_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_Y_c_454_n 0.0138068f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.217
cc_85 VPB N_Y_c_455_n 0.00173134f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.19
cc_86 VPB N_Y_c_456_n 0.0034184f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_Y_c_457_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_Y_c_458_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_Y_c_459_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_460_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_Y_c_461_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB Y 0.00762934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB Y 0.0187691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 N_C_M1023_g N_B_M1009_g 0.0243494f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_95 N_C_c_104_n N_B_c_183_n 0.0231619f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_C_c_100_n N_B_c_181_n 0.0243494f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_97 C B 0.00794911f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_98 N_C_c_100_n B 9.44011e-19 $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_99 N_C_c_101_n N_VPWR_c_342_n 0.00871449f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_100 C N_VPWR_c_342_n 0.0190812f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_101 N_C_c_99_n N_VPWR_c_342_n 0.0053674f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C_c_101_n N_VPWR_c_343_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_103 N_C_c_102_n N_VPWR_c_343_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_104 N_C_c_102_n N_VPWR_c_344_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_105 N_C_c_103_n N_VPWR_c_344_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_106 N_C_c_103_n N_VPWR_c_345_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_107 N_C_c_104_n N_VPWR_c_345_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C_c_104_n N_VPWR_c_346_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_109 N_C_c_101_n N_VPWR_c_340_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_C_c_102_n N_VPWR_c_340_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_C_c_103_n N_VPWR_c_340_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_112 N_C_c_104_n N_VPWR_c_340_n 0.011869f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_113 N_C_c_101_n N_Y_c_450_n 0.0046976f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_102_n N_Y_c_450_n 0.00116723f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_115 C N_Y_c_450_n 0.0305808f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_116 N_C_c_100_n N_Y_c_450_n 0.0074788f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_117 N_C_c_101_n N_Y_c_468_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_118 N_C_c_102_n N_Y_c_468_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_119 N_C_c_103_n N_Y_c_468_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_120 N_C_c_102_n N_Y_c_451_n 0.0153933f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_121 N_C_c_103_n N_Y_c_451_n 0.0113962f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_122 C N_Y_c_451_n 0.040258f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_123 N_C_c_100_n N_Y_c_451_n 0.00725062f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_124 N_C_c_102_n N_Y_c_475_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_125 N_C_c_103_n N_Y_c_475_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_C_c_104_n N_Y_c_475_n 0.0106251f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_127 N_C_c_104_n N_Y_c_452_n 0.017118f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 C N_Y_c_452_n 0.00101487f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_129 N_C_c_100_n N_Y_c_452_n 3.62813e-19 $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_130 N_C_c_104_n N_Y_c_481_n 6.48386e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C_c_103_n N_Y_c_457_n 0.00292783f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C_c_104_n N_Y_c_457_n 0.00116723f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 C N_Y_c_457_n 0.0305808f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_134 N_C_c_100_n N_Y_c_457_n 0.0074788f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_135 N_C_M1002_g N_A_27_47#_c_605_n 0.0108433f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_136 N_C_M1017_g N_A_27_47#_c_605_n 0.0060427f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_137 C N_A_27_47#_c_605_n 0.0396411f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_138 N_C_c_100_n N_A_27_47#_c_605_n 0.00375198f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_139 C N_A_27_47#_c_606_n 0.0255512f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_140 N_C_c_99_n N_A_27_47#_c_606_n 0.00756929f $X=0.395 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C_M1002_g N_A_27_47#_c_620_n 5.85252e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_142 N_C_M1017_g N_A_27_47#_c_620_n 0.00864756f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_143 N_C_M1017_g N_A_27_47#_c_607_n 0.00266283f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_144 C N_A_27_47#_c_607_n 0.030512f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_145 N_C_c_100_n N_A_27_47#_c_607_n 0.00332f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_146 N_C_M1018_g N_A_27_47#_c_608_n 0.0107068f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_147 N_C_M1023_g N_A_27_47#_c_608_n 0.00687942f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_148 C N_A_27_47#_c_608_n 0.0345087f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_149 N_C_c_100_n N_A_27_47#_c_608_n 0.0031956f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_150 N_C_M1018_g N_A_27_47#_c_609_n 2.65385e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_151 N_C_M1023_g N_A_27_47#_c_609_n 0.00711615f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_152 N_C_M1002_g N_VGND_c_684_n 0.00276126f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_153 N_C_M1017_g N_VGND_c_684_n 0.00361688f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_154 N_C_M1017_g N_VGND_c_685_n 0.00397237f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_155 N_C_M1018_g N_VGND_c_685_n 0.00439206f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_156 N_C_M1018_g N_VGND_c_686_n 0.00276126f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_157 N_C_M1023_g N_VGND_c_686_n 0.00615f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_158 N_C_M1023_g N_VGND_c_687_n 0.00433241f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_159 N_C_M1002_g N_VGND_c_688_n 0.00703713f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_160 N_C_M1017_g N_VGND_c_688_n 0.00582631f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_161 N_C_M1018_g N_VGND_c_688_n 0.00616524f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_162 N_C_M1023_g N_VGND_c_688_n 0.00612841f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_163 N_C_M1002_g N_VGND_c_689_n 0.00439206f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_164 N_C_M1023_g N_A_485_47#_c_755_n 7.03111e-19 $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_165 N_B_c_181_n N_A_c_266_n 0.00741568f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_166 B N_A_c_266_n 7.55054e-19 $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_167 N_B_c_181_n A 6.88356e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_168 B A 0.0152145f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_169 N_B_c_183_n N_VPWR_c_346_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_c_184_n N_VPWR_c_347_n 0.0052072f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B_c_185_n N_VPWR_c_347_n 0.004751f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_c_186_n N_VPWR_c_348_n 0.00825342f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B_c_183_n N_VPWR_c_351_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B_c_184_n N_VPWR_c_351_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B_c_185_n N_VPWR_c_357_n 0.00597712f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_186_n N_VPWR_c_357_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B_c_183_n N_VPWR_c_340_n 0.0100198f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B_c_184_n N_VPWR_c_340_n 0.0118438f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_185_n N_VPWR_c_340_n 0.00999457f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_186_n N_VPWR_c_340_n 0.0131262f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B_c_183_n N_Y_c_475_n 6.24674e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B_c_183_n N_Y_c_452_n 0.0113403f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B_c_181_n N_Y_c_452_n 3.10838e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_184 B N_Y_c_452_n 0.00840447f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_185 N_B_c_183_n N_Y_c_481_n 0.0130707f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_184_n N_Y_c_481_n 0.0106251f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_185_n N_Y_c_481_n 6.24674e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_184_n N_Y_c_453_n 0.0153933f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B_c_185_n N_Y_c_453_n 0.0113962f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_181_n N_Y_c_453_n 0.00725062f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_191 B N_Y_c_453_n 0.040258f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_192 N_B_c_184_n N_Y_c_497_n 6.48386e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_c_185_n N_Y_c_497_n 0.0130707f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B_c_186_n N_Y_c_497_n 0.0153658f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B_c_186_n N_Y_c_454_n 0.0179883f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_181_n N_Y_c_454_n 3.10838e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_197 B N_Y_c_454_n 0.0227895f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_198 N_B_c_183_n N_Y_c_458_n 0.00292783f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_184_n N_Y_c_458_n 0.00116723f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_181_n N_Y_c_458_n 0.0074788f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_201 B N_Y_c_458_n 0.0305808f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_202 N_B_c_185_n N_Y_c_459_n 0.00292783f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_186_n N_Y_c_459_n 0.00116723f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_181_n N_Y_c_459_n 0.00723098f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_205 B N_Y_c_459_n 0.0305808f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_206 N_B_M1009_g N_A_27_47#_c_609_n 0.00322747f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_207 N_B_M1013_g N_A_27_47#_c_609_n 2.40584e-19 $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_208 B N_A_27_47#_c_609_n 0.12623f $X=3.93 $Y=1.19 $X2=0 $Y2=0
cc_209 N_B_M1009_g N_A_27_47#_c_610_n 0.00853013f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_210 N_B_M1013_g N_A_27_47#_c_610_n 0.00773532f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_211 N_B_c_181_n N_A_27_47#_c_610_n 0.0031956f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_212 N_B_M1009_g N_A_27_47#_c_611_n 2.40584e-19 $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_213 N_B_M1013_g N_A_27_47#_c_611_n 0.00298321f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_214 N_B_M1019_g N_A_27_47#_c_611_n 0.00300245f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B_M1020_g N_A_27_47#_c_611_n 2.42175e-19 $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_216 N_B_c_181_n N_A_27_47#_c_611_n 0.00322716f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_217 N_B_M1019_g N_A_27_47#_c_612_n 2.65832e-19 $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_218 N_B_M1020_g N_A_27_47#_c_612_n 0.00556724f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_219 N_B_M1019_g N_A_27_47#_c_613_n 0.00799428f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_220 N_B_M1020_g N_A_27_47#_c_613_n 0.00568546f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_221 N_B_c_181_n N_A_27_47#_c_613_n 0.00433688f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_222 N_B_M1009_g N_VGND_c_687_n 0.00420703f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_223 N_B_M1013_g N_VGND_c_687_n 0.00357877f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_224 N_B_M1019_g N_VGND_c_687_n 0.00357877f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_225 N_B_M1020_g N_VGND_c_687_n 0.00357877f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_226 N_B_M1009_g N_VGND_c_688_n 0.00602822f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_227 N_B_M1013_g N_VGND_c_688_n 0.00548399f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_228 N_B_M1019_g N_VGND_c_688_n 0.00559933f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_229 N_B_M1020_g N_VGND_c_688_n 0.00684455f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_230 N_B_M1009_g N_A_485_47#_c_755_n 0.00518064f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_231 N_B_M1013_g N_A_485_47#_c_755_n 0.0099669f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_232 N_B_M1019_g N_A_485_47#_c_755_n 0.0099669f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_233 N_B_M1020_g N_A_485_47#_c_755_n 0.0122603f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_234 N_A_c_269_n N_VPWR_c_348_n 0.00762417f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_270_n N_VPWR_c_349_n 0.0052072f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_c_271_n N_VPWR_c_349_n 0.004751f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_c_272_n N_VPWR_c_350_n 0.00728278f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A_c_269_n N_VPWR_c_353_n 0.00597712f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_270_n N_VPWR_c_353_n 0.00673617f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_c_271_n N_VPWR_c_355_n 0.00597712f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_c_272_n N_VPWR_c_355_n 0.00673617f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_c_269_n N_VPWR_c_340_n 0.0112769f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_c_270_n N_VPWR_c_340_n 0.0118438f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_c_271_n N_VPWR_c_340_n 0.00999457f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_c_272_n N_VPWR_c_340_n 0.0129051f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_269_n N_Y_c_454_n 0.0139912f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_266_n N_Y_c_454_n 0.00729564f $X=4.675 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_267_n N_Y_c_454_n 2.73568e-19 $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_249 A N_Y_c_454_n 0.0401373f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_250 N_A_M1004_g N_Y_c_447_n 0.00863645f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A_M1006_g N_Y_c_447_n 0.0111698f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A_M1011_g N_Y_c_447_n 0.0111698f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_253 N_A_M1016_g N_Y_c_447_n 0.0134479f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_c_267_n N_Y_c_447_n 0.00968149f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_255 A N_Y_c_447_n 0.115822f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_256 N_A_c_269_n N_Y_c_521_n 0.0178402f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_c_270_n N_Y_c_521_n 0.0106251f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_271_n N_Y_c_521_n 6.24674e-19 $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_c_270_n N_Y_c_455_n 0.0153933f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_271_n N_Y_c_455_n 0.0113962f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_267_n N_Y_c_455_n 0.00725062f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_262 A N_Y_c_455_n 0.040258f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_263 N_A_c_270_n N_Y_c_528_n 6.48386e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_271_n N_Y_c_528_n 0.0130707f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_272_n N_Y_c_528_n 0.0153658f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_c_272_n N_Y_c_456_n 0.0176391f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_c_267_n N_Y_c_456_n 3.10838e-19 $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_268 A N_Y_c_456_n 0.0185134f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_269 N_A_c_269_n N_Y_c_460_n 0.00292783f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_c_270_n N_Y_c_460_n 0.00116723f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_c_267_n N_Y_c_460_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_272 A N_Y_c_460_n 0.0305808f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_273 N_A_c_271_n N_Y_c_461_n 0.00292783f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_c_272_n N_Y_c_461_n 0.00116723f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_267_n N_Y_c_461_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_276 A N_Y_c_461_n 0.0305808f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_277 N_A_c_272_n Y 0.00109426f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_M1016_g Y 0.00575311f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_c_267_n Y 0.00571229f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_280 A Y 0.0160804f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_281 N_A_M1004_g N_A_27_47#_c_612_n 0.00400917f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_M1004_g N_VGND_c_687_n 0.00357877f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_M1006_g N_VGND_c_687_n 0.00357877f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_M1011_g N_VGND_c_687_n 0.00357877f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_M1016_g N_VGND_c_687_n 0.00357877f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_M1004_g N_VGND_c_688_n 0.00668309f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_M1006_g N_VGND_c_688_n 0.00548399f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_M1011_g N_VGND_c_688_n 0.00548399f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_M1016_g N_VGND_c_688_n 0.00646571f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_M1004_g N_A_485_47#_c_755_n 0.0105253f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_M1006_g N_A_485_47#_c_755_n 0.00958923f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_M1011_g N_A_485_47#_c_755_n 0.00958923f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_M1016_g N_A_485_47#_c_755_n 0.00958923f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_294 N_A_c_266_n N_A_485_47#_c_755_n 0.00630022f $X=4.675 $Y=1.16 $X2=0 $Y2=0
cc_295 A N_A_485_47#_c_755_n 0.0145371f $X=6.235 $Y=1.19 $X2=0 $Y2=0
cc_296 N_VPWR_c_340_n N_Y_M1001_s 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_340_n N_Y_M1015_s 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_c_340_n N_Y_M1000_s 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_340_n N_Y_M1008_s 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_340_n N_Y_M1003_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_340_n N_Y_M1014_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_342_n N_Y_c_450_n 0.0178509f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_303 N_VPWR_c_342_n N_Y_c_468_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_304 N_VPWR_c_343_n N_Y_c_468_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_305 N_VPWR_c_344_n N_Y_c_468_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_306 N_VPWR_c_340_n N_Y_c_468_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_307 N_VPWR_M1010_d N_Y_c_451_n 0.00180012f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_308 N_VPWR_c_344_n N_Y_c_451_n 0.0139097f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_309 N_VPWR_c_344_n N_Y_c_475_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_310 N_VPWR_c_345_n N_Y_c_475_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_311 N_VPWR_c_346_n N_Y_c_475_n 0.0385613f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_312 N_VPWR_c_340_n N_Y_c_475_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_313 N_VPWR_M1021_d N_Y_c_452_n 0.00180012f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_314 N_VPWR_c_346_n N_Y_c_452_n 0.0139097f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_315 N_VPWR_c_346_n N_Y_c_481_n 0.0470327f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_316 N_VPWR_c_347_n N_Y_c_481_n 0.0385613f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_317 N_VPWR_c_351_n N_Y_c_481_n 0.0223557f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_340_n N_Y_c_481_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_M1005_d N_Y_c_453_n 0.00180012f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_320 N_VPWR_c_347_n N_Y_c_453_n 0.0139097f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_321 N_VPWR_c_347_n N_Y_c_497_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_322 N_VPWR_c_348_n N_Y_c_497_n 0.0429581f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_323 N_VPWR_c_357_n N_Y_c_497_n 0.0223557f $X=3.935 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_340_n N_Y_c_497_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_325 N_VPWR_M1012_d N_Y_c_454_n 0.00313113f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_326 N_VPWR_M1003_s N_Y_c_454_n 0.00313113f $X=4.415 $Y=1.485 $X2=0 $Y2=0
cc_327 N_VPWR_c_348_n N_Y_c_454_n 0.0578207f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_328 N_VPWR_c_348_n N_Y_c_521_n 0.0523533f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_329 N_VPWR_c_349_n N_Y_c_521_n 0.0385613f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_330 N_VPWR_c_353_n N_Y_c_521_n 0.0223557f $X=5.395 $Y=2.72 $X2=0 $Y2=0
cc_331 N_VPWR_c_340_n N_Y_c_521_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_332 N_VPWR_M1007_s N_Y_c_455_n 0.00180012f $X=5.335 $Y=1.485 $X2=0 $Y2=0
cc_333 N_VPWR_c_349_n N_Y_c_455_n 0.0139097f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_334 N_VPWR_c_349_n N_Y_c_528_n 0.0470327f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_335 N_VPWR_c_350_n N_Y_c_528_n 0.0398607f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_336 N_VPWR_c_355_n N_Y_c_528_n 0.0223557f $X=6.335 $Y=2.72 $X2=0 $Y2=0
cc_337 N_VPWR_c_340_n N_Y_c_528_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_338 N_VPWR_M1022_s N_Y_c_456_n 0.00331674f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_339 N_VPWR_c_350_n N_Y_c_456_n 0.0180943f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_340 N_VPWR_c_350_n Y 0.004029f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_341 N_VPWR_c_342_n N_A_27_47#_c_606_n 7.91944e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_342 N_Y_c_452_n N_A_27_47#_c_608_n 0.0138466f $X=2.395 $Y=1.555 $X2=0 $Y2=0
cc_343 N_Y_c_454_n N_A_27_47#_c_612_n 0.00567975f $X=4.795 $Y=1.555 $X2=0 $Y2=0
cc_344 N_Y_c_447_n N_A_27_47#_c_612_n 0.00823418f $X=6.555 $Y=0.78 $X2=0 $Y2=0
cc_345 N_Y_c_449_n N_VGND_c_687_n 0.00360587f $X=6.67 $Y=0.905 $X2=0 $Y2=0
cc_346 N_Y_M1004_s N_VGND_c_688_n 0.00256987f $X=4.875 $Y=0.235 $X2=0 $Y2=0
cc_347 N_Y_M1011_s N_VGND_c_688_n 0.00256987f $X=5.815 $Y=0.235 $X2=0 $Y2=0
cc_348 N_Y_c_449_n N_VGND_c_688_n 0.00559591f $X=6.67 $Y=0.905 $X2=0 $Y2=0
cc_349 N_Y_c_447_n N_A_485_47#_M1006_d 0.00214463f $X=6.555 $Y=0.78 $X2=0 $Y2=0
cc_350 N_Y_c_447_n N_A_485_47#_M1016_d 0.00333519f $X=6.555 $Y=0.78 $X2=0 $Y2=0
cc_351 N_Y_M1004_s N_A_485_47#_c_755_n 0.00401739f $X=4.875 $Y=0.235 $X2=0 $Y2=0
cc_352 N_Y_M1011_s N_A_485_47#_c_755_n 0.00401739f $X=5.815 $Y=0.235 $X2=0 $Y2=0
cc_353 N_Y_c_447_n N_A_485_47#_c_755_n 0.0962868f $X=6.555 $Y=0.78 $X2=0 $Y2=0
cc_354 N_Y_c_449_n N_A_485_47#_c_755_n 0.00368247f $X=6.67 $Y=0.905 $X2=0 $Y2=0
cc_355 N_A_27_47#_c_605_n N_VGND_M1002_s 0.00251598f $X=0.985 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_356 N_A_27_47#_c_608_n N_VGND_M1018_s 0.00251598f $X=1.925 $Y=0.78 $X2=0
+ $Y2=0
cc_357 N_A_27_47#_c_605_n N_VGND_c_684_n 0.0127122f $X=0.985 $Y=0.82 $X2=0 $Y2=0
cc_358 N_A_27_47#_c_620_n N_VGND_c_684_n 0.0231432f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_359 N_A_27_47#_c_605_n N_VGND_c_685_n 0.00194552f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_360 N_A_27_47#_c_620_n N_VGND_c_685_n 0.023074f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_361 N_A_27_47#_c_608_n N_VGND_c_685_n 0.00248202f $X=1.925 $Y=0.78 $X2=0
+ $Y2=0
cc_362 N_A_27_47#_c_608_n N_VGND_c_686_n 0.0127122f $X=1.925 $Y=0.78 $X2=0 $Y2=0
cc_363 N_A_27_47#_c_608_n N_VGND_c_687_n 0.00194552f $X=1.925 $Y=0.78 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_609_n N_VGND_c_687_n 0.00548985f $X=2.305 $Y=0.78 $X2=0
+ $Y2=0
cc_365 N_A_27_47#_c_610_n N_VGND_c_687_n 0.00117399f $X=2.865 $Y=0.78 $X2=0
+ $Y2=0
cc_366 N_A_27_47#_M1002_d N_VGND_c_688_n 0.00259235f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_27_47#_M1017_d N_VGND_c_688_n 0.00264276f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_27_47#_M1023_d N_VGND_c_688_n 0.00323135f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_369 N_A_27_47#_M1013_d N_VGND_c_688_n 0.00256987f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_370 N_A_27_47#_M1020_d N_VGND_c_688_n 0.00210147f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_371 N_A_27_47#_c_604_n N_VGND_c_688_n 0.0128092f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_372 N_A_27_47#_c_605_n N_VGND_c_688_n 0.00966112f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_373 N_A_27_47#_c_620_n N_VGND_c_688_n 0.0141066f $X=1.2 $Y=0.4 $X2=0 $Y2=0
cc_374 N_A_27_47#_c_608_n N_VGND_c_688_n 0.00966112f $X=1.925 $Y=0.78 $X2=0
+ $Y2=0
cc_375 N_A_27_47#_c_609_n N_VGND_c_688_n 0.0101904f $X=2.305 $Y=0.78 $X2=0 $Y2=0
cc_376 N_A_27_47#_c_610_n N_VGND_c_688_n 0.00294408f $X=2.865 $Y=0.78 $X2=0
+ $Y2=0
cc_377 N_A_27_47#_c_604_n N_VGND_c_689_n 0.0221535f $X=0.26 $Y=0.4 $X2=0 $Y2=0
cc_378 N_A_27_47#_c_605_n N_VGND_c_689_n 0.00248202f $X=0.985 $Y=0.82 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_610_n N_A_485_47#_M1009_s 0.00253128f $X=2.865 $Y=0.78
+ $X2=-0.19 $Y2=-0.24
cc_380 N_A_27_47#_c_613_n N_A_485_47#_M1019_s 0.00322814f $X=3.805 $Y=0.78 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_M1013_d N_A_485_47#_c_755_n 0.00401739f $X=2.895 $Y=0.235
+ $X2=0 $Y2=0
cc_382 N_A_27_47#_M1020_d N_A_485_47#_c_755_n 0.00511748f $X=3.885 $Y=0.235
+ $X2=0 $Y2=0
cc_383 N_A_27_47#_c_610_n N_A_485_47#_c_755_n 0.0175415f $X=2.865 $Y=0.78 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_611_n N_A_485_47#_c_755_n 0.0190148f $X=3.245 $Y=0.78 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_612_n N_A_485_47#_c_755_n 0.0232109f $X=4.02 $Y=0.74 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_613_n N_A_485_47#_c_755_n 0.0219645f $X=3.805 $Y=0.78 $X2=0
+ $Y2=0
cc_387 N_VGND_c_688_n N_A_485_47#_M1009_s 0.00255381f $X=6.67 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_388 N_VGND_c_688_n N_A_485_47#_M1019_s 0.00295535f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_688_n N_A_485_47#_M1004_d 0.00250339f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_688_n N_A_485_47#_M1006_d 0.00255381f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_688_n N_A_485_47#_M1016_d 0.00217543f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_686_n N_A_485_47#_c_755_n 0.00620687f $X=1.67 $Y=0.4 $X2=0 $Y2=0
cc_393 N_VGND_c_687_n N_A_485_47#_c_755_n 0.244926f $X=6.67 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_688_n N_A_485_47#_c_755_n 0.152161f $X=6.67 $Y=0 $X2=0 $Y2=0
