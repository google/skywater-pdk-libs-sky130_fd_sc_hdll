# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb4to1_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  25.76000 BY  2.720000 ;
  SITE unithd ;
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.395000 1.055000 1.785000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.095000 1.055000 12.485000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.275000 1.055000 14.665000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.975000 1.055000 25.365000 1.325000 ;
    END
  END D[3]
  PIN S[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 0.995000 6.355000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.525000 0.995000 7.120000 1.325000 ;
    END
  END S[1]
  PIN S[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.640000 0.995000 19.235000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 19.405000 0.995000 20.000000 1.325000 ;
    END
  END S[3]
  PIN Z
    ANTENNADIFFAREA  1.992000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  2.985000 1.755000  3.275000 1.800000 ;
        RECT  2.985000 1.800000 22.775000 1.940000 ;
        RECT  2.985000 1.940000  3.275000 1.985000 ;
        RECT  3.925000 1.755000  4.215000 1.800000 ;
        RECT  3.925000 1.940000  4.215000 1.985000 ;
        RECT  8.665000 1.755000  8.955000 1.800000 ;
        RECT  8.665000 1.940000  8.955000 1.985000 ;
        RECT  9.605000 1.755000  9.895000 1.800000 ;
        RECT  9.605000 1.940000  9.895000 1.985000 ;
        RECT 15.865000 1.755000 16.155000 1.800000 ;
        RECT 15.865000 1.940000 16.155000 1.985000 ;
        RECT 16.805000 1.755000 17.095000 1.800000 ;
        RECT 16.805000 1.940000 17.095000 1.985000 ;
        RECT 21.545000 1.755000 21.835000 1.800000 ;
        RECT 21.545000 1.940000 21.835000 1.985000 ;
        RECT 22.485000 1.755000 22.775000 1.800000 ;
        RECT 22.485000 1.940000 22.775000 1.985000 ;
    END
  END Z
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 25.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 25.760000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 25.760000 0.085000 ;
      RECT  0.000000  2.635000 25.760000 2.805000 ;
      RECT  0.125000  1.495000  0.395000 2.635000 ;
      RECT  0.145000  0.085000  0.395000 0.885000 ;
      RECT  0.565000  0.255000  0.895000 0.715000 ;
      RECT  0.565000  0.715000  2.695000 0.885000 ;
      RECT  0.565000  1.495000  2.795000 1.665000 ;
      RECT  0.565000  1.665000  0.895000 2.465000 ;
      RECT  1.065000  0.085000  1.335000 0.545000 ;
      RECT  1.065000  1.835000  1.335000 2.635000 ;
      RECT  1.505000  0.255000  1.835000 0.715000 ;
      RECT  1.505000  1.665000  1.835000 2.465000 ;
      RECT  2.005000  0.085000  2.255000 0.545000 ;
      RECT  2.005000  1.835000  2.275000 2.635000 ;
      RECT  2.425000  0.255000  4.455000 0.425000 ;
      RECT  2.425000  0.425000  2.695000 0.715000 ;
      RECT  2.495000  1.665000  2.795000 2.295000 ;
      RECT  2.495000  2.295000  4.705000 2.465000 ;
      RECT  2.865000  0.595000  3.195000 0.885000 ;
      RECT  2.965000  0.885000  3.195000 1.065000 ;
      RECT  2.965000  1.065000  4.235000 1.365000 ;
      RECT  2.965000  1.365000  3.295000 2.125000 ;
      RECT  3.365000  0.425000  3.535000 0.770000 ;
      RECT  3.465000  1.535000  3.735000 2.295000 ;
      RECT  3.705000  0.595000  4.035000 1.065000 ;
      RECT  3.905000  1.365000  4.235000 2.125000 ;
      RECT  4.205000  0.425000  4.455000 0.770000 ;
      RECT  4.405000  1.065000  5.590000 1.395000 ;
      RECT  4.405000  1.565000  4.705000 2.295000 ;
      RECT  4.950000  1.605000  5.225000 2.635000 ;
      RECT  4.960000  0.085000  5.250000 0.610000 ;
      RECT  5.420000  0.280000  5.670000 0.825000 ;
      RECT  5.420000  0.825000  5.590000 1.065000 ;
      RECT  5.420000  1.395000  5.590000 1.605000 ;
      RECT  5.420000  1.605000  5.750000 2.465000 ;
      RECT  5.880000  0.085000  6.170000 0.610000 ;
      RECT  5.920000  1.605000  6.220000 2.635000 ;
      RECT  6.660000  1.605000  6.960000 2.635000 ;
      RECT  6.710000  0.085000  7.000000 0.610000 ;
      RECT  7.130000  1.605000  7.460000 2.465000 ;
      RECT  7.210000  0.280000  7.460000 0.825000 ;
      RECT  7.290000  0.825000  7.460000 1.065000 ;
      RECT  7.290000  1.065000  8.475000 1.395000 ;
      RECT  7.290000  1.395000  7.460000 1.605000 ;
      RECT  7.630000  0.085000  7.920000 0.610000 ;
      RECT  7.655000  1.605000  7.930000 2.635000 ;
      RECT  8.175000  1.565000  8.475000 2.295000 ;
      RECT  8.175000  2.295000 10.385000 2.465000 ;
      RECT  8.425000  0.255000 10.455000 0.425000 ;
      RECT  8.425000  0.425000  8.675000 0.770000 ;
      RECT  8.645000  1.065000  9.915000 1.365000 ;
      RECT  8.645000  1.365000  8.975000 2.125000 ;
      RECT  8.845000  0.595000  9.175000 1.065000 ;
      RECT  9.145000  1.535000  9.415000 2.295000 ;
      RECT  9.345000  0.425000  9.515000 0.770000 ;
      RECT  9.585000  1.365000  9.915000 2.125000 ;
      RECT  9.685000  0.595000 10.015000 0.885000 ;
      RECT  9.685000  0.885000  9.915000 1.065000 ;
      RECT 10.085000  1.495000 12.315000 1.665000 ;
      RECT 10.085000  1.665000 10.385000 2.295000 ;
      RECT 10.185000  0.425000 10.455000 0.715000 ;
      RECT 10.185000  0.715000 12.315000 0.885000 ;
      RECT 10.605000  1.835000 10.875000 2.635000 ;
      RECT 10.625000  0.085000 10.875000 0.545000 ;
      RECT 11.045000  0.255000 11.375000 0.715000 ;
      RECT 11.045000  1.665000 11.375000 2.465000 ;
      RECT 11.545000  0.085000 11.815000 0.545000 ;
      RECT 11.545000  1.835000 11.815000 2.635000 ;
      RECT 11.985000  0.255000 12.315000 0.715000 ;
      RECT 11.985000  1.665000 12.315000 2.465000 ;
      RECT 12.485000  0.085000 12.735000 0.885000 ;
      RECT 12.485000  1.495000 12.755000 2.635000 ;
      RECT 13.005000  1.495000 13.275000 2.635000 ;
      RECT 13.025000  0.085000 13.275000 0.885000 ;
      RECT 13.445000  0.255000 13.775000 0.715000 ;
      RECT 13.445000  0.715000 15.575000 0.885000 ;
      RECT 13.445000  1.495000 15.675000 1.665000 ;
      RECT 13.445000  1.665000 13.775000 2.465000 ;
      RECT 13.945000  0.085000 14.215000 0.545000 ;
      RECT 13.945000  1.835000 14.215000 2.635000 ;
      RECT 14.385000  0.255000 14.715000 0.715000 ;
      RECT 14.385000  1.665000 14.715000 2.465000 ;
      RECT 14.885000  0.085000 15.135000 0.545000 ;
      RECT 14.885000  1.835000 15.155000 2.635000 ;
      RECT 15.305000  0.255000 17.335000 0.425000 ;
      RECT 15.305000  0.425000 15.575000 0.715000 ;
      RECT 15.375000  1.665000 15.675000 2.295000 ;
      RECT 15.375000  2.295000 17.585000 2.465000 ;
      RECT 15.745000  0.595000 16.075000 0.885000 ;
      RECT 15.845000  0.885000 16.075000 1.065000 ;
      RECT 15.845000  1.065000 17.115000 1.365000 ;
      RECT 15.845000  1.365000 16.175000 2.125000 ;
      RECT 16.245000  0.425000 16.415000 0.770000 ;
      RECT 16.345000  1.535000 16.615000 2.295000 ;
      RECT 16.585000  0.595000 16.915000 1.065000 ;
      RECT 16.785000  1.365000 17.115000 2.125000 ;
      RECT 17.085000  0.425000 17.335000 0.770000 ;
      RECT 17.285000  1.065000 18.470000 1.395000 ;
      RECT 17.285000  1.565000 17.585000 2.295000 ;
      RECT 17.830000  1.605000 18.105000 2.635000 ;
      RECT 17.840000  0.085000 18.130000 0.610000 ;
      RECT 18.300000  0.280000 18.550000 0.825000 ;
      RECT 18.300000  0.825000 18.470000 1.065000 ;
      RECT 18.300000  1.395000 18.470000 1.605000 ;
      RECT 18.300000  1.605000 18.630000 2.465000 ;
      RECT 18.760000  0.085000 19.050000 0.610000 ;
      RECT 18.800000  1.605000 19.100000 2.635000 ;
      RECT 19.540000  1.605000 19.840000 2.635000 ;
      RECT 19.590000  0.085000 19.880000 0.610000 ;
      RECT 20.010000  1.605000 20.340000 2.465000 ;
      RECT 20.090000  0.280000 20.340000 0.825000 ;
      RECT 20.170000  0.825000 20.340000 1.065000 ;
      RECT 20.170000  1.065000 21.355000 1.395000 ;
      RECT 20.170000  1.395000 20.340000 1.605000 ;
      RECT 20.510000  0.085000 20.800000 0.610000 ;
      RECT 20.535000  1.605000 20.810000 2.635000 ;
      RECT 21.055000  1.565000 21.355000 2.295000 ;
      RECT 21.055000  2.295000 23.265000 2.465000 ;
      RECT 21.305000  0.255000 23.335000 0.425000 ;
      RECT 21.305000  0.425000 21.555000 0.770000 ;
      RECT 21.525000  1.065000 22.795000 1.365000 ;
      RECT 21.525000  1.365000 21.855000 2.125000 ;
      RECT 21.725000  0.595000 22.055000 1.065000 ;
      RECT 22.025000  1.535000 22.295000 2.295000 ;
      RECT 22.225000  0.425000 22.395000 0.770000 ;
      RECT 22.465000  1.365000 22.795000 2.125000 ;
      RECT 22.565000  0.595000 22.895000 0.885000 ;
      RECT 22.565000  0.885000 22.795000 1.065000 ;
      RECT 22.965000  1.495000 25.195000 1.665000 ;
      RECT 22.965000  1.665000 23.265000 2.295000 ;
      RECT 23.065000  0.425000 23.335000 0.715000 ;
      RECT 23.065000  0.715000 25.195000 0.885000 ;
      RECT 23.485000  1.835000 23.755000 2.635000 ;
      RECT 23.505000  0.085000 23.755000 0.545000 ;
      RECT 23.925000  0.255000 24.255000 0.715000 ;
      RECT 23.925000  1.665000 24.255000 2.465000 ;
      RECT 24.425000  0.085000 24.695000 0.545000 ;
      RECT 24.425000  1.835000 24.695000 2.635000 ;
      RECT 24.865000  0.255000 25.195000 0.715000 ;
      RECT 24.865000  1.665000 25.195000 2.465000 ;
      RECT 25.365000  0.085000 25.615000 0.885000 ;
      RECT 25.365000  1.495000 25.635000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.045000  1.785000  3.215000 1.955000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  3.985000  1.785000  4.155000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.725000  1.785000  8.895000 1.955000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.665000  1.785000  9.835000 1.955000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
      RECT 15.785000 -0.085000 15.955000 0.085000 ;
      RECT 15.785000  2.635000 15.955000 2.805000 ;
      RECT 15.925000  1.785000 16.095000 1.955000 ;
      RECT 16.245000 -0.085000 16.415000 0.085000 ;
      RECT 16.245000  2.635000 16.415000 2.805000 ;
      RECT 16.705000 -0.085000 16.875000 0.085000 ;
      RECT 16.705000  2.635000 16.875000 2.805000 ;
      RECT 16.865000  1.785000 17.035000 1.955000 ;
      RECT 17.165000 -0.085000 17.335000 0.085000 ;
      RECT 17.165000  2.635000 17.335000 2.805000 ;
      RECT 17.625000 -0.085000 17.795000 0.085000 ;
      RECT 17.625000  2.635000 17.795000 2.805000 ;
      RECT 18.085000 -0.085000 18.255000 0.085000 ;
      RECT 18.085000  2.635000 18.255000 2.805000 ;
      RECT 18.545000 -0.085000 18.715000 0.085000 ;
      RECT 18.545000  2.635000 18.715000 2.805000 ;
      RECT 19.005000 -0.085000 19.175000 0.085000 ;
      RECT 19.005000  2.635000 19.175000 2.805000 ;
      RECT 19.465000 -0.085000 19.635000 0.085000 ;
      RECT 19.465000  2.635000 19.635000 2.805000 ;
      RECT 19.925000 -0.085000 20.095000 0.085000 ;
      RECT 19.925000  2.635000 20.095000 2.805000 ;
      RECT 20.385000 -0.085000 20.555000 0.085000 ;
      RECT 20.385000  2.635000 20.555000 2.805000 ;
      RECT 20.845000 -0.085000 21.015000 0.085000 ;
      RECT 20.845000  2.635000 21.015000 2.805000 ;
      RECT 21.305000 -0.085000 21.475000 0.085000 ;
      RECT 21.305000  2.635000 21.475000 2.805000 ;
      RECT 21.605000  1.785000 21.775000 1.955000 ;
      RECT 21.765000 -0.085000 21.935000 0.085000 ;
      RECT 21.765000  2.635000 21.935000 2.805000 ;
      RECT 22.225000 -0.085000 22.395000 0.085000 ;
      RECT 22.225000  2.635000 22.395000 2.805000 ;
      RECT 22.545000  1.785000 22.715000 1.955000 ;
      RECT 22.685000 -0.085000 22.855000 0.085000 ;
      RECT 22.685000  2.635000 22.855000 2.805000 ;
      RECT 23.145000 -0.085000 23.315000 0.085000 ;
      RECT 23.145000  2.635000 23.315000 2.805000 ;
      RECT 23.605000 -0.085000 23.775000 0.085000 ;
      RECT 23.605000  2.635000 23.775000 2.805000 ;
      RECT 24.065000 -0.085000 24.235000 0.085000 ;
      RECT 24.065000  2.635000 24.235000 2.805000 ;
      RECT 24.525000 -0.085000 24.695000 0.085000 ;
      RECT 24.525000  2.635000 24.695000 2.805000 ;
      RECT 24.985000 -0.085000 25.155000 0.085000 ;
      RECT 24.985000  2.635000 25.155000 2.805000 ;
      RECT 25.445000 -0.085000 25.615000 0.085000 ;
      RECT 25.445000  2.635000 25.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_4
END LIBRARY
