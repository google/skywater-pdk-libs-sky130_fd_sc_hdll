* File: sky130_fd_sc_hdll__or4_4.pxi.spice
* Created: Thu Aug 27 19:25:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4_4%D N_D_c_79_n N_D_M1014_g N_D_c_76_n N_D_M1013_g D
+ D N_D_c_78_n PM_SKY130_FD_SC_HDLL__OR4_4%D
x_PM_SKY130_FD_SC_HDLL__OR4_4%C N_C_c_107_n N_C_M1008_g N_C_c_108_n N_C_M1006_g
+ N_C_c_109_n C C C PM_SKY130_FD_SC_HDLL__OR4_4%C
x_PM_SKY130_FD_SC_HDLL__OR4_4%B N_B_c_150_n N_B_M1001_g N_B_c_151_n N_B_M1005_g
+ N_B_c_152_n B B PM_SKY130_FD_SC_HDLL__OR4_4%B
x_PM_SKY130_FD_SC_HDLL__OR4_4%A N_A_c_188_n N_A_M1003_g N_A_c_189_n N_A_M1010_g
+ A N_A_c_190_n A PM_SKY130_FD_SC_HDLL__OR4_4%A
x_PM_SKY130_FD_SC_HDLL__OR4_4%A_32_297# N_A_32_297#_M1013_d N_A_32_297#_M1005_d
+ N_A_32_297#_M1014_s N_A_32_297#_c_227_n N_A_32_297#_M1002_g
+ N_A_32_297#_c_235_n N_A_32_297#_M1000_g N_A_32_297#_c_228_n
+ N_A_32_297#_M1004_g N_A_32_297#_c_236_n N_A_32_297#_M1009_g
+ N_A_32_297#_c_229_n N_A_32_297#_M1007_g N_A_32_297#_c_237_n
+ N_A_32_297#_M1012_g N_A_32_297#_c_238_n N_A_32_297#_M1015_g
+ N_A_32_297#_c_230_n N_A_32_297#_M1011_g N_A_32_297#_c_239_n
+ N_A_32_297#_c_231_n N_A_32_297#_c_247_n N_A_32_297#_c_256_n
+ N_A_32_297#_c_248_n N_A_32_297#_c_347_p N_A_32_297#_c_268_n
+ N_A_32_297#_c_232_n N_A_32_297#_c_233_n N_A_32_297#_c_297_p
+ N_A_32_297#_c_263_n N_A_32_297#_c_234_n PM_SKY130_FD_SC_HDLL__OR4_4%A_32_297#
x_PM_SKY130_FD_SC_HDLL__OR4_4%VPWR N_VPWR_M1010_d N_VPWR_M1009_s N_VPWR_M1015_s
+ N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n VPWR N_VPWR_c_384_n
+ N_VPWR_c_375_n VPWR PM_SKY130_FD_SC_HDLL__OR4_4%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4_4%X N_X_M1002_d N_X_M1007_d N_X_M1000_d N_X_M1012_d
+ N_X_c_436_n N_X_c_480_n N_X_c_445_n N_X_c_437_n N_X_c_430_n N_X_c_431_n
+ N_X_c_463_n N_X_c_484_n N_X_c_438_n N_X_c_432_n N_X_c_433_n N_X_c_439_n X
+ N_X_c_435_n PM_SKY130_FD_SC_HDLL__OR4_4%X
x_PM_SKY130_FD_SC_HDLL__OR4_4%VGND N_VGND_M1013_s N_VGND_M1006_d N_VGND_M1003_d
+ N_VGND_M1004_s N_VGND_M1011_s N_VGND_c_509_n N_VGND_c_510_n N_VGND_c_511_n
+ N_VGND_c_512_n N_VGND_c_513_n N_VGND_c_514_n N_VGND_c_515_n N_VGND_c_516_n
+ N_VGND_c_517_n N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n VGND
+ N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n VGND
+ PM_SKY130_FD_SC_HDLL__OR4_4%VGND
cc_1 VNB N_D_c_76_n 0.0201074f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_2 VNB D 0.0218021f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=0.765
cc_3 VNB N_D_c_78_n 0.0397829f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_4 VNB N_C_c_107_n 0.0260391f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_5 VNB N_C_c_108_n 0.0176935f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_6 VNB N_C_c_109_n 0.00111747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_150_n 0.0216949f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_8 VNB N_B_c_151_n 0.01695f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_9 VNB N_B_c_152_n 0.00629304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_188_n 0.0177853f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.41
cc_11 VNB N_A_c_189_n 0.0260553f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_12 VNB N_A_c_190_n 0.00110961f $X=-0.19 $Y=-0.24 $X2=0.285 $Y2=1.16
cc_13 VNB N_A_32_297#_c_227_n 0.0171624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_32_297#_c_228_n 0.0167557f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_15 VNB N_A_32_297#_c_229_n 0.0171987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_32_297#_c_230_n 0.0200831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_32_297#_c_231_n 0.00303358f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_32_297#_c_232_n 0.0016277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_32_297#_c_233_n 0.00376665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_32_297#_c_234_n 0.0762306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_375_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_430_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_431_n 0.0017592f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_432_n 0.00123315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_433_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.0211332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_435_n 0.00911365f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_509_n 0.0106918f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=0.85
cc_29 VNB N_VGND_c_510_n 0.0185321f $X=-0.19 $Y=-0.24 $X2=0.227 $Y2=1.16
cc_30 VNB N_VGND_c_511_n 0.0195679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_512_n 0.00226425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_513_n 0.00260546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_514_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_515_n 0.0129152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_516_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_517_n 0.0173964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_518_n 0.00609289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_519_n 0.0178379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_520_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_521_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_522_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_523_n 0.239263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_D_c_79_n 0.0215949f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_44 VPB D 0.00425673f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=0.765
cc_45 VPB N_D_c_78_n 0.017203f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_46 VPB N_C_c_107_n 0.02828f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_47 VPB N_C_c_109_n 0.0010374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_B_c_150_n 0.0249345f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.41
cc_49 VPB N_B_c_152_n 0.00576121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB B 2.10939e-19 $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_51 VPB N_A_c_189_n 0.0263982f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=0.995
cc_52 VPB N_A_c_190_n 0.00184998f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_53 VPB A 0.00416191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_32_297#_c_235_n 0.0171649f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_55 VPB N_A_32_297#_c_236_n 0.0159743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_32_297#_c_237_n 0.0159556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_32_297#_c_238_n 0.0191486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_32_297#_c_239_n 0.0310345f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_32_297#_c_231_n 0.00869004f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_32_297#_c_234_n 0.0467455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_376_n 0.00519418f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_62 VPB N_VPWR_c_377_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=0.85
cc_63 VPB N_VPWR_c_378_n 0.0136825f $X=-0.19 $Y=1.305 $X2=0.227 $Y2=1.16
cc_64 VPB N_VPWR_c_379_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_380_n 0.0632257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_381_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_382_n 0.0213107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_383_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_384_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_375_n 0.0490581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_X_c_436_n 0.00190706f $X=-0.19 $Y=1.305 $X2=0.285 $Y2=1.16
cc_72 VPB N_X_c_437_n 0.00206401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_X_c_438_n 0.0122447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_X_c_439_n 0.00161374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB X 0.00789266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 N_D_c_79_n N_C_c_107_n 0.0335457f $X=0.52 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_77 N_D_c_78_n N_C_c_107_n 0.0180828f $X=0.52 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_78 N_D_c_76_n N_C_c_108_n 0.0203545f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_79 N_D_c_79_n N_C_c_109_n 6.27534e-19 $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_80 N_D_c_78_n N_C_c_109_n 5.11753e-19 $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_81 N_D_c_79_n C 0.00616947f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_82 N_D_c_79_n N_A_32_297#_c_239_n 0.0142367f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_83 N_D_c_79_n N_A_32_297#_c_231_n 0.0214918f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_84 N_D_c_76_n N_A_32_297#_c_231_n 0.00440389f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_85 D N_A_32_297#_c_231_n 0.0564286f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_86 N_D_c_78_n N_A_32_297#_c_231_n 0.0167795f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_87 N_D_c_76_n N_A_32_297#_c_247_n 0.00446123f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_88 N_D_c_76_n N_A_32_297#_c_248_n 0.0109239f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_89 D N_A_32_297#_c_248_n 0.00562567f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_90 N_D_c_79_n N_VPWR_c_380_n 0.00674013f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_91 N_D_c_79_n N_VPWR_c_375_n 0.0132274f $X=0.52 $Y=1.41 $X2=0 $Y2=0
cc_92 D N_VGND_M1013_s 0.00399065f $X=0.14 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_93 D N_VGND_c_509_n 5.41347e-19 $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_94 N_D_c_76_n N_VGND_c_510_n 0.00707235f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_95 D N_VGND_c_510_n 0.0214679f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_96 N_D_c_78_n N_VGND_c_510_n 0.00100535f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_97 N_D_c_76_n N_VGND_c_511_n 0.00501458f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_98 N_D_c_76_n N_VGND_c_512_n 0.0013206f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_99 N_D_c_76_n N_VGND_c_523_n 0.00951998f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_100 D N_VGND_c_523_n 0.00197281f $X=0.14 $Y=0.765 $X2=0 $Y2=0
cc_101 N_C_c_107_n N_B_c_150_n 0.0738038f $X=1.1 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_102 N_C_c_109_n N_B_c_150_n 9.93623e-19 $X=1.015 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_103 C N_B_c_150_n 0.0049168f $X=1.11 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_104 N_C_c_108_n N_B_c_151_n 0.0215326f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C_c_107_n N_B_c_152_n 0.00326052f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_106 N_C_c_109_n N_B_c_152_n 0.0239913f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_107 N_C_c_107_n B 0.00134972f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C_c_109_n B 0.00594195f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_109 C B 0.029771f $X=1.11 $Y=1.785 $X2=0 $Y2=0
cc_110 C B 0.029771f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_111 N_C_c_107_n N_A_32_297#_c_239_n 9.88251e-19 $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_112 C N_A_32_297#_c_239_n 0.0250465f $X=1.11 $Y=1.785 $X2=0 $Y2=0
cc_113 N_C_c_107_n N_A_32_297#_c_231_n 0.00330726f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_108_n N_A_32_297#_c_231_n 0.00340748f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_115 N_C_c_109_n N_A_32_297#_c_231_n 0.0509163f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_116 N_C_c_108_n N_A_32_297#_c_247_n 0.00540738f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_c_107_n N_A_32_297#_c_256_n 7.10472e-19 $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_118 N_C_c_108_n N_A_32_297#_c_256_n 0.0150804f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_119 N_C_c_109_n N_A_32_297#_c_256_n 0.0110068f $X=1.015 $Y=1.16 $X2=0 $Y2=0
cc_120 N_C_c_107_n N_A_32_297#_c_248_n 0.00189854f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_121 N_C_c_109_n A_122_297# 0.00117691f $X=1.015 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_122 C A_122_297# 0.00260417f $X=1.11 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_123 C A_122_297# 0.00813819f $X=1.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_124 C A_238_297# 0.00540645f $X=1.11 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_125 C A_238_297# 0.00569444f $X=1.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_126 N_C_c_107_n N_VPWR_c_380_n 0.00450951f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_127 C N_VPWR_c_380_n 0.0149389f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_128 N_C_c_107_n N_VPWR_c_375_n 0.00647188f $X=1.1 $Y=1.41 $X2=0 $Y2=0
cc_129 C N_VPWR_c_375_n 0.0137424f $X=1.145 $Y=1.87 $X2=0 $Y2=0
cc_130 N_C_c_108_n N_VGND_c_511_n 0.00199015f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_131 N_C_c_108_n N_VGND_c_512_n 0.0117441f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_132 N_C_c_108_n N_VGND_c_523_n 0.00304119f $X=1.125 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_151_n N_A_c_188_n 0.0249402f $X=1.595 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 N_B_c_150_n N_A_c_189_n 0.0741097f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_135 N_B_c_152_n N_A_c_189_n 0.00309823f $X=1.545 $Y=1.16 $X2=0 $Y2=0
cc_136 B N_A_c_189_n 0.0098765f $X=1.67 $Y=1.785 $X2=0 $Y2=0
cc_137 N_B_c_150_n N_A_c_190_n 5.80057e-19 $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_138 N_B_c_152_n N_A_c_190_n 0.0341568f $X=1.545 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B_c_150_n A 2.07758e-19 $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_152_n A 0.00792632f $X=1.545 $Y=1.16 $X2=0 $Y2=0
cc_141 N_B_c_150_n N_A_32_297#_c_256_n 6.47027e-19 $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_151_n N_A_32_297#_c_256_n 0.01167f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B_c_152_n N_A_32_297#_c_256_n 0.0222059f $X=1.545 $Y=1.16 $X2=0 $Y2=0
cc_144 N_B_c_152_n N_A_32_297#_c_263_n 0.00316818f $X=1.545 $Y=1.16 $X2=0 $Y2=0
cc_145 B A_332_297# 0.0103992f $X=1.67 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_146 B A_332_297# 0.0068829f $X=1.67 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_147 B N_VPWR_c_376_n 0.0278745f $X=1.67 $Y=1.785 $X2=0 $Y2=0
cc_148 N_B_c_150_n N_VPWR_c_380_n 0.00480294f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_149 B N_VPWR_c_380_n 0.0147961f $X=1.67 $Y=2.125 $X2=0 $Y2=0
cc_150 N_B_c_150_n N_VPWR_c_375_n 0.00699328f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_151 B N_VPWR_c_375_n 0.0127233f $X=1.67 $Y=2.125 $X2=0 $Y2=0
cc_152 N_B_c_151_n N_VGND_c_512_n 0.00176556f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B_c_151_n N_VGND_c_517_n 0.00428022f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B_c_151_n N_VGND_c_523_n 0.00585784f $X=1.595 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_188_n N_A_32_297#_c_227_n 0.0169356f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_189_n N_A_32_297#_c_235_n 0.0300132f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_190_n N_A_32_297#_c_235_n 6.97767e-19 $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_158 A N_A_32_297#_c_235_n 0.00138427f $X=2.27 $Y=1.53 $X2=0 $Y2=0
cc_159 N_A_c_188_n N_A_32_297#_c_268_n 0.0121667f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_c_189_n N_A_32_297#_c_268_n 0.00208416f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_190_n N_A_32_297#_c_268_n 0.0179369f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_162 A N_A_32_297#_c_268_n 0.00496743f $X=2.27 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A_c_188_n N_A_32_297#_c_232_n 0.00323346f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_189_n N_A_32_297#_c_232_n 5.19892e-19 $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_190_n N_A_32_297#_c_232_n 0.00588362f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_c_189_n N_A_32_297#_c_233_n 0.00127183f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_190_n N_A_32_297#_c_233_n 0.0141416f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_168 A N_A_32_297#_c_233_n 0.00707041f $X=2.27 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_c_189_n N_A_32_297#_c_234_n 0.0187825f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_190_n N_A_32_297#_c_234_n 0.00248787f $X=2.075 $Y=1.16 $X2=0 $Y2=0
cc_171 A N_VPWR_M1010_d 0.00517956f $X=2.27 $Y=1.53 $X2=-0.19 $Y2=-0.24
cc_172 N_A_c_189_n N_VPWR_c_376_n 0.0121442f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_173 A N_VPWR_c_376_n 0.0193325f $X=2.27 $Y=1.53 $X2=0 $Y2=0
cc_174 N_A_c_189_n N_VPWR_c_380_n 0.00702461f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_189_n N_VPWR_c_375_n 0.0130026f $X=2.04 $Y=1.41 $X2=0 $Y2=0
cc_176 A N_X_c_436_n 0.00200305f $X=2.27 $Y=1.53 $X2=0 $Y2=0
cc_177 N_A_c_188_n N_VGND_c_513_n 0.00473127f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_188_n N_VGND_c_517_n 0.00428022f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_188_n N_VGND_c_523_n 0.00626581f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_32_297#_c_231_n A_122_297# 0.00564644f $X=0.65 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_181 N_A_32_297#_c_235_n N_VPWR_c_376_n 0.0101706f $X=2.62 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_32_297#_c_236_n N_VPWR_c_377_n 0.00300743f $X=3.09 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_32_297#_c_237_n N_VPWR_c_377_n 0.00300743f $X=3.56 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_32_297#_c_238_n N_VPWR_c_379_n 0.00479105f $X=4.03 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_32_297#_c_239_n N_VPWR_c_380_n 0.0195512f $X=0.285 $Y=2.34 $X2=0
+ $Y2=0
cc_186 N_A_32_297#_c_235_n N_VPWR_c_382_n 0.00702461f $X=2.62 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_32_297#_c_236_n N_VPWR_c_382_n 0.00702461f $X=3.09 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_32_297#_c_237_n N_VPWR_c_384_n 0.00702461f $X=3.56 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_32_297#_c_238_n N_VPWR_c_384_n 0.00702461f $X=4.03 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_32_297#_M1014_s N_VPWR_c_375_n 0.00218082f $X=0.16 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_32_297#_c_235_n N_VPWR_c_375_n 0.0128986f $X=2.62 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_32_297#_c_236_n N_VPWR_c_375_n 0.0124092f $X=3.09 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_32_297#_c_237_n N_VPWR_c_375_n 0.0124092f $X=3.56 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_32_297#_c_238_n N_VPWR_c_375_n 0.0133833f $X=4.03 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_32_297#_c_239_n N_VPWR_c_375_n 0.0125731f $X=0.285 $Y=2.34 $X2=0
+ $Y2=0
cc_196 N_A_32_297#_c_235_n N_X_c_436_n 3.19638e-19 $X=2.62 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_32_297#_c_297_p N_X_c_436_n 0.0172229f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A_32_297#_c_234_n N_X_c_436_n 0.00674235f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A_32_297#_c_227_n N_X_c_445_n 0.00489827f $X=2.595 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_32_297#_c_228_n N_X_c_445_n 0.00766092f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_32_297#_c_229_n N_X_c_445_n 5.47877e-19 $X=3.535 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_32_297#_c_268_n N_X_c_445_n 0.00459795f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_203 N_A_32_297#_c_236_n N_X_c_437_n 0.0158555f $X=3.09 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_32_297#_c_237_n N_X_c_437_n 0.0159162f $X=3.56 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_32_297#_c_297_p N_X_c_437_n 0.0406907f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_32_297#_c_234_n N_X_c_437_n 0.00881912f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_207 N_A_32_297#_c_228_n N_X_c_430_n 0.00901745f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_32_297#_c_229_n N_X_c_430_n 0.00895898f $X=3.535 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_32_297#_c_297_p N_X_c_430_n 0.0392656f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_210 N_A_32_297#_c_234_n N_X_c_430_n 0.00345541f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_211 N_A_32_297#_c_227_n N_X_c_431_n 0.00157721f $X=2.595 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_32_297#_c_228_n N_X_c_431_n 0.00270583f $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_32_297#_c_268_n N_X_c_431_n 0.00715387f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_214 N_A_32_297#_c_232_n N_X_c_431_n 0.00518689f $X=2.465 $Y=1.075 $X2=0 $Y2=0
cc_215 N_A_32_297#_c_297_p N_X_c_431_n 0.0199589f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_32_297#_c_234_n N_X_c_431_n 0.0033272f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A_32_297#_c_228_n N_X_c_463_n 5.24597e-19 $X=3.065 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_32_297#_c_229_n N_X_c_463_n 0.00651696f $X=3.535 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_32_297#_c_238_n N_X_c_438_n 0.0186965f $X=4.03 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_32_297#_c_297_p N_X_c_438_n 0.00405064f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_32_297#_c_234_n N_X_c_438_n 9.44246e-19 $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_222 N_A_32_297#_c_230_n N_X_c_432_n 0.0139406f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_32_297#_c_297_p N_X_c_432_n 0.00208021f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_32_297#_c_229_n N_X_c_433_n 0.00119564f $X=3.535 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_32_297#_c_297_p N_X_c_433_n 0.0304076f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_32_297#_c_234_n N_X_c_433_n 0.00486271f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_227 N_A_32_297#_c_297_p N_X_c_439_n 0.0172229f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_32_297#_c_234_n N_X_c_439_n 0.0065364f $X=4.03 $Y=1.202 $X2=0 $Y2=0
cc_229 N_A_32_297#_c_238_n X 0.00177528f $X=4.03 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_32_297#_c_230_n X 0.019947f $X=4.055 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_32_297#_c_297_p X 0.0114448f $X=3.825 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_32_297#_c_256_n N_VGND_M1006_d 0.0075965f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_233 N_A_32_297#_c_268_n N_VGND_M1003_d 0.00762812f $X=2.38 $Y=0.74 $X2=0
+ $Y2=0
cc_234 N_A_32_297#_c_232_n N_VGND_M1003_d 7.52091e-19 $X=2.465 $Y=1.075 $X2=0
+ $Y2=0
cc_235 N_A_32_297#_c_247_n N_VGND_c_510_n 0.011573f $X=0.835 $Y=0.49 $X2=0 $Y2=0
cc_236 N_A_32_297#_c_247_n N_VGND_c_511_n 0.00852533f $X=0.835 $Y=0.49 $X2=0
+ $Y2=0
cc_237 N_A_32_297#_c_248_n N_VGND_c_511_n 0.00586573f $X=0.92 $Y=0.74 $X2=0
+ $Y2=0
cc_238 N_A_32_297#_c_247_n N_VGND_c_512_n 0.0118543f $X=0.835 $Y=0.49 $X2=0
+ $Y2=0
cc_239 N_A_32_297#_c_256_n N_VGND_c_512_n 0.0214497f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_240 N_A_32_297#_c_227_n N_VGND_c_513_n 0.00816884f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_32_297#_c_228_n N_VGND_c_513_n 0.00115121f $X=3.065 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_32_297#_c_268_n N_VGND_c_513_n 0.0252021f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_243 N_A_32_297#_c_228_n N_VGND_c_514_n 0.00379224f $X=3.065 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_32_297#_c_229_n N_VGND_c_514_n 0.00276126f $X=3.535 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_32_297#_c_230_n N_VGND_c_516_n 0.00438629f $X=4.055 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_32_297#_c_256_n N_VGND_c_517_n 0.0029785f $X=1.72 $Y=0.74 $X2=0 $Y2=0
cc_247 N_A_32_297#_c_347_p N_VGND_c_517_n 0.00846569f $X=1.805 $Y=0.49 $X2=0
+ $Y2=0
cc_248 N_A_32_297#_c_268_n N_VGND_c_517_n 0.0035399f $X=2.38 $Y=0.74 $X2=0 $Y2=0
cc_249 N_A_32_297#_c_227_n N_VGND_c_519_n 0.00496106f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_250 N_A_32_297#_c_228_n N_VGND_c_519_n 0.00423334f $X=3.065 $Y=0.995 $X2=0
+ $Y2=0
cc_251 N_A_32_297#_c_229_n N_VGND_c_521_n 0.00423334f $X=3.535 $Y=0.995 $X2=0
+ $Y2=0
cc_252 N_A_32_297#_c_230_n N_VGND_c_521_n 0.00437852f $X=4.055 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_32_297#_M1013_d N_VGND_c_523_n 0.00454252f $X=0.62 $Y=0.235 $X2=0
+ $Y2=0
cc_254 N_A_32_297#_M1005_d N_VGND_c_523_n 0.00256656f $X=1.67 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_A_32_297#_c_227_n N_VGND_c_523_n 0.0083553f $X=2.595 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_A_32_297#_c_228_n N_VGND_c_523_n 0.00613677f $X=3.065 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_32_297#_c_229_n N_VGND_c_523_n 0.00608558f $X=3.535 $Y=0.995 $X2=0
+ $Y2=0
cc_258 N_A_32_297#_c_230_n N_VGND_c_523_n 0.0071478f $X=4.055 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_32_297#_c_247_n N_VGND_c_523_n 0.00618681f $X=0.835 $Y=0.49 $X2=0
+ $Y2=0
cc_260 N_A_32_297#_c_256_n N_VGND_c_523_n 0.00691826f $X=1.72 $Y=0.74 $X2=0
+ $Y2=0
cc_261 N_A_32_297#_c_248_n N_VGND_c_523_n 0.0107733f $X=0.92 $Y=0.74 $X2=0 $Y2=0
cc_262 N_A_32_297#_c_347_p N_VGND_c_523_n 0.00625722f $X=1.805 $Y=0.49 $X2=0
+ $Y2=0
cc_263 N_A_32_297#_c_268_n N_VGND_c_523_n 0.00878037f $X=2.38 $Y=0.74 $X2=0
+ $Y2=0
cc_264 A_122_297# N_VPWR_c_375_n 0.0143816f $X=0.61 $Y=1.485 $X2=0 $Y2=0
cc_265 A_238_297# N_VPWR_c_375_n 0.00761629f $X=1.19 $Y=1.485 $X2=0 $Y2=0
cc_266 A_332_297# N_VPWR_c_375_n 0.00520913f $X=1.66 $Y=1.485 $X2=0 $Y2=0
cc_267 N_VPWR_c_375_n N_X_M1000_d 0.00370124f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_c_375_n N_X_M1012_d 0.00370124f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_382_n N_X_c_480_n 0.0149311f $X=3.2 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_375_n N_X_c_480_n 0.00955092f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_M1009_s N_X_c_437_n 0.00187091f $X=3.18 $Y=1.485 $X2=0 $Y2=0
cc_272 N_VPWR_c_377_n N_X_c_437_n 0.0143191f $X=3.325 $Y=1.96 $X2=0 $Y2=0
cc_273 N_VPWR_c_384_n N_X_c_484_n 0.0149311f $X=4.14 $Y=2.72 $X2=0 $Y2=0
cc_274 N_VPWR_c_375_n N_X_c_484_n 0.00955092f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_M1015_s N_X_c_438_n 0.00359214f $X=4.12 $Y=1.485 $X2=0 $Y2=0
cc_276 N_VPWR_c_379_n N_X_c_438_n 0.0187873f $X=4.265 $Y=1.96 $X2=0 $Y2=0
cc_277 N_X_c_430_n N_VGND_M1004_s 0.00251047f $X=3.58 $Y=0.815 $X2=0 $Y2=0
cc_278 N_X_c_432_n N_VGND_M1011_s 2.28588e-19 $X=4.21 $Y=0.815 $X2=0 $Y2=0
cc_279 N_X_c_435_n N_VGND_M1011_s 0.00344973f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_280 N_X_c_445_n N_VGND_c_513_n 0.0140037f $X=2.855 $Y=0.485 $X2=0 $Y2=0
cc_281 N_X_c_445_n N_VGND_c_514_n 0.0177813f $X=2.855 $Y=0.485 $X2=0 $Y2=0
cc_282 N_X_c_430_n N_VGND_c_514_n 0.0127273f $X=3.58 $Y=0.815 $X2=0 $Y2=0
cc_283 N_X_c_435_n N_VGND_c_515_n 0.00225104f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_284 N_X_c_432_n N_VGND_c_516_n 0.00177288f $X=4.21 $Y=0.815 $X2=0 $Y2=0
cc_285 N_X_c_435_n N_VGND_c_516_n 0.0120207f $X=4.347 $Y=0.905 $X2=0 $Y2=0
cc_286 N_X_c_445_n N_VGND_c_519_n 0.0153475f $X=2.855 $Y=0.485 $X2=0 $Y2=0
cc_287 N_X_c_430_n N_VGND_c_519_n 0.00266636f $X=3.58 $Y=0.815 $X2=0 $Y2=0
cc_288 N_X_c_430_n N_VGND_c_521_n 0.00198695f $X=3.58 $Y=0.815 $X2=0 $Y2=0
cc_289 N_X_c_463_n N_VGND_c_521_n 0.0231806f $X=3.795 $Y=0.39 $X2=0 $Y2=0
cc_290 N_X_c_432_n N_VGND_c_521_n 0.00254521f $X=4.21 $Y=0.815 $X2=0 $Y2=0
cc_291 N_X_M1002_d N_VGND_c_523_n 0.00607585f $X=2.67 $Y=0.235 $X2=0 $Y2=0
cc_292 N_X_M1007_d N_VGND_c_523_n 0.00304143f $X=3.61 $Y=0.235 $X2=0 $Y2=0
cc_293 N_X_c_445_n N_VGND_c_523_n 0.00940698f $X=2.855 $Y=0.485 $X2=0 $Y2=0
cc_294 N_X_c_430_n N_VGND_c_523_n 0.00972452f $X=3.58 $Y=0.815 $X2=0 $Y2=0
cc_295 N_X_c_463_n N_VGND_c_523_n 0.0143352f $X=3.795 $Y=0.39 $X2=0 $Y2=0
cc_296 N_X_c_432_n N_VGND_c_523_n 0.00509281f $X=4.21 $Y=0.815 $X2=0 $Y2=0
cc_297 N_X_c_435_n N_VGND_c_523_n 0.00444357f $X=4.347 $Y=0.905 $X2=0 $Y2=0
