* File: sky130_fd_sc_hdll__and2b_4.spice
* Created: Thu Aug 27 18:57:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2b_4.pex.spice"
.subckt sky130_fd_sc_hdll__and2b_4  VNB VPB B A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* B	B
* VPB	VPB
* VNB	VNB
MM1008 A_119_47# N_A_33_199#_M1008_g N_A_27_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.2015 PD=0.86 PS=1.92 NRD=9.228 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B_M1003_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.156
+ AS=0.06825 PD=1.13 PS=0.86 NRD=23.076 NRS=9.228 M=1 R=4.33333 SA=75000.6
+ SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1003_d N_A_27_47#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.156 AS=0.10725 PD=1.13 PS=0.98 NRD=13.836 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_27_47#_M1004_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=8.304 NRS=0.912 M=1 R=4.33333
+ SA=75001.7 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1004_d N_A_27_47#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.1235 PD=0.98 PS=1.03 NRD=0.912 NRS=9.228 M=1 R=4.33333
+ SA=75002.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_27_47#_M1012_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.142453 AS=0.1235 PD=1.28178 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333
+ SA=75002.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_A_33_199#_M1006_d N_A_N_M1006_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0920467 PD=1.46 PS=0.828224 NRD=11.424 NRS=46.896 M=1 R=2.8
+ SA=75003.3 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1005 N_A_27_47#_M1005_d N_A_33_199#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_B_M1000_g N_A_27_47#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.195 AS=0.145 PD=1.39 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1000_d N_A_27_47#_M1001_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.195 AS=0.16 PD=1.39 PS=1.32 NRD=9.8303 NRS=6.8753 M=1 R=5.55556
+ SA=90001.2 SB=90001.9 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_27_47#_M1007_g N_X_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.16 PD=1.29 PS=1.32 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.7 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1007_d N_A_27_47#_M1011_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.2 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1013_d N_A_27_47#_M1013_g N_X_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.229366 AS=0.145 PD=1.93662 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.7 SB=90000.4 A=0.18 P=2.36 MULT=1
MM1010 N_A_33_199#_M1010_d N_A_N_M1010_g N_VPWR_M1013_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1344 AS=0.0963338 PD=1.48 PS=0.81338 NRD=25.7873 NRS=81.7747 M=1
+ R=2.33333 SA=90003.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__and2b_4.pxi.spice"
*
.ends
*
*
