* File: sky130_fd_sc_hdll__mux2_4.pex.spice
* Created: Wed Sep  2 08:34:37 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%S 1 3 4 6 9 11 12 14 16 17 18 20 25 27 32
+ 33
r94 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.51
+ $Y=1.16 $X2=3.51 $Y2=1.16
r95 27 34 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.965 $Y=1.16 $X2=3.05
+ $Y2=1.16
r96 27 33 15.6453 $w=3.28e-07 $l=4.48e-07 $layer=LI1_cond $X=3.062 $Y=1.16
+ $X2=3.51 $Y2=1.16
r97 27 34 0.41907 $w=3.28e-07 $l=1.2e-08 $layer=LI1_cond $X=3.062 $Y=1.16
+ $X2=3.05 $Y2=1.16
r98 22 25 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=1.16
+ $X2=0.705 $Y2=1.16
r99 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r100 20 27 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.995
+ $X2=2.965 $Y2=1.16
r101 19 20 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=2.965 $Y=0.805
+ $X2=2.965 $Y2=0.995
r102 17 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.88 $Y=0.72
+ $X2=2.965 $Y2=0.805
r103 17 18 136.353 $w=1.68e-07 $l=2.09e-06 $layer=LI1_cond $X=2.88 $Y=0.72
+ $X2=0.79 $Y2=0.72
r104 16 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.705 $Y=0.995
+ $X2=0.705 $Y2=1.16
r105 15 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.705 $Y=0.805
+ $X2=0.79 $Y2=0.72
r106 15 16 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.705 $Y=0.805
+ $X2=0.705 $Y2=0.995
r107 12 32 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.595 $Y2=1.202
r108 12 14 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.62 $Y=0.995
+ $X2=3.62 $Y2=0.56
r109 9 32 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.595 $Y=1.41
+ $X2=3.595 $Y2=1.202
r110 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.595 $Y=1.41
+ $X2=3.595 $Y2=1.985
r111 4 23 38.578 $w=2.95e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.54 $Y2=1.16
r112 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r113 1 23 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.54 $Y2=1.16
r114 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A_27_47# 1 2 7 9 10 12 14 17 19 23 27 30
c50 23 0 1.19188e-19 $X=1.045 $Y=1.16
r51 27 29 8.74048 $w=2.53e-07 $l=1.65e-07 $layer=LI1_cond $X=0.217 $Y=0.46
+ $X2=0.217 $Y2=0.625
r52 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.045
+ $Y=1.16 $X2=1.045 $Y2=1.16
r53 21 23 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.07 $Y=1.495
+ $X2=1.07 $Y2=1.16
r54 20 30 2.15711 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.58
+ $X2=0.217 $Y2=1.58
r55 19 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.96 $Y=1.58
+ $X2=1.07 $Y2=1.495
r56 19 20 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=0.96 $Y=1.58
+ $X2=0.345 $Y2=1.58
r57 15 30 4.27425 $w=2.12e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.58
r58 15 17 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=1.665
+ $X2=0.217 $Y2=1.96
r59 14 30 4.27425 $w=2.12e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.175 $Y=1.495
+ $X2=0.217 $Y2=1.58
r60 14 29 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=0.175 $Y=1.495
+ $X2=0.175 $Y2=0.625
r61 10 24 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.07 $Y2=1.16
r62 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r63 7 24 48.1208 $w=2.95e-07 $l=2.73861e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.07 $Y2=1.16
r64 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41 $X2=1.02
+ $Y2=1.985
r65 2 17 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
r66 1 27 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A0 1 3 4 6 7 8 9 10 15
c33 15 0 1.43803e-19 $X=1.71 $Y=1.16
r34 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.71
+ $Y=1.16 $X2=1.71 $Y2=1.16
r35 9 10 11.3574 $w=3.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.622 $Y=1.19
+ $X2=1.622 $Y2=1.53
r36 9 15 1.00212 $w=3.43e-07 $l=3e-08 $layer=LI1_cond $X=1.622 $Y=1.19 $X2=1.622
+ $Y2=1.16
r37 7 14 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=1.93 $Y=1.16 $X2=1.71
+ $Y2=1.16
r38 7 8 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.93 $Y=1.16
+ $X2=2.03 $Y2=1.202
r39 4 8 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.055 $Y=0.995
+ $X2=2.03 $Y2=1.202
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.055 $Y=0.995
+ $X2=2.055 $Y2=0.56
r41 1 8 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.03 $Y=1.41
+ $X2=2.03 $Y2=1.202
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.03 $Y=1.41 $X2=2.03
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A1 1 3 4 6 7 11 13
c31 1 0 1.43803e-19 $X=2.55 $Y=1.41
r32 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5
+ $Y=1.16 $X2=2.5 $Y2=1.16
r33 7 11 15.0167 $w=3.28e-07 $l=4.3e-07 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=2.5
+ $Y2=1.16
r34 7 13 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=1.16 $X2=2.065
+ $Y2=1.16
r35 4 10 38.578 $w=2.95e-07 $l=1.88348e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.525 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.575 $Y=0.995
+ $X2=2.575 $Y2=0.56
r37 1 10 48.1208 $w=2.95e-07 $l=2.62202e-07 $layer=POLY_cond $X=2.55 $Y=1.41
+ $X2=2.525 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.55 $Y=1.41 $X2=2.55
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A_424_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 35 40 41 42 44 46 52 55 64
c136 64 0 1.54761e-19 $X=5.475 $Y=1.202
r137 64 65 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.202
+ $X2=5.5 $Y2=1.202
r138 61 62 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=5.005 $Y=1.202
+ $X2=5.03 $Y2=1.202
r139 60 61 58.1274 $w=3.69e-07 $l=4.45e-07 $layer=POLY_cond $X=4.56 $Y=1.202
+ $X2=5.005 $Y2=1.202
r140 59 60 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.535 $Y=1.202
+ $X2=4.56 $Y2=1.202
r141 56 57 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=4.065 $Y=1.202
+ $X2=4.09 $Y2=1.202
r142 53 64 27.4309 $w=3.69e-07 $l=2.1e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.475 $Y2=1.202
r143 53 62 30.6965 $w=3.69e-07 $l=2.35e-07 $layer=POLY_cond $X=5.265 $Y=1.202
+ $X2=5.03 $Y2=1.202
r144 52 53 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.265
+ $Y=1.16 $X2=5.265 $Y2=1.16
r145 50 59 57.4743 $w=3.69e-07 $l=4.4e-07 $layer=POLY_cond $X=4.095 $Y=1.202
+ $X2=4.535 $Y2=1.202
r146 50 57 0.653117 $w=3.69e-07 $l=5e-09 $layer=POLY_cond $X=4.095 $Y=1.202
+ $X2=4.09 $Y2=1.202
r147 49 52 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.095 $Y=1.16
+ $X2=5.265 $Y2=1.16
r148 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.095
+ $Y=1.16 $X2=4.095 $Y2=1.16
r149 47 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=1.16
+ $X2=3.9 $Y2=1.16
r150 47 49 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.985 $Y=1.16
+ $X2=4.095 $Y2=1.16
r151 45 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=1.245 $X2=3.9
+ $Y2=1.16
r152 45 46 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=3.9 $Y=1.245
+ $X2=3.9 $Y2=1.595
r153 44 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.9 $Y=1.075 $X2=3.9
+ $Y2=1.16
r154 43 44 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.9 $Y=0.825
+ $X2=3.9 $Y2=1.075
r155 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=0.74
+ $X2=3.9 $Y2=0.825
r156 41 42 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.815 $Y=0.74
+ $X2=3.43 $Y2=0.74
r157 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.345 $Y=0.655
+ $X2=3.43 $Y2=0.74
r158 39 40 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.345 $Y=0.465
+ $X2=3.345 $Y2=0.655
r159 35 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.815 $Y=1.68
+ $X2=3.9 $Y2=1.595
r160 35 37 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=3.815 $Y=1.68
+ $X2=2.295 $Y2=1.68
r161 31 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.26 $Y=0.38
+ $X2=3.345 $Y2=0.465
r162 31 33 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.26 $Y=0.38
+ $X2=2.29 $Y2=0.38
r163 28 65 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.5 $Y=0.995
+ $X2=5.5 $Y2=1.202
r164 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.5 $Y=0.995
+ $X2=5.5 $Y2=0.56
r165 25 64 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.202
r166 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.985
r167 22 62 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.03 $Y2=1.202
r168 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.03 $Y2=0.56
r169 19 61 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.202
r170 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.985
r171 16 60 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.56 $Y=0.995
+ $X2=4.56 $Y2=1.202
r172 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.56 $Y=0.995
+ $X2=4.56 $Y2=0.56
r173 13 59 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.202
r174 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.535 $Y=1.41
+ $X2=4.535 $Y2=1.985
r175 10 57 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=1.202
r176 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.09 $Y=0.995
+ $X2=4.09 $Y2=0.56
r177 7 56 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.065 $Y=1.41
+ $X2=4.065 $Y2=1.202
r178 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.065 $Y=1.41
+ $X2=4.065 $Y2=1.985
r179 2 37 600 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=2.12
+ $Y=1.485 $X2=2.295 $Y2=1.68
r180 1 33 182 $w=1.7e-07 $l=2.20907e-07 $layer=licon1_NDIFF $count=1 $X=2.13
+ $Y=0.235 $X2=2.29 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%VPWR 1 2 3 4 15 19 21 23 25 27 32 40 45 51
+ 54 61 65
r83 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r84 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r85 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r86 54 57 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.805 $Y=2.34
+ $X2=3.805 $Y2=2.72
r87 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 49 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r89 49 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r91 46 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=4.745 $Y2=2.72
r92 46 48 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.935 $Y=2.72
+ $X2=5.29 $Y2=2.72
r93 45 64 5.23377 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.737 $Y2=2.72
r94 45 48 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=2.72
+ $X2=5.29 $Y2=2.72
r95 44 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r96 44 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r98 41 57 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.995 $Y=2.72
+ $X2=3.805 $Y2=2.72
r99 41 43 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.995 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 40 61 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.745 $Y2=2.72
r101 40 43 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.37 $Y2=2.72
r102 39 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r103 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 36 39 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r105 36 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r106 35 38 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r108 33 51 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.692 $Y2=2.72
r109 33 35 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=1.15 $Y2=2.72
r110 32 57 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.805 $Y2=2.72
r111 32 38 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=2.72
+ $X2=3.45 $Y2=2.72
r112 27 51 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.692 $Y2=2.72
r113 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r114 25 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r116 21 64 2.96292 $w=3.8e-07 $l=1.07912e-07 $layer=LI1_cond $X=5.685 $Y=2.635
+ $X2=5.737 $Y2=2.72
r117 21 23 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=5.685 $Y=2.635
+ $X2=5.685 $Y2=2
r118 17 61 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.745 $Y=2.635
+ $X2=4.745 $Y2=2.72
r119 17 19 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.745 $Y=2.635
+ $X2=4.745 $Y2=2
r120 13 51 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.692 $Y=2.635
+ $X2=0.692 $Y2=2.72
r121 13 15 20.6141 $w=3.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.692 $Y=2.635
+ $X2=0.692 $Y2=2
r122 4 23 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2
r123 3 19 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=2
r124 2 54 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.685
+ $Y=1.485 $X2=3.83 $Y2=2.34
r125 1 15 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A_222_297# 1 2 9 12
c23 1 0 1.19188e-19 $X=1.11 $Y=1.485
r24 12 14 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.24 $Y=2.02
+ $X2=1.24 $Y2=2.36
r25 7 14 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=1.44 $Y=2.36 $X2=1.24
+ $Y2=2.36
r26 7 9 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.44 $Y=2.36
+ $X2=2.805 $Y2=2.36
r27 2 9 600 $w=1.7e-07 $l=9.53939e-07 $layer=licon1_PDIFF $count=1 $X=2.64
+ $Y=1.485 $X2=2.805 $Y2=2.36
r28 1 12 300 $w=1.7e-07 $l=6.11964e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.485 $X2=1.275 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%A_334_297# 1 2 7 13
r24 11 13 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.36 $Y=2.105
+ $X2=3.36 $Y2=2.3
r25 7 11 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.275 $Y=2.02
+ $X2=3.36 $Y2=2.105
r26 7 9 96.5562 $w=1.68e-07 $l=1.48e-06 $layer=LI1_cond $X=3.275 $Y=2.02
+ $X2=1.795 $Y2=2.02
r27 2 13 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=3.235
+ $Y=1.485 $X2=3.36 $Y2=2.3
r28 1 9 600 $w=1.7e-07 $l=5.94222e-07 $layer=licon1_PDIFF $count=1 $X=1.67
+ $Y=1.485 $X2=1.795 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35 37
+ 38 39 40 41 47 48 50 56
r76 48 56 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.765 $Y=1.575
+ $X2=5.765 $Y2=1.53
r77 47 50 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=5.765 $Y=0.805
+ $X2=5.765 $Y2=0.85
r78 41 48 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.765 $Y=1.66
+ $X2=5.765 $Y2=1.575
r79 41 56 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=5.765 $Y=1.51
+ $X2=5.765 $Y2=1.53
r80 40 41 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.765 $Y=1.19
+ $X2=5.765 $Y2=1.51
r81 39 47 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.765 $Y=0.72
+ $X2=5.765 $Y2=0.805
r82 39 40 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=5.765 $Y=0.87
+ $X2=5.765 $Y2=1.19
r83 39 50 1.00212 $w=2.28e-07 $l=2e-08 $layer=LI1_cond $X=5.765 $Y=0.87
+ $X2=5.765 $Y2=0.85
r84 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=1.66
+ $X2=5.24 $Y2=1.66
r85 35 41 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.65 $Y=1.66
+ $X2=5.765 $Y2=1.66
r86 35 36 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.65 $Y=1.66
+ $X2=5.325 $Y2=1.66
r87 34 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.325 $Y=0.72
+ $X2=5.24 $Y2=0.72
r88 33 39 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.65 $Y=0.72
+ $X2=5.765 $Y2=0.72
r89 33 34 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=5.65 $Y=0.72
+ $X2=5.325 $Y2=0.72
r90 29 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=1.745
+ $X2=5.24 $Y2=1.66
r91 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.24 $Y=1.745
+ $X2=5.24 $Y2=1.96
r92 25 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.635
+ $X2=5.24 $Y2=0.72
r93 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.24 $Y=0.635
+ $X2=5.24 $Y2=0.42
r94 23 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=1.66
+ $X2=5.24 $Y2=1.66
r95 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.155 $Y=1.66
+ $X2=4.385 $Y2=1.66
r96 21 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.155 $Y=0.72
+ $X2=5.24 $Y2=0.72
r97 21 22 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.155 $Y=0.72
+ $X2=4.385 $Y2=0.72
r98 17 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.3 $Y=1.745
+ $X2=4.385 $Y2=1.66
r99 17 19 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.3 $Y=1.745
+ $X2=4.3 $Y2=1.96
r100 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.3 $Y=0.635
+ $X2=4.385 $Y2=0.72
r101 13 15 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.3 $Y=0.635
+ $X2=4.3 $Y2=0.42
r102 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=1.485 $X2=5.24 $Y2=1.96
r103 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.155
+ $Y=1.485 $X2=4.3 $Y2=1.96
r104 2 27 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.235 $X2=5.24 $Y2=0.42
r105 1 15 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.165
+ $Y=0.235 $X2=4.3 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_4%VGND 1 2 3 4 13 15 20 28 33 40 47 54 60 61
c82 47 0 1.54761e-19 $X=3.91 $Y=0
r83 60 63 11.2524 $w=4.12e-07 $l=3.8e-07 $layer=LI1_cond $X=5.737 $Y=0 $X2=5.737
+ $Y2=0.38
r84 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r85 54 57 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.745 $Y=0 $X2=4.745
+ $Y2=0.38
r86 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r87 47 50 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.805
+ $Y2=0.38
r88 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r89 40 43 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r90 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r91 37 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r92 37 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.83
+ $Y2=0
r93 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r94 34 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=4.745
+ $Y2=0
r95 34 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=4.935 $Y=0 $X2=5.29
+ $Y2=0
r96 33 60 5.95845 $w=1.7e-07 $l=2.42e-07 $layer=LI1_cond $X=5.495 $Y=0 $X2=5.737
+ $Y2=0
r97 33 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.495 $Y=0 $X2=5.29
+ $Y2=0
r98 32 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r99 32 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r100 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r101 29 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.805
+ $Y2=0
r102 29 31 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.995 $Y=0
+ $X2=4.37 $Y2=0
r103 28 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.555 $Y=0 $X2=4.745
+ $Y2=0
r104 28 31 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=0
+ $X2=4.37 $Y2=0
r105 27 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r106 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r107 24 27 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r108 24 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r109 23 26 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.45
+ $Y2=0
r110 23 24 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r111 21 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r112 21 23 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r113 20 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.615 $Y=0 $X2=3.805
+ $Y2=0
r114 20 26 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.615 $Y=0
+ $X2=3.45 $Y2=0
r115 15 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r116 15 17 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r117 13 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r118 13 17 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r119 4 63 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.38
r120 3 57 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=0.235 $X2=4.77 $Y2=0.38
r121 2 50 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.235 $X2=3.83 $Y2=0.38
r122 1 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

