* File: sky130_fd_sc_hdll__dlygate4sd3_1.spice
* Created: Thu Aug 27 19:06:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dlygate4sd3_1.pex.spice"
.subckt sky130_fd_sc_hdll__dlygate4sd3_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_27_47#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0588 AS=0.126 PD=0.7 PS=1.44 NRD=1.428 NRS=9.996 M=1 R=2.8 SA=75000.2
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1003 N_A_273_47#_M1003_d N_A_27_47#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.5
+ W=0.42 AD=0.1092 AS=0.0588 PD=1.36 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1006 N_VGND_M1006_d N_A_273_47#_M1006_g N_A_379_93#_M1006_s VNB NSHORT L=0.5
+ W=0.42 AD=0.0965607 AS=0.1092 PD=0.828224 PS=1.36 NRD=49.968 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1005 N_X_M1005_d N_A_379_93#_M1005_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.149439 PD=1.84 PS=1.28178 NRD=0.912 NRS=11.988 M=1 R=4.33333
+ SA=75000.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0588 AS=0.1134 PD=0.7 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1007 N_A_273_47#_M1007_d N_A_27_47#_M1007_g N_VPWR_M1002_d VPB PHIGHVT L=0.5
+ W=0.42 AD=0.1092 AS=0.0588 PD=1.36 PS=0.7 NRD=0 NRS=0 M=1 R=0.84 SA=250000
+ SB=250000 A=0.21 P=1.84 MULT=1
MM1000 N_VPWR_M1000_d N_A_273_47#_M1000_g N_A_379_93#_M1000_s VPB PHIGHVT L=0.5
+ W=0.42 AD=0.0980493 AS=0.1092 PD=0.81338 PS=1.36 NRD=28.1316 NRS=0 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1001 N_X_M1001_d N_A_379_93#_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.233451 PD=2.54 PS=1.93662 NRD=0.9653 NRS=6.8753 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_61 VPB 0 1.21278e-19 $X=0.14 $Y=2.635
*
.include "sky130_fd_sc_hdll__dlygate4sd3_1.pxi.spice"
*
.ends
*
*
