# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand3b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.430000 1.075000 0.830000 1.275000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.150000 1.075000 3.440000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.890000 1.275000 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA  0.429500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.630000  0.085000 0.940000 0.905000 ;
        RECT 1.710000  0.085000 1.960000 0.545000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.465700 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.630000 1.835000 0.940000 2.635000 ;
        RECT 1.710000 2.175000 1.880000 2.635000 ;
        RECT 2.650000 2.175000 2.900000 2.635000 ;
        RECT 3.090000 2.175000 3.390000 2.635000 ;
        RECT 4.160000 2.175000 4.450000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.110500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.110000 1.785000 4.490000 1.955000 ;
        RECT 1.110000 1.955000 2.430000 2.005000 ;
        RECT 1.110000 2.005000 1.490000 2.465000 ;
        RECT 2.050000 2.005000 2.430000 2.465000 ;
        RECT 3.560000 0.635000 4.490000 0.905000 ;
        RECT 3.560000 1.955000 4.490000 2.005000 ;
        RECT 3.560000 2.005000 3.860000 2.465000 ;
        RECT 4.250000 0.905000 4.490000 1.785000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.410000 0.655000 ;
      RECT 0.090000 0.655000 0.260000 1.445000 ;
      RECT 0.090000 1.445000 4.000000 1.615000 ;
      RECT 0.090000 1.615000 0.260000 2.065000 ;
      RECT 0.090000 2.065000 0.410000 2.465000 ;
      RECT 1.110000 0.255000 1.490000 0.715000 ;
      RECT 1.110000 0.715000 3.000000 0.905000 ;
      RECT 2.200000 0.255000 4.450000 0.465000 ;
      RECT 2.200000 0.635000 3.000000 0.715000 ;
      RECT 3.220000 0.465000 3.390000 0.905000 ;
      RECT 3.670000 1.075000 4.000000 1.445000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3b_2
