* File: sky130_fd_sc_hdll__sdlclkp_4.pex.spice
* Created: Wed Sep  2 08:52:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%SCE 2 3 5 8 10 11 19
c30 8 0 1.073e-19 $X=0.52 $Y=0.445
c31 3 0 1.54309e-19 $X=0.495 $Y=1.77
r32 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r33 15 18 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r34 10 11 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=0.215 $Y=1.16
+ $X2=0.215 $Y2=1.53
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r36 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r37 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r38 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r39 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r40 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r41 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GATE 2 3 5 8 10 11 16 17
c46 17 0 3.16691e-19 $X=0.99 $Y=1.16
c47 16 0 9.53816e-20 $X=0.99 $Y=1.16
c48 10 0 1.54309e-19 $X=1.155 $Y=1.53
c49 3 0 1.23918e-19 $X=0.905 $Y=1.77
r50 16 18 37.8338 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=1.16
+ $X2=0.99 $Y2=1.325
r51 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=1.16 $X2=0.99 $Y2=1.16
r52 10 11 9.0076 $w=4.33e-07 $l=3.4e-07 $layer=LI1_cond $X=1.122 $Y=1.53
+ $X2=1.122 $Y2=1.87
r53 10 17 7.20187 $w=5.58e-07 $l=2.85e-07 $layer=LI1_cond $X=1.1 $Y=1.445
+ $X2=1.1 $Y2=1.16
r54 6 16 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.16
r55 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.99 $Y=0.995 $X2=0.99
+ $Y2=0.445
r56 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=2.165
r57 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.905 $Y=1.67 $X2=0.905
+ $Y2=1.77
r58 2 18 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.905 $Y=1.67
+ $X2=0.905 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_280_21# 1 2 9 11 13 14 17 20 25 26 28
+ 34 36 39 41 43 47 48 53 54 57 60
c172 57 0 1.562e-19 $X=1.765 $Y=1.53
c173 54 0 1.83164e-19 $X=1.91 $Y=1.53
c174 47 0 1.91701e-19 $X=1.74 $Y=1.325
c175 34 0 1.88819e-19 $X=4.677 $Y=1.495
c176 25 0 3.03377e-20 $X=1.565 $Y=0.87
c177 9 0 2.22956e-20 $X=1.475 $Y=0.415
r178 68 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.74 $X2=1.93 $Y2=1.74
r179 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.745 $Y=1.53
+ $X2=4.745 $Y2=1.53
r180 57 69 4.97379 $w=5.03e-07 $l=2.1e-07 $layer=LI1_cond $X=1.762 $Y=1.53
+ $X2=1.762 $Y2=1.74
r181 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.765 $Y=1.53
+ $X2=1.765 $Y2=1.53
r182 54 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.91 $Y=1.53
+ $X2=1.765 $Y2=1.53
r183 53 60 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.6 $Y=1.53
+ $X2=4.745 $Y2=1.53
r184 53 54 3.3292 $w=1.4e-07 $l=2.69e-06 $layer=MET1_cond $X=4.6 $Y=1.53
+ $X2=1.91 $Y2=1.53
r185 47 57 4.85537 $w=5.03e-07 $l=2.05e-07 $layer=LI1_cond $X=1.762 $Y=1.325
+ $X2=1.762 $Y2=1.53
r186 46 47 3.4935 $w=5.03e-07 $l=1.2e-07 $layer=LI1_cond $X=1.74 $Y=1.205
+ $X2=1.74 $Y2=1.325
r187 41 43 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=5.12 $Y=0.615
+ $X2=5.12 $Y2=0.465
r188 37 61 3.79964 $w=2.5e-07 $l=1.53e-07 $layer=LI1_cond $X=4.83 $Y=1.62
+ $X2=4.677 $Y2=1.62
r189 37 39 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.83 $Y=1.62
+ $X2=5.21 $Y2=1.62
r190 36 48 3.17288 $w=2.97e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.685 $Y=1.105
+ $X2=4.677 $Y2=1.19
r191 35 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.685 $Y=0.7
+ $X2=5.12 $Y2=0.7
r192 35 36 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=4.685 $Y=0.785
+ $X2=4.685 $Y2=1.105
r193 34 61 3.10428 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=4.677 $Y=1.495
+ $X2=4.677 $Y2=1.62
r194 33 48 3.17288 $w=2.97e-07 $l=8.5e-08 $layer=LI1_cond $X=4.677 $Y=1.275
+ $X2=4.677 $Y2=1.19
r195 33 34 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=4.677 $Y=1.275
+ $X2=4.677 $Y2=1.495
r196 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.4
+ $Y=1.19 $X2=4.4 $Y2=1.19
r197 28 48 3.41642 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.525 $Y=1.19
+ $X2=4.677 $Y2=1.19
r198 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.525 $Y=1.19
+ $X2=4.4 $Y2=1.19
r199 26 63 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=1.565 $Y=0.87
+ $X2=1.475 $Y2=0.87
r200 25 46 9.89919 $w=3.88e-07 $l=3.35e-07 $layer=LI1_cond $X=1.66 $Y=0.87
+ $X2=1.66 $Y2=1.205
r201 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=0.87 $X2=1.565 $Y2=0.87
r202 18 31 34.1407 $w=3.26e-07 $l=1.46969e-07 $layer=POLY_cond $X=4.4 $Y=1.055
+ $X2=4.425 $Y2=1.19
r203 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.4 $Y=1.055
+ $X2=4.4 $Y2=0.445
r204 14 31 46.5577 $w=3.26e-07 $l=2.73861e-07 $layer=POLY_cond $X=4.375 $Y=1.44
+ $X2=4.425 $Y2=1.19
r205 14 17 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.375 $Y=1.44
+ $X2=4.375 $Y2=1.835
r206 11 68 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.015 $Y=1.99
+ $X2=1.955 $Y2=1.74
r207 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.015 $Y=1.99
+ $X2=2.015 $Y2=2.275
r208 7 63 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.475 $Y=0.735
+ $X2=1.475 $Y2=0.87
r209 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.475 $Y=0.735
+ $X2=1.475 $Y2=0.415
r210 2 39 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.065
+ $Y=1.515 $X2=5.21 $Y2=1.66
r211 1 43 182 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_NDIFF $count=1 $X=4.945
+ $Y=0.235 $X2=5.08 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_277_243# 1 2 8 9 11 12 13 16 18 21 24
+ 28 30 31 37 38 41 42 43
c124 42 0 2.22956e-20 $X=2.11 $Y=0.87
c125 37 0 5.69068e-21 $X=4.235 $Y=0.85
c126 28 0 1.17835e-19 $X=4.14 $Y=1.66
c127 18 0 2.62261e-20 $X=2.075 $Y=1.215
c128 8 0 3.27168e-20 $X=1.485 $Y=1.89
r129 41 44 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=0.87
+ $X2=2.135 $Y2=1.035
r130 41 43 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.135 $Y=0.87
+ $X2=2.135 $Y2=0.705
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.11
+ $Y=0.87 $X2=2.11 $Y2=0.87
r132 38 50 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=4.107 $Y=0.85
+ $X2=4.107 $Y2=0.935
r133 38 49 2.91128 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=4.107 $Y=0.85
+ $X2=4.107 $Y2=0.765
r134 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.235 $Y=0.85
+ $X2=4.235 $Y2=0.85
r135 33 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.275 $Y=0.85
+ $X2=2.275 $Y2=0.85
r136 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.42 $Y=0.85
+ $X2=2.275 $Y2=0.85
r137 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.09 $Y=0.85
+ $X2=4.235 $Y2=0.85
r138 30 31 2.06683 $w=1.4e-07 $l=1.67e-06 $layer=MET1_cond $X=4.09 $Y=0.85
+ $X2=2.42 $Y2=0.85
r139 25 28 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.98 $Y=1.66
+ $X2=4.14 $Y2=1.66
r140 24 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.98 $Y=1.575
+ $X2=3.98 $Y2=1.66
r141 24 50 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.98 $Y=1.575
+ $X2=3.98 $Y2=0.935
r142 21 49 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=4.06 $Y=0.465
+ $X2=4.06 $Y2=0.765
r143 18 44 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=2.075 $Y=1.215
+ $X2=2.075 $Y2=1.035
r144 16 43 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.05 $Y=0.415
+ $X2=2.05 $Y2=0.705
r145 12 18 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=1.975 $Y=1.29
+ $X2=2.075 $Y2=1.215
r146 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=1.975 $Y=1.29
+ $X2=1.585 $Y2=1.29
r147 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.99
+ $X2=1.485 $Y2=2.275
r148 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.485 $Y=1.89 $X2=1.485
+ $Y2=1.99
r149 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=1.485 $Y=1.365
+ $X2=1.585 $Y2=1.29
r150 7 8 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=1.485 $Y=1.365
+ $X2=1.485 $Y2=1.89
r151 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=4.015
+ $Y=1.515 $X2=4.14 $Y2=1.66
r152 1 21 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.14 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_505_315# 1 2 7 9 12 14 16 17 19 20 24
+ 28 30 34 41 42
c122 30 0 5.88603e-20 $X=5.565 $Y=2
c123 12 0 1.28601e-19 $X=2.76 $Y=0.445
r124 38 41 5.12956 $w=3.28e-07 $l=1.35e-07 $layer=LI1_cond $X=2.66 $Y=1.74
+ $X2=2.795 $Y2=1.74
r125 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.74 $X2=2.66 $Y2=1.74
r126 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.79
+ $Y=1.16 $X2=5.79 $Y2=1.16
r127 32 34 24.8598 $w=3.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.74 $Y=1.915
+ $X2=5.74 $Y2=1.16
r128 31 42 3.05 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.705 $Y=2
+ $X2=3.595 $Y2=1.86
r129 30 32 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.565 $Y=2
+ $X2=5.74 $Y2=1.915
r130 30 31 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=5.565 $Y=2
+ $X2=3.705 $Y2=2
r131 26 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.595 $Y=2.085
+ $X2=3.595 $Y2=1.86
r132 26 28 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.595 $Y=2.085
+ $X2=3.595 $Y2=2.205
r133 22 42 3.05 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.595 $Y=1.635
+ $X2=3.595 $Y2=1.86
r134 22 24 63.6463 $w=2.18e-07 $l=1.215e-06 $layer=LI1_cond $X=3.595 $Y=1.635
+ $X2=3.595 $Y2=0.42
r135 20 42 3.05 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.485 $Y=1.77
+ $X2=3.595 $Y2=1.86
r136 20 41 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.485 $Y=1.77
+ $X2=2.795 $Y2=1.77
r137 17 35 39.2524 $w=3.82e-07 $l=2.24332e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=5.87 $Y2=1.16
r138 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.01 $Y=0.995
+ $X2=6.01 $Y2=0.56
r139 14 35 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=5.985 $Y=1.41
+ $X2=5.87 $Y2=1.16
r140 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.985 $Y=1.41
+ $X2=5.985 $Y2=1.985
r141 10 39 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.76 $Y=1.575
+ $X2=2.68 $Y2=1.74
r142 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.76 $Y=1.575
+ $X2=2.76 $Y2=0.445
r143 7 39 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=2.625 $Y=1.99
+ $X2=2.68 $Y2=1.74
r144 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.625 $Y=1.99
+ $X2=2.625 $Y2=2.275
r145 2 28 600 $w=1.7e-07 $l=7.89177e-07 $layer=licon1_PDIFF $count=1 $X=3.475
+ $Y=1.485 $X2=3.62 $Y2=2.205
r146 1 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.235 $X2=3.62 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_310_47# 1 2 7 9 10 12 13 17 22 24 25
+ 27
c93 25 0 3.27168e-20 $X=2.7 $Y=1.185
c94 24 0 3.03377e-20 $X=2.615 $Y=0.995
r95 30 31 14.6301 $w=2.46e-07 $l=2.95e-07 $layer=LI1_cond $X=2.32 $Y=1.205
+ $X2=2.615 $Y2=1.205
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.18
+ $Y=1.16 $X2=3.18 $Y2=1.16
r97 25 31 4.2431 $w=3.8e-07 $l=9.44722e-08 $layer=LI1_cond $X=2.7 $Y=1.185
+ $X2=2.615 $Y2=1.205
r98 25 27 14.5572 $w=3.78e-07 $l=4.8e-07 $layer=LI1_cond $X=2.7 $Y=1.185
+ $X2=3.18 $Y2=1.185
r99 24 31 2.90119 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=2.615 $Y=0.995
+ $X2=2.615 $Y2=1.205
r100 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.615 $Y=0.535
+ $X2=2.615 $Y2=0.995
r101 21 30 2.90119 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.32 $Y=1.375
+ $X2=2.32 $Y2=1.205
r102 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.32 $Y=1.375
+ $X2=2.32 $Y2=2.125
r103 17 22 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.235 $Y=2.295
+ $X2=2.32 $Y2=2.125
r104 17 19 16.4393 $w=3.38e-07 $l=4.85e-07 $layer=LI1_cond $X=2.235 $Y=2.295
+ $X2=1.75 $Y2=2.295
r105 13 23 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.53 $Y=0.395
+ $X2=2.615 $Y2=0.535
r106 13 15 30.6632 $w=2.78e-07 $l=7.45e-07 $layer=LI1_cond $X=2.53 $Y=0.395
+ $X2=1.785 $Y2=0.395
r107 10 28 39.3952 $w=3.9e-07 $l=2.26164e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.265 $Y2=1.16
r108 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.56
r109 7 28 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.265 $Y2=1.16
r110 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.385 $Y=1.41
+ $X2=3.385 $Y2=1.985
r111 2 19 600 $w=1.7e-07 $l=3.2596e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=2.065 $X2=1.75 $Y2=2.315
r112 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.235 $X2=1.785 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%CLK 1 3 4 7 8 10 11 13 15 16 18 21 25 28
+ 39
c94 11 0 5.88603e-20 $X=6.455 $Y=1.41
c95 8 0 1.23841e-19 $X=6.37 $Y=0.995
c96 7 0 1.17835e-19 $X=4.975 $Y=1.835
c97 4 0 5.69068e-21 $X=4.975 $Y=1.44
r98 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.43
+ $Y=1.16 $X2=6.43 $Y2=1.16
r99 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.21
+ $Y=1.16 $X2=5.21 $Y2=1.16
r100 21 39 0.0224562 $w=2.3e-07 $l=3.5e-08 $layer=MET1_cond $X=5.16 $Y=1.19
+ $X2=5.125 $Y2=1.19
r101 21 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.2 $Y=1.19 $X2=5.2
+ $Y2=1.19
r102 19 28 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.245 $Y=1.16
+ $X2=6.43 $Y2=1.16
r103 18 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.245 $Y=1.19
+ $X2=6.245 $Y2=1.19
r104 16 21 0.141131 $w=2.3e-07 $l=1.85e-07 $layer=MET1_cond $X=5.345 $Y=1.19
+ $X2=5.16 $Y2=1.19
r105 15 18 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.1 $Y=1.19
+ $X2=6.245 $Y2=1.19
r106 15 16 0.934404 $w=1.4e-07 $l=7.55e-07 $layer=MET1_cond $X=6.1 $Y=1.19
+ $X2=5.345 $Y2=1.19
r107 11 27 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.455 $Y=1.41
+ $X2=6.455 $Y2=1.16
r108 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.455 $Y=1.41
+ $X2=6.455 $Y2=1.985
r109 8 27 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=6.37 $Y=0.995
+ $X2=6.455 $Y2=1.16
r110 8 10 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.37 $Y=0.995
+ $X2=6.37 $Y2=0.56
r111 4 24 47.9649 $w=4.43e-07 $l=3.24037e-07 $layer=POLY_cond $X=4.975 $Y=1.44
+ $X2=5.07 $Y2=1.16
r112 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.975 $Y=1.44
+ $X2=4.975 $Y2=1.835
r113 1 24 69.3486 $w=4.43e-07 $l=5.20481e-07 $layer=POLY_cond $X=4.87 $Y=0.73
+ $X2=5.07 $Y2=1.16
r114 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.87 $Y=0.73 $X2=4.87
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_1125_47# 1 2 9 11 13 16 18 20 23 25 27
+ 28 29 30 32 35 37 38 40 44 46 47 52 58 60
c155 60 0 5.46563e-20 $X=6.825 $Y=1.185
c156 35 0 1.27609e-19 $X=8.55 $Y=0.56
c157 29 0 1.64127e-19 $X=8.02 $Y=1.16
r158 66 67 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.895 $Y=1.217
+ $X2=7.92 $Y2=1.217
r159 65 66 64.997 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=7.45 $Y=1.217
+ $X2=7.895 $Y2=1.217
r160 64 65 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=7.425 $Y=1.217
+ $X2=7.45 $Y2=1.217
r161 61 62 3.65152 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=6.955 $Y=1.217
+ $X2=6.98 $Y2=1.217
r162 56 58 12.2649 $w=5.88e-07 $l=6.05e-07 $layer=LI1_cond $X=6.22 $Y=1.79
+ $X2=6.825 $Y2=1.79
r163 52 54 6.58539 $w=4.18e-07 $l=2.4e-07 $layer=LI1_cond $X=5.625 $Y=0.46
+ $X2=5.625 $Y2=0.7
r164 50 64 55.503 $w=3.3e-07 $l=3.8e-07 $layer=POLY_cond $X=7.045 $Y=1.217
+ $X2=7.425 $Y2=1.217
r165 50 62 9.49394 $w=3.3e-07 $l=6.5e-08 $layer=POLY_cond $X=7.045 $Y=1.217
+ $X2=6.98 $Y2=1.217
r166 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.045
+ $Y=1.16 $X2=7.045 $Y2=1.16
r167 47 60 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.91 $Y=1.185
+ $X2=6.825 $Y2=1.185
r168 47 49 6.33462 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=6.91 $Y=1.185
+ $X2=7.045 $Y2=1.185
r169 46 58 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.825 $Y=1.495
+ $X2=6.825 $Y2=1.79
r170 45 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=1.315
+ $X2=6.825 $Y2=1.185
r171 45 46 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.825 $Y=1.315
+ $X2=6.825 $Y2=1.495
r172 44 60 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.825 $Y=1.055
+ $X2=6.825 $Y2=1.185
r173 43 44 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.825 $Y=0.785
+ $X2=6.825 $Y2=1.055
r174 40 56 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.22 $Y=2.085
+ $X2=6.22 $Y2=1.79
r175 40 42 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=6.22 $Y=2.085 $X2=6.22
+ $Y2=2.125
r176 39 54 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.835 $Y=0.7
+ $X2=5.625 $Y2=0.7
r177 38 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.74 $Y=0.7
+ $X2=6.825 $Y2=0.785
r178 38 39 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.74 $Y=0.7
+ $X2=5.835 $Y2=0.7
r179 33 37 30.0832 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=8.55 $Y=1.025
+ $X2=8.525 $Y2=1.217
r180 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.55 $Y=1.025
+ $X2=8.55 $Y2=0.56
r181 30 37 30.0832 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=8.525 $Y=1.41
+ $X2=8.525 $Y2=1.217
r182 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.525 $Y=1.41
+ $X2=8.525 $Y2=1.985
r183 29 67 16.3418 $w=3.3e-07 $l=1.253e-07 $layer=POLY_cond $X=8.02 $Y=1.16
+ $X2=7.92 $Y2=1.217
r184 28 37 1.40033 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=8.425 $Y=1.16
+ $X2=8.525 $Y2=1.217
r185 28 29 89.9803 $w=2.7e-07 $l=4.05e-07 $layer=POLY_cond $X=8.425 $Y=1.16
+ $X2=8.02 $Y2=1.16
r186 25 67 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.92 $Y=1.41
+ $X2=7.92 $Y2=1.217
r187 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.92 $Y=1.41
+ $X2=7.92 $Y2=1.985
r188 21 66 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.895 $Y=1.025
+ $X2=7.895 $Y2=1.217
r189 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.895 $Y=1.025
+ $X2=7.895 $Y2=0.56
r190 18 65 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.45 $Y=1.41
+ $X2=7.45 $Y2=1.217
r191 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.45 $Y=1.41
+ $X2=7.45 $Y2=1.985
r192 14 64 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.425 $Y=1.025
+ $X2=7.425 $Y2=1.217
r193 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.425 $Y=1.025
+ $X2=7.425 $Y2=0.56
r194 11 62 16.9318 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.98 $Y=1.41
+ $X2=6.98 $Y2=1.217
r195 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.98 $Y=1.41
+ $X2=6.98 $Y2=1.985
r196 7 61 21.2229 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.955 $Y=1.025
+ $X2=6.955 $Y2=1.217
r197 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.955 $Y=1.025
+ $X2=6.955 $Y2=0.56
r198 2 42 600 $w=1.7e-07 $l=7.08802e-07 $layer=licon1_PDIFF $count=1 $X=6.075
+ $Y=1.485 $X2=6.22 $Y2=2.125
r199 1 52 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.625
+ $Y=0.235 $X2=5.75 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VPWR 1 2 3 4 5 6 7 22 24 30 34 36 38 43
+ 44 45 55 56 62 71 81 84 88 93 95 99
r118 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r119 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 90 93 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.75 $Y=2.53
+ $X2=5.915 $Y2=2.53
r121 90 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r122 86 88 6.56995 $w=5.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=3.895 $Y2=2.53
r123 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 84 88 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.265 $Y=2.72
+ $X2=3.895 $Y2=2.72
r125 83 84 11.8978 $w=7.28e-07 $l=2.2e-07 $layer=LI1_cond $X=3.045 $Y=2.44
+ $X2=3.265 $Y2=2.44
r126 80 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 79 83 0.901155 $w=7.28e-07 $l=5.5e-08 $layer=LI1_cond $X=2.99 $Y=2.44
+ $X2=3.045 $Y2=2.44
r128 79 81 15.0928 $w=7.28e-07 $l=4.15e-07 $layer=LI1_cond $X=2.99 $Y=2.44
+ $X2=2.575 $Y2=2.44
r129 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r130 74 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.97 $Y2=2.72
r131 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r132 71 98 4.11661 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=8.765 $Y=2.72
+ $X2=8.982 $Y2=2.72
r133 71 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.765 $Y=2.72
+ $X2=8.51 $Y2=2.72
r134 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r135 70 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r136 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r137 67 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.885 $Y=2.72
+ $X2=6.72 $Y2=2.72
r138 67 69 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=6.885 $Y=2.72
+ $X2=7.59 $Y2=2.72
r139 66 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r140 66 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r141 65 93 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=5.915 $Y2=2.72
r142 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r143 62 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.72 $Y2=2.72
r144 62 65 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.21 $Y2=2.72
r145 59 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.75 $Y2=2.72
r146 59 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 58 61 6.6328 $w=5.48e-07 $l=3.05e-07 $layer=LI1_cond $X=4.37 $Y=2.53
+ $X2=4.675 $Y2=2.53
r148 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r149 56 86 5.65419 $w=5.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.17 $Y=2.53
+ $X2=3.91 $Y2=2.53
r150 56 58 4.34938 $w=5.48e-07 $l=2e-07 $layer=LI1_cond $X=4.17 $Y=2.53 $X2=4.37
+ $Y2=2.53
r151 55 90 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.64 $Y=2.53
+ $X2=5.75 $Y2=2.53
r152 55 61 20.9857 $w=5.48e-07 $l=9.65e-07 $layer=LI1_cond $X=5.64 $Y=2.53
+ $X2=4.675 $Y2=2.53
r153 54 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r154 53 81 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=2.575 $Y2=2.72
r155 53 54 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r156 51 54 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r157 50 53 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r158 50 51 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r159 48 76 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r160 48 50 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r161 45 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r162 45 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r163 43 69 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.6 $Y=2.72 $X2=7.59
+ $Y2=2.72
r164 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.6 $Y=2.72
+ $X2=7.725 $Y2=2.72
r165 42 73 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.85 $Y=2.72
+ $X2=8.51 $Y2=2.72
r166 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.85 $Y=2.72
+ $X2=7.725 $Y2=2.72
r167 38 41 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.9 $Y=1.66 $X2=8.9
+ $Y2=2.34
r168 36 98 3.16808 $w=2.7e-07 $l=1.19143e-07 $layer=LI1_cond $X=8.9 $Y=2.635
+ $X2=8.982 $Y2=2.72
r169 36 41 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.9 $Y=2.635
+ $X2=8.9 $Y2=2.34
r170 32 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=2.635
+ $X2=7.725 $Y2=2.72
r171 32 34 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.725 $Y=2.635
+ $X2=7.725 $Y2=2
r172 28 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.72 $Y=2.635
+ $X2=6.72 $Y2=2.72
r173 28 30 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.72 $Y=2.635
+ $X2=6.72 $Y2=2.36
r174 22 76 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r175 22 24 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r176 7 41 400 $w=1.7e-07 $l=9.65376e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=1.485 $X2=8.85 $Y2=2.34
r177 7 38 400 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=8.615
+ $Y=1.485 $X2=8.85 $Y2=1.66
r178 6 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.54
+ $Y=1.485 $X2=7.685 $Y2=2
r179 5 30 600 $w=1.7e-07 $l=9.58514e-07 $layer=licon1_PDIFF $count=1 $X=6.545
+ $Y=1.485 $X2=6.72 $Y2=2.36
r180 4 90 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=5.605
+ $Y=1.485 $X2=5.75 $Y2=2.36
r181 3 61 600 $w=1.7e-07 $l=9.24054e-07 $layer=licon1_PDIFF $count=1 $X=4.465
+ $Y=1.515 $X2=4.675 $Y2=2.34
r182 2 83 600 $w=1.7e-07 $l=4.54148e-07 $layer=licon1_PDIFF $count=1 $X=2.715
+ $Y=2.065 $X2=3.045 $Y2=2.36
r183 1 24 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%A_27_47# 1 2 3 12 15 16 17 18 20 24
r52 22 24 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.205 $Y=0.615
+ $X2=1.205 $Y2=0.42
r53 18 20 15.5919 $w=3.38e-07 $l=4.6e-07 $layer=LI1_cond $X=0.735 $Y=2.295
+ $X2=1.195 $Y2=2.295
r54 16 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=1.205 $Y2=0.615
r55 16 17 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=0.735 $Y2=0.7
r56 15 18 7.23167 $w=3.4e-07 $l=2.18174e-07 $layer=LI1_cond $X=0.625 $Y=2.125
+ $X2=0.735 $Y2=2.295
r57 14 17 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.625 $Y=0.7
+ $X2=0.735 $Y2=0.7
r58 14 15 70.1943 $w=2.18e-07 $l=1.34e-06 $layer=LI1_cond $X=0.625 $Y=0.785
+ $X2=0.625 $Y2=2.125
r59 10 14 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.625 $Y2=0.7
r60 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r61 3 20 600 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.845 $X2=1.195 $Y2=2.29
r62 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.42
r63 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%GCLK 1 2 3 4 14 17 19 20 21 22 24 26 28
+ 32 33 34 35 36 37 38 39 48 53
c89 32 0 1.23116e-19 $X=7.735 $Y=1.185
c90 28 0 2.87968e-19 $X=7.215 $Y=0.36
c91 19 0 1.27609e-19 $X=7.65 $Y=0.8
r92 37 38 10.0469 $w=3.88e-07 $l=3.4e-07 $layer=LI1_cond $X=8.4 $Y=1.87 $X2=8.4
+ $Y2=2.21
r93 37 61 1.62524 $w=3.88e-07 $l=5.5e-08 $layer=LI1_cond $X=8.4 $Y=1.87 $X2=8.4
+ $Y2=1.815
r94 36 61 8.4217 $w=3.88e-07 $l=2.85e-07 $layer=LI1_cond $X=8.4 $Y=1.53 $X2=8.4
+ $Y2=1.815
r95 36 57 6.35321 $w=3.88e-07 $l=2.15e-07 $layer=LI1_cond $X=8.4 $Y=1.53 $X2=8.4
+ $Y2=1.315
r96 35 51 4.06667 $w=3.9e-07 $l=1.3e-07 $layer=LI1_cond $X=8.4 $Y=1.185 $X2=8.4
+ $Y2=1.055
r97 35 57 4.06667 $w=3.9e-07 $l=1.3e-07 $layer=LI1_cond $X=8.4 $Y=1.185 $X2=8.4
+ $Y2=1.315
r98 35 48 9.15 $w=2.6e-07 $l=1.95e-07 $layer=LI1_cond $X=8.4 $Y=1.185 $X2=8.205
+ $Y2=1.185
r99 35 39 11.8382 $w=4.28e-07 $l=3.75e-07 $layer=LI1_cond $X=8.595 $Y=1.185
+ $X2=8.97 $Y2=1.185
r100 34 51 6.05771 $w=3.88e-07 $l=2.05e-07 $layer=LI1_cond $X=8.4 $Y=0.85
+ $X2=8.4 $Y2=1.055
r101 34 53 12.7064 $w=3.88e-07 $l=4.3e-07 $layer=LI1_cond $X=8.4 $Y=0.85 $X2=8.4
+ $Y2=0.42
r102 33 48 6.87033 $w=2.58e-07 $l=1.55e-07 $layer=LI1_cond $X=8.05 $Y=1.185
+ $X2=8.205 $Y2=1.185
r103 31 33 10.1947 $w=2.58e-07 $l=2.3e-07 $layer=LI1_cond $X=7.82 $Y=1.185
+ $X2=8.05 $Y2=1.185
r104 31 32 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.82 $Y=1.185
+ $X2=7.735 $Y2=1.185
r105 25 32 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.735 $Y=1.315
+ $X2=7.735 $Y2=1.185
r106 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.735 $Y=1.315
+ $X2=7.735 $Y2=1.485
r107 24 32 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.735 $Y=1.055
+ $X2=7.735 $Y2=1.185
r108 23 24 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.735 $Y=0.885
+ $X2=7.735 $Y2=1.055
r109 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.65 $Y=1.57
+ $X2=7.735 $Y2=1.485
r110 21 22 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=1.57
+ $X2=7.38 $Y2=1.57
r111 19 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.65 $Y=0.8
+ $X2=7.735 $Y2=0.885
r112 19 20 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.65 $Y=0.8 $X2=7.38
+ $Y2=0.8
r113 15 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.255 $Y=1.655
+ $X2=7.38 $Y2=1.57
r114 15 17 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=7.255 $Y=1.655
+ $X2=7.255 $Y2=1.815
r115 14 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.255 $Y=0.715
+ $X2=7.38 $Y2=0.8
r116 14 28 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=7.255 $Y=0.715
+ $X2=7.255 $Y2=0.445
r117 4 61 300 $w=1.7e-07 $l=4.48665e-07 $layer=licon1_PDIFF $count=2 $X=8.01
+ $Y=1.485 $X2=8.29 $Y2=1.815
r118 3 17 300 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=2 $X=7.07
+ $Y=1.485 $X2=7.215 $Y2=1.815
r119 2 53 182 $w=1.7e-07 $l=4.01995e-07 $layer=licon1_NDIFF $count=1 $X=7.97
+ $Y=0.235 $X2=8.29 $Y2=0.42
r120 1 28 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.03
+ $Y=0.235 $X2=7.215 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_4%VGND 1 2 3 4 5 6 21 25 27 29 31 32 39 40
+ 41 43 48 71 77 83 88 94 97
r131 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r132 92 94 9.59153 $w=5.28e-07 $l=1.6e-07 $layer=LI1_cond $X=6.67 $Y=0.18
+ $X2=6.83 $Y2=0.18
r133 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r134 90 92 0.112838 $w=5.28e-07 $l=5e-09 $layer=LI1_cond $X=6.665 $Y=0.18
+ $X2=6.67 $Y2=0.18
r135 87 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r136 86 90 10.2682 $w=5.28e-07 $l=4.55e-07 $layer=LI1_cond $X=6.21 $Y=0.18
+ $X2=6.665 $Y2=0.18
r137 86 88 10.6071 $w=5.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.21 $Y=0.18
+ $X2=6.005 $Y2=0.18
r138 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r139 83 84 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r140 77 80 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.36
r141 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r142 74 97 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r143 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r144 71 96 4.11661 $w=1.7e-07 $l=2.17e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.982 $Y2=0
r145 71 73 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.51 $Y2=0
r146 70 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.51
+ $Y2=0
r147 70 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=6.67
+ $Y2=0
r148 69 94 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.59 $Y=0 $X2=6.83
+ $Y2=0
r149 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r150 66 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r151 65 88 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=6.005 $Y2=0
r152 65 66 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r153 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r154 62 65 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r155 62 63 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r156 59 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r157 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r158 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r159 56 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r160 55 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r161 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r162 53 83 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=3.092 $Y2=0
r163 53 55 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=3.265 $Y=0
+ $X2=3.45 $Y2=0
r164 52 84 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r165 52 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r166 51 52 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r167 49 77 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r168 49 51 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r169 48 83 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.92 $Y=0 $X2=3.092
+ $Y2=0
r170 48 51 115.476 $w=1.68e-07 $l=1.77e-06 $layer=LI1_cond $X=2.92 $Y=0 $X2=1.15
+ $Y2=0
r171 43 77 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r172 43 45 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r173 41 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r174 41 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r175 39 69 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=7.6 $Y=0 $X2=7.59
+ $Y2=0
r176 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.6 $Y=0 $X2=7.725
+ $Y2=0
r177 38 73 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=7.85 $Y=0 $X2=8.51
+ $Y2=0
r178 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.85 $Y=0 $X2=7.725
+ $Y2=0
r179 34 62 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.83
+ $Y2=0
r180 32 58 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.37
+ $Y2=0
r181 31 36 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.585 $Y=0
+ $X2=4.585 $Y2=0.36
r182 31 34 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.775
+ $Y2=0
r183 31 32 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.585 $Y=0 $X2=4.395
+ $Y2=0
r184 27 96 3.16808 $w=2.7e-07 $l=1.19143e-07 $layer=LI1_cond $X=8.9 $Y=0.085
+ $X2=8.982 $Y2=0
r185 27 29 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.9 $Y=0.085
+ $X2=8.9 $Y2=0.38
r186 23 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.725 $Y=0.085
+ $X2=7.725 $Y2=0
r187 23 25 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=7.725 $Y=0.085
+ $X2=7.725 $Y2=0.38
r188 19 83 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.092 $Y=0.085
+ $X2=3.092 $Y2=0
r189 19 21 14.1968 $w=3.43e-07 $l=4.25e-07 $layer=LI1_cond $X=3.092 $Y=0.085
+ $X2=3.092 $Y2=0.51
r190 6 29 91 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_NDIFF $count=2 $X=8.625
+ $Y=0.235 $X2=8.85 $Y2=0.38
r191 5 25 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.5
+ $Y=0.235 $X2=7.685 $Y2=0.38
r192 4 90 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=6.445
+ $Y=0.235 $X2=6.665 $Y2=0.36
r193 3 36 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.235 $X2=4.61 $Y2=0.36
r194 2 21 182 $w=1.7e-07 $l=3.72659e-07 $layer=licon1_NDIFF $count=1 $X=2.835
+ $Y=0.235 $X2=3.065 $Y2=0.51
r195 1 80 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

