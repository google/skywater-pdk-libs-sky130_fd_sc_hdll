* File: sky130_fd_sc_hdll__mux2i_1.pxi.spice
* Created: Wed Sep  2 08:34:52 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A0 N_A0_c_67_n N_A0_M1000_g N_A0_c_64_n
+ N_A0_M1005_g A0 N_A0_c_66_n PM_SKY130_FD_SC_HDLL__MUX2I_1%A0
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A1 N_A1_c_91_n N_A1_M1002_g N_A1_c_92_n
+ N_A1_M1007_g N_A1_c_93_n A1 A1 PM_SKY130_FD_SC_HDLL__MUX2I_1%A1
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A_303_205# N_A_303_205#_M1003_s
+ N_A_303_205#_M1004_s N_A_303_205#_c_131_n N_A_303_205#_M1006_g
+ N_A_303_205#_M1008_g N_A_303_205#_c_127_n N_A_303_205#_c_128_n
+ N_A_303_205#_c_129_n N_A_303_205#_c_134_n N_A_303_205#_c_130_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%A_303_205#
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%S N_S_M1009_g N_S_c_199_n N_S_M1001_g
+ N_S_c_194_n N_S_c_195_n N_S_M1004_g N_S_c_196_n N_S_M1003_g N_S_c_197_n S S S
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%S
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_297# N_A_27_297#_M1000_s
+ N_A_27_297#_M1001_d N_A_27_297#_c_250_n N_A_27_297#_c_251_n
+ N_A_27_297#_c_259_n N_A_27_297#_c_264_n N_A_27_297#_c_252_n
+ N_A_27_297#_c_253_n N_A_27_297#_c_254_n N_A_27_297#_c_255_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%Y N_Y_M1005_d N_Y_M1000_d Y Y N_Y_c_295_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%Y
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%VPWR N_VPWR_M1006_d N_VPWR_M1004_d
+ N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n N_VPWR_c_323_n VPWR
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_319_n N_VPWR_c_327_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1008_s
+ N_A_27_47#_c_359_n N_A_27_47#_c_373_p N_A_27_47#_c_360_n N_A_27_47#_c_361_n
+ N_A_27_47#_c_367_n PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%A_207_47# N_A_207_47#_M1002_d
+ N_A_207_47#_M1009_d N_A_207_47#_c_386_n N_A_207_47#_c_387_n
+ N_A_207_47#_c_388_n N_A_207_47#_c_398_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%A_207_47#
x_PM_SKY130_FD_SC_HDLL__MUX2I_1%VGND N_VGND_M1008_d N_VGND_M1003_d
+ N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n N_VGND_c_425_n VGND
+ N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n
+ PM_SKY130_FD_SC_HDLL__MUX2I_1%VGND
cc_1 VNB N_A0_c_64_n 0.0215747f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB A0 0.00925368f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A0_c_66_n 0.0412594f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_4 VNB N_A1_c_91_n 0.02219f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_A1_c_92_n 0.0277352f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_6 VNB N_A1_c_93_n 0.00468622f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_7 VNB N_A_303_205#_M1008_g 0.0240599f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_8 VNB N_A_303_205#_c_127_n 0.0156054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_303_205#_c_128_n 0.0365721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_303_205#_c_129_n 0.0108388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_303_205#_c_130_n 5.41669e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_S_M1009_g 0.0304312f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_13 VNB N_S_c_194_n 0.0338928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_S_c_195_n 0.0354084f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_15 VNB N_S_c_196_n 0.0228128f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_16 VNB N_S_c_197_n 0.004855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB S 0.0210425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_295_n 0.00330557f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_319_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_359_n 0.0176849f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_21 VNB N_A_27_47#_c_360_n 0.00649749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_361_n 0.00921644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_207_47#_c_386_n 0.00316787f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_24 VNB N_A_207_47#_c_387_n 0.00419053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_207_47#_c_388_n 0.0111518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_422_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_27 VNB N_VGND_c_423_n 0.016033f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_28 VNB N_VGND_c_424_n 0.0357301f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_425_n 0.00420404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_426_n 0.0489331f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_427_n 0.0149861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_428_n 0.243602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_429_n 0.00323881f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A0_c_67_n 0.0204286f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_35 VPB N_A0_c_66_n 0.0179842f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_36 VPB N_A1_c_92_n 0.0286995f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_37 VPB A1 0.00164497f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_38 VPB N_A_303_205#_c_131_n 0.0190683f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_39 VPB N_A_303_205#_c_127_n 0.00570321f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_303_205#_c_128_n 0.00783497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_303_205#_c_134_n 0.0106045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_S_c_199_n 0.0212794f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.56
cc_43 VPB N_S_c_194_n 0.0316061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_S_c_195_n 0.038033f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_45 VPB N_S_c_197_n 0.00733532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB S 0.01231f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_297#_c_250_n 0.00712721f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_48 VPB N_A_27_297#_c_251_n 0.0334885f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_49 VPB N_A_27_297#_c_252_n 0.0040699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_297#_c_253_n 2.7441e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_254_n 0.00349529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_255_n 0.00803767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB Y 0.00254915f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_54 VPB N_Y_c_295_n 0.0015013f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_320_n 0.00536298f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_56 VPB N_VPWR_c_321_n 0.0313134f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_57 VPB N_VPWR_c_322_n 0.0355085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_323_n 0.00564836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_324_n 0.0468849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_325_n 0.0139174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_319_n 0.0660902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_327_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 N_A0_c_64_n N_A1_c_91_n 0.0227443f $X=0.54 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_64 N_A0_c_67_n N_A1_c_92_n 0.0235943f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A0_c_66_n N_A1_c_92_n 0.0227443f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_66 N_A0_c_66_n N_A1_c_93_n 2.44243e-19 $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_67 N_A0_c_67_n N_A_27_297#_c_251_n 7.43495e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_68 A0 N_A_27_297#_c_251_n 0.0246129f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_69 N_A0_c_66_n N_A_27_297#_c_251_n 0.0071827f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_70 N_A0_c_67_n N_A_27_297#_c_259_n 0.0143148f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A0_c_67_n N_Y_c_295_n 0.00146642f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A0_c_64_n N_Y_c_295_n 0.00893972f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_73 A0 N_Y_c_295_n 0.0153721f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A0_c_66_n N_Y_c_295_n 0.0154028f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_75 N_A0_c_67_n N_VPWR_c_324_n 0.00429453f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A0_c_67_n N_VPWR_c_319_n 0.00702073f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A0_c_64_n N_A_27_47#_c_359_n 0.0112573f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_78 A0 N_A_27_47#_c_359_n 0.0197608f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_79 N_A0_c_66_n N_A_27_47#_c_359_n 0.00590828f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_80 A0 N_A_27_47#_c_361_n 0.00188679f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_A0_c_66_n N_A_27_47#_c_361_n 0.00161682f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_82 N_A0_c_64_n N_A_27_47#_c_367_n 0.0154935f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A0_c_64_n N_VGND_c_426_n 0.00357877f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A0_c_64_n N_VGND_c_428_n 0.00634625f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A1_c_92_n N_A_303_205#_c_131_n 0.0284749f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_86 A1 N_A_303_205#_c_131_n 0.0037694f $X=1.095 $Y=1.445 $X2=0 $Y2=0
cc_87 N_A1_c_92_n N_A_303_205#_M1008_g 4.39614e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A1_c_93_n N_A_303_205#_M1008_g 4.74514e-19 $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A1_c_92_n N_A_303_205#_c_127_n 9.43845e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A1_c_93_n N_A_303_205#_c_127_n 0.0168965f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A1_c_92_n N_A_303_205#_c_128_n 0.0158241f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A1_c_93_n N_A_303_205#_c_128_n 0.00394642f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A1_c_92_n N_A_27_297#_c_259_n 0.0168954f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_94 A1 N_A_27_297#_c_259_n 0.009947f $X=1.095 $Y=1.445 $X2=0 $Y2=0
cc_95 A1 N_A_27_297#_c_253_n 0.00507385f $X=1.095 $Y=1.445 $X2=0 $Y2=0
cc_96 N_A1_c_92_n Y 2.54491e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_97 A1 Y 0.0233929f $X=1.095 $Y=1.445 $X2=0 $Y2=0
cc_98 N_A1_c_91_n N_Y_c_295_n 0.00611657f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A1_c_92_n N_Y_c_295_n 3.67561e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A1_c_93_n N_Y_c_295_n 0.0249375f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_101 A1 N_Y_c_295_n 0.00760459f $X=1.095 $Y=1.445 $X2=0 $Y2=0
cc_102 A1 A_215_297# 0.0079464f $X=1.095 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_103 N_A1_c_92_n N_VPWR_c_324_n 0.00429453f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A1_c_92_n N_VPWR_c_319_n 0.00650299f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A1_c_91_n N_A_27_47#_c_367_n 0.0153854f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A1_c_91_n N_A_207_47#_c_388_n 0.00260151f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A1_c_92_n N_A_207_47#_c_388_n 0.00131673f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_93_n N_A_207_47#_c_388_n 0.017945f $X=1.09 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A1_c_91_n N_VGND_c_426_n 0.00357877f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A1_c_91_n N_VGND_c_428_n 0.00666937f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_303_205#_M1008_g N_S_M1009_g 0.0214782f $X=1.9 $Y=0.56 $X2=0 $Y2=0
cc_112 N_A_303_205#_c_127_n N_S_M1009_g 0.00656427f $X=2.93 $Y=1.192 $X2=0 $Y2=0
cc_113 N_A_303_205#_c_129_n N_S_M1009_g 0.00526495f $X=3.11 $Y=0.42 $X2=0 $Y2=0
cc_114 N_A_303_205#_c_131_n N_S_c_199_n 0.0200311f $X=1.615 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_303_205#_c_134_n N_S_c_199_n 0.00325818f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_116 N_A_303_205#_c_127_n N_S_c_194_n 0.0225281f $X=2.93 $Y=1.192 $X2=0 $Y2=0
cc_117 N_A_303_205#_c_134_n N_S_c_194_n 0.00854395f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_118 N_A_303_205#_c_130_n N_S_c_194_n 0.0138834f $X=3.062 $Y=1.192 $X2=0 $Y2=0
cc_119 N_A_303_205#_c_134_n N_S_c_195_n 0.0160079f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_120 N_A_303_205#_c_130_n N_S_c_195_n 0.00233064f $X=3.062 $Y=1.192 $X2=0
+ $Y2=0
cc_121 N_A_303_205#_c_129_n N_S_c_196_n 0.0215846f $X=3.11 $Y=0.42 $X2=0 $Y2=0
cc_122 N_A_303_205#_c_127_n N_S_c_197_n 0.00705723f $X=2.93 $Y=1.192 $X2=0 $Y2=0
cc_123 N_A_303_205#_c_128_n N_S_c_197_n 0.0248443f $X=1.68 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_303_205#_c_134_n N_S_c_197_n 0.00151238f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_125 N_A_303_205#_c_129_n S 0.0245223f $X=3.11 $Y=0.42 $X2=0 $Y2=0
cc_126 N_A_303_205#_c_134_n S 0.0236642f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_127 N_A_303_205#_c_130_n S 0.0193755f $X=3.062 $Y=1.192 $X2=0 $Y2=0
cc_128 N_A_303_205#_c_131_n N_A_27_297#_c_259_n 0.00867534f $X=1.615 $Y=1.41
+ $X2=0 $Y2=0
cc_129 N_A_303_205#_c_131_n N_A_27_297#_c_264_n 0.0207367f $X=1.615 $Y=1.41
+ $X2=0 $Y2=0
cc_130 N_A_303_205#_c_127_n N_A_27_297#_c_252_n 0.0484467f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_131 N_A_303_205#_c_128_n N_A_27_297#_c_252_n 0.00167684f $X=1.68 $Y=1.16
+ $X2=0 $Y2=0
cc_132 N_A_303_205#_c_131_n N_A_27_297#_c_253_n 0.00971925f $X=1.615 $Y=1.41
+ $X2=0 $Y2=0
cc_133 N_A_303_205#_c_127_n N_A_27_297#_c_253_n 0.0173997f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_134 N_A_303_205#_c_128_n N_A_27_297#_c_253_n 6.18809e-19 $X=1.68 $Y=1.16
+ $X2=0 $Y2=0
cc_135 N_A_303_205#_c_127_n N_A_27_297#_c_254_n 0.0309672f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_136 N_A_303_205#_c_134_n N_A_27_297#_c_254_n 0.0120199f $X=3.11 $Y=1.96 $X2=0
+ $Y2=0
cc_137 N_A_303_205#_c_131_n N_A_27_297#_c_255_n 2.85809e-19 $X=1.615 $Y=1.41
+ $X2=0 $Y2=0
cc_138 N_A_303_205#_c_134_n N_A_27_297#_c_255_n 0.0547824f $X=3.11 $Y=1.96 $X2=0
+ $Y2=0
cc_139 N_A_303_205#_c_131_n N_VPWR_c_320_n 0.00538702f $X=1.615 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_303_205#_c_134_n N_VPWR_c_322_n 0.015687f $X=3.11 $Y=1.96 $X2=0 $Y2=0
cc_141 N_A_303_205#_c_131_n N_VPWR_c_324_n 0.00429201f $X=1.615 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_303_205#_M1004_s N_VPWR_c_319_n 0.00519837f $X=2.975 $Y=1.485 $X2=0
+ $Y2=0
cc_143 N_A_303_205#_c_131_n N_VPWR_c_319_n 0.00701728f $X=1.615 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_303_205#_c_134_n N_VPWR_c_319_n 0.00858812f $X=3.11 $Y=1.96 $X2=0
+ $Y2=0
cc_145 N_A_303_205#_M1008_g N_A_27_47#_c_360_n 0.00292079f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_146 N_A_303_205#_M1008_g N_A_207_47#_c_386_n 0.013723f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_147 N_A_303_205#_c_127_n N_A_207_47#_c_386_n 0.0182513f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_148 N_A_303_205#_c_129_n N_A_207_47#_c_386_n 0.011974f $X=3.11 $Y=0.42 $X2=0
+ $Y2=0
cc_149 N_A_303_205#_c_129_n N_A_207_47#_c_387_n 0.0296971f $X=3.11 $Y=0.42 $X2=0
+ $Y2=0
cc_150 N_A_303_205#_c_127_n N_A_207_47#_c_388_n 0.00502436f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_151 N_A_303_205#_c_128_n N_A_207_47#_c_388_n 0.0015462f $X=1.68 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_303_205#_M1008_g N_A_207_47#_c_398_n 0.00268976f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_153 N_A_303_205#_c_127_n N_A_207_47#_c_398_n 0.0519644f $X=2.93 $Y=1.192
+ $X2=0 $Y2=0
cc_154 N_A_303_205#_c_128_n N_A_207_47#_c_398_n 0.00618549f $X=1.68 $Y=1.16
+ $X2=0 $Y2=0
cc_155 N_A_303_205#_M1008_g N_VGND_c_422_n 0.00268723f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_156 N_A_303_205#_c_129_n N_VGND_c_424_n 0.0185411f $X=3.11 $Y=0.42 $X2=0
+ $Y2=0
cc_157 N_A_303_205#_M1008_g N_VGND_c_426_n 0.00420765f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_158 N_A_303_205#_M1003_s N_VGND_c_428_n 0.00703964f $X=2.965 $Y=0.235 $X2=0
+ $Y2=0
cc_159 N_A_303_205#_M1008_g N_VGND_c_428_n 0.00705894f $X=1.9 $Y=0.56 $X2=0
+ $Y2=0
cc_160 N_A_303_205#_c_129_n N_VGND_c_428_n 0.0101286f $X=3.11 $Y=0.42 $X2=0
+ $Y2=0
cc_161 N_S_c_199_n N_A_27_297#_c_252_n 0.0110989f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_162 N_S_c_197_n N_A_27_297#_c_252_n 2.964e-19 $X=2.345 $Y=1.287 $X2=0 $Y2=0
cc_163 N_S_c_199_n N_A_27_297#_c_254_n 0.00211974f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_164 N_S_c_194_n N_A_27_297#_c_254_n 0.00679421f $X=3.265 $Y=1.257 $X2=0 $Y2=0
cc_165 N_S_c_197_n N_A_27_297#_c_254_n 3.07171e-19 $X=2.345 $Y=1.287 $X2=0 $Y2=0
cc_166 N_S_c_199_n N_A_27_297#_c_255_n 0.0143694f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_167 S N_VPWR_M1004_d 0.00313909f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_168 N_S_c_199_n N_VPWR_c_320_n 0.010235f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_169 N_S_c_195_n N_VPWR_c_321_n 0.00585219f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_170 S N_VPWR_c_321_n 0.0180155f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_171 N_S_c_199_n N_VPWR_c_322_n 0.00597712f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_172 N_S_c_195_n N_VPWR_c_322_n 0.00702461f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_173 N_S_c_199_n N_VPWR_c_319_n 0.0119454f $X=2.345 $Y=1.41 $X2=0 $Y2=0
cc_174 N_S_c_195_n N_VPWR_c_319_n 0.014779f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_175 N_S_M1009_g N_A_207_47#_c_386_n 0.0129919f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_176 N_S_c_194_n N_A_207_47#_c_386_n 0.00134749f $X=3.265 $Y=1.257 $X2=0 $Y2=0
cc_177 N_S_M1009_g N_A_207_47#_c_387_n 0.00700894f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_178 S N_VGND_M1003_d 0.00265397f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_179 N_S_M1009_g N_VGND_c_422_n 0.00268723f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_180 N_S_c_195_n N_VGND_c_423_n 9.95348e-19 $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_181 N_S_c_196_n N_VGND_c_423_n 0.0044587f $X=3.39 $Y=0.99 $X2=0 $Y2=0
cc_182 S N_VGND_c_423_n 0.0150646f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_183 N_S_M1009_g N_VGND_c_424_n 0.00436487f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_184 N_S_c_196_n N_VGND_c_424_n 0.00491017f $X=3.39 $Y=0.99 $X2=0 $Y2=0
cc_185 S N_VGND_c_424_n 0.00170758f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_186 S N_VGND_c_427_n 2.1649e-19 $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_187 N_S_M1009_g N_VGND_c_428_n 0.00731071f $X=2.32 $Y=0.56 $X2=0 $Y2=0
cc_188 N_S_c_196_n N_VGND_c_428_n 0.0101019f $X=3.39 $Y=0.99 $X2=0 $Y2=0
cc_189 S N_VGND_c_428_n 0.00497188f $X=3.515 $Y=0.765 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_259_n N_Y_M1000_d 0.00352392f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_251_n Y 0.0267271f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_192 N_A_27_297#_c_259_n Y 0.0134101f $X=1.505 $Y=2.38 $X2=0 $Y2=0
cc_193 N_A_27_297#_c_259_n A_215_297# 0.0132306f $X=1.505 $Y=2.38 $X2=-0.19
+ $Y2=1.305
cc_194 N_A_27_297#_c_252_n N_VPWR_M1006_d 0.0108115f $X=2.365 $Y=1.565 $X2=-0.19
+ $Y2=1.305
cc_195 N_A_27_297#_c_252_n N_VPWR_c_320_n 0.0212328f $X=2.365 $Y=1.565 $X2=0
+ $Y2=0
cc_196 N_A_27_297#_c_255_n N_VPWR_c_320_n 0.044794f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_255_n N_VPWR_c_322_n 0.0244686f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_198 N_A_27_297#_c_250_n N_VPWR_c_324_n 0.0193052f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_259_n N_VPWR_c_324_n 0.0757804f $X=1.505 $Y=2.38 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_M1000_s N_VPWR_c_319_n 0.00230701f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_M1001_d N_VPWR_c_319_n 0.00217517f $X=2.435 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_27_297#_c_250_n N_VPWR_c_319_n 0.0115483f $X=0.27 $Y=2.295 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_259_n N_VPWR_c_319_n 0.0463457f $X=1.505 $Y=2.38 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_255_n N_VPWR_c_319_n 0.0141694f $X=2.58 $Y=2.32 $X2=0 $Y2=0
cc_205 N_Y_M1000_d N_VPWR_c_319_n 0.00232092f $X=0.605 $Y=1.485 $X2=0 $Y2=0
cc_206 N_Y_c_295_n N_A_27_47#_c_359_n 0.0155375f $X=0.75 $Y=0.76 $X2=0 $Y2=0
cc_207 N_Y_M1005_d N_A_27_47#_c_367_n 0.00312348f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_208 N_Y_c_295_n N_A_27_47#_c_367_n 0.0124912f $X=0.75 $Y=0.76 $X2=0 $Y2=0
cc_209 N_Y_M1005_d N_VGND_c_428_n 0.00216833f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_210 A_215_297# N_VPWR_c_319_n 0.00362899f $X=1.075 $Y=1.485 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_373_p N_A_207_47#_M1002_d 0.00430243f $X=1.275 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_212 N_A_27_47#_c_360_n N_A_207_47#_M1002_d 6.11981e-19 $X=1.69 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_213 N_A_27_47#_M1008_s N_A_207_47#_c_386_n 3.55274e-19 $X=1.565 $Y=0.235
+ $X2=0 $Y2=0
cc_214 N_A_27_47#_c_360_n N_A_207_47#_c_386_n 0.00225424f $X=1.69 $Y=0.38 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_M1008_s N_A_207_47#_c_388_n 2.69323e-19 $X=1.565 $Y=0.235
+ $X2=0 $Y2=0
cc_216 N_A_27_47#_c_373_p N_A_207_47#_c_388_n 0.0214613f $X=1.275 $Y=0.36 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_367_n N_A_207_47#_c_388_n 0.0014352f $X=1.065 $Y=0.36 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_M1008_s N_A_207_47#_c_398_n 0.00619419f $X=1.565 $Y=0.235
+ $X2=0 $Y2=0
cc_219 N_A_27_47#_c_360_n N_A_207_47#_c_398_n 0.0214613f $X=1.69 $Y=0.38 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_c_361_n N_VGND_c_426_n 0.10479f $X=0.44 $Y=0.36 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1005_s N_VGND_c_428_n 0.0026754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_222 N_A_27_47#_M1008_s N_VGND_c_428_n 0.00209344f $X=1.565 $Y=0.235 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_361_n N_VGND_c_428_n 0.0645352f $X=0.44 $Y=0.36 $X2=0 $Y2=0
cc_224 N_A_207_47#_c_386_n N_VGND_M1008_d 0.00343381f $X=2.465 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_225 N_A_207_47#_c_386_n N_VGND_c_422_n 0.0110546f $X=2.465 $Y=0.8 $X2=0 $Y2=0
cc_226 N_A_207_47#_c_386_n N_VGND_c_424_n 0.00307482f $X=2.465 $Y=0.8 $X2=0
+ $Y2=0
cc_227 N_A_207_47#_c_387_n N_VGND_c_424_n 0.0163122f $X=2.56 $Y=0.55 $X2=0 $Y2=0
cc_228 N_A_207_47#_c_386_n N_VGND_c_426_n 0.00203142f $X=2.465 $Y=0.8 $X2=0
+ $Y2=0
cc_229 N_A_207_47#_M1002_d N_VGND_c_428_n 0.00210147f $X=1.035 $Y=0.235 $X2=0
+ $Y2=0
cc_230 N_A_207_47#_M1009_d N_VGND_c_428_n 0.00267671f $X=2.395 $Y=0.235 $X2=0
+ $Y2=0
cc_231 N_A_207_47#_c_386_n N_VGND_c_428_n 0.0111916f $X=2.465 $Y=0.8 $X2=0 $Y2=0
cc_232 N_A_207_47#_c_387_n N_VGND_c_428_n 0.00895528f $X=2.56 $Y=0.55 $X2=0
+ $Y2=0
