* NGSPICE file created from sky130_fd_sc_hdll__muxb8to1_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__muxb8to1_2 D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[7]
+ S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
M1000 VPWR D[2] a_1315_297# VPB phighvt w=1e+06u l=180000u
+  ad=3.76e+12p pd=3.152e+07u as=8.211e+11p ps=7.41e+06u
M1001 VPWR D[3] a_2112_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.211e+11p ps=7.41e+06u
M1002 VPWR S[4] a_2854_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1003 a_27_297# D[0] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1004 Z a_1566_265# a_1315_297# VPB phighvt w=820000u l=180000u
+  ad=1.9024e+12p pd=1.776e+07u as=0p ps=0u
M1005 Z a_1989_47# a_2112_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# a_278_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_4565_47# S[7] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=1.9656e+12p ps=2.104e+07u
M1008 VPWR S[0] a_278_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1009 a_1989_47# S[3] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1010 Z S[5] a_3421_69# VNB nshort w=520000u l=150000u
+  ad=1.1232e+12p pd=1.264e+07u as=5.6745e+11p ps=5.52e+06u
M1011 a_4709_69# D[7] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1012 a_2133_69# D[3] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1013 Z a_278_265# a_27_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_2603_297# D[4] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1015 a_845_69# S[1] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1016 a_2603_297# a_2854_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_47# S[0] Z VNB nshort w=520000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1018 Z S[1] a_845_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_27_47# D[0] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 Z S[0] a_27_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 Z S[4] a_2603_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1022 a_824_333# D[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1023 a_1989_47# S[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1024 a_3400_333# a_3277_47# Z VPB phighvt w=820000u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1025 a_3400_333# D[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_3421_69# S[5] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VGND D[7] a_4709_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_3277_47# S[5] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1029 a_3891_297# D[6] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1030 a_4688_333# D[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.211e+11p pd=7.41e+06u as=0p ps=0u
M1031 VGND D[4] a_2603_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND S[4] a_2854_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1033 a_3891_297# a_4142_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VPWR D[0] a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1035 a_701_47# S[1] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1036 VGND D[1] a_845_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1037 VPWR D[4] a_2603_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1038 VPWR D[5] a_3400_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VPWR S[6] a_4142_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1040 a_824_333# a_701_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1041 Z a_2854_265# a_2603_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1042 Z a_3277_47# a_3400_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1043 VGND S[0] a_278_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1044 a_2603_47# S[4] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1045 a_701_47# S[1] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1046 Z a_4142_265# a_3891_297# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1047 VGND D[5] a_3421_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1048 a_2603_47# D[4] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1049 VPWR D[1] a_824_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1050 a_3277_47# S[5] VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1051 a_845_69# D[1] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1052 Z S[3] a_2133_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1053 VGND D[0] a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1054 a_3421_69# D[5] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1055 Z S[7] a_4709_69# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1056 Z a_701_47# a_824_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1057 a_1315_47# D[2] VGND VNB nshort w=650000u l=150000u
+  ad=5.6745e+11p pd=5.52e+06u as=0p ps=0u
M1058 Z S[2] a_1315_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1059 Z S[6] a_3891_47# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=5.6745e+11p ps=5.52e+06u
M1060 a_1315_297# D[2] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1061 a_1315_297# a_1566_265# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1062 a_2112_333# a_1989_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1063 VGND D[2] a_1315_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1064 a_4688_333# a_4565_47# Z VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1065 a_2133_69# S[3] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1066 a_4565_47# S[7] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1067 VPWR S[2] a_1566_265# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1068 a_2112_333# D[3] VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1069 VPWR D[7] a_4688_333# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1070 VGND D[6] a_3891_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1071 a_4709_69# S[7] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1072 VPWR D[6] a_3891_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1073 Z a_4565_47# a_4688_333# VPB phighvt w=820000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1074 a_3891_47# S[6] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1075 VGND S[6] a_4142_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1076 a_1315_47# S[2] Z VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1077 VGND S[2] a_1566_265# VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=1.352e+11p ps=1.56e+06u
M1078 VGND D[3] a_2133_69# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1079 a_3891_47# D[6] VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

