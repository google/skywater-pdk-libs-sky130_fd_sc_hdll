* File: sky130_fd_sc_hdll__and3_4.pex.spice
* Created: Thu Aug 27 18:58:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3_4%A 1 3 4 6 7 8 9 10 11 19 20
r31 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.74
+ $Y=1.16 $X2=0.74 $Y2=1.16
r32 11 19 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=0.64 $Y=1.167 $X2=0.74
+ $Y2=1.167
r33 11 25 10.3553 $w=3.43e-07 $l=3.1e-07 $layer=LI1_cond $X=0.64 $Y=1.167
+ $X2=0.33 $Y2=1.167
r34 9 10 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=2.21
r35 8 9 18.2247 $w=2.13e-07 $l=3.4e-07 $layer=LI1_cond $X=0.222 $Y=1.53
+ $X2=0.222 $Y2=1.87
r36 8 20 10.1844 $w=2.13e-07 $l=1.9e-07 $layer=LI1_cond $X=0.222 $Y=1.53
+ $X2=0.222 $Y2=1.34
r37 7 20 4.49766 $w=2.15e-07 $l=1.73e-07 $layer=LI1_cond $X=0.222 $Y=1.167
+ $X2=0.222 $Y2=1.34
r38 7 25 2.80779 $w=3.45e-07 $l=1.08e-07 $layer=LI1_cond $X=0.222 $Y=1.167
+ $X2=0.33 $Y2=1.167
r39 4 18 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.85 $Y=0.995
+ $X2=0.765 $Y2=1.16
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.85 $Y=0.995 $X2=0.85
+ $Y2=0.56
r41 1 18 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.825 $Y=1.41
+ $X2=0.765 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.825 $Y=1.41
+ $X2=0.825 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%B 1 3 4 6 7 8
c31 7 0 1.93824e-19 $X=1.115 $Y=0.765
r32 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r33 8 13 1.11527 $w=3.08e-07 $l=3e-08 $layer=LI1_cond $X=1.2 $Y=1.19 $X2=1.2
+ $Y2=1.16
r34 7 13 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=1.2 $Y=0.85 $X2=1.2
+ $Y2=1.16
r35 4 12 39.3227 $w=3.86e-07 $l=2.25433e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.352 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r37 1 12 45.0491 $w=3.86e-07 $l=3.03315e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.352 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.41 $X2=1.47
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%C 1 3 4 6 7 11 13
c39 4 0 3.89502e-19 $X=1.95 $Y=1.41
r40 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.16 $X2=1.915 $Y2=1.16
r41 7 11 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.71 $Y=1.16
+ $X2=1.915 $Y2=1.16
r42 7 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=1.16 $X2=1.61
+ $Y2=1.16
r43 4 10 48.1208 $w=2.95e-07 $l=2.54951e-07 $layer=POLY_cond $X=1.95 $Y=1.41
+ $X2=1.94 $Y2=1.16
r44 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.95 $Y=1.41 $X2=1.95
+ $Y2=1.985
r45 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.94 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%A_85_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 38 40 41 42 46 49 50 52 53 55 57 63 67 68 69 78
c143 78 0 1.13405e-19 $X=3.945 $Y=1.202
c144 55 0 1.95678e-19 $X=2.325 $Y=1.02
r145 78 79 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.945 $Y=1.202
+ $X2=3.97 $Y2=1.202
r146 75 76 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.465 $Y2=1.202
r147 74 75 59.1132 $w=3.71e-07 $l=4.55e-07 $layer=POLY_cond $X=2.985 $Y=1.202
+ $X2=3.44 $Y2=1.202
r148 73 74 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.96 $Y=1.202
+ $X2=2.985 $Y2=1.202
r149 70 71 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.48 $Y=1.202
+ $X2=2.505 $Y2=1.202
r150 64 78 26.6334 $w=3.71e-07 $l=2.05e-07 $layer=POLY_cond $X=3.74 $Y=1.202
+ $X2=3.945 $Y2=1.202
r151 64 76 35.7278 $w=3.71e-07 $l=2.75e-07 $layer=POLY_cond $X=3.74 $Y=1.202
+ $X2=3.465 $Y2=1.202
r152 63 64 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.74
+ $Y=1.16 $X2=3.74 $Y2=1.16
r153 61 73 50.6685 $w=3.71e-07 $l=3.9e-07 $layer=POLY_cond $X=2.57 $Y=1.202
+ $X2=2.96 $Y2=1.202
r154 61 71 8.44474 $w=3.71e-07 $l=6.5e-08 $layer=POLY_cond $X=2.57 $Y=1.202
+ $X2=2.505 $Y2=1.202
r155 60 63 40.2495 $w=3.33e-07 $l=1.17e-06 $layer=LI1_cond $X=2.57 $Y=1.187
+ $X2=3.74 $Y2=1.187
r156 60 61 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.57
+ $Y=1.16 $X2=2.57 $Y2=1.16
r157 58 69 0.271299 $w=3.35e-07 $l=1.05e-07 $layer=LI1_cond $X=2.43 $Y=1.187
+ $X2=2.325 $Y2=1.187
r158 58 60 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=2.43 $Y=1.187
+ $X2=2.57 $Y2=1.187
r159 56 69 7.47207 $w=2.1e-07 $l=1.68e-07 $layer=LI1_cond $X=2.325 $Y=1.355
+ $X2=2.325 $Y2=1.187
r160 56 57 11.8831 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=2.325 $Y=1.355
+ $X2=2.325 $Y2=1.58
r161 55 69 7.47207 $w=2.1e-07 $l=1.67e-07 $layer=LI1_cond $X=2.325 $Y=1.02
+ $X2=2.325 $Y2=1.187
r162 54 55 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=2.325 $Y=0.805
+ $X2=2.325 $Y2=1.02
r163 52 54 6.83868 $w=1.9e-07 $l=1.44914e-07 $layer=LI1_cond $X=2.22 $Y=0.71
+ $X2=2.325 $Y2=0.805
r164 52 53 23.0574 $w=1.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.22 $Y=0.71
+ $X2=1.825 $Y2=0.71
r165 51 68 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.8 $Y=1.665 $X2=1.71
+ $Y2=1.665
r166 50 57 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=2.325 $Y2=1.58
r167 50 51 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=2.22 $Y=1.665
+ $X2=1.8 $Y2=1.665
r168 49 53 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=1.73 $Y=0.615
+ $X2=1.825 $Y2=0.71
r169 48 49 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=1.73 $Y=0.445
+ $X2=1.73 $Y2=0.615
r170 44 68 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=1.75
+ $X2=1.71 $Y2=1.665
r171 44 46 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=1.71 $Y=1.75
+ $X2=1.71 $Y2=1.96
r172 43 67 4.80081 $w=1.9e-07 $l=1.68e-07 $layer=LI1_cond $X=0.8 $Y=0.35
+ $X2=0.632 $Y2=0.35
r173 42 48 6.81649 $w=1.9e-07 $l=1.3435e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=1.73 $Y2=0.445
r174 42 43 48.7416 $w=1.88e-07 $l=8.35e-07 $layer=LI1_cond $X=1.635 $Y=0.35
+ $X2=0.8 $Y2=0.35
r175 40 68 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=1.62 $Y=1.665 $X2=1.71
+ $Y2=1.665
r176 40 41 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.62 $Y=1.665
+ $X2=0.68 $Y2=1.665
r177 36 41 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.59 $Y=1.75
+ $X2=0.68 $Y2=1.665
r178 36 38 12.9394 $w=1.78e-07 $l=2.1e-07 $layer=LI1_cond $X=0.59 $Y=1.75
+ $X2=0.59 $Y2=1.96
r179 31 79 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.97 $Y=0.995
+ $X2=3.97 $Y2=1.202
r180 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.97 $Y=0.995
+ $X2=3.97 $Y2=0.56
r181 28 78 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.945 $Y=1.41
+ $X2=3.945 $Y2=1.202
r182 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.945 $Y=1.41
+ $X2=3.945 $Y2=1.985
r183 25 76 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.202
r184 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.465 $Y=1.41
+ $X2=3.465 $Y2=1.985
r185 22 75 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=1.202
r186 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=0.56
r187 19 74 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.202
r188 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.985
r189 16 73 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=2.96 $Y2=1.202
r190 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=2.96 $Y2=0.56
r191 13 71 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.202
r192 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.985
r193 10 70 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.48 $Y2=1.202
r194 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.48 $Y2=0.56
r195 3 46 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=1.485 $X2=1.71 $Y2=1.96
r196 2 38 300 $w=1.7e-07 $l=5.51362e-07 $layer=licon1_PDIFF $count=2 $X=0.425
+ $Y=1.485 $X2=0.59 $Y2=1.96
r197 1 67 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.47
+ $Y=0.235 $X2=0.635 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%VPWR 1 2 3 4 15 17 21 25 27 29 32 33 34 36
+ 45 50 53 57
r64 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r65 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r66 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 48 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 45 56 4.91801 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=3.97 $Y=2.72
+ $X2=4.285 $Y2=2.72
r71 45 47 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=2.72 $X2=3.91
+ $Y2=2.72
r72 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r73 44 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r74 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r75 41 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.39 $Y=2.72
+ $X2=2.225 $Y2=2.72
r76 41 43 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.39 $Y=2.72 $X2=2.99
+ $Y2=2.72
r77 39 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r78 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 36 50 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.145 $Y2=2.72
r80 36 38 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.69 $Y2=2.72
r81 34 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r82 32 43 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=2.72 $X2=2.99
+ $Y2=2.72
r83 32 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.01 $Y=2.72 $X2=3.2
+ $Y2=2.72
r84 31 47 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=3.91 $Y2=2.72
r85 31 33 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.39 $Y=2.72 $X2=3.2
+ $Y2=2.72
r86 27 56 3.27868 $w=3.8e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.285 $Y2=2.72
r87 27 29 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=4.16 $Y=2.635
+ $X2=4.16 $Y2=2.02
r88 23 33 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.2 $Y=2.635 $X2=3.2
+ $Y2=2.72
r89 23 25 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=3.2 $Y=2.635
+ $X2=3.2 $Y2=2.02
r90 19 53 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.72
r91 19 21 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.225 $Y=2.635
+ $X2=2.225 $Y2=2.02
r92 18 50 11.2921 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.395 $Y=2.72
+ $X2=1.145 $Y2=2.72
r93 17 53 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=2.225 $Y2=2.72
r94 17 18 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=1.395 $Y2=2.72
r95 13 50 2.07448 $w=5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.72
r96 13 15 14.7118 $w=4.98e-07 $l=6.15e-07 $layer=LI1_cond $X=1.145 $Y=2.635
+ $X2=1.145 $Y2=2.02
r97 4 29 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.485 $X2=4.185 $Y2=2.02
r98 3 25 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.485 $X2=3.225 $Y2=2.02
r99 2 21 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=1.485 $X2=2.225 $Y2=2.02
r100 1 15 300 $w=1.7e-07 $l=6.54217e-07 $layer=licon1_PDIFF $count=2 $X=0.915
+ $Y=1.485 $X2=1.18 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%X 1 2 3 4 15 17 19 20 23 27 29 31 36 38 40
+ 42 45 47
c60 29 0 1.13405e-19 $X=4.21 $Y=0.73
r61 45 47 0.205793 $w=2.78e-07 $l=5e-09 $layer=LI1_cond $X=4.35 $Y=0.845
+ $X2=4.35 $Y2=0.85
r62 42 45 3.11269 $w=2.8e-07 $l=1.15e-07 $layer=LI1_cond $X=4.35 $Y=0.73
+ $X2=4.35 $Y2=0.845
r63 42 47 1.64635 $w=2.78e-07 $l=4e-08 $layer=LI1_cond $X=4.35 $Y=0.89 $X2=4.35
+ $Y2=0.85
r64 41 42 26.5473 $w=2.78e-07 $l=6.45e-07 $layer=LI1_cond $X=4.35 $Y=1.535
+ $X2=4.35 $Y2=0.89
r65 34 36 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.745 $Y=0.68
+ $X2=2.84 $Y2=0.68
r66 32 40 4.43576 $w=2.27e-07 $l=9.5e-08 $layer=LI1_cond $X=3.8 $Y=1.65
+ $X2=3.705 $Y2=1.65
r67 31 41 6.90206 $w=2.3e-07 $l=1.88944e-07 $layer=LI1_cond $X=4.21 $Y=1.65
+ $X2=4.35 $Y2=1.535
r68 31 32 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.21 $Y=1.65 $X2=3.8
+ $Y2=1.65
r69 30 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.8 $Y=0.73 $X2=3.705
+ $Y2=0.73
r70 29 42 3.78936 $w=2.3e-07 $l=1.4e-07 $layer=LI1_cond $X=4.21 $Y=0.73 $X2=4.35
+ $Y2=0.73
r71 29 30 20.5435 $w=2.28e-07 $l=4.1e-07 $layer=LI1_cond $X=4.21 $Y=0.73 $X2=3.8
+ $Y2=0.73
r72 25 40 1.99853 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=1.65
r73 25 27 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.705 $Y=1.765
+ $X2=3.705 $Y2=1.96
r74 21 38 2.03875 $w=1.9e-07 $l=1.15e-07 $layer=LI1_cond $X=3.705 $Y=0.615
+ $X2=3.705 $Y2=0.73
r75 21 23 11.3828 $w=1.88e-07 $l=1.95e-07 $layer=LI1_cond $X=3.705 $Y=0.615
+ $X2=3.705 $Y2=0.42
r76 19 40 4.43576 $w=2.27e-07 $l=9.64883e-08 $layer=LI1_cond $X=3.61 $Y=1.647
+ $X2=3.705 $Y2=1.65
r77 19 20 39.4392 $w=2.23e-07 $l=7.7e-07 $layer=LI1_cond $X=3.61 $Y=1.647
+ $X2=2.84 $Y2=1.647
r78 17 38 4.39427 $w=2.3e-07 $l=9.5e-08 $layer=LI1_cond $X=3.61 $Y=0.73
+ $X2=3.705 $Y2=0.73
r79 17 36 38.5818 $w=2.28e-07 $l=7.7e-07 $layer=LI1_cond $X=3.61 $Y=0.73
+ $X2=2.84 $Y2=0.73
r80 13 20 6.87974 $w=2.25e-07 $l=1.5331e-07 $layer=LI1_cond $X=2.745 $Y=1.76
+ $X2=2.84 $Y2=1.647
r81 13 15 11.6746 $w=1.88e-07 $l=2e-07 $layer=LI1_cond $X=2.745 $Y=1.76
+ $X2=2.745 $Y2=1.96
r82 4 40 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=3.555
+ $Y=1.485 $X2=3.705 $Y2=1.62
r83 4 27 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=3.555
+ $Y=1.485 $X2=3.705 $Y2=1.96
r84 3 15 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.485 $X2=2.745 $Y2=1.96
r85 2 38 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.705 $Y2=0.76
r86 2 23 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=3.515
+ $Y=0.235 $X2=3.705 $Y2=0.42
r87 1 34 182 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.745 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3_4%VGND 1 2 3 12 14 15 21 23 32 37 40 41
r65 40 43 9.54783 $w=4.6e-07 $l=3.6e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.285
+ $Y2=0.36
r66 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r67 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r68 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r70 32 40 6.6364 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.285
+ $Y2=0
r71 32 34 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.91
+ $Y2=0
r72 31 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r73 31 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r74 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r75 28 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.22
+ $Y2=0
r76 28 30 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=2.385 $Y=0 $X2=2.99
+ $Y2=0
r77 23 37 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.22
+ $Y2=0
r78 23 25 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=0.23 $Y2=0
r79 21 38 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r80 21 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r81 17 34 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=0 $X2=3.91
+ $Y2=0
r82 15 30 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.99
+ $Y2=0
r83 14 19 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.2
+ $Y2=0.36
r84 14 17 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.39
+ $Y2=0
r85 14 15 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.2 $Y=0 $X2=3.01
+ $Y2=0
r86 10 37 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0
r87 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.22 $Y=0.085
+ $X2=2.22 $Y2=0.36
r88 3 43 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=4.045
+ $Y=0.235 $X2=4.185 $Y2=0.36
r89 2 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.235 $X2=3.225 $Y2=0.36
r90 1 12 182 $w=1.7e-07 $l=3.46915e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.22 $Y2=0.36
.ends

