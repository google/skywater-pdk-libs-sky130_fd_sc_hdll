* File: sky130_fd_sc_hdll__einvp_1.pxi.spice
* Created: Wed Sep  2 08:31:33 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVP_1%TE N_TE_M1003_g N_TE_c_42_n N_TE_c_47_n
+ N_TE_c_48_n N_TE_M1001_g N_TE_c_43_n N_TE_c_44_n N_TE_M1005_g TE TE
+ N_TE_c_45_n PM_SKY130_FD_SC_HDLL__EINVP_1%TE
x_PM_SKY130_FD_SC_HDLL__EINVP_1%A_27_47# N_A_27_47#_M1003_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_74_n N_A_27_47#_M1000_g N_A_27_47#_c_75_n N_A_27_47#_c_80_n
+ N_A_27_47#_c_76_n N_A_27_47#_c_77_n N_A_27_47#_c_81_n N_A_27_47#_c_82_n
+ N_A_27_47#_c_78_n PM_SKY130_FD_SC_HDLL__EINVP_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVP_1%A N_A_c_132_n N_A_M1002_g N_A_c_135_n
+ N_A_M1004_g A A A N_A_c_134_n PM_SKY130_FD_SC_HDLL__EINVP_1%A
x_PM_SKY130_FD_SC_HDLL__EINVP_1%VPWR N_VPWR_M1001_d N_VPWR_c_162_n
+ N_VPWR_c_163_n VPWR N_VPWR_c_164_n N_VPWR_c_161_n N_VPWR_c_166_n
+ N_VPWR_c_167_n PM_SKY130_FD_SC_HDLL__EINVP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVP_1%Z N_Z_M1002_d N_Z_M1004_d N_Z_c_196_n
+ N_Z_c_203_n Z Z Z Z PM_SKY130_FD_SC_HDLL__EINVP_1%Z
x_PM_SKY130_FD_SC_HDLL__EINVP_1%VGND N_VGND_M1003_d VGND N_VGND_c_230_n
+ N_VGND_c_231_n N_VGND_c_232_n N_VGND_c_233_n
+ PM_SKY130_FD_SC_HDLL__EINVP_1%VGND
cc_1 VNB N_TE_M1003_g 0.0344245f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_TE_c_42_n 0.0270103f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_3 VNB N_TE_c_43_n 0.0287017f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.035
cc_4 VNB N_TE_c_44_n 0.0163246f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.96
cc_5 VNB N_TE_c_45_n 0.0157585f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_6 VNB N_A_27_47#_c_74_n 0.032401f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_7 VNB N_A_27_47#_c_75_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.96
cc_8 VNB N_A_27_47#_c_76_n 0.00290698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_77_n 0.0100644f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.035
cc_10 VNB N_A_27_47#_c_78_n 0.00464834f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.19
cc_11 VNB N_A_c_132_n 0.0254329f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.96
cc_12 VNB A 0.0141935f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_13 VNB N_A_c_134_n 0.0399523f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_14 VNB N_VPWR_c_161_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Z_c_196_n 0.00354501f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_16 VNB Z 0.0239154f $X=-0.19 $Y=-0.24 $X2=0.87 $Y2=1.035
cc_17 VNB N_VGND_c_230_n 0.0352237f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_18 VNB N_VGND_c_231_n 0.163936f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_232_n 0.0143174f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_20 VNB N_VGND_c_233_n 0.0187033f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_TE_c_42_n 0.00361987f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_22 VPB N_TE_c_47_n 0.0442496f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_23 VPB N_TE_c_48_n 0.0303777f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_24 VPB N_TE_c_45_n 0.0208919f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_25 VPB N_A_27_47#_c_74_n 0.0297645f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_26 VPB N_A_27_47#_c_80_n 0.0155207f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_27 VPB N_A_27_47#_c_81_n 0.00442449f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_28 VPB N_A_27_47#_c_82_n 0.0101173f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_29 VPB N_A_27_47#_c_78_n 0.00588859f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.19
cc_30 VPB N_A_c_135_n 0.019994f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB A 0.025575f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_32 VPB N_A_c_134_n 0.0184221f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_33 VPB N_VPWR_c_162_n 0.0143812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_163_n 0.00443975f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_35 VPB N_VPWR_c_164_n 0.0277791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_161_n 0.0456683f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_166_n 0.0143174f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_38 VPB N_VPWR_c_167_n 0.00572156f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.53
cc_39 VPB N_Z_c_196_n 0.00139111f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_40 VPB Z 0.0151105f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.035
cc_41 N_TE_c_43_n N_A_27_47#_c_74_n 0.00267339f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_42 N_TE_c_48_n N_A_27_47#_c_80_n 0.00465345f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_43 N_TE_M1003_g N_A_27_47#_c_76_n 0.0133165f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_44 N_TE_c_42_n N_A_27_47#_c_76_n 3.50292e-19 $X=0.495 $Y=1.325 $X2=0 $Y2=0
cc_45 N_TE_c_43_n N_A_27_47#_c_76_n 0.00460481f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_46 N_TE_c_44_n N_A_27_47#_c_76_n 0.0108703f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_47 N_TE_c_45_n N_A_27_47#_c_76_n 0.019301f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_48 N_TE_c_45_n N_A_27_47#_c_77_n 0.0238604f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_49 N_TE_c_48_n N_A_27_47#_c_81_n 0.017012f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_50 N_TE_c_45_n N_A_27_47#_c_81_n 0.0193441f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_51 N_TE_c_45_n N_A_27_47#_c_82_n 0.0239512f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_52 N_TE_M1003_g N_A_27_47#_c_78_n 0.00353276f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_53 N_TE_c_42_n N_A_27_47#_c_78_n 0.0203673f $X=0.495 $Y=1.325 $X2=0 $Y2=0
cc_54 N_TE_c_43_n N_A_27_47#_c_78_n 0.0163163f $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_55 N_TE_c_44_n N_A_27_47#_c_78_n 0.0059842f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_56 N_TE_c_45_n N_A_27_47#_c_78_n 0.0621966f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_57 N_TE_c_48_n N_VPWR_c_163_n 0.0129436f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_58 N_TE_c_48_n N_VPWR_c_161_n 0.00472246f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_59 N_TE_c_48_n N_VPWR_c_166_n 0.00316478f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_60 N_TE_M1003_g N_VGND_c_231_n 0.00500115f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_61 N_TE_M1003_g N_VGND_c_232_n 0.00341689f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_62 N_TE_M1003_g N_VGND_c_233_n 0.00891715f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_63 N_TE_c_43_n N_VGND_c_233_n 2.84564e-19 $X=0.87 $Y=1.035 $X2=0 $Y2=0
cc_64 N_TE_c_44_n N_VGND_c_233_n 0.0204061f $X=0.945 $Y=0.96 $X2=0 $Y2=0
cc_65 N_A_27_47#_c_76_n N_A_c_132_n 9.90876e-19 $X=0.765 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_27_47#_c_78_n N_A_c_132_n 9.9219e-19 $X=1.605 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_27_47#_c_74_n N_A_c_135_n 0.0273887f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_78_n N_A_c_135_n 5.49191e-19 $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_27_47#_c_74_n N_A_c_134_n 0.0119509f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_27_47#_c_78_n N_A_c_134_n 6.49022e-19 $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_81_n N_VPWR_M1001_d 0.0165297f $X=0.765 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_27_47#_c_78_n N_VPWR_M1001_d 0.0162533f $X=1.605 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_27_47#_c_80_n N_VPWR_c_163_n 0.0185477f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_81_n N_VPWR_c_163_n 0.085954f $X=0.765 $Y=1.98 $X2=0 $Y2=0
cc_75 N_A_27_47#_M1001_s N_VPWR_c_161_n 0.00241145f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_76 N_A_27_47#_c_80_n N_VPWR_c_161_n 0.00989054f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_81_n N_VPWR_c_161_n 0.00966156f $X=0.765 $Y=1.98 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_80_n N_VPWR_c_166_n 0.0179755f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_81_n N_VPWR_c_166_n 0.00275296f $X=0.765 $Y=1.98 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_74_n N_VPWR_c_167_n 0.0248548f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_74_n N_Z_c_196_n 0.00620124f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_76_n N_Z_c_196_n 0.0010987f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_78_n N_Z_c_196_n 0.046658f $X=1.605 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_74_n N_Z_c_203_n 0.00358172f $X=1.57 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_76_n Z 0.00900095f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_76_n N_VGND_M1003_d 0.0040323f $X=0.765 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_27_47#_c_78_n N_VGND_M1003_d 8.38854e-19 $X=1.605 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_27_47#_c_76_n N_VGND_c_230_n 0.0035086f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_89 N_A_27_47#_M1003_s N_VGND_c_231_n 0.00229009f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_c_75_n N_VGND_c_231_n 0.00989054f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_76_n N_VGND_c_231_n 0.014355f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_75_n N_VGND_c_232_n 0.0177719f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_76_n N_VGND_c_232_n 0.00273399f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_76_n N_VGND_c_233_n 0.0680352f $X=0.765 $Y=0.74 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_76_n A_204_47# 0.0144983f $X=0.765 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_27_47#_c_78_n A_204_47# 0.00100307f $X=1.605 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_c_135_n N_VPWR_c_164_n 0.00429397f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_135_n N_VPWR_c_161_n 0.00740777f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_135_n N_VPWR_c_167_n 0.00304135f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_100 A N_Z_M1004_d 0.0110954f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_101 N_A_c_132_n N_Z_c_196_n 0.0108246f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_c_135_n N_Z_c_196_n 0.022237f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_103 A N_Z_c_196_n 0.0555592f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A_c_134_n N_Z_c_196_n 0.0120508f $X=2.205 $Y=1.202 $X2=0 $Y2=0
cc_105 N_A_c_135_n N_Z_c_203_n 0.00517799f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_c_132_n Z 0.0234059f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_107 A Z 0.021531f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A_c_134_n Z 0.00600202f $X=2.205 $Y=1.202 $X2=0 $Y2=0
cc_109 N_A_c_135_n Z 0.0121935f $X=2.205 $Y=1.41 $X2=0 $Y2=0
cc_110 A Z 0.0197866f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_111 N_A_c_132_n N_VGND_c_230_n 0.00357877f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_c_132_n N_VGND_c_231_n 0.00764649f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A_c_132_n N_VGND_c_233_n 0.00355303f $X=2.18 $Y=0.995 $X2=0 $Y2=0
cc_114 N_VPWR_c_161_n A_332_297# 0.0113589f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_115 N_VPWR_c_167_n A_332_297# 0.00382754f $X=1.74 $Y=2.52 $X2=-0.19 $Y2=-0.24
cc_116 N_VPWR_c_161_n N_Z_M1004_d 0.00225742f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_117 N_VPWR_c_164_n N_Z_c_203_n 0.0101671f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_118 N_VPWR_c_161_n N_Z_c_203_n 0.00654677f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_119 N_VPWR_c_167_n N_Z_c_203_n 0.0159044f $X=1.74 $Y=2.52 $X2=0 $Y2=0
cc_120 N_VPWR_c_164_n Z 0.0291486f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_121 N_VPWR_c_161_n Z 0.01706f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_122 A_332_297# N_Z_c_196_n 0.00718748f $X=1.66 $Y=1.485 $X2=0.15 $Y2=2.635
cc_123 A_332_297# N_Z_c_203_n 0.00485573f $X=1.66 $Y=1.485 $X2=0 $Y2=0
cc_124 Z N_VGND_c_230_n 0.0402646f $X=2.4 $Y=0.425 $X2=0 $Y2=0
cc_125 N_Z_M1002_d N_VGND_c_231_n 0.00258538f $X=2.255 $Y=0.235 $X2=0 $Y2=0
cc_126 Z N_VGND_c_231_n 0.0239314f $X=2.4 $Y=0.425 $X2=0 $Y2=0
cc_127 Z N_VGND_c_233_n 0.00945052f $X=2.4 $Y=0.425 $X2=0 $Y2=0
cc_128 N_Z_c_196_n A_204_47# 0.00128538f $X=2.067 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_129 Z A_204_47# 0.0148409f $X=2.4 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_130 N_VGND_c_231_n A_204_47# 0.0157178f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_131 N_VGND_c_233_n A_204_47# 0.0128716f $X=1.5 $Y=0.2 $X2=-0.19 $Y2=-0.24
