* File: sky130_fd_sc_hdll__or2b_2.spice
* Created: Thu Aug 27 19:23:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or2b_2.pex.spice"
.subckt sky130_fd_sc_hdll__or2b_2  VNB VPB B_N A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_B_N_M1000_g N_A_27_53#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.16695 AS=0.1302 PD=1.215 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.8 A=0.063 P=1.14 MULT=1
MM1001 N_A_228_297#_M1001_d N_A_27_53#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.16695 PD=0.69 PS=1.215 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75001.2 SB=75001.9 A=0.063 P=1.14 MULT=1
MM1009 N_VGND_M1009_d N_A_M1009_g N_A_228_297#_M1001_d VNB NSHORT L=0.15 W=0.42
+ AD=0.100977 AS=0.0567 PD=0.855701 PS=0.69 NRD=27.132 NRS=0 M=1 R=2.8
+ SA=75001.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1009_d N_A_228_297#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.156273 AS=0.16575 PD=1.3243 PS=1.16 NRD=11.988 NRS=34.152 M=1 R=4.33333
+ SA=75001.5 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_228_297#_M1007_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.16575 PD=1.87 PS=1.16 NRD=3.684 NRS=8.304 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_53#_M1003_d N_B_N_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1004 A_318_297# N_A_27_53#_M1004_g N_A_228_297#_M1004_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0483 AS=0.1134 PD=0.65 PS=1.38 NRD=28.1316 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g A_318_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0483 PD=0.804507 PS=0.65 NRD=76.83 NRS=28.1316 M=1 R=2.33333
+ SA=90000.6 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1005_d N_A_228_297#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.218803 AS=0.24 PD=1.91549 PS=1.48 NRD=1.9503 NRS=38.3953 M=1 R=5.55556
+ SA=90000.6 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_228_297#_M1008_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.24 PD=2.59 PS=1.48 NRD=5.91 NRS=0.9653 M=1 R=5.55556 SA=90001.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_62 VPB 0 8.49032e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or2b_2.pxi.spice"
*
.ends
*
*
