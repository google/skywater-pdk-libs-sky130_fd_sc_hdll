* File: sky130_fd_sc_hdll__xor2_2.pex.spice
* Created: Wed Sep  2 08:54:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 26 28 29 31 38 40 41 42 47 52
c126 52 0 1.92034e-19 $X=3.355 $Y=1.202
c127 38 0 1.47612e-19 $X=0.84 $Y=1.175
c128 26 0 1.61073e-19 $X=0.84 $Y=1.445
r129 52 53 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=3.355 $Y=1.202
+ $X2=3.38 $Y2=1.202
r130 49 50 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=2.91 $Y=1.202
+ $X2=2.935 $Y2=1.202
r131 47 48 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.202
+ $X2=1.005 $Y2=1.202
r132 44 45 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.485 $Y=1.202
+ $X2=0.51 $Y2=1.202
r133 41 42 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.86 $Y=1.53
+ $X2=1.15 $Y2=1.53
r134 40 42 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.925 $Y=1.53
+ $X2=1.15 $Y2=1.53
r135 36 47 27.9053 $w=3.8e-07 $l=2.2e-07 $layer=POLY_cond $X=0.76 $Y=1.202
+ $X2=0.98 $Y2=1.202
r136 36 45 31.7105 $w=3.8e-07 $l=2.5e-07 $layer=POLY_cond $X=0.76 $Y=1.202
+ $X2=0.51 $Y2=1.202
r137 35 38 4.43636 $w=1.98e-07 $l=8e-08 $layer=LI1_cond $X=0.76 $Y=1.175
+ $X2=0.84 $Y2=1.175
r138 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.76
+ $Y=1.16 $X2=0.76 $Y2=1.16
r139 32 52 5.11406 $w=3.77e-07 $l=4e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.355 $Y2=1.202
r140 32 50 48.5836 $w=3.77e-07 $l=3.8e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=2.935 $Y2=1.202
r141 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.315
+ $Y=1.16 $X2=3.315 $Y2=1.16
r142 29 31 68.4864 $w=1.98e-07 $l=1.235e-06 $layer=LI1_cond $X=2.08 $Y=1.175
+ $X2=3.315 $Y2=1.175
r143 28 41 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.97 $Y=1.445
+ $X2=1.86 $Y2=1.53
r144 27 29 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=1.97 $Y=1.275
+ $X2=2.08 $Y2=1.175
r145 27 28 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=1.97 $Y=1.275
+ $X2=1.97 $Y2=1.445
r146 26 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.84 $Y=1.445
+ $X2=0.925 $Y2=1.53
r147 25 38 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.84 $Y=1.275 $X2=0.84
+ $Y2=1.175
r148 25 26 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.84 $Y=1.275
+ $X2=0.84 $Y2=1.445
r149 22 53 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.202
r150 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r151 19 52 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.355 $Y=0.995
+ $X2=3.355 $Y2=1.202
r152 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.355 $Y=0.995
+ $X2=3.355 $Y2=0.56
r153 16 50 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.935 $Y2=1.202
r154 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.935 $Y=0.995
+ $X2=2.935 $Y2=0.56
r155 13 49 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.202
r156 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.985
r157 10 48 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r158 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r159 7 47 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.202
r160 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r161 4 45 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.202
r162 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.985
r163 1 44 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=1.202
r164 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.485 $Y=0.995
+ $X2=0.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 31 36 37 43 44
c116 37 0 1.47612e-19 $X=1.92 $Y=1.202
c117 31 0 1.92034e-19 $X=3.91 $Y=1.19
c118 1 0 1.61073e-19 $X=1.45 $Y=1.41
r119 44 45 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=4.375 $Y=1.202
+ $X2=4.4 $Y2=1.202
r120 43 51 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=4.275 $Y=1.175
+ $X2=3.91 $Y2=1.175
r121 42 44 12.8191 $w=3.76e-07 $l=1e-07 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.375 $Y2=1.202
r122 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.275
+ $Y=1.16 $X2=4.275 $Y2=1.16
r123 40 42 54.4814 $w=3.76e-07 $l=4.25e-07 $layer=POLY_cond $X=3.85 $Y=1.202
+ $X2=4.275 $Y2=1.202
r124 39 40 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=3.825 $Y=1.202
+ $X2=3.85 $Y2=1.202
r125 37 38 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.92 $Y=1.202
+ $X2=1.945 $Y2=1.202
r126 35 37 56.4447 $w=3.8e-07 $l=4.45e-07 $layer=POLY_cond $X=1.475 $Y=1.202
+ $X2=1.92 $Y2=1.202
r127 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.475
+ $Y=1.16 $X2=1.475 $Y2=1.16
r128 33 35 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.45 $Y=1.202
+ $X2=1.475 $Y2=1.202
r129 31 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=1.19
+ $X2=3.91 $Y2=1.19
r130 29 36 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=1.25 $Y=1.175
+ $X2=1.475 $Y2=1.175
r131 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.25 $Y=1.19
+ $X2=1.25 $Y2=1.19
r132 26 28 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.395 $Y=1.19
+ $X2=1.25 $Y2=1.19
r133 25 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.765 $Y=1.19
+ $X2=3.91 $Y2=1.19
r134 25 26 2.93316 $w=1.4e-07 $l=2.37e-06 $layer=MET1_cond $X=3.765 $Y=1.19
+ $X2=1.395 $Y2=1.19
r135 22 45 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.4 $Y=0.995
+ $X2=4.4 $Y2=1.202
r136 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.4 $Y=0.995
+ $X2=4.4 $Y2=0.56
r137 19 44 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.202
r138 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.375 $Y=1.41
+ $X2=4.375 $Y2=1.985
r139 16 40 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.202
r140 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.85 $Y2=1.985
r141 13 39 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.825 $Y=0.995
+ $X2=3.825 $Y2=1.202
r142 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.825 $Y=0.995
+ $X2=3.825 $Y2=0.56
r143 10 38 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=1.202
r144 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.945 $Y=0.995
+ $X2=1.945 $Y2=0.56
r145 7 37 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.202
r146 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.92 $Y=1.41
+ $X2=1.92 $Y2=1.985
r147 4 35 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=1.202
r148 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.475 $Y=0.995
+ $X2=1.475 $Y2=0.56
r149 1 33 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.202
r150 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.45 $Y=1.41
+ $X2=1.45 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%A_112_47# 1 2 3 10 12 13 15 16 18 19 21 23
+ 24 25 26 27 30 32 36 38 41 42 43 45 46 48 51 52 60
c165 16 0 1.72656e-19 $X=5.835 $Y=1.41
r166 60 61 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.835 $Y=1.202
+ $X2=5.86 $Y2=1.202
r167 57 58 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.34 $Y=1.202
+ $X2=5.365 $Y2=1.202
r168 52 55 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.685 $Y=1.87
+ $X2=1.685 $Y2=1.96
r169 49 60 34.8816 $w=3.8e-07 $l=2.75e-07 $layer=POLY_cond $X=5.56 $Y=1.202
+ $X2=5.835 $Y2=1.202
r170 49 58 24.7342 $w=3.8e-07 $l=1.95e-07 $layer=POLY_cond $X=5.56 $Y=1.202
+ $X2=5.365 $Y2=1.202
r171 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.56
+ $Y=1.16 $X2=5.56 $Y2=1.16
r172 46 48 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.185 $Y=1.16
+ $X2=5.56 $Y2=1.16
r173 44 46 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.1 $Y=1.245
+ $X2=5.185 $Y2=1.16
r174 44 45 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=5.1 $Y=1.245 $X2=5.1
+ $Y2=1.445
r175 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.015 $Y=1.53
+ $X2=5.1 $Y2=1.445
r176 42 43 169.299 $w=1.68e-07 $l=2.595e-06 $layer=LI1_cond $X=5.015 $Y=1.53
+ $X2=2.42 $Y2=1.53
r177 40 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=1.615
+ $X2=2.42 $Y2=1.53
r178 40 41 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.335 $Y=1.615
+ $X2=2.335 $Y2=1.785
r179 39 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.81 $Y=1.87
+ $X2=1.685 $Y2=1.87
r180 38 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.25 $Y=1.87
+ $X2=2.335 $Y2=1.785
r181 38 39 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.25 $Y=1.87
+ $X2=1.81 $Y2=1.87
r182 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.66 $Y=0.725
+ $X2=1.66 $Y2=0.39
r183 33 51 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.91 $Y=0.815
+ $X2=0.72 $Y2=0.815
r184 32 34 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=1.47 $Y=0.815
+ $X2=1.66 $Y2=0.725
r185 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.47 $Y=0.815
+ $X2=0.91 $Y2=0.815
r186 28 51 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=0.72 $Y=0.725 $X2=0.72
+ $Y2=0.815
r187 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.72 $Y=0.725
+ $X2=0.72 $Y2=0.39
r188 26 52 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.56 $Y=1.87
+ $X2=1.685 $Y2=1.87
r189 26 27 82.8556 $w=1.68e-07 $l=1.27e-06 $layer=LI1_cond $X=1.56 $Y=1.87
+ $X2=0.29 $Y2=1.87
r190 24 51 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.53 $Y=0.815
+ $X2=0.72 $Y2=0.815
r191 24 25 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=0.53 $Y=0.815
+ $X2=0.29 $Y2=0.815
r192 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.205 $Y=1.785
+ $X2=0.29 $Y2=1.87
r193 22 25 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.29 $Y2=0.815
r194 22 23 57.4118 $w=1.68e-07 $l=8.8e-07 $layer=LI1_cond $X=0.205 $Y=0.905
+ $X2=0.205 $Y2=1.785
r195 19 61 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.86 $Y=0.995
+ $X2=5.86 $Y2=1.202
r196 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.86 $Y=0.995
+ $X2=5.86 $Y2=0.56
r197 16 60 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.835 $Y=1.41
+ $X2=5.835 $Y2=1.202
r198 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.835 $Y=1.41
+ $X2=5.835 $Y2=1.985
r199 13 58 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.202
r200 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.985
r201 10 57 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=1.202
r202 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=0.56
r203 3 55 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.54
+ $Y=1.485 $X2=1.685 $Y2=1.96
r204 2 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=1.55
+ $Y=0.235 $X2=1.685 $Y2=0.39
r205 1 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.56
+ $Y=0.235 $X2=0.745 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%A_27_297# 1 2 3 10 13 17 18 21 24 25
c56 24 0 1.9698e-19 $X=1.25 $Y=2.21
r57 25 31 8.39676 $w=2.47e-07 $l=1.7e-07 $layer=LI1_cond $X=1.215 $Y=2.21
+ $X2=1.215 $Y2=2.38
r58 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.25 $Y=2.21
+ $X2=1.25 $Y2=2.21
r59 20 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.21
+ $X2=0.23 $Y2=2.21
r60 18 20 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.375 $Y=2.21
+ $X2=0.23 $Y2=2.21
r61 17 24 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.105 $Y=2.21
+ $X2=1.25 $Y2=2.21
r62 17 18 0.903464 $w=1.4e-07 $l=7.3e-07 $layer=MET1_cond $X=1.105 $Y=2.21
+ $X2=0.375 $Y2=2.21
r63 13 15 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.155 $Y=2.3 $X2=2.155
+ $Y2=2.38
r64 11 31 2.92482 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.34 $Y=2.38
+ $X2=1.215 $Y2=2.38
r65 10 15 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.03 $Y=2.38
+ $X2=2.155 $Y2=2.38
r66 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.03 $Y=2.38 $X2=1.34
+ $Y2=2.38
r67 3 13 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.01
+ $Y=1.485 $X2=2.155 $Y2=2.3
r68 2 25 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.07
+ $Y=1.485 $X2=1.215 $Y2=2.3
r69 1 21 600 $w=1.7e-07 $l=8.82227e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%VPWR 1 2 3 14 18 22 25 26 28 29 30 46 47 50
c88 25 0 1.9698e-19 $X=3.02 $Y=2.72
r89 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r90 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r91 44 47 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r92 43 46 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r93 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r94 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r95 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 38 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r98 35 38 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r99 35 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 34 37 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r101 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 32 50 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=0.745 $Y2=2.72
r103 32 34 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.87 $Y=2.72
+ $X2=1.15 $Y2=2.72
r104 30 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 28 40 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=3.96 $Y=2.72 $X2=3.91
+ $Y2=2.72
r106 28 29 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.96 $Y=2.72
+ $X2=4.112 $Y2=2.72
r107 27 43 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.37 $Y2=2.72
r108 27 29 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.265 $Y=2.72
+ $X2=4.112 $Y2=2.72
r109 25 37 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.02 $Y=2.72 $X2=2.99
+ $Y2=2.72
r110 25 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=3.145 $Y2=2.72
r111 24 40 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 24 26 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=3.145 $Y2=2.72
r113 20 29 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.112 $Y=2.635
+ $X2=4.112 $Y2=2.72
r114 20 22 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=4.112 $Y=2.635
+ $X2=4.112 $Y2=2.3
r115 16 26 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2.72
r116 16 18 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.145 $Y=2.635
+ $X2=3.145 $Y2=2.3
r117 12 50 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r118 12 14 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.3
r119 3 22 600 $w=1.7e-07 $l=9.09519e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.485 $X2=4.14 $Y2=2.3
r120 2 18 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3
+ $Y=1.485 $X2=3.145 $Y2=2.3
r121 1 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.745 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_297# 1 2 3 4 5 19 20 21 24 28 32 35
+ 38 41 44
r47 43 44 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=5.13 $Y=2.125
+ $X2=5.255 $Y2=2.125
r48 40 43 9.14648 $w=6.78e-07 $l=5.2e-07 $layer=LI1_cond $X=4.61 $Y=2.125
+ $X2=5.13 $Y2=2.125
r49 40 41 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=4.61 $Y=2.125
+ $X2=4.485 $Y2=2.125
r50 35 36 7.68595 $w=3.13e-07 $l=1.75e-07 $layer=LI1_cond $X=2.642 $Y=2.3
+ $X2=2.642 $Y2=2.125
r51 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.07 $Y=2.295
+ $X2=6.07 $Y2=1.96
r52 28 30 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.945 $Y=2.38
+ $X2=6.07 $Y2=2.295
r53 28 44 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.945 $Y=2.38
+ $X2=5.255 $Y2=2.38
r54 27 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.74 $Y=1.87
+ $X2=3.615 $Y2=1.87
r55 27 41 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.74 $Y=1.87
+ $X2=4.485 $Y2=1.87
r56 22 38 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.955
+ $X2=3.615 $Y2=1.87
r57 22 24 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=3.615 $Y=1.955
+ $X2=3.615 $Y2=1.96
r58 20 38 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.49 $Y=1.87
+ $X2=3.615 $Y2=1.87
r59 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.49 $Y=1.87 $X2=2.8
+ $Y2=1.87
r60 19 36 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.695 $Y=1.96
+ $X2=2.695 $Y2=2.125
r61 16 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.695 $Y=1.955
+ $X2=2.8 $Y2=1.87
r62 16 19 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=2.695 $Y=1.955
+ $X2=2.695 $Y2=1.96
r63 5 32 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.925
+ $Y=1.485 $X2=6.07 $Y2=1.96
r64 4 43 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=5.005
+ $Y=1.485 $X2=5.13 $Y2=1.96
r65 3 40 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.465
+ $Y=1.485 $X2=4.61 $Y2=1.96
r66 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.47
+ $Y=1.485 $X2=3.615 $Y2=1.96
r67 1 35 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.485 $X2=2.675 $Y2=2.3
r68 1 19 600 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=1 $X=2.55
+ $Y=1.485 $X2=2.675 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%X 1 2 3 14 16 19 23 26 27 29 30
c54 19 0 1.72656e-19 $X=6.167 $Y=1.415
r55 25 27 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=5.6 $Y=0.775
+ $X2=5.765 $Y2=0.775
r56 25 26 10.6316 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=5.6 $Y=0.775
+ $X2=5.385 $Y2=0.775
r57 23 26 66.5455 $w=1.78e-07 $l=1.08e-06 $layer=LI1_cond $X=4.305 $Y=0.815
+ $X2=5.385 $Y2=0.815
r58 21 23 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.14 $Y=0.775
+ $X2=4.305 $Y2=0.775
r59 19 30 2.73707 $w=3.65e-07 $l=1.05e-07 $layer=LI1_cond $X=6.167 $Y=1.415
+ $X2=6.167 $Y2=1.52
r60 18 19 16.1026 $w=3.63e-07 $l=5.1e-07 $layer=LI1_cond $X=6.167 $Y=0.905
+ $X2=6.167 $Y2=1.415
r61 16 18 7.89155 $w=1.8e-07 $l=2.22495e-07 $layer=LI1_cond $X=5.985 $Y=0.815
+ $X2=6.167 $Y2=0.905
r62 16 27 13.5556 $w=1.78e-07 $l=2.2e-07 $layer=LI1_cond $X=5.985 $Y=0.815
+ $X2=5.765 $Y2=0.815
r63 15 29 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.725 $Y=1.52
+ $X2=5.6 $Y2=1.52
r64 14 30 4.74426 $w=2.1e-07 $l=1.82e-07 $layer=LI1_cond $X=5.985 $Y=1.52
+ $X2=6.167 $Y2=1.52
r65 14 15 13.7316 $w=2.08e-07 $l=2.6e-07 $layer=LI1_cond $X=5.985 $Y=1.52
+ $X2=5.725 $Y2=1.52
r66 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.455
+ $Y=1.485 $X2=5.6 $Y2=1.62
r67 2 25 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.6 $Y2=0.73
r68 1 21 182 $w=1.7e-07 $l=6.03179e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.14 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%VGND 1 2 3 4 5 6 19 21 23 27 29 33 37 41 45
+ 48 49 51 52 53 54 55 56 73 78 81
r102 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r103 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r104 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r105 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r106 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r107 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r108 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r109 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r110 64 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.83 $Y2=0
r111 63 66 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r112 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r113 61 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r114 61 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r115 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r116 58 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.155
+ $Y2=0
r117 58 60 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.24 $Y=0 $X2=2.99
+ $Y2=0
r118 56 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r119 56 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 54 69 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=5.985 $Y=0
+ $X2=5.75 $Y2=0
r121 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=0 $X2=6.07
+ $Y2=0
r122 53 72 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.21
+ $Y2=0
r123 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.155 $Y=0 $X2=6.07
+ $Y2=0
r124 51 66 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=4.83 $Y2=0
r125 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0 $X2=5.13
+ $Y2=0
r126 50 69 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=5.215 $Y=0
+ $X2=5.75 $Y2=0
r127 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.215 $Y=0 $X2=5.13
+ $Y2=0
r128 48 60 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=2.99
+ $Y2=0
r129 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=0 $X2=3.145
+ $Y2=0
r130 47 63 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.45
+ $Y2=0
r131 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.23 $Y=0 $X2=3.145
+ $Y2=0
r132 43 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0
r133 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.07 $Y=0.085
+ $X2=6.07 $Y2=0.39
r134 39 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.13 $Y=0.085
+ $X2=5.13 $Y2=0
r135 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.13 $Y=0.085
+ $X2=5.13 $Y2=0.39
r136 35 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0
r137 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0.39
r138 31 81 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0
r139 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.155 $Y=0.085
+ $X2=2.155 $Y2=0.39
r140 30 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0 $X2=1.215
+ $Y2=0
r141 29 81 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.155
+ $Y2=0
r142 29 30 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.3
+ $Y2=0
r143 25 78 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0
r144 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.215 $Y=0.085
+ $X2=1.215 $Y2=0.39
r145 24 75 3.40825 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r146 23 78 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.215
+ $Y2=0
r147 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.36
+ $Y2=0
r148 19 75 3.40825 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.18 $Y2=0
r149 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.39
r150 6 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.935
+ $Y=0.235 $X2=6.07 $Y2=0.39
r151 5 41 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.005
+ $Y=0.235 $X2=5.13 $Y2=0.39
r152 4 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.01
+ $Y=0.235 $X2=3.145 $Y2=0.39
r153 3 33 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.02
+ $Y=0.235 $X2=2.155 $Y2=0.39
r154 2 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.215 $Y2=0.39
r155 1 21 182 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.275 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR2_2%A_510_47# 1 2 3 12 14 15 19 20 22
r45 20 22 47.6692 $w=2.18e-07 $l=9.1e-07 $layer=LI1_cond $X=3.7 $Y=0.365
+ $X2=4.61 $Y2=0.365
r46 17 19 7.10673 $w=2.98e-07 $l=1.85e-07 $layer=LI1_cond $X=3.55 $Y=0.725
+ $X2=3.55 $Y2=0.54
r47 16 20 7.02845 $w=2.2e-07 $l=1.97484e-07 $layer=LI1_cond $X=3.55 $Y=0.475
+ $X2=3.7 $Y2=0.365
r48 16 19 2.49696 $w=2.98e-07 $l=6.5e-08 $layer=LI1_cond $X=3.55 $Y=0.475
+ $X2=3.55 $Y2=0.54
r49 14 17 7.38573 $w=1.8e-07 $l=1.89737e-07 $layer=LI1_cond $X=3.4 $Y=0.815
+ $X2=3.55 $Y2=0.725
r50 14 15 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.4 $Y=0.815
+ $X2=2.84 $Y2=0.815
r51 10 15 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=2.675 $Y=0.725
+ $X2=2.84 $Y2=0.815
r52 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.675 $Y=0.725
+ $X2=2.675 $Y2=0.39
r53 3 22 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.475
+ $Y=0.235 $X2=4.61 $Y2=0.39
r54 2 19 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.615 $Y2=0.54
r55 1 12 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=2.55
+ $Y=0.235 $X2=2.675 $Y2=0.39
.ends

