* File: sky130_fd_sc_hdll__clkbuf_8.pex.spice
* Created: Thu Aug 27 19:02:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_8%A 1 3 6 8 10 13 15 16 26
c39 15 0 1.46759e-19 $X=0.23 $Y=0.85
r40 25 26 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.155
+ $X2=1.005 $Y2=1.155
r41 24 25 47.733 $w=5.1e-07 $l=4.55e-07 $layer=POLY_cond $X=0.525 $Y=1.155
+ $X2=0.98 $Y2=1.155
r42 23 24 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=0.5 $Y=1.155
+ $X2=0.525 $Y2=1.155
r43 20 23 24.1288 $w=5.1e-07 $l=2.3e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.5 $Y2=1.155
r44 16 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r45 15 16 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r46 11 26 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.005 $Y=0.9
+ $X2=1.005 $Y2=1.155
r47 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.005 $Y=0.9
+ $X2=1.005 $Y2=0.445
r48 8 25 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.155
r49 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r50 4 24 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.525 $Y=0.9
+ $X2=0.525 $Y2=1.155
r51 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.525 $Y=0.9
+ $X2=0.525 $Y2=0.445
r52 1 23 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.155
r53 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_8%A_118_297# 1 2 9 11 13 16 18 20 23 25 27
+ 30 32 34 37 39 41 44 46 48 51 53 55 56 58 61 65 69 76 79 96
r145 96 97 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=4.82 $Y=1.18
+ $X2=4.845 $Y2=1.18
r146 95 96 56.0194 $w=4.13e-07 $l=4.8e-07 $layer=POLY_cond $X=4.34 $Y=1.18
+ $X2=4.82 $Y2=1.18
r147 94 95 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=4.315 $Y=1.18
+ $X2=4.34 $Y2=1.18
r148 93 94 53.1017 $w=4.13e-07 $l=4.55e-07 $layer=POLY_cond $X=3.86 $Y=1.18
+ $X2=4.315 $Y2=1.18
r149 92 93 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.18
+ $X2=3.86 $Y2=1.18
r150 89 90 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=3.355 $Y=1.18
+ $X2=3.38 $Y2=1.18
r151 88 89 53.1017 $w=4.13e-07 $l=4.55e-07 $layer=POLY_cond $X=2.9 $Y=1.18
+ $X2=3.355 $Y2=1.18
r152 87 88 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=2.875 $Y=1.18
+ $X2=2.9 $Y2=1.18
r153 86 87 53.1017 $w=4.13e-07 $l=4.55e-07 $layer=POLY_cond $X=2.42 $Y=1.18
+ $X2=2.875 $Y2=1.18
r154 85 86 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=2.395 $Y=1.18
+ $X2=2.42 $Y2=1.18
r155 84 85 53.1017 $w=4.13e-07 $l=4.55e-07 $layer=POLY_cond $X=1.94 $Y=1.18
+ $X2=2.395 $Y2=1.18
r156 83 84 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=1.915 $Y=1.18
+ $X2=1.94 $Y2=1.18
r157 80 81 2.91768 $w=4.13e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.18
+ $X2=1.46 $Y2=1.18
r158 77 92 28.0097 $w=4.13e-07 $l=2.4e-07 $layer=POLY_cond $X=3.595 $Y=1.18
+ $X2=3.835 $Y2=1.18
r159 77 90 25.092 $w=4.13e-07 $l=2.15e-07 $layer=POLY_cond $X=3.595 $Y=1.18
+ $X2=3.38 $Y2=1.18
r160 76 77 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.595
+ $Y=1.16 $X2=3.595 $Y2=1.16
r161 74 83 25.6755 $w=4.13e-07 $l=2.2e-07 $layer=POLY_cond $X=1.695 $Y=1.18
+ $X2=1.915 $Y2=1.18
r162 74 81 27.4261 $w=4.13e-07 $l=2.35e-07 $layer=POLY_cond $X=1.695 $Y=1.18
+ $X2=1.46 $Y2=1.18
r163 73 76 87.5857 $w=2.48e-07 $l=1.9e-06 $layer=LI1_cond $X=1.695 $Y=1.2
+ $X2=3.595 $Y2=1.2
r164 73 74 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=1.695
+ $Y=1.16 $X2=1.695 $Y2=1.16
r165 71 79 1.34256 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.87 $Y=1.2
+ $X2=0.745 $Y2=1.2
r166 71 73 38.0306 $w=2.48e-07 $l=8.25e-07 $layer=LI1_cond $X=0.87 $Y=1.2
+ $X2=1.695 $Y2=1.2
r167 67 79 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.325
+ $X2=0.745 $Y2=1.2
r168 67 69 16.8257 $w=2.48e-07 $l=3.65e-07 $layer=LI1_cond $X=0.745 $Y=1.325
+ $X2=0.745 $Y2=1.69
r169 63 79 5.16603 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.075
+ $X2=0.745 $Y2=1.2
r170 63 65 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.745 $Y=1.075
+ $X2=0.745 $Y2=0.445
r171 59 97 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.845 $Y=0.95
+ $X2=4.845 $Y2=1.18
r172 59 61 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.845 $Y=0.95
+ $X2=4.845 $Y2=0.445
r173 56 96 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.18
r174 56 58 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.985
r175 53 95 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.18
r176 53 55 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.985
r177 49 94 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.315 $Y=0.95
+ $X2=4.315 $Y2=1.18
r178 49 51 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.315 $Y=0.95
+ $X2=4.315 $Y2=0.445
r179 46 93 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.18
r180 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.985
r181 42 92 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.835 $Y=0.95
+ $X2=3.835 $Y2=1.18
r182 42 44 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.835 $Y=0.95
+ $X2=3.835 $Y2=0.445
r183 39 90 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.18
r184 39 41 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r185 35 89 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.355 $Y=0.95
+ $X2=3.355 $Y2=1.18
r186 35 37 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.355 $Y=0.95
+ $X2=3.355 $Y2=0.445
r187 32 88 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.9 $Y=1.41 $X2=2.9
+ $Y2=1.18
r188 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.9 $Y=1.41
+ $X2=2.9 $Y2=1.985
r189 28 87 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.875 $Y=0.95
+ $X2=2.875 $Y2=1.18
r190 28 30 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.875 $Y=0.95
+ $X2=2.875 $Y2=0.445
r191 25 86 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.18
r192 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.985
r193 21 85 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.395 $Y=0.95
+ $X2=2.395 $Y2=1.18
r194 21 23 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.395 $Y=0.95
+ $X2=2.395 $Y2=0.445
r195 18 84 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.18
r196 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.985
r197 14 83 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.915 $Y=0.95
+ $X2=1.915 $Y2=1.18
r198 14 16 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.915 $Y=0.95
+ $X2=1.915 $Y2=0.445
r199 11 81 22.226 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.18
r200 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.985
r201 7 80 26.6457 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=1.435 $Y=0.95
+ $X2=1.435 $Y2=1.18
r202 7 9 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=1.435 $Y=0.95
+ $X2=1.435 $Y2=0.445
r203 2 69 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.69
r204 1 65 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_8%VPWR 1 2 3 4 5 6 19 21 23 27 29 33 37 41
+ 45 48 49 51 52 54 55 56 69 70 76 79
c79 6 0 4.2343e-20 $X=4.91 $Y=1.485
c80 5 0 1.26981e-19 $X=3.95 $Y=1.485
r81 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r82 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r83 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r84 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r85 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r86 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r87 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r88 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r89 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r90 61 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r91 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r92 58 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.31 $Y=2.72 $X2=2.18
+ $Y2=2.72
r93 58 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=2.72
+ $X2=2.99 $Y2=2.72
r94 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 56 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 54 66 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.93 $Y=2.72 $X2=4.83
+ $Y2=2.72
r97 54 55 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=4.93 $Y=2.72
+ $X2=5.077 $Y2=2.72
r98 53 69 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.29 $Y2=2.72
r99 53 55 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=5.225 $Y=2.72
+ $X2=5.077 $Y2=2.72
r100 51 63 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=2.72 $X2=3.91
+ $Y2=2.72
r101 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.97 $Y=2.72 $X2=4.1
+ $Y2=2.72
r102 50 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.23 $Y=2.72 $X2=4.83
+ $Y2=2.72
r103 50 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.23 $Y=2.72 $X2=4.1
+ $Y2=2.72
r104 48 60 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=2.72 $X2=2.99
+ $Y2=2.72
r105 48 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.01 $Y=2.72
+ $X2=3.14 $Y2=2.72
r106 47 63 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=3.91 $Y2=2.72
r107 47 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.27 $Y=2.72
+ $X2=3.14 $Y2=2.72
r108 43 55 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=5.077 $Y=2.635
+ $X2=5.077 $Y2=2.72
r109 43 45 16.2123 $w=2.93e-07 $l=4.15e-07 $layer=LI1_cond $X=5.077 $Y=2.635
+ $X2=5.077 $Y2=2.22
r110 39 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.635
+ $X2=4.1 $Y2=2.72
r111 39 41 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=4.1 $Y=2.635
+ $X2=4.1 $Y2=2.22
r112 35 49 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=2.635
+ $X2=3.14 $Y2=2.72
r113 35 37 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=3.14 $Y=2.635
+ $X2=3.14 $Y2=2.22
r114 31 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=2.635
+ $X2=2.18 $Y2=2.72
r115 31 33 18.3948 $w=2.58e-07 $l=4.15e-07 $layer=LI1_cond $X=2.18 $Y=2.635
+ $X2=2.18 $Y2=2.22
r116 30 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=1.22 $Y2=2.72
r117 29 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.05 $Y=2.72
+ $X2=2.18 $Y2=2.72
r118 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.05 $Y=2.72 $X2=1.35
+ $Y2=2.72
r119 25 76 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r120 25 27 41.8869 $w=2.58e-07 $l=9.45e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=1.69
r121 24 73 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r122 23 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=1.22 $Y2=2.72
r123 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=2.72 $X2=0.39
+ $Y2=2.72
r124 19 73 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.195 $Y2=2.72
r125 19 21 36.9172 $w=2.93e-07 $l=9.45e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.69
r126 6 45 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.485 $X2=5.06 $Y2=2.22
r127 5 41 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.485 $X2=4.1 $Y2=2.22
r128 4 37 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.485 $X2=3.14 $Y2=2.22
r129 3 33 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.485 $X2=2.18 $Y2=2.22
r130 2 27 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.22 $Y2=1.69
r131 1 21 300 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.69
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_8%X 1 2 3 4 5 6 7 8 27 31 32 33 37 41 43 47
+ 51 53 57 62 63 65 66 68 69 70 71
c115 69 0 1.69324e-19 $X=4.835 $Y=0.85
r116 71 86 2.07573 $w=6.65e-07 $l=1.2e-07 $layer=LI1_cond $X=4.695 $Y=1.615
+ $X2=4.695 $Y2=1.495
r117 71 86 0.285047 $w=1.068e-06 $l=2.5e-08 $layer=LI1_cond $X=4.695 $Y=1.47
+ $X2=4.695 $Y2=1.495
r118 70 71 3.19252 $w=1.068e-06 $l=2.8e-07 $layer=LI1_cond $X=4.695 $Y=1.19
+ $X2=4.695 $Y2=1.47
r119 69 85 1.49612 $w=6.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=0.82
+ $X2=4.695 $Y2=0.905
r120 69 70 3.0785 $w=1.068e-06 $l=2.7e-07 $layer=LI1_cond $X=4.695 $Y=0.92
+ $X2=4.695 $Y2=1.19
r121 69 85 0.171028 $w=1.068e-06 $l=1.5e-08 $layer=LI1_cond $X=4.695 $Y=0.92
+ $X2=4.695 $Y2=0.905
r122 55 69 1.49612 $w=6.65e-07 $l=1.51658e-07 $layer=LI1_cond $X=4.58 $Y=0.735
+ $X2=4.695 $Y2=0.82
r123 55 57 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.58 $Y=0.735
+ $X2=4.58 $Y2=0.445
r124 54 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.75 $Y=1.615
+ $X2=3.62 $Y2=1.615
r125 53 71 5.17024 $w=2.4e-07 $l=5.35e-07 $layer=LI1_cond $X=4.16 $Y=1.615
+ $X2=4.695 $Y2=1.615
r126 53 54 19.6876 $w=2.38e-07 $l=4.1e-07 $layer=LI1_cond $X=4.16 $Y=1.615
+ $X2=3.75 $Y2=1.615
r127 52 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.75 $Y=0.82
+ $X2=3.62 $Y2=0.82
r128 51 69 6.49904 $w=1.7e-07 $l=5.35e-07 $layer=LI1_cond $X=4.16 $Y=0.82
+ $X2=4.695 $Y2=0.82
r129 51 52 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=4.16 $Y=0.82
+ $X2=3.75 $Y2=0.82
r130 45 66 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.82
r131 45 47 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.445
r132 44 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.79 $Y=1.615
+ $X2=2.66 $Y2=1.615
r133 43 68 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.49 $Y=1.615
+ $X2=3.62 $Y2=1.615
r134 43 44 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=3.49 $Y=1.615
+ $X2=2.79 $Y2=1.615
r135 42 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.79 $Y=0.82
+ $X2=2.66 $Y2=0.82
r136 41 66 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.49 $Y=0.82
+ $X2=3.62 $Y2=0.82
r137 41 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.49 $Y=0.82 $X2=2.79
+ $Y2=0.82
r138 35 63 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.735
+ $X2=2.66 $Y2=0.82
r139 35 37 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.66 $Y=0.735
+ $X2=2.66 $Y2=0.445
r140 34 62 3.55196 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=1.83 $Y=1.615
+ $X2=1.7 $Y2=1.615
r141 33 65 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.53 $Y=1.615
+ $X2=2.66 $Y2=1.615
r142 33 34 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=2.53 $Y=1.615
+ $X2=1.83 $Y2=1.615
r143 31 63 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.53 $Y=0.82
+ $X2=2.66 $Y2=0.82
r144 31 32 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.53 $Y=0.82 $X2=1.83
+ $Y2=0.82
r145 25 32 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.7 $Y=0.735
+ $X2=1.83 $Y2=0.82
r146 25 27 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=1.7 $Y=0.735
+ $X2=1.7 $Y2=0.445
r147 8 71 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.58 $Y2=1.69
r148 7 68 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=3.47
+ $Y=1.485 $X2=3.62 $Y2=1.69
r149 6 65 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=1.485 $X2=2.66 $Y2=1.69
r150 5 62 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=1.55
+ $Y=1.485 $X2=1.7 $Y2=1.69
r151 4 57 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.235 $X2=4.58 $Y2=0.445
r152 3 47 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.62 $Y2=0.445
r153 2 37 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.66 $Y2=0.445
r154 1 27 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.235 $X2=1.7 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_8%VGND 1 2 3 4 5 6 19 21 23 27 29 33 37 41
+ 45 48 49 51 52 54 55 56 69 70 76 79
c84 23 0 1.46759e-19 $X=1.09 $Y=0
r85 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r86 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r87 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r88 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r89 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r90 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r91 64 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r92 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r93 61 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r94 61 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r95 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r96 58 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.18
+ $Y2=0
r97 58 60 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.99
+ $Y2=0
r98 56 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r99 56 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r100 54 66 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.83
+ $Y2=0
r101 54 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.08
+ $Y2=0
r102 53 69 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.29
+ $Y2=0
r103 53 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.08
+ $Y2=0
r104 51 63 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.91
+ $Y2=0
r105 51 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.1
+ $Y2=0
r106 50 66 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.83
+ $Y2=0
r107 50 52 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.1
+ $Y2=0
r108 48 60 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.99
+ $Y2=0
r109 48 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=3.14
+ $Y2=0
r110 47 63 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.91
+ $Y2=0
r111 47 49 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.14
+ $Y2=0
r112 43 55 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.08 $Y=0.085
+ $X2=5.08 $Y2=0
r113 43 45 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=5.08 $Y=0.085
+ $X2=5.08 $Y2=0.4
r114 39 52 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0.085
+ $X2=4.1 $Y2=0
r115 39 41 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=4.1 $Y=0.085
+ $X2=4.1 $Y2=0.4
r116 35 49 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r117 35 37 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.4
r118 31 79 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r119 31 33 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.4
r120 30 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.22
+ $Y2=0
r121 29 79 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.18
+ $Y2=0
r122 29 30 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.35
+ $Y2=0
r123 25 76 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r124 25 27 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.445
r125 24 73 3.93884 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r126 23 76 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.22
+ $Y2=0
r127 23 24 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.39
+ $Y2=0
r128 19 73 3.17127 $w=2.45e-07 $l=1.15521e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.195 $Y2=0
r129 19 21 13.8764 $w=2.43e-07 $l=2.95e-07 $layer=LI1_cond $X=0.267 $Y=0.085
+ $X2=0.267 $Y2=0.38
r130 6 45 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=4.92
+ $Y=0.235 $X2=5.065 $Y2=0.4
r131 5 41 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=0.235 $X2=4.1 $Y2=0.4
r132 4 37 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.235 $X2=3.14 $Y2=0.4
r133 3 33 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.235 $X2=2.18 $Y2=0.4
r134 2 27 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.445
r135 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

