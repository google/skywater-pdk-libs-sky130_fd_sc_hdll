* File: sky130_fd_sc_hdll__o2bb2ai_4.spice
* Created: Thu Aug 27 19:22:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o2bb2ai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o2bb2ai_4  VNB VPB A2_N A1_N B2 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* B2	B2
* A1_N	A1_N
* A2_N	A2_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_27_47#_M1003_d N_A2_N_M1003_g N_A_113_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.182 AS=0.104 PD=1.86 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1021 N_A_27_47#_M1021_d N_A2_N_M1021_g N_A_113_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1022 N_A_27_47#_M1021_d N_A2_N_M1022_g N_A_113_47#_M1022_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1037 N_A_27_47#_M1037_d N_A2_N_M1037_g N_A_113_47#_M1022_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1015_d N_A1_N_M1015_g N_A_27_47#_M1037_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1017 N_VGND_M1015_d N_A1_N_M1017_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1031 N_VGND_M1031_d N_A1_N_M1031_g N_A_27_47#_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1038 N_VGND_M1031_d N_A1_N_M1038_g N_A_27_47#_M1038_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_113_47#_M1006_g N_A_887_47#_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1008 N_Y_M1006_d N_A_113_47#_M1008_g N_A_887_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1028 N_Y_M1028_d N_A_113_47#_M1028_g N_A_887_47#_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75005 A=0.0975 P=1.6 MULT=1
MM1033 N_Y_M1028_d N_A_113_47#_M1033_g N_A_887_47#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.247 PD=1.02 PS=1.41 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_B2_M1000_g N_A_887_47#_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.247 PD=0.97 PS=1.41 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1000_d N_B2_M1013_g N_A_887_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_B2_M1016_g N_A_887_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.5
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1034 N_VGND_M1016_d N_B2_M1034_g N_A_887_47#_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_B1_M1009_g N_A_887_47#_M1034_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1009_d N_B1_M1012_g N_A_887_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.9
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1026_d N_B1_M1026_g N_A_887_47#_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1026_d N_B1_M1027_g N_A_887_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_113_47#_M1002_d N_A2_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90005.8 A=0.18 P=2.36 MULT=1
MM1010 N_A_113_47#_M1002_d N_A2_N_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1018 N_A_113_47#_M1018_d N_A2_N_M1018_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1029 N_A_113_47#_M1018_d N_A2_N_M1029_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1001 N_A_113_47#_M1001_d N_A1_N_M1001_g N_VPWR_M1029_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90004 A=0.18 P=2.36 MULT=1
MM1023 N_A_113_47#_M1001_d N_A1_N_M1023_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1035 N_A_113_47#_M1035_d N_A1_N_M1035_g N_VPWR_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1039 N_A_113_47#_M1035_d N_A1_N_M1039_g N_VPWR_M1039_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.39 PD=1.29 PS=1.78 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1039_s N_A_113_47#_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.39 AS=0.145 PD=1.78 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_113_47#_M1007_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1007_d N_A_113_47#_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1036 N_VPWR_M1036_d N_A_113_47#_M1036_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1011_d N_B2_M1011_g N_A_1361_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1024 N_Y_M1011_d N_B2_M1024_g N_A_1361_297#_M1024_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1030 N_Y_M1030_d N_B2_M1030_g N_A_1361_297#_M1024_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1032 N_Y_M1030_d N_B2_M1032_g N_A_1361_297#_M1032_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_B1_M1005_g N_A_1361_297#_M1032_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1005_d N_B1_M1014_g N_A_1361_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_B1_M1020_g N_A_1361_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1020_d N_B1_M1025_g N_A_1361_297#_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=18.3291 P=26.05
pX41_noxref noxref_14 A2_N A2_N PROBETYPE=1
pX42_noxref noxref_15 A1_N A1_N PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o2bb2ai_4.pxi.spice"
*
.ends
*
*
