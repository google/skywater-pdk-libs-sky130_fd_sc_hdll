* File: sky130_fd_sc_hdll__clkinv_4.pxi.spice
* Created: Wed Sep  2 08:26:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_4%A N_A_c_87_n N_A_M1000_g N_A_M1001_g N_A_c_88_n
+ N_A_M1003_g N_A_c_74_n N_A_M1002_g N_A_c_89_n N_A_M1004_g N_A_c_76_n
+ N_A_M1006_g N_A_c_90_n N_A_M1005_g N_A_c_78_n N_A_M1008_g N_A_c_91_n
+ N_A_M1007_g N_A_c_92_n N_A_M1009_g N_A_c_80_n N_A_c_81_n N_A_c_82_n N_A_c_83_n
+ N_A_c_84_n N_A_c_85_n N_A_c_86_n A A A A A A A A A A
+ PM_SKY130_FD_SC_HDLL__CLKINV_4%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_4%VPWR N_VPWR_M1000_d N_VPWR_M1003_d
+ N_VPWR_M1005_d N_VPWR_M1009_d N_VPWR_c_182_n N_VPWR_c_183_n N_VPWR_c_184_n
+ N_VPWR_c_185_n N_VPWR_c_186_n N_VPWR_c_187_n N_VPWR_c_188_n N_VPWR_c_189_n
+ N_VPWR_c_190_n VPWR N_VPWR_c_191_n N_VPWR_c_192_n N_VPWR_c_181_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_4%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_4%Y N_Y_M1001_d N_Y_M1006_d N_Y_M1000_s
+ N_Y_M1004_s N_Y_M1007_s N_Y_c_233_n N_Y_c_234_n N_Y_c_235_n N_Y_c_245_n
+ N_Y_c_246_n N_Y_c_314_n N_Y_c_247_n N_Y_c_236_n N_Y_c_237_n N_Y_c_318_n
+ N_Y_c_248_n N_Y_c_238_n N_Y_c_239_n N_Y_c_322_n N_Y_c_249_n N_Y_c_250_n
+ N_Y_c_240_n N_Y_c_251_n N_Y_c_241_n N_Y_c_252_n Y Y Y N_Y_c_243_n N_Y_c_254_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_4%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_4%VGND N_VGND_M1001_s N_VGND_M1002_s
+ N_VGND_M1008_s N_VGND_c_350_n N_VGND_c_351_n N_VGND_c_352_n N_VGND_c_353_n
+ N_VGND_c_354_n N_VGND_c_355_n VGND N_VGND_c_356_n N_VGND_c_357_n
+ N_VGND_c_358_n N_VGND_c_359_n N_VGND_c_360_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_4%VGND
cc_1 VNB N_A_M1001_g 0.0380238f $X=-0.19 $Y=-0.24 $X2=0.995 $Y2=0.445
cc_2 VNB N_A_c_74_n 0.0183247f $X=-0.19 $Y=-0.24 $X2=1.4 $Y2=1.16
cc_3 VNB N_A_M1002_g 0.0299271f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=0.445
cc_4 VNB N_A_c_76_n 0.0183228f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_5 VNB N_A_M1006_g 0.029927f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=0.445
cc_6 VNB N_A_c_78_n 0.0183247f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=1.16
cc_7 VNB N_A_M1008_g 0.0401409f $X=-0.19 $Y=-0.24 $X2=2.435 $Y2=0.445
cc_8 VNB N_A_c_80_n 0.0184882f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=1.16
cc_9 VNB N_A_c_81_n 0.0209725f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_10 VNB N_A_c_82_n 0.00629246f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.217
cc_11 VNB N_A_c_83_n 0.00629259f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.217
cc_12 VNB N_A_c_84_n 0.00629259f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=1.217
cc_13 VNB N_A_c_85_n 0.00755835f $X=-0.19 $Y=-0.24 $X2=2.46 $Y2=1.217
cc_14 VNB N_A_c_86_n 0.0397617f $X=-0.19 $Y=-0.24 $X2=2.84 $Y2=1.16
cc_15 VNB N_VPWR_c_181_n 0.155873f $X=-0.19 $Y=-0.24 $X2=2.185 $Y2=1.105
cc_16 VNB N_Y_c_233_n 0.0202092f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.41
cc_17 VNB N_Y_c_234_n 0.0164024f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.985
cc_18 VNB N_Y_c_235_n 0.0104981f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.985
cc_19 VNB N_Y_c_236_n 0.0013073f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=1.16
cc_20 VNB N_Y_c_237_n 0.00732848f $X=-0.19 $Y=-0.24 $X2=2.435 $Y2=0.445
cc_21 VNB N_Y_c_238_n 0.00130439f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.16
cc_22 VNB N_Y_c_239_n 0.0194357f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.217
cc_23 VNB N_Y_c_240_n 0.00191689f $X=-0.19 $Y=-0.24 $X2=2.695 $Y2=1.105
cc_24 VNB N_Y_c_241_n 0.00187002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB Y 0.0267466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_Y_c_243_n 0.0132373f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.177
cc_27 VNB N_VGND_c_350_n 0.00571301f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=1.16
cc_28 VNB N_VGND_c_351_n 0.0182484f $X=-0.19 $Y=-0.24 $X2=1.475 $Y2=0.445
cc_29 VNB N_VGND_c_352_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=1.5 $Y2=1.985
cc_30 VNB N_VGND_c_353_n 0.00546241f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.025
cc_31 VNB N_VGND_c_354_n 0.0181341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_355_n 0.00574268f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=1.41
cc_33 VNB N_VGND_c_356_n 0.0184172f $X=-0.19 $Y=-0.24 $X2=2.36 $Y2=1.16
cc_34 VNB N_VGND_c_357_n 0.025462f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.985
cc_35 VNB N_VGND_c_358_n 0.213527f $X=-0.19 $Y=-0.24 $X2=2.94 $Y2=1.985
cc_36 VNB N_VGND_c_359_n 0.00660796f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.217
cc_37 VNB N_VGND_c_360_n 0.00497354f $X=-0.19 $Y=-0.24 $X2=2.56 $Y2=1.16
cc_38 VPB N_A_c_87_n 0.0192616f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.41
cc_39 VPB N_A_c_88_n 0.0161615f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.41
cc_40 VPB N_A_c_89_n 0.0161805f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.41
cc_41 VPB N_A_c_90_n 0.0161805f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.41
cc_42 VPB N_A_c_91_n 0.0161805f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=1.41
cc_43 VPB N_A_c_92_n 0.0193091f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.41
cc_44 VPB N_A_c_80_n 0.00693507f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=1.16
cc_45 VPB N_A_c_82_n 0.00639463f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.217
cc_46 VPB N_A_c_83_n 0.00639603f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.217
cc_47 VPB N_A_c_84_n 0.00639603f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.217
cc_48 VPB N_A_c_85_n 0.00638057f $X=-0.19 $Y=1.305 $X2=2.46 $Y2=1.217
cc_49 VPB N_A_c_86_n 0.00703453f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.16
cc_50 VPB N_VPWR_c_182_n 0.0115225f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=1.025
cc_51 VPB N_VPWR_c_183_n 0.0335458f $X=-0.19 $Y=1.305 $X2=1.475 $Y2=0.445
cc_52 VPB N_VPWR_c_184_n 0.0199672f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.41
cc_53 VPB N_VPWR_c_185_n 0.00522213f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_54 VPB N_VPWR_c_186_n 0.00522213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_187_n 0.0173956f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.985
cc_56 VPB N_VPWR_c_188_n 0.0335277f $X=-0.19 $Y=1.305 $X2=2.36 $Y2=1.16
cc_57 VPB N_VPWR_c_189_n 0.0199672f $X=-0.19 $Y=1.305 $X2=2.435 $Y2=0.445
cc_58 VPB N_VPWR_c_190_n 0.00497514f $X=-0.19 $Y=1.305 $X2=2.435 $Y2=0.445
cc_59 VPB N_VPWR_c_191_n 0.0199228f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.985
cc_60 VPB N_VPWR_c_192_n 0.00497514f $X=-0.19 $Y=1.305 $X2=2.84 $Y2=1.16
cc_61 VPB N_VPWR_c_181_n 0.0488761f $X=-0.19 $Y=1.305 $X2=2.185 $Y2=1.105
cc_62 VPB N_Y_c_233_n 0.00767241f $X=-0.19 $Y=1.305 $X2=1.5 $Y2=1.41
cc_63 VPB N_Y_c_245_n 0.00244569f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_64 VPB N_Y_c_246_n 0.00750725f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.16
cc_65 VPB N_Y_c_247_n 0.00204767f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=1.41
cc_66 VPB N_Y_c_248_n 0.0020177f $X=-0.19 $Y=1.305 $X2=2.94 $Y2=1.41
cc_67 VPB N_Y_c_249_n 0.00336463f $X=-0.19 $Y=1.305 $X2=1.165 $Y2=1.105
cc_68 VPB N_Y_c_250_n 0.00156219f $X=-0.19 $Y=1.305 $X2=2.185 $Y2=1.105
cc_69 VPB N_Y_c_251_n 0.00156219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_252_n 0.00159282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB Y 0.00903212f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_Y_c_254_n 0.0141507f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 N_A_c_87_n N_VPWR_c_183_n 0.00489113f $X=0.54 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_87_n N_VPWR_c_184_n 0.00702461f $X=0.54 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_88_n N_VPWR_c_184_n 0.00702461f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_88_n N_VPWR_c_185_n 0.00303578f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_89_n N_VPWR_c_185_n 0.00303578f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_90_n N_VPWR_c_186_n 0.00303578f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_91_n N_VPWR_c_186_n 0.00303578f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_92_n N_VPWR_c_188_n 0.00492609f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_VPWR_c_189_n 0.00702461f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_90_n N_VPWR_c_189_n 0.00702461f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_91_n N_VPWR_c_191_n 0.00702461f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_92_n N_VPWR_c_191_n 0.00702461f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_c_87_n N_VPWR_c_181_n 0.0134641f $X=0.54 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_88_n N_VPWR_c_181_n 0.0125388f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_89_n N_VPWR_c_181_n 0.0125388f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_90_n N_VPWR_c_181_n 0.0125388f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_c_91_n N_VPWR_c_181_n 0.0125388f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_92_n N_VPWR_c_181_n 0.0135862f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_87_n N_Y_c_233_n 0.00170353f $X=0.54 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_M1001_g N_Y_c_233_n 0.00270363f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_c_80_n N_Y_c_233_n 0.0119622f $X=0.64 $Y=1.16 $X2=0 $Y2=0
cc_94 A N_Y_c_233_n 0.0178211f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_95 N_A_M1001_g N_Y_c_234_n 0.0145702f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_96 N_A_c_80_n N_Y_c_234_n 0.0117529f $X=0.64 $Y=1.16 $X2=0 $Y2=0
cc_97 A N_Y_c_234_n 0.0493103f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_98 N_A_c_87_n N_Y_c_245_n 0.0188912f $X=0.54 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_80_n N_Y_c_245_n 5.58945e-19 $X=0.64 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_c_81_n N_Y_c_245_n 3.02991e-19 $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_101 A N_Y_c_245_n 0.0145864f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A_c_88_n N_Y_c_247_n 0.0175259f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_74_n N_Y_c_247_n 0.00664449f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A_c_89_n N_Y_c_247_n 0.0175259f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_76_n N_Y_c_247_n 3.71188e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_c_82_n N_Y_c_247_n 6.07109e-19 $X=1.02 $Y=1.217 $X2=0 $Y2=0
cc_107 N_A_c_83_n N_Y_c_247_n 6.07109e-19 $X=1.5 $Y=1.217 $X2=0 $Y2=0
cc_108 A N_Y_c_247_n 0.0499117f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_109 N_A_M1001_g N_Y_c_236_n 0.00510542f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_M1002_g N_Y_c_236_n 0.00200232f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_M1002_g N_Y_c_237_n 0.012818f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_c_76_n N_Y_c_237_n 0.00338337f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_M1006_g N_Y_c_237_n 0.012818f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_114 A N_Y_c_237_n 0.0497753f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A_c_76_n N_Y_c_248_n 2.38621e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_90_n N_Y_c_248_n 0.0175259f $X=1.98 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_78_n N_Y_c_248_n 0.00664449f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_c_91_n N_Y_c_248_n 0.0175259f $X=2.46 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_84_n N_Y_c_248_n 6.07109e-19 $X=1.98 $Y=1.217 $X2=0 $Y2=0
cc_120 N_A_c_85_n N_Y_c_248_n 5.70451e-19 $X=2.46 $Y=1.217 $X2=0 $Y2=0
cc_121 A N_Y_c_248_n 0.0495466f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_M1006_g N_Y_c_238_n 0.0050845f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_123 N_A_M1008_g N_Y_c_238_n 0.00198218f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_124 N_A_M1008_g N_Y_c_239_n 0.0145702f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_125 N_A_c_85_n N_Y_c_239_n 0.0136433f $X=2.46 $Y=1.217 $X2=0 $Y2=0
cc_126 A N_Y_c_239_n 0.0405478f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_c_92_n N_Y_c_249_n 0.0203908f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_86_n N_Y_c_249_n 7.78878e-19 $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_129 A N_Y_c_249_n 0.00554358f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A_c_81_n N_Y_c_250_n 0.00574389f $X=0.92 $Y=1.16 $X2=0 $Y2=0
cc_131 A N_Y_c_250_n 0.0209566f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_c_74_n N_Y_c_240_n 0.00350792f $X=1.4 $Y=1.16 $X2=0 $Y2=0
cc_133 A N_Y_c_240_n 0.0211887f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_76_n N_Y_c_251_n 0.00625592f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_135 A N_Y_c_251_n 0.0209566f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_c_78_n N_Y_c_241_n 0.00350792f $X=2.36 $Y=1.16 $X2=0 $Y2=0
cc_137 A N_Y_c_241_n 0.0207812f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_c_86_n N_Y_c_252_n 0.00585652f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_139 A N_Y_c_252_n 0.0213675f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A_c_92_n Y 0.00169878f $X=2.94 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_86_n Y 0.012036f $X=2.84 $Y=1.16 $X2=0 $Y2=0
cc_142 A Y 0.0105775f $X=2.695 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_M1001_g N_VGND_c_350_n 0.00492552f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_144 N_A_M1001_g N_VGND_c_351_n 0.00437852f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_145 N_A_M1002_g N_VGND_c_351_n 0.00437852f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_M1002_g N_VGND_c_352_n 0.00480861f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_M1006_g N_VGND_c_352_n 0.00313102f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_148 N_A_M1008_g N_VGND_c_353_n 0.0045088f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_149 N_A_M1006_g N_VGND_c_354_n 0.00437852f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_M1008_g N_VGND_c_354_n 0.00437852f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_151 N_A_M1001_g N_VGND_c_358_n 0.0073136f $X=0.995 $Y=0.445 $X2=0 $Y2=0
cc_152 N_A_M1002_g N_VGND_c_358_n 0.00626392f $X=1.475 $Y=0.445 $X2=0 $Y2=0
cc_153 N_A_M1006_g N_VGND_c_358_n 0.00613846f $X=1.955 $Y=0.445 $X2=0 $Y2=0
cc_154 N_A_M1008_g N_VGND_c_358_n 0.00742651f $X=2.435 $Y=0.445 $X2=0 $Y2=0
cc_155 N_VPWR_c_181_n N_Y_M1000_s 0.00405474f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_181_n N_Y_M1004_s 0.00405474f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_181_n N_Y_M1007_s 0.00388144f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_M1000_d N_Y_c_245_n 0.00124373f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_159 N_VPWR_c_183_n N_Y_c_245_n 0.00956383f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_160 N_VPWR_M1000_d N_Y_c_246_n 0.00263276f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_161 N_VPWR_c_183_n N_Y_c_246_n 0.0153867f $X=0.3 $Y=1.965 $X2=0 $Y2=0
cc_162 N_VPWR_c_184_n N_Y_c_314_n 0.0129843f $X=1.13 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_181_n N_Y_c_314_n 0.00960102f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_M1003_d N_Y_c_247_n 0.00197722f $X=1.11 $Y=1.485 $X2=0 $Y2=0
cc_165 N_VPWR_c_185_n N_Y_c_247_n 0.0151327f $X=1.26 $Y=1.965 $X2=0 $Y2=0
cc_166 N_VPWR_c_189_n N_Y_c_318_n 0.0129843f $X=2.09 $Y=2.72 $X2=0 $Y2=0
cc_167 N_VPWR_c_181_n N_Y_c_318_n 0.00960102f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_168 N_VPWR_M1005_d N_Y_c_248_n 0.00197722f $X=2.07 $Y=1.485 $X2=0 $Y2=0
cc_169 N_VPWR_c_186_n N_Y_c_248_n 0.0151327f $X=2.22 $Y=1.965 $X2=0 $Y2=0
cc_170 N_VPWR_c_191_n N_Y_c_322_n 0.0131352f $X=3.05 $Y=2.72 $X2=0 $Y2=0
cc_171 N_VPWR_c_181_n N_Y_c_322_n 0.00979076f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_172 N_VPWR_M1009_d N_Y_c_249_n 0.00240495f $X=3.03 $Y=1.485 $X2=0 $Y2=0
cc_173 N_VPWR_c_188_n N_Y_c_249_n 0.0148521f $X=3.18 $Y=1.965 $X2=0 $Y2=0
cc_174 N_VPWR_M1009_d N_Y_c_254_n 0.00219558f $X=3.03 $Y=1.485 $X2=0 $Y2=0
cc_175 N_VPWR_c_188_n N_Y_c_254_n 0.0149598f $X=3.18 $Y=1.965 $X2=0 $Y2=0
cc_176 N_Y_c_234_n N_VGND_c_350_n 0.0252244f $X=1.13 $Y=0.81 $X2=0 $Y2=0
cc_177 N_Y_c_234_n N_VGND_c_351_n 0.00305995f $X=1.13 $Y=0.81 $X2=0 $Y2=0
cc_178 N_Y_c_236_n N_VGND_c_351_n 0.0141727f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_179 N_Y_c_237_n N_VGND_c_351_n 0.00305995f $X=2.09 $Y=0.81 $X2=0 $Y2=0
cc_180 N_Y_c_237_n N_VGND_c_352_n 0.0184664f $X=2.09 $Y=0.81 $X2=0 $Y2=0
cc_181 N_Y_c_239_n N_VGND_c_353_n 0.0236483f $X=3.27 $Y=0.81 $X2=0 $Y2=0
cc_182 N_Y_c_237_n N_VGND_c_354_n 0.00305995f $X=2.09 $Y=0.81 $X2=0 $Y2=0
cc_183 N_Y_c_238_n N_VGND_c_354_n 0.0140179f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_184 N_Y_c_239_n N_VGND_c_354_n 0.00305995f $X=3.27 $Y=0.81 $X2=0 $Y2=0
cc_185 N_Y_c_234_n N_VGND_c_356_n 0.00440462f $X=1.13 $Y=0.81 $X2=0 $Y2=0
cc_186 N_Y_c_235_n N_VGND_c_356_n 0.00289403f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_187 N_Y_c_239_n N_VGND_c_357_n 0.00615732f $X=3.27 $Y=0.81 $X2=0 $Y2=0
cc_188 N_Y_c_243_n N_VGND_c_357_n 0.00510712f $X=3.42 $Y=0.895 $X2=0 $Y2=0
cc_189 N_Y_M1001_d N_VGND_c_358_n 0.00299282f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_190 N_Y_M1006_d N_VGND_c_358_n 0.00301747f $X=2.03 $Y=0.235 $X2=0 $Y2=0
cc_191 N_Y_c_234_n N_VGND_c_358_n 0.0140191f $X=1.13 $Y=0.81 $X2=0 $Y2=0
cc_192 N_Y_c_235_n N_VGND_c_358_n 0.00478629f $X=0.275 $Y=0.81 $X2=0 $Y2=0
cc_193 N_Y_c_236_n N_VGND_c_358_n 0.00978777f $X=1.26 $Y=0.445 $X2=0 $Y2=0
cc_194 N_Y_c_237_n N_VGND_c_358_n 0.0110611f $X=2.09 $Y=0.81 $X2=0 $Y2=0
cc_195 N_Y_c_238_n N_VGND_c_358_n 0.00959809f $X=2.22 $Y=0.445 $X2=0 $Y2=0
cc_196 N_Y_c_239_n N_VGND_c_358_n 0.0168867f $X=3.27 $Y=0.81 $X2=0 $Y2=0
cc_197 N_Y_c_243_n N_VGND_c_358_n 0.0084464f $X=3.42 $Y=0.895 $X2=0 $Y2=0
