* NGSPICE file created from sky130_fd_sc_hdll__fill_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__fill_1 VGND VNB VPB VPWR
.ends

