* File: sky130_fd_sc_hdll__sdfxbp_1.pex.spice
* Created: Wed Sep  2 08:52:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%CLK 1 2 3 5 6 8 13
c40 1 0 2.71124e-20 $X=0.31 $Y=1.325
r41 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r42 6 16 86.4067 $w=2.69e-07 $l=5.05816e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.355 $Y2=1.16
r43 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r44 3 9 94.8617 $w=1.5e-07 $l=1.85e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.31 $Y2=1.665
r45 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r46 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r47 1 16 38.9235 $w=2.69e-07 $l=1.86145e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.355 $Y2=1.16
r48 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_27_47# 1 2 8 9 11 14 18 20 21 23 24 26
+ 28 29 31 32 36 40 44 45 46 50 51 53 56 57 58 59 60 61 68 70 76 81 85
c244 85 0 5.22246e-20 $X=7.2 $Y=1.41
c245 68 0 1.55016e-19 $X=5.7 $Y=1.87
c246 61 0 1.98979e-19 $X=5.845 $Y=1.87
c247 53 0 1.8505e-19 $X=0.81 $Y=1.235
c248 51 0 1.77499e-19 $X=0.78 $Y=1.795
c249 46 0 1.03679e-19 $X=0.665 $Y=1.88
r250 84 86 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.225 $Y=1.41
+ $X2=7.225 $Y2=1.575
r251 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.2
+ $Y=1.41 $X2=7.2 $Y2=1.41
r252 81 84 16.2293 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=7.225 $Y=1.32
+ $X2=7.225 $Y2=1.41
r253 79 80 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.5
+ $Y=1.74 $X2=5.5 $Y2=1.74
r254 75 76 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r255 71 85 22.0885 $w=2.38e-07 $l=4.6e-07 $layer=LI1_cond $X=7.235 $Y=1.87
+ $X2=7.235 $Y2=1.41
r256 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.26 $Y=1.87
+ $X2=7.26 $Y2=1.87
r257 68 80 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=5.7 $Y=1.832 $X2=5.5
+ $Y2=1.832
r258 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.7 $Y=1.87 $X2=5.7
+ $Y2=1.87
r259 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.78 $Y=1.87
+ $X2=0.78 $Y2=1.87
r260 61 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.845 $Y=1.87
+ $X2=5.7 $Y2=1.87
r261 60 70 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.115 $Y=1.87
+ $X2=7.26 $Y2=1.87
r262 60 61 1.57178 $w=1.4e-07 $l=1.27e-06 $layer=MET1_cond $X=7.115 $Y=1.87
+ $X2=5.845 $Y2=1.87
r263 59 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.925 $Y=1.87
+ $X2=0.78 $Y2=1.87
r264 58 67 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.555 $Y=1.87
+ $X2=5.7 $Y2=1.87
r265 58 59 5.73019 $w=1.4e-07 $l=4.63e-06 $layer=MET1_cond $X=5.555 $Y=1.87
+ $X2=0.925 $Y2=1.87
r266 54 75 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.965 $Y2=1.235
r267 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r268 51 64 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.88
r269 51 53 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.235
r270 50 57 6.0623 $w=2.28e-07 $l=1.15e-07 $layer=LI1_cond $X=0.78 $Y=1.085
+ $X2=0.78 $Y2=0.97
r271 50 53 7.51593 $w=2.28e-07 $l=1.5e-07 $layer=LI1_cond $X=0.78 $Y=1.085
+ $X2=0.78 $Y2=1.235
r272 48 57 9.38461 $w=1.93e-07 $l=1.65e-07 $layer=LI1_cond $X=0.762 $Y=0.805
+ $X2=0.762 $Y2=0.97
r273 47 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r274 46 64 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.78 $Y2=1.88
r275 46 47 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.345 $Y2=1.88
r276 44 48 6.85817 $w=1.7e-07 $l=1.32868e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.762 $Y2=0.805
r277 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.345 $Y2=0.72
r278 38 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r279 38 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r280 34 36 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=8 $Y=1.245 $X2=8
+ $Y2=0.415
r281 33 81 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.385 $Y=1.32
+ $X2=7.225 $Y2=1.32
r282 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.925 $Y=1.32
+ $X2=8 $Y2=1.245
r283 32 33 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.925 $Y=1.32
+ $X2=7.385 $Y2=1.32
r284 29 31 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.23 $Y=1.99
+ $X2=7.23 $Y2=2.275
r285 28 29 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.23 $Y=1.89 $X2=7.23
+ $Y2=1.99
r286 28 86 104.447 $w=2e-07 $l=3.15e-07 $layer=POLY_cond $X=7.23 $Y=1.89
+ $X2=7.23 $Y2=1.575
r287 24 79 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.465 $Y=1.99
+ $X2=5.525 $Y2=1.74
r288 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.465 $Y=1.99
+ $X2=5.465 $Y2=2.275
r289 23 79 31.9848 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.465 $Y=1.575
+ $X2=5.525 $Y2=1.74
r290 22 23 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=5.465 $Y=1.395
+ $X2=5.465 $Y2=1.575
r291 20 22 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=5.365 $Y=1.32
+ $X2=5.465 $Y2=1.395
r292 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.365 $Y=1.32
+ $X2=5.005 $Y2=1.32
r293 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.93 $Y=1.245
+ $X2=5.005 $Y2=1.32
r294 16 18 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.93 $Y=1.245
+ $X2=4.93 $Y2=0.415
r295 12 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r296 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r297 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r298 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r299 7 75 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r300 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r301 2 56 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r302 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_319_47# 1 2 9 11 13 15 18 20 23 24 26
+ 29 32 36 38 39 41 47
c120 41 0 1.77453e-19 $X=3.42 $Y=1.52
c121 23 0 1.68628e-19 $X=2.335 $Y=1.86
r122 41 44 8.82014 $w=2.18e-07 $l=1.65e-07 $layer=LI1_cond $X=3.445 $Y=1.52
+ $X2=3.445 $Y2=1.685
r123 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=1.52 $X2=3.42 $Y2=1.52
r124 33 36 7.88038 $w=1.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.605 $Y=0.35
+ $X2=1.74 $Y2=0.35
r125 32 44 9.95338 $w=1.93e-07 $l=1.75e-07 $layer=LI1_cond $X=3.432 $Y=1.86
+ $X2=3.432 $Y2=1.685
r126 30 39 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.42 $Y=1.967
+ $X2=2.335 $Y2=1.967
r127 29 32 6.83761 $w=2.15e-07 $l=1.47743e-07 $layer=LI1_cond $X=3.335 $Y=1.967
+ $X2=3.432 $Y2=1.86
r128 29 30 49.0458 $w=2.13e-07 $l=9.15e-07 $layer=LI1_cond $X=3.335 $Y=1.967
+ $X2=2.42 $Y2=1.967
r129 27 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=2.48 $Y=1.04 $X2=2.57
+ $Y2=1.04
r130 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.48
+ $Y=1.04 $X2=2.48 $Y2=1.04
r131 24 26 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=2.42 $Y=1.04 $X2=2.48
+ $Y2=1.04
r132 23 39 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.335 $Y=1.86
+ $X2=2.335 $Y2=1.967
r133 22 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.335 $Y=1.125
+ $X2=2.42 $Y2=1.04
r134 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.335 $Y=1.125
+ $X2=2.335 $Y2=1.86
r135 21 38 1.54683 $w=2.15e-07 $l=1.43e-07 $layer=LI1_cond $X=1.805 $Y=1.967
+ $X2=1.662 $Y2=1.967
r136 20 39 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=1.967
+ $X2=2.335 $Y2=1.967
r137 20 21 23.8529 $w=2.13e-07 $l=4.45e-07 $layer=LI1_cond $X=2.25 $Y=1.967
+ $X2=1.805 $Y2=1.967
r138 16 38 4.92743 $w=2.27e-07 $l=1.08e-07 $layer=LI1_cond $X=1.662 $Y=2.075
+ $X2=1.662 $Y2=1.967
r139 16 18 4.04366 $w=2.83e-07 $l=1e-07 $layer=LI1_cond $X=1.662 $Y=2.075
+ $X2=1.662 $Y2=2.175
r140 15 38 4.92743 $w=2.27e-07 $l=1.32469e-07 $layer=LI1_cond $X=1.605 $Y=1.86
+ $X2=1.662 $Y2=1.967
r141 14 33 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=0.35
r142 14 15 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.605 $Y=0.445
+ $X2=1.605 $Y2=1.86
r143 11 42 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.4 $Y=1.77
+ $X2=3.445 $Y2=1.52
r144 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.4 $Y=1.77
+ $X2=3.4 $Y2=2.165
r145 7 47 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.57 $Y=0.905
+ $X2=2.57 $Y2=1.04
r146 7 9 235.872 $w=1.5e-07 $l=4.6e-07 $layer=POLY_cond $X=2.57 $Y=0.905
+ $X2=2.57 $Y2=0.445
r147 2 18 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=2.175
r148 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.74 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%SCE 1 3 6 8 10 12 15 17 21 24 25 26 35 37
+ 39
c103 37 0 1.62494e-19 $X=3.425 $Y=0.785
r104 37 39 3.40495 $w=2.18e-07 $l=6.5e-08 $layer=LI1_cond $X=3.425 $Y=0.785
+ $X2=3.425 $Y2=0.85
r105 32 35 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.4 $Y=0.95
+ $X2=3.51 $Y2=0.95
r106 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.4
+ $Y=0.95 $X2=3.4 $Y2=0.95
r107 26 37 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.425 $Y=0.7
+ $X2=3.425 $Y2=0.785
r108 26 33 4.71454 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=3.425 $Y=0.86
+ $X2=3.425 $Y2=0.95
r109 26 39 0.523838 $w=2.18e-07 $l=1e-08 $layer=LI1_cond $X=3.425 $Y=0.86
+ $X2=3.425 $Y2=0.85
r110 24 26 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.315 $Y=0.7
+ $X2=3.425 $Y2=0.7
r111 24 25 83.8342 $w=1.68e-07 $l=1.285e-06 $layer=LI1_cond $X=3.315 $Y=0.7
+ $X2=2.03 $Y2=0.7
r112 22 30 8.87117 $w=3.26e-07 $l=6e-08 $layer=POLY_cond $X=1.97 $Y=1.52
+ $X2=1.97 $Y2=1.58
r113 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.945
+ $Y=1.52 $X2=1.945 $Y2=1.52
r114 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.945 $Y=0.785
+ $X2=2.03 $Y2=0.7
r115 19 21 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.945 $Y=0.785
+ $X2=1.945 $Y2=1.52
r116 13 35 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.51 $Y=0.785
+ $X2=3.51 $Y2=0.95
r117 13 15 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.51 $Y=0.785
+ $X2=3.51 $Y2=0.445
r118 10 17 63.8074 $w=2e-07 $l=1.9e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=1.58
r119 10 12 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r120 9 30 20.933 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=2.16 $Y=1.58 $X2=1.97
+ $Y2=1.58
r121 8 17 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=2.325 $Y=1.58
+ $X2=2.425 $Y2=1.58
r122 8 9 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.325 $Y=1.58
+ $X2=2.16 $Y2=1.58
r123 4 22 34.1407 $w=3.26e-07 $l=1.39911e-07 $layer=POLY_cond $X=1.98 $Y=1.385
+ $X2=1.97 $Y2=1.52
r124 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.98 $Y=1.385 $X2=1.98
+ $Y2=0.445
r125 1 30 37.6865 $w=3.26e-07 $l=1.97358e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.97 $Y2=1.58
r126 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%D 1 3 6 8 16
r37 8 16 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.89 $Y=1.52
+ $X2=2.975 $Y2=1.52
r38 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.89
+ $Y=1.52 $X2=2.89 $Y2=1.52
r39 4 11 38.578 $w=2.95e-07 $l=1.94808e-07 $layer=POLY_cond $X=2.98 $Y=1.355
+ $X2=2.915 $Y2=1.52
r40 4 6 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=2.98 $Y=1.355 $X2=2.98
+ $Y2=0.445
r41 1 11 48.1208 $w=2.95e-07 $l=2.57391e-07 $layer=POLY_cond $X=2.93 $Y=1.77
+ $X2=2.915 $Y2=1.52
r42 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.93 $Y=1.77 $X2=2.93
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%SCD 3 6 7 9 10 13
c50 3 0 1.62494e-19 $X=3.89 $Y=0.445
r51 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.355
+ $X2=3.975 $Y2=1.52
r52 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.975 $Y=1.355
+ $X2=3.975 $Y2=1.19
r53 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.95
+ $Y=1.355 $X2=3.95 $Y2=1.355
r54 10 14 3.72364 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.08 $Y=1.19
+ $X2=4.08 $Y2=1.355
r55 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.915 $Y=1.77
+ $X2=3.915 $Y2=2.165
r56 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.915 $Y=1.67 $X2=3.915
+ $Y2=1.77
r57 6 16 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.915 $Y=1.67 $X2=3.915
+ $Y2=1.52
r58 3 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.89 $Y=0.445
+ $X2=3.89 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_211_363# 1 2 7 9 10 12 13 15 16 18 21
+ 25 26 30 33 34 36 37 38 41 47 49 57 62
c205 37 0 5.22246e-20 $X=7.125 $Y=0.85
c206 36 0 1.41526e-19 $X=5.215 $Y=0.735
c207 21 0 1.98979e-19 $X=4.94 $Y=1.74
r208 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.48
+ $Y=0.87 $X2=7.48 $Y2=0.87
r209 59 62 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.335 $Y=0.87
+ $X2=7.48 $Y2=0.87
r210 54 57 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.4 $Y=0.87
+ $X2=5.51 $Y2=0.87
r211 50 63 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=7.27 $Y=0.87
+ $X2=7.48 $Y2=0.87
r212 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.27 $Y=0.85
+ $X2=7.27 $Y2=0.85
r213 47 75 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=5.29 $Y=0.87 $X2=5
+ $Y2=0.87
r214 47 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.4
+ $Y=0.87 $X2=5.4 $Y2=0.87
r215 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0.85
+ $X2=5.29 $Y2=0.85
r216 43 46 0.0481203 $w=2.3e-07 $l=7.5e-08 $layer=MET1_cond $X=5.215 $Y=0.85
+ $X2=5.29 $Y2=0.85
r217 41 70 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=1.2 $Y=0.51
+ $X2=1.2 $Y2=1.96
r218 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=0.51 $X2=1.2
+ $Y2=0.51
r219 38 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=0.85
+ $X2=5.29 $Y2=0.85
r220 37 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.125 $Y=0.85
+ $X2=7.27 $Y2=0.85
r221 37 38 2.09158 $w=1.4e-07 $l=1.69e-06 $layer=MET1_cond $X=7.125 $Y=0.85
+ $X2=5.435 $Y2=0.85
r222 36 43 0.0373109 $w=1.4e-07 $l=1.15e-07 $layer=MET1_cond $X=5.215 $Y=0.735
+ $X2=5.215 $Y2=0.85
r223 35 36 0.191831 $w=1.4e-07 $l=1.55e-07 $layer=MET1_cond $X=5.215 $Y=0.58
+ $X2=5.215 $Y2=0.735
r224 34 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=0.51
+ $X2=1.2 $Y2=0.51
r225 33 35 0.0698411 $w=1.4e-07 $l=9.89949e-08 $layer=MET1_cond $X=5.145 $Y=0.51
+ $X2=5.215 $Y2=0.58
r226 33 34 4.70296 $w=1.4e-07 $l=3.8e-06 $layer=MET1_cond $X=5.145 $Y=0.51
+ $X2=1.345 $Y2=0.51
r227 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.76
+ $Y=1.74 $X2=7.76 $Y2=1.74
r228 27 30 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.62 $Y=1.74
+ $X2=7.76 $Y2=1.74
r229 26 63 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.525 $Y=0.87
+ $X2=7.48 $Y2=0.87
r230 25 27 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.62 $Y=1.575
+ $X2=7.62 $Y2=1.74
r231 24 26 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.62 $Y=1.035
+ $X2=7.525 $Y2=0.87
r232 24 25 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.62 $Y=1.035
+ $X2=7.62 $Y2=1.575
r233 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.94
+ $Y=1.74 $X2=4.94 $Y2=1.74
r234 19 75 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5 $Y=1.035 $X2=5
+ $Y2=0.87
r235 19 21 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5 $Y=1.035 $X2=5
+ $Y2=1.74
r236 16 31 46.5577 $w=3.26e-07 $l=2.89396e-07 $layer=POLY_cond $X=7.7 $Y=1.99
+ $X2=7.785 $Y2=1.74
r237 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.7 $Y=1.99
+ $X2=7.7 $Y2=2.275
r238 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.335 $Y=0.705
+ $X2=7.335 $Y2=0.87
r239 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.335 $Y=0.705
+ $X2=7.335 $Y2=0.415
r240 10 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.51 $Y=0.705
+ $X2=5.51 $Y2=0.87
r241 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.51 $Y=0.705
+ $X2=5.51 $Y2=0.415
r242 7 22 46.5577 $w=3.26e-07 $l=2.57391e-07 $layer=POLY_cond $X=4.95 $Y=1.99
+ $X2=4.965 $Y2=1.74
r243 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.95 $Y=1.99
+ $X2=4.95 $Y2=2.275
r244 2 70 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r245 1 41 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_1179_183# 1 2 8 9 11 14 16 19 22 24 30
+ 31 33 34 37
c100 37 0 1.19883e-19 $X=6 $Y=0.93
c101 9 0 1.55016e-19 $X=5.995 $Y=1.99
r102 36 37 0.919847 $w=2.62e-07 $l=5e-09 $layer=POLY_cond $X=5.995 $Y=0.93 $X2=6
+ $Y2=0.93
r103 33 34 7.18001 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=2.3
+ $X2=6.875 $Y2=2.135
r104 28 37 33.1145 $w=2.62e-07 $l=1.8e-07 $layer=POLY_cond $X=6.18 $Y=0.93 $X2=6
+ $Y2=0.93
r105 27 30 3.0866 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=0.93
+ $X2=6.265 $Y2=0.93
r106 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.18
+ $Y=0.93 $X2=6.18 $Y2=0.93
r107 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.945 $Y=0.45
+ $X2=7.07 $Y2=0.45
r108 20 31 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=1.065
+ $X2=6.835 $Y2=0.915
r109 20 34 56.0506 $w=2.18e-07 $l=1.07e-06 $layer=LI1_cond $X=6.835 $Y=1.065
+ $X2=6.835 $Y2=2.135
r110 19 31 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=0.765
+ $X2=6.835 $Y2=0.915
r111 18 22 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.835 $Y=0.535
+ $X2=6.945 $Y2=0.45
r112 18 19 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=6.835 $Y=0.535
+ $X2=6.835 $Y2=0.765
r113 16 31 0.253446 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.725 $Y=0.915
+ $X2=6.835 $Y2=0.915
r114 16 30 17.6708 $w=2.98e-07 $l=4.6e-07 $layer=LI1_cond $X=6.725 $Y=0.915
+ $X2=6.265 $Y2=0.915
r115 12 37 15.8058 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6 $Y=0.795 $X2=6
+ $Y2=0.93
r116 12 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6 $Y=0.795 $X2=6
+ $Y2=0.445
r117 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.995 $Y=1.99
+ $X2=5.995 $Y2=2.275
r118 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.995 $Y=1.89 $X2=5.995
+ $Y2=1.99
r119 7 36 9.16944 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=5.995 $Y=1.065
+ $X2=5.995 $Y2=0.93
r120 7 8 273.551 $w=2e-07 $l=8.25e-07 $layer=POLY_cond $X=5.995 $Y=1.065
+ $X2=5.995 $Y2=1.89
r121 2 33 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.735 $X2=6.94 $Y2=2.3
r122 1 24 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.905
+ $Y=0.235 $X2=7.07 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_1001_47# 1 2 8 9 11 14 15 16 17 18 19
+ 23 28 30 32
c116 28 0 2.90402e-19 $X=5.79 $Y=1.315
r117 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.47
+ $Y=1.41 $X2=6.47 $Y2=1.41
r118 32 34 18.3251 $w=2.43e-07 $l=3.65e-07 $layer=LI1_cond $X=6.105 $Y=1.41
+ $X2=6.47 $Y2=1.41
r119 29 32 1.31576 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.105 $Y=1.575
+ $X2=6.105 $Y2=1.41
r120 29 30 32.216 $w=2.18e-07 $l=6.15e-07 $layer=LI1_cond $X=6.105 $Y=1.575
+ $X2=6.105 $Y2=2.19
r121 28 32 15.8148 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=5.79 $Y=1.41
+ $X2=6.105 $Y2=1.41
r122 27 28 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=5.79 $Y=0.535
+ $X2=5.79 $Y2=1.315
r123 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.705 $Y=0.45
+ $X2=5.79 $Y2=0.535
r124 23 25 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.705 $Y=0.45
+ $X2=5.25 $Y2=0.45
r125 19 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=5.995 $Y=2.275
+ $X2=6.105 $Y2=2.19
r126 19 21 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=5.995 $Y=2.275
+ $X2=5.21 $Y2=2.275
r127 17 35 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.47 $Y2=1.41
r128 17 18 0.448535 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.705 $Y2=1.467
r129 15 16 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.755 $Y=0.95
+ $X2=6.755 $Y2=1.1
r130 14 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.83 $Y=0.555
+ $X2=6.83 $Y2=0.95
r131 9 18 27.0491 $w=1.9e-07 $l=1.93e-07 $layer=POLY_cond $X=6.705 $Y=1.66
+ $X2=6.705 $Y2=1.467
r132 9 11 120.5 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.705 $Y=1.66
+ $X2=6.705 $Y2=2.11
r133 8 18 27.0491 $w=1.9e-07 $l=1.92e-07 $layer=POLY_cond $X=6.705 $Y=1.275
+ $X2=6.705 $Y2=1.467
r134 8 16 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=6.705 $Y=1.275
+ $X2=6.705 $Y2=1.1
r135 2 21 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=5.04
+ $Y=2.065 $X2=5.21 $Y2=2.275
r136 1 25 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=5.005
+ $Y=0.235 $X2=5.25 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_1653_315# 1 2 7 9 12 14 16 17 19 20 22
+ 23 24 26 27 29 31 38 42 45 47 50 51 53 54 55
c115 51 0 3.89057e-19 $X=9.915 $Y=1.16
r116 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.915
+ $Y=1.16 $X2=9.915 $Y2=1.16
r117 48 55 0.63164 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=9.4 $Y=1.16
+ $X2=9.307 $Y2=1.16
r118 48 50 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=9.4 $Y=1.16
+ $X2=9.915 $Y2=1.16
r119 47 54 6.72893 $w=2.37e-07 $l=1.89222e-07 $layer=LI1_cond $X=9.307 $Y=1.575
+ $X2=9.255 $Y2=1.74
r120 46 55 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=9.307 $Y=1.325
+ $X2=9.307 $Y2=1.16
r121 46 47 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=9.307 $Y=1.325
+ $X2=9.307 $Y2=1.575
r122 45 55 8.10876 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=9.307 $Y=0.995
+ $X2=9.307 $Y2=1.16
r123 45 53 10.1916 $w=1.83e-07 $l=1.7e-07 $layer=LI1_cond $X=9.307 $Y=0.995
+ $X2=9.307 $Y2=0.825
r124 40 54 6.72893 $w=2.37e-07 $l=1.65e-07 $layer=LI1_cond $X=9.255 $Y=1.905
+ $X2=9.255 $Y2=1.74
r125 40 42 1.78827 $w=2.88e-07 $l=4.5e-08 $layer=LI1_cond $X=9.255 $Y=1.905
+ $X2=9.255 $Y2=1.95
r126 36 53 7.96936 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=9.235 $Y=0.66
+ $X2=9.235 $Y2=0.825
r127 36 38 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=9.235 $Y=0.66
+ $X2=9.235 $Y2=0.385
r128 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.57
+ $Y=1.74 $X2=8.57 $Y2=1.74
r129 31 54 0.189605 $w=3.3e-07 $l=1.45e-07 $layer=LI1_cond $X=9.11 $Y=1.74
+ $X2=9.255 $Y2=1.74
r130 31 33 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.11 $Y=1.74
+ $X2=8.57 $Y2=1.74
r131 27 29 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=10.955 $Y=0.73
+ $X2=10.955 $Y2=0.445
r132 24 26 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=10.93 $Y=1.77
+ $X2=10.93 $Y2=2.165
r133 23 24 52.9784 $w=2.32e-07 $l=2.92276e-07 $layer=POLY_cond $X=10.85 $Y=1.515
+ $X2=10.93 $Y2=1.77
r134 22 23 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=10.85 $Y=1.325
+ $X2=10.85 $Y2=1.515
r135 21 51 3.90195 $w=3.3e-07 $l=3.32415e-07 $layer=POLY_cond $X=10.04 $Y=1.16
+ $X2=9.78 $Y2=0.995
r136 20 22 46.3768 $w=1.76e-07 $l=1.89222e-07 $layer=POLY_cond $X=10.902 $Y=1.16
+ $X2=10.85 $Y2=1.325
r137 20 27 118.951 $w=1.76e-07 $l=4.5573e-07 $layer=POLY_cond $X=10.902 $Y=1.16
+ $X2=10.955 $Y2=0.73
r138 20 21 128.523 $w=3.3e-07 $l=7.35e-07 $layer=POLY_cond $X=10.775 $Y=1.16
+ $X2=10.04 $Y2=1.16
r139 17 51 34.7346 $w=1.65e-07 $l=1.85e-07 $layer=POLY_cond $X=9.965 $Y=0.995
+ $X2=9.78 $Y2=0.995
r140 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.965 $Y=0.995
+ $X2=9.965 $Y2=0.56
r141 14 51 34.7346 $w=1.65e-07 $l=4.88493e-07 $layer=POLY_cond $X=9.94 $Y=1.41
+ $X2=9.78 $Y2=0.995
r142 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.94 $Y=1.41
+ $X2=9.94 $Y2=1.985
r143 10 34 39.3952 $w=3.9e-07 $l=1.74714e-07 $layer=POLY_cond $X=8.505 $Y=1.575
+ $X2=8.485 $Y2=1.74
r144 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=8.505 $Y=1.575
+ $X2=8.505 $Y2=0.445
r145 7 34 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=8.365 $Y=1.99
+ $X2=8.485 $Y2=1.74
r146 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.365 $Y=1.99
+ $X2=8.365 $Y2=2.275
r147 2 42 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=9.11
+ $Y=1.485 $X2=9.235 $Y2=1.95
r148 1 38 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=9.11
+ $Y=0.235 $X2=9.235 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_1464_413# 1 2 7 9 10 12 13 14 15 19 26
+ 29 32 33
c85 14 0 1.12604e-19 $X=9.47 $Y=1.202
r86 32 34 11.1226 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=8.11 $Y=1.16
+ $X2=8.11 $Y2=1.405
r87 32 33 7.01492 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.11 $Y=1.16
+ $X2=8.11 $Y2=0.995
r88 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.96
+ $Y=1.16 $X2=8.96 $Y2=1.16
r89 27 32 1.07274 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=8.285 $Y=1.16
+ $X2=8.11 $Y2=1.16
r90 27 29 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.285 $Y=1.16
+ $X2=8.96 $Y2=1.16
r91 26 34 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.2 $Y=2.165 $X2=8.2
+ $Y2=1.405
r92 23 33 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=8.045 $Y=0.535
+ $X2=8.045 $Y2=0.995
r93 19 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.935 $Y=0.45
+ $X2=8.045 $Y2=0.535
r94 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.935 $Y=0.45
+ $X2=7.68 $Y2=0.45
r95 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.115 $Y=2.25
+ $X2=8.2 $Y2=2.165
r96 15 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.115 $Y=2.25
+ $X2=7.465 $Y2=2.25
r97 13 30 71.6931 $w=3.3e-07 $l=4.1e-07 $layer=POLY_cond $X=9.37 $Y=1.16
+ $X2=8.96 $Y2=1.16
r98 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=9.37 $Y=1.16
+ $X2=9.47 $Y2=1.202
r99 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=9.495 $Y=0.995
+ $X2=9.47 $Y2=1.202
r100 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.495 $Y=0.995
+ $X2=9.495 $Y2=0.56
r101 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=9.47 $Y=1.41
+ $X2=9.47 $Y2=1.202
r102 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.47 $Y=1.41
+ $X2=9.47 $Y2=1.985
r103 2 17 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.32
+ $Y=2.065 $X2=7.465 $Y2=2.25
r104 1 21 182 $w=1.7e-07 $l=3.6187e-07 $layer=licon1_NDIFF $count=1 $X=7.41
+ $Y=0.235 $X2=7.68 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_2114_47# 1 2 7 9 10 12 15 19 23 26
r44 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.355
+ $Y=1.16 $X2=11.355 $Y2=1.16
r45 21 26 0.364692 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=10.86 $Y=1.16
+ $X2=10.735 $Y2=1.16
r46 21 23 17.2866 $w=3.28e-07 $l=4.95e-07 $layer=LI1_cond $X=10.86 $Y=1.16
+ $X2=11.355 $Y2=1.16
r47 17 26 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.735 $Y=1.325
+ $X2=10.735 $Y2=1.16
r48 17 19 37.5696 $w=2.48e-07 $l=8.15e-07 $layer=LI1_cond $X=10.735 $Y=1.325
+ $X2=10.735 $Y2=2.14
r49 13 26 6.46576 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=10.735 $Y=0.995
+ $X2=10.735 $Y2=1.16
r50 13 15 22.3574 $w=2.48e-07 $l=4.85e-07 $layer=LI1_cond $X=10.735 $Y=0.995
+ $X2=10.735 $Y2=0.51
r51 10 24 38.5363 $w=3.15e-07 $l=2.08315e-07 $layer=POLY_cond $X=11.49 $Y=0.995
+ $X2=11.392 $Y2=1.16
r52 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.49 $Y=0.995
+ $X2=11.49 $Y2=0.56
r53 7 24 47.0331 $w=3.15e-07 $l=2.84165e-07 $layer=POLY_cond $X=11.465 $Y=1.41
+ $X2=11.392 $Y2=1.16
r54 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.465 $Y=1.41
+ $X2=11.465 $Y2=1.985
r55 2 19 600 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_PDIFF $count=1 $X=10.57
+ $Y=1.845 $X2=10.695 $Y2=2.14
r56 1 15 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=10.57
+ $Y=0.235 $X2=10.695 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 48
+ 53 54 56 57 59 60 62 63 64 66 71 98 107 108 111 114 117
c177 108 0 1.77499e-19 $X=11.73 $Y=2.72
c178 44 0 1.94529e-19 $X=9.705 $Y=1.79
c179 2 0 1.68628e-19 $X=2.045 $Y=1.845
c180 1 0 1.03679e-19 $X=0.585 $Y=1.815
r181 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r182 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r183 111 112 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r184 108 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r185 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r186 105 117 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=11.395 $Y=2.72
+ $X2=11.242 $Y2=2.72
r187 105 107 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.395 $Y=2.72
+ $X2=11.73 $Y2=2.72
r188 104 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r189 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r190 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r191 100 103 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r192 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r193 98 117 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.09 $Y=2.72
+ $X2=11.242 $Y2=2.72
r194 98 103 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=11.09 $Y=2.72
+ $X2=10.81 $Y2=2.72
r195 97 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r196 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r197 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r198 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r199 91 94 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r200 90 93 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r201 90 91 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r202 88 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r203 87 88 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r204 85 88 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r205 84 87 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r206 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r207 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r208 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r209 79 82 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r210 79 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r211 78 81 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r212 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r213 76 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.165 $Y2=2.72
r214 76 78 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=2.72
+ $X2=2.53 $Y2=2.72
r215 75 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r216 75 112 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r217 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r218 72 111 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r219 72 74 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r220 71 114 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.165 $Y2=2.72
r221 71 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r222 66 111 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r223 66 68 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r224 64 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r225 64 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r226 62 96 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.43 $Y2=2.72
r227 62 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.62 $Y=2.72
+ $X2=9.705 $Y2=2.72
r228 61 100 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=9.79 $Y=2.72
+ $X2=9.89 $Y2=2.72
r229 61 63 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=2.72
+ $X2=9.705 $Y2=2.72
r230 59 93 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.515 $Y=2.72
+ $X2=8.51 $Y2=2.72
r231 59 60 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.515 $Y=2.72
+ $X2=8.667 $Y2=2.72
r232 58 96 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.82 $Y=2.72
+ $X2=9.43 $Y2=2.72
r233 58 60 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.82 $Y=2.72
+ $X2=8.667 $Y2=2.72
r234 56 87 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.21 $Y2=2.72
r235 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.47 $Y2=2.72
r236 55 90 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.67 $Y2=2.72
r237 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.47 $Y2=2.72
r238 53 81 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.09 $Y=2.72
+ $X2=3.91 $Y2=2.72
r239 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=2.72
+ $X2=4.175 $Y2=2.72
r240 52 84 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.26 $Y=2.72
+ $X2=4.37 $Y2=2.72
r241 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=2.72
+ $X2=4.175 $Y2=2.72
r242 48 51 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=11.242 $Y=1.66
+ $X2=11.242 $Y2=2
r243 46 117 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.242 $Y=2.635
+ $X2=11.242 $Y2=2.72
r244 46 51 23.9935 $w=3.03e-07 $l=6.35e-07 $layer=LI1_cond $X=11.242 $Y=2.635
+ $X2=11.242 $Y2=2
r245 42 63 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.705 $Y=2.635
+ $X2=9.705 $Y2=2.72
r246 42 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.705 $Y=2.635
+ $X2=9.705 $Y2=1.79
r247 38 60 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.667 $Y=2.635
+ $X2=8.667 $Y2=2.72
r248 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.667 $Y=2.635
+ $X2=8.667 $Y2=2.3
r249 34 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2.72
r250 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2
r251 30 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=2.635
+ $X2=4.175 $Y2=2.72
r252 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.175 $Y=2.635
+ $X2=4.175 $Y2=2.33
r253 26 114 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.165 $Y=2.635
+ $X2=2.165 $Y2=2.72
r254 26 28 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.165 $Y=2.635
+ $X2=2.165 $Y2=2.33
r255 22 111 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r256 22 24 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r257 7 51 300 $w=1.7e-07 $l=2.76857e-07 $layer=licon1_PDIFF $count=2 $X=11.02
+ $Y=1.845 $X2=11.23 $Y2=2
r258 7 48 600 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_PDIFF $count=1 $X=11.02
+ $Y=1.845 $X2=11.23 $Y2=1.66
r259 6 44 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=9.56
+ $Y=1.485 $X2=9.705 $Y2=1.79
r260 5 40 600 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_PDIFF $count=1 $X=8.455
+ $Y=2.065 $X2=8.71 $Y2=2.3
r261 4 36 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.085
+ $Y=2.065 $X2=6.47 $Y2=2
r262 3 32 600 $w=1.7e-07 $l=5.63627e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.845 $X2=4.175 $Y2=2.33
r263 2 28 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2.33
r264 1 24 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%A_604_369# 1 2 3 4 13 17 22 24 25 26 27
+ 28 30 32 36 38 39
c118 13 0 1.77453e-19 $X=3.7 $Y=2.33
r119 39 41 18.6318 $w=2.39e-07 $l=3.65e-07 $layer=LI1_cond $X=4.657 $Y=1.91
+ $X2=4.657 $Y2=2.275
r120 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.6 $Y=0.45 $X2=4.7
+ $Y2=0.45
r121 32 39 5.37298 $w=2.39e-07 $l=1.09864e-07 $layer=LI1_cond $X=4.6 $Y=1.825
+ $X2=4.657 $Y2=1.91
r122 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.885 $X2=4.6
+ $Y2=0.8
r123 31 32 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.6 $Y=0.885
+ $X2=4.6 $Y2=1.825
r124 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.715 $X2=4.6
+ $Y2=0.8
r125 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.6 $Y=0.535
+ $X2=4.6 $Y2=0.45
r126 29 30 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.6 $Y=0.535
+ $X2=4.6 $Y2=0.715
r127 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.515 $Y=0.8 $X2=4.6
+ $Y2=0.8
r128 27 28 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=4.515 $Y=0.8
+ $X2=3.875 $Y2=0.8
r129 25 39 2.73298 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=4.515 $Y=1.91
+ $X2=4.657 $Y2=1.91
r130 25 26 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.515 $Y=1.91
+ $X2=3.87 $Y2=1.91
r131 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=0.715
+ $X2=3.875 $Y2=0.8
r132 23 24 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=3.79 $Y=0.445
+ $X2=3.79 $Y2=0.715
r133 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.785 $Y=1.995
+ $X2=3.87 $Y2=1.91
r134 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.785 $Y=1.995
+ $X2=3.785 $Y2=2.245
r135 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.705 $Y=0.36
+ $X2=3.79 $Y2=0.445
r136 17 19 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.705 $Y=0.36
+ $X2=3.245 $Y2=0.36
r137 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.7 $Y=2.33
+ $X2=3.785 $Y2=2.245
r138 13 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.7 $Y=2.33
+ $X2=3.165 $Y2=2.33
r139 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=2.065 $X2=4.715 $Y2=2.275
r140 3 15 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=3.02
+ $Y=1.845 $X2=3.165 $Y2=2.33
r141 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.575
+ $Y=0.235 $X2=4.7 $Y2=0.45
r142 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.055
+ $Y=0.235 $X2=3.245 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%Q 1 2 12 13 14 17
c36 13 0 1.12604e-19 $X=10.21 $Y=1.505
r37 14 21 11.3935 $w=4.78e-07 $l=3.15e-07 $layer=LI1_cond $X=10.2 $Y=0.51
+ $X2=10.2 $Y2=0.825
r38 14 17 2.8656 $w=4.78e-07 $l=1.15e-07 $layer=LI1_cond $X=10.2 $Y=0.51
+ $X2=10.2 $Y2=0.395
r39 13 21 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=10.33 $Y=1.505
+ $X2=10.33 $Y2=0.825
r40 12 13 7.56008 $w=4.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.21 $Y=1.67
+ $X2=10.21 $Y2=1.505
r41 2 12 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=10.03
+ $Y=1.485 $X2=10.175 $Y2=1.67
r42 1 17 91 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_NDIFF $count=2 $X=10.04
+ $Y=0.235 $X2=10.175 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%Q_N 1 2 7 10
r12 7 15 13.1062 $w=2.53e-07 $l=2.9e-07 $layer=LI1_cond $X=11.742 $Y=1.53
+ $X2=11.742 $Y2=1.82
r13 7 10 40.6745 $w=2.53e-07 $l=9e-07 $layer=LI1_cond $X=11.742 $Y=1.53
+ $X2=11.742 $Y2=0.63
r14 2 15 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=11.555
+ $Y=1.485 $X2=11.7 $Y2=1.82
r15 1 10 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=11.565
+ $Y=0.235 $X2=11.7 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXBP_1%VGND 1 2 3 4 5 6 7 24 28 32 36 40 44 47
+ 48 50 51 53 54 55 57 75 79 91 100 101 105 111 114 117
c168 101 0 1.46995e-19 $X=11.73 $Y=0
c169 40 0 1.94529e-19 $X=9.705 $Y=0.53
r170 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r171 114 115 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r172 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r173 105 108 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r174 105 106 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r175 101 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r176 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r177 98 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.395 $Y=0
+ $X2=11.23 $Y2=0
r178 98 100 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=11.395 $Y=0
+ $X2=11.73 $Y2=0
r179 97 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r180 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r181 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r182 93 96 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=9.89 $Y=0 $X2=10.81
+ $Y2=0
r183 93 94 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r184 91 117 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.065 $Y=0
+ $X2=11.23 $Y2=0
r185 91 96 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.065 $Y=0
+ $X2=10.81 $Y2=0
r186 90 94 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=9.89
+ $Y2=0
r187 90 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.51 $Y2=0
r188 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r189 87 114 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.8 $Y=0 $X2=8.59
+ $Y2=0
r190 87 89 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=8.8 $Y=0 $X2=9.43
+ $Y2=0
r191 86 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.51 $Y2=0
r192 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r193 83 86 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r194 83 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r195 82 85 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=0 $X2=8.05
+ $Y2=0
r196 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r197 80 111 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.36 $Y2=0
r198 80 82 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=0
+ $X2=6.67 $Y2=0
r199 79 114 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.38 $Y=0 $X2=8.59
+ $Y2=0
r200 79 85 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=8.38 $Y=0 $X2=8.05
+ $Y2=0
r201 78 112 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.21 $Y2=0
r202 77 78 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r203 75 111 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.175 $Y=0
+ $X2=6.36 $Y2=0
r204 75 77 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=6.175 $Y=0
+ $X2=4.37 $Y2=0
r205 74 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r206 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r207 71 74 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r208 70 73 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r209 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r210 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r211 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r212 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r213 65 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r214 64 67 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r215 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r216 62 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r217 62 64 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r218 57 105 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r219 57 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r220 55 106 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r221 55 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r222 53 89 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=9.62 $Y=0 $X2=9.43
+ $Y2=0
r223 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.62 $Y=0 $X2=9.705
+ $Y2=0
r224 52 93 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=9.79 $Y=0 $X2=9.89
+ $Y2=0
r225 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.79 $Y=0 $X2=9.705
+ $Y2=0
r226 50 73 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=0
+ $X2=3.91 $Y2=0
r227 50 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.095 $Y=0 $X2=4.195
+ $Y2=0
r228 49 77 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.37
+ $Y2=0
r229 49 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.295 $Y=0 $X2=4.195
+ $Y2=0
r230 47 67 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.07
+ $Y2=0
r231 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.31
+ $Y2=0
r232 46 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.53
+ $Y2=0
r233 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.31
+ $Y2=0
r234 42 117 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0
r235 42 44 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.23 $Y=0.085
+ $X2=11.23 $Y2=0.38
r236 38 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.705 $Y=0.085
+ $X2=9.705 $Y2=0
r237 38 40 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.705 $Y=0.085
+ $X2=9.705 $Y2=0.53
r238 34 114 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.59 $Y=0.085
+ $X2=8.59 $Y2=0
r239 34 36 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=8.59 $Y=0.085
+ $X2=8.59 $Y2=0.45
r240 30 111 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0
r241 30 32 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.36 $Y=0.085
+ $X2=6.36 $Y2=0.42
r242 26 51 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=0.085
+ $X2=4.195 $Y2=0
r243 26 28 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=4.195 $Y=0.085
+ $X2=4.195 $Y2=0.38
r244 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=0.085
+ $X2=2.31 $Y2=0
r245 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.31 $Y=0.085
+ $X2=2.31 $Y2=0.36
r246 7 44 91 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_NDIFF $count=2 $X=11.03
+ $Y=0.235 $X2=11.23 $Y2=0.38
r247 6 40 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=9.57
+ $Y=0.235 $X2=9.705 $Y2=0.53
r248 5 36 182 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_NDIFF $count=1 $X=8.58
+ $Y=0.235 $X2=8.715 $Y2=0.45
r249 4 32 182 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_NDIFF $count=1 $X=6.075
+ $Y=0.235 $X2=6.43 $Y2=0.42
r250 3 28 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=3.965
+ $Y=0.235 $X2=4.18 $Y2=0.38
r251 2 24 182 $w=1.7e-07 $l=3.11288e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.31 $Y2=0.36
r252 1 108 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

