* File: sky130_fd_sc_hdll__clkbuf_1.spice
* Created: Thu Aug 27 19:01:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_1.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_1  VNB VPB A X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A	A
* VPB	VPB
* VNB	VNB
MM1003 N_VGND_M1003_d N_A_75_212#_M1003_g N_X_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.169 AS=0.1612 PD=1.17 PS=1.66 NRD=1.152 NRS=10.38 M=1 R=3.46667
+ SA=75000.2 SB=75001 A=0.078 P=1.34 MULT=1
MM1001 N_A_75_212#_M1001_d N_A_M1001_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.52
+ AD=0.1404 AS=0.169 PD=1.58 PS=1.17 NRD=1.152 NRS=5.76 M=1 R=3.46667 SA=75001
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1000 N_VPWR_M1000_d N_A_75_212#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=0.79
+ AD=0.26465 AS=0.2133 PD=1.46 PS=2.12 NRD=3.7233 NRS=1.2411 M=1 R=4.38889
+ SA=90000.2 SB=90001 A=0.1422 P=1.94 MULT=1
MM1002 N_A_75_212#_M1002_d N_A_M1002_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=0.79
+ AD=0.2133 AS=0.26465 PD=2.12 PS=1.46 NRD=1.2411 NRS=8.7271 M=1 R=4.38889
+ SA=90001 SB=90000.2 A=0.1422 P=1.94 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.5631 P=7.65
pX5_noxref noxref_8 VGND VGND PROBETYPE=1
pX6_noxref noxref_9 VPWR VPWR PROBETYPE=1
*
.include "sky130_fd_sc_hdll__clkbuf_1.pxi.spice"
*
.ends
*
*
