* File: sky130_fd_sc_hdll__nor4bb_2.spice
* Created: Thu Aug 27 19:17:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor4bb_2.pex.spice"
.subckt sky130_fd_sc_hdll__nor4bb_2  VNB VPB D_N C_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* C_N	C_N
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1019 N_VGND_M1019_d N_D_N_M1019_g N_A_27_93#_M1019_s VNB NSHORT L=0.15 W=0.42
+ AD=0.08085 AS=0.1092 PD=0.805 PS=1.36 NRD=24.276 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_216_93#_M1002_d N_C_N_M1002_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1197 AS=0.08085 PD=1.41 PS=0.805 NRD=5.712 NRS=5.712 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_Y_M1000_d N_A_216_93#_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2535 PD=0.97 PS=2.08 NRD=0 NRS=23.076 M=1 R=4.33333 SA=75000.3
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1012 N_Y_M1000_d N_A_216_93#_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1012_s N_A_27_93#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1010_d N_A_27_93#_M1010_g N_Y_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_B_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65 AD=0.182
+ AS=0.12025 PD=1.86 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2 SB=75001.7
+ A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_B_M1016_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1005 N_Y_M1005_d N_A_M1005_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1005_d N_A_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.17875 PD=1.02 PS=1.85 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_D_N_M1008_g N_A_27_93#_M1008_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.126812 AS=0.1134 PD=1.34 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1013 N_A_216_93#_M1013_d N_C_N_M1013_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.126812 PD=1.38 PS=1.34 NRD=2.3443 NRS=115.816 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1003 N_A_433_297#_M1003_d N_A_216_93#_M1003_g N_A_343_297#_M1003_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1018 N_A_433_297#_M1003_d N_A_216_93#_M1018_g N_A_343_297#_M1018_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 N_A_343_297#_M1018_s N_A_27_93#_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1017 N_A_343_297#_M1017_d N_A_27_93#_M1017_g N_Y_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1009 N_A_823_297#_M1009_d N_B_M1009_g N_A_433_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 N_A_823_297#_M1015_d N_B_M1015_g N_A_433_297#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_A_823_297#_M1015_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1007 N_A_823_297#_M1007_d N_A_M1007_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.285 AS=0.145 PD=2.57 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__nor4bb_2.pxi.spice"
*
.ends
*
*
