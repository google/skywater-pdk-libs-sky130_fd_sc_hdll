* File: sky130_fd_sc_hdll__and4bb_2.pex.spice
* Created: Thu Aug 27 18:59:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%A_N 2 3 5 8 10 11 19
r32 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r33 15 18 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r34 10 11 22.798 $w=1.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.24 $Y=1.16 $X2=0.24
+ $Y2=1.53
r35 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r36 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r37 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r38 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r39 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r40 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r41 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%A_184_21# 1 2 3 10 12 13 15 16 18 19 21
+ 24 27 28 31 33 34 37 39 40 43 54
c113 39 0 1.28225e-19 $X=3.545 $Y=2
r114 53 54 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.465 $Y=1.202
+ $X2=1.49 $Y2=1.202
r115 52 53 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=1.02 $Y=1.202
+ $X2=1.465 $Y2=1.202
r116 51 52 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=0.995 $Y=1.202
+ $X2=1.02 $Y2=1.202
r117 41 43 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.63 $Y=2.085
+ $X2=3.63 $Y2=2.3
r118 40 50 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2 $X2=2.68
+ $Y2=2
r119 39 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.545 $Y=2
+ $X2=3.63 $Y2=2.085
r120 39 40 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.545 $Y=2
+ $X2=2.765 $Y2=2
r121 35 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.68 $Y=2.085
+ $X2=2.68 $Y2=2
r122 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.68 $Y=2.085
+ $X2=2.68 $Y2=2.3
r123 34 50 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.495 $Y=2
+ $X2=2.68 $Y2=2
r124 33 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.495 $Y=0.72
+ $X2=2.23 $Y2=0.72
r125 33 34 58.146 $w=2.18e-07 $l=1.11e-06 $layer=LI1_cond $X=2.495 $Y=0.805
+ $X2=2.495 $Y2=1.915
r126 29 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.635
+ $X2=2.23 $Y2=0.72
r127 29 31 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.23 $Y=0.635
+ $X2=2.23 $Y2=0.42
r128 27 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=0.72
+ $X2=2.23 $Y2=0.72
r129 27 28 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=2.145 $Y=0.72
+ $X2=1.735 $Y2=0.72
r130 25 54 14.2911 $w=3.71e-07 $l=1.1e-07 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=1.49 $Y2=1.202
r131 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r132 22 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.625 $Y=0.805
+ $X2=1.735 $Y2=0.72
r133 22 24 18.5962 $w=2.18e-07 $l=3.55e-07 $layer=LI1_cond $X=1.625 $Y=0.805
+ $X2=1.625 $Y2=1.16
r134 19 54 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.202
r135 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.985
r136 16 53 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=1.202
r137 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=0.56
r138 13 52 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.202
r139 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r140 10 51 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=1.202
r141 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=0.56
r142 3 43 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=3.485
+ $Y=2.065 $X2=3.63 $Y2=2.3
r143 2 37 600 $w=1.7e-07 $l=3.10403e-07 $layer=licon1_PDIFF $count=1 $X=2.505
+ $Y=2.065 $X2=2.68 $Y2=2.3
r144 1 31 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.105
+ $Y=0.235 $X2=2.23 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%A_27_47# 1 2 8 9 11 14 18 22 24 25 26 27
+ 29 40 46
r95 45 46 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=2.415 $Y=1.16
+ $X2=2.44 $Y2=1.16
r96 41 45 49.8355 $w=3.3e-07 $l=2.85e-07 $layer=POLY_cond $X=2.13 $Y=1.16
+ $X2=2.415 $Y2=1.16
r97 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.13
+ $Y=1.16 $X2=2.13 $Y2=1.16
r98 37 40 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.99 $Y=1.16
+ $X2=2.13 $Y2=1.16
r99 28 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.99 $Y=1.325
+ $X2=1.99 $Y2=1.16
r100 28 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.99 $Y=1.325
+ $X2=1.99 $Y2=1.885
r101 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.905 $Y=1.97
+ $X2=1.99 $Y2=1.885
r102 26 27 77.3102 $w=1.68e-07 $l=1.185e-06 $layer=LI1_cond $X=1.905 $Y=1.97
+ $X2=0.72 $Y2=1.97
r103 25 27 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=0.61 $Y=1.97
+ $X2=0.72 $Y2=1.97
r104 25 34 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.61 $Y=1.97
+ $X2=0.26 $Y2=1.97
r105 24 30 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=0.61 $Y=0.72
+ $X2=0.26 $Y2=0.72
r106 24 25 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=0.61 $Y=0.805
+ $X2=0.61 $Y2=1.885
r107 20 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.055
+ $X2=0.26 $Y2=1.97
r108 20 22 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=2.055
+ $X2=0.26 $Y2=2.3
r109 16 30 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.72
r110 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r111 12 46 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.44 $Y=0.995
+ $X2=2.44 $Y2=1.16
r112 12 14 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.44 $Y=0.995
+ $X2=2.44 $Y2=0.445
r113 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.415 $Y=1.99
+ $X2=2.415 $Y2=2.275
r114 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.415 $Y=1.89 $X2=2.415
+ $Y2=1.99
r115 7 45 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.415 $Y=1.325
+ $X2=2.415 $Y2=1.16
r116 7 8 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.415 $Y=1.325
+ $X2=2.415 $Y2=1.89
r117 2 22 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r118 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%A_545_280# 1 2 8 9 11 14 16 19 20 21 24
+ 27 29 30 37 39
c74 30 0 1.28225e-19 $X=2.88 $Y=1.565
c75 21 0 1.24949e-19 $X=4.105 $Y=2
r76 35 37 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=4.74 $Y=0.42 $X2=4.83
+ $Y2=0.42
r77 30 42 39.9599 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.565
+ $X2=2.87 $Y2=1.73
r78 30 41 48.0588 $w=2.9e-07 $l=1.65e-07 $layer=POLY_cond $X=2.87 $Y=1.565
+ $X2=2.87 $Y2=1.4
r79 29 32 4.97646 $w=2.18e-07 $l=9.5e-08 $layer=LI1_cond $X=2.905 $Y=1.565
+ $X2=2.905 $Y2=1.66
r80 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.88
+ $Y=1.565 $X2=2.88 $Y2=1.565
r81 27 39 4.23118 $w=2.15e-07 $l=1.05119e-07 $layer=LI1_cond $X=4.83 $Y=1.915
+ $X2=4.785 $Y2=2
r82 26 37 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.83 $Y=0.585
+ $X2=4.83 $Y2=0.42
r83 26 27 86.7701 $w=1.68e-07 $l=1.33e-06 $layer=LI1_cond $X=4.83 $Y=0.585
+ $X2=4.83 $Y2=1.915
r84 22 39 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=4.785 $Y=2.085
+ $X2=4.785 $Y2=2
r85 22 24 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=4.785 $Y=2.085
+ $X2=4.785 $Y2=2.3
r86 20 39 2.20034 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.655 $Y=2 $X2=4.785
+ $Y2=2
r87 20 21 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=4.655 $Y=2 $X2=4.105
+ $Y2=2
r88 19 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.995 $Y=1.915
+ $X2=4.105 $Y2=2
r89 18 19 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.995 $Y=1.745
+ $X2=3.995 $Y2=1.915
r90 17 32 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.015 $Y=1.66
+ $X2=2.905 $Y2=1.66
r91 16 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.885 $Y=1.66
+ $X2=3.995 $Y2=1.745
r92 16 17 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=3.885 $Y=1.66
+ $X2=3.015 $Y2=1.66
r93 14 41 489.691 $w=1.5e-07 $l=9.55e-07 $layer=POLY_cond $X=2.935 $Y=0.445
+ $X2=2.935 $Y2=1.4
r94 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.915 $Y=1.99
+ $X2=2.915 $Y2=2.275
r95 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.915 $Y=1.89 $X2=2.915
+ $Y2=1.99
r96 8 42 53.0523 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=2.915 $Y=1.89 $X2=2.915
+ $Y2=1.73
r97 2 24 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.595
+ $Y=2.065 $X2=4.74 $Y2=2.3
r98 1 35 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.605
+ $Y=0.235 $X2=4.74 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%C 2 3 5 8 9 10 11 16 18
c40 3 0 1.24949e-19 $X=3.395 $Y=1.99
r41 16 19 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=0.94
+ $X2=3.36 $Y2=1.105
r42 16 18 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.36 $Y=0.94
+ $X2=3.36 $Y2=0.775
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.36
+ $Y=0.94 $X2=3.36 $Y2=0.94
r44 11 17 10.8721 $w=2.63e-07 $l=2.5e-07 $layer=LI1_cond $X=3.402 $Y=1.19
+ $X2=3.402 $Y2=0.94
r45 10 17 3.91396 $w=2.63e-07 $l=9e-08 $layer=LI1_cond $X=3.402 $Y=0.85
+ $X2=3.402 $Y2=0.94
r46 9 10 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=3.402 $Y=0.51
+ $X2=3.402 $Y2=0.85
r47 8 18 106.04 $w=1.5e-07 $l=3.3e-07 $layer=POLY_cond $X=3.42 $Y=0.445 $X2=3.42
+ $Y2=0.775
r48 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.395 $Y=1.99
+ $X2=3.395 $Y2=2.275
r49 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.395 $Y=1.89 $X2=3.395
+ $Y2=1.99
r50 2 19 260.288 $w=2e-07 $l=7.85e-07 $layer=POLY_cond $X=3.395 $Y=1.89
+ $X2=3.395 $Y2=1.105
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%D 3 6 7 9 10 11 12 17
r47 17 20 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.24 $X2=3.9
+ $Y2=1.405
r48 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.9 $Y=1.24 $X2=3.9
+ $Y2=1.075
r49 12 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.9
+ $Y=1.24 $X2=3.9 $Y2=1.24
r50 11 12 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.855 $Y=0.85
+ $X2=3.855 $Y2=1.19
r51 10 11 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=3.855 $Y=0.51
+ $X2=3.855 $Y2=0.85
r52 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.865 $Y=1.99
+ $X2=3.865 $Y2=2.275
r53 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.865 $Y=1.89 $X2=3.865
+ $Y2=1.99
r54 6 20 160.815 $w=2e-07 $l=4.85e-07 $layer=POLY_cond $X=3.865 $Y=1.89
+ $X2=3.865 $Y2=1.405
r55 3 19 323.043 $w=1.5e-07 $l=6.3e-07 $layer=POLY_cond $X=3.84 $Y=0.445
+ $X2=3.84 $Y2=1.075
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%B_N 2 3 5 8 9 10 14 16 21
c35 14 0 1.38925e-19 $X=4.44 $Y=0.93
r36 15 21 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=4.35 $Y=0.93 $X2=4.35
+ $Y2=0.89
r37 14 17 39.6736 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=0.93
+ $X2=4.455 $Y2=1.095
r38 14 16 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=4.455 $Y=0.93
+ $X2=4.455 $Y2=0.765
r39 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.44
+ $Y=0.93 $X2=4.44 $Y2=0.93
r40 10 15 8.56101 $w=3.48e-07 $l=2.6e-07 $layer=LI1_cond $X=4.35 $Y=1.19
+ $X2=4.35 $Y2=0.93
r41 9 21 1.31708 $w=3.48e-07 $l=4e-08 $layer=LI1_cond $X=4.35 $Y=0.85 $X2=4.35
+ $Y2=0.89
r42 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.53 $Y=0.445
+ $X2=4.53 $Y2=0.765
r43 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.505 $Y=1.99
+ $X2=4.505 $Y2=2.275
r44 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.505 $Y=1.89 $X2=4.505
+ $Y2=1.99
r45 2 17 263.604 $w=2e-07 $l=7.95e-07 $layer=POLY_cond $X=4.505 $Y=1.89
+ $X2=4.505 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%VPWR 1 2 3 4 13 17 20 21 22 24 39 40 43
+ 52 55 57
r80 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r81 57 60 11.2289 $w=3.88e-07 $l=3.8e-07 $layer=LI1_cond $X=3.13 $Y=2.34
+ $X2=3.13 $Y2=2.72
r82 54 55 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.145 $Y=2.53
+ $X2=2.31 $Y2=2.53
r83 51 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r84 50 54 1.63102 $w=5.48e-07 $l=7.5e-08 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=2.145 $Y2=2.53
r85 50 52 15.5949 $w=5.48e-07 $l=4.3e-07 $layer=LI1_cond $X=2.07 $Y=2.53
+ $X2=1.64 $Y2=2.53
r86 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r87 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 43 46 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=2.34
+ $X2=0.705 $Y2=2.72
r89 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r91 37 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r92 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r93 34 60 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.13 $Y2=2.72
r94 34 36 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.91 $Y2=2.72
r95 33 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r96 33 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r97 32 52 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=1.61 $Y=2.72 $X2=1.64
+ $Y2=2.72
r98 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r99 30 46 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r100 30 32 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r101 24 46 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r102 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r103 22 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r104 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r105 20 36 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 20 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.27 $Y2=2.72
r107 19 39 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 19 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.27 $Y2=2.72
r109 15 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=2.635
+ $X2=4.27 $Y2=2.72
r110 15 17 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=4.27 $Y=2.635
+ $X2=4.27 $Y2=2.34
r111 13 60 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=2.935 $Y=2.72
+ $X2=3.13 $Y2=2.72
r112 13 55 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.935 $Y=2.72
+ $X2=2.31 $Y2=2.72
r113 4 17 600 $w=1.7e-07 $l=4.31103e-07 $layer=licon1_PDIFF $count=1 $X=3.955
+ $Y=2.065 $X2=4.27 $Y2=2.34
r114 3 57 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=2.065 $X2=3.15 $Y2=2.34
r115 2 54 300 $w=1.7e-07 $l=1.10186e-06 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.485 $X2=2.145 $Y2=2.34
r116 1 43 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%X 1 2 7 8 9 16 26
r23 26 29 0.628605 $w=2.73e-07 $l=1.5e-08 $layer=LI1_cond $X=1.202 $Y=1.53
+ $X2=1.202 $Y2=1.545
r24 9 29 1.75177 $w=3.53e-07 $l=3.5e-08 $layer=LI1_cond $X=1.242 $Y=1.58
+ $X2=1.242 $Y2=1.545
r25 9 26 1.46675 $w=2.73e-07 $l=3.5e-08 $layer=LI1_cond $X=1.202 $Y=1.495
+ $X2=1.202 $Y2=1.53
r26 8 9 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=1.202 $Y=1.19
+ $X2=1.202 $Y2=1.495
r27 7 8 14.2484 $w=2.73e-07 $l=3.4e-07 $layer=LI1_cond $X=1.202 $Y=0.85
+ $X2=1.202 $Y2=1.19
r28 7 16 18.02 $w=2.73e-07 $l=4.3e-07 $layer=LI1_cond $X=1.202 $Y=0.85 $X2=1.202
+ $Y2=0.42
r29 2 9 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.485 $X2=1.255 $Y2=1.63
r30 1 16 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.255 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4BB_2%VGND 1 2 3 12 15 16 17 19 24 37 38 42 49
c74 37 0 1.38925e-19 $X=4.83 $Y=0
r75 49 52 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.7
+ $Y2=0.38
r76 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r77 42 45 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r78 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r79 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r80 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r81 34 35 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r82 32 35 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r83 32 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r84 31 34 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r85 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r86 29 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.7
+ $Y2=0
r87 29 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.07
+ $Y2=0
r88 28 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r89 28 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r90 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r91 25 42 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r92 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r93 24 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.7
+ $Y2=0
r94 24 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r95 19 42 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r96 19 21 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r97 17 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r98 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r99 15 34 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=3.91
+ $Y2=0
r100 15 16 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.31
+ $Y2=0
r101 14 37 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.83 $Y2=0
r102 14 16 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0 $X2=4.31
+ $Y2=0
r103 10 16 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0
r104 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0.42
r105 3 12 182 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_NDIFF $count=1 $X=3.915
+ $Y=0.235 $X2=4.27 $Y2=0.42
r106 2 52 182 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.71 $Y2=0.38
r107 1 45 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

