* File: sky130_fd_sc_hdll__sdfxtp_4.pxi.spice
* Created: Wed Sep  2 08:52:36 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%CLK N_CLK_c_218_n N_CLK_c_222_n N_CLK_c_219_n
+ N_CLK_M1035_g N_CLK_c_223_n N_CLK_M1001_g CLK
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%CLK
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_27_47# N_A_27_47#_M1035_s N_A_27_47#_M1001_s
+ N_A_27_47#_M1009_g N_A_27_47#_c_268_n N_A_27_47#_c_269_n N_A_27_47#_M1026_g
+ N_A_27_47#_M1034_g N_A_27_47#_c_258_n N_A_27_47#_c_259_n N_A_27_47#_c_272_n
+ N_A_27_47#_c_273_n N_A_27_47#_M1013_g N_A_27_47#_c_274_n N_A_27_47#_c_275_n
+ N_A_27_47#_M1003_g N_A_27_47#_c_260_n N_A_27_47#_M1027_g N_A_27_47#_c_482_p
+ N_A_27_47#_c_262_n N_A_27_47#_c_263_n N_A_27_47#_c_277_n N_A_27_47#_c_384_p
+ N_A_27_47#_c_264_n N_A_27_47#_c_279_n N_A_27_47#_c_280_n N_A_27_47#_c_281_n
+ N_A_27_47#_c_282_n N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_285_n
+ N_A_27_47#_c_265_n N_A_27_47#_c_266_n N_A_27_47#_c_267_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCE N_SCE_c_500_n N_SCE_M1012_g N_SCE_M1016_g
+ N_SCE_c_502_n N_SCE_M1008_g N_SCE_M1036_g N_SCE_c_496_n N_SCE_c_497_n SCE
+ N_SCE_c_503_n N_SCE_c_498_n N_SCE_c_517_p SCE
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCE
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_319_47# N_A_319_47#_M1016_s
+ N_A_319_47#_M1012_s N_A_319_47#_M1020_g N_A_319_47#_c_600_n
+ N_A_319_47#_M1031_g N_A_319_47#_c_595_n N_A_319_47#_c_602_n
+ N_A_319_47#_c_608_n N_A_319_47#_c_596_n N_A_319_47#_c_610_n
+ N_A_319_47#_c_604_n N_A_319_47#_c_597_n N_A_319_47#_c_605_n
+ N_A_319_47#_c_598_n N_A_319_47#_c_599_n N_A_319_47#_c_615_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_319_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%D N_D_c_713_n N_D_M1037_g N_D_M1002_g D D
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%D
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCD N_SCD_M1029_g N_SCD_c_754_n N_SCD_c_755_n
+ N_SCD_M1028_g SCD N_SCD_c_753_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%SCD
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_203_47# N_A_203_47#_M1009_d
+ N_A_203_47#_M1026_d N_A_203_47#_c_818_n N_A_203_47#_M1024_g
+ N_A_203_47#_c_804_n N_A_203_47#_M1021_g N_A_203_47#_c_805_n
+ N_A_203_47#_M1014_g N_A_203_47#_c_819_n N_A_203_47#_M1033_g
+ N_A_203_47#_c_806_n N_A_203_47#_c_807_n N_A_203_47#_c_808_n
+ N_A_203_47#_c_822_n N_A_203_47#_c_809_n N_A_203_47#_c_810_n
+ N_A_203_47#_c_811_n N_A_203_47#_c_812_n N_A_203_47#_c_813_n
+ N_A_203_47#_c_814_n N_A_203_47#_c_815_n N_A_203_47#_c_816_n
+ N_A_203_47#_c_817_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_203_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1189_183# N_A_1189_183#_M1032_d
+ N_A_1189_183#_M1022_d N_A_1189_183#_c_1009_n N_A_1189_183#_c_1016_n
+ N_A_1189_183#_M1000_g N_A_1189_183#_M1007_g N_A_1189_183#_c_1011_n
+ N_A_1189_183#_c_1040_n N_A_1189_183#_c_1059_p N_A_1189_183#_c_1041_n
+ N_A_1189_183#_c_1012_n N_A_1189_183#_c_1026_n N_A_1189_183#_c_1013_n
+ N_A_1189_183#_c_1014_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1189_183#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1011_47# N_A_1011_47#_M1034_d
+ N_A_1011_47#_M1024_d N_A_1011_47#_c_1107_n N_A_1011_47#_c_1115_n
+ N_A_1011_47#_M1022_g N_A_1011_47#_M1032_g N_A_1011_47#_c_1108_n
+ N_A_1011_47#_c_1109_n N_A_1011_47#_c_1110_n N_A_1011_47#_c_1111_n
+ N_A_1011_47#_c_1131_n N_A_1011_47#_c_1135_n N_A_1011_47#_c_1112_n
+ N_A_1011_47#_c_1118_n N_A_1011_47#_c_1113_n N_A_1011_47#_c_1114_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1011_47#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1667_315# N_A_1667_315#_M1019_s
+ N_A_1667_315#_M1030_s N_A_1667_315#_c_1233_n N_A_1667_315#_M1010_g
+ N_A_1667_315#_M1005_g N_A_1667_315#_c_1225_n N_A_1667_315#_M1006_g
+ N_A_1667_315#_c_1235_n N_A_1667_315#_M1004_g N_A_1667_315#_c_1226_n
+ N_A_1667_315#_M1011_g N_A_1667_315#_c_1236_n N_A_1667_315#_M1018_g
+ N_A_1667_315#_c_1227_n N_A_1667_315#_M1015_g N_A_1667_315#_c_1237_n
+ N_A_1667_315#_M1023_g N_A_1667_315#_c_1238_n N_A_1667_315#_M1025_g
+ N_A_1667_315#_c_1228_n N_A_1667_315#_M1017_g N_A_1667_315#_c_1239_n
+ N_A_1667_315#_c_1247_p N_A_1667_315#_c_1229_n N_A_1667_315#_c_1240_n
+ N_A_1667_315#_c_1230_n N_A_1667_315#_c_1231_n N_A_1667_315#_c_1249_p
+ N_A_1667_315#_c_1258_p N_A_1667_315#_c_1232_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1667_315#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1474_413# N_A_1474_413#_M1014_d
+ N_A_1474_413#_M1003_d N_A_1474_413#_c_1369_n N_A_1474_413#_M1030_g
+ N_A_1474_413#_c_1363_n N_A_1474_413#_M1019_g N_A_1474_413#_c_1364_n
+ N_A_1474_413#_c_1365_n N_A_1474_413#_c_1375_n N_A_1474_413#_c_1379_n
+ N_A_1474_413#_c_1372_n N_A_1474_413#_c_1366_n N_A_1474_413#_c_1367_n
+ N_A_1474_413#_c_1368_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_1474_413#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%VPWR N_VPWR_M1001_d N_VPWR_M1012_d
+ N_VPWR_M1028_d N_VPWR_M1000_d N_VPWR_M1010_d N_VPWR_M1030_d N_VPWR_M1018_d
+ N_VPWR_M1025_d N_VPWR_c_1453_n N_VPWR_c_1454_n N_VPWR_c_1455_n N_VPWR_c_1456_n
+ N_VPWR_c_1457_n N_VPWR_c_1458_n N_VPWR_c_1459_n N_VPWR_c_1460_n
+ N_VPWR_c_1461_n N_VPWR_c_1462_n N_VPWR_c_1463_n N_VPWR_c_1464_n
+ N_VPWR_c_1465_n N_VPWR_c_1466_n N_VPWR_c_1467_n N_VPWR_c_1468_n
+ N_VPWR_c_1469_n N_VPWR_c_1470_n N_VPWR_c_1471_n VPWR N_VPWR_c_1472_n
+ N_VPWR_c_1473_n N_VPWR_c_1474_n N_VPWR_c_1475_n N_VPWR_c_1476_n
+ N_VPWR_c_1452_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_608_369# N_A_608_369#_M1002_d
+ N_A_608_369#_M1034_s N_A_608_369#_M1037_d N_A_608_369#_M1024_s
+ N_A_608_369#_c_1640_n N_A_608_369#_c_1652_n N_A_608_369#_c_1664_n
+ N_A_608_369#_c_1629_n N_A_608_369#_c_1636_n N_A_608_369#_c_1637_n
+ N_A_608_369#_c_1630_n N_A_608_369#_c_1631_n N_A_608_369#_c_1632_n
+ N_A_608_369#_c_1633_n N_A_608_369#_c_1634_n N_A_608_369#_c_1635_n
+ N_A_608_369#_c_1639_n PM_SKY130_FD_SC_HDLL__SDFXTP_4%A_608_369#
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%Q N_Q_M1006_s N_Q_M1015_s N_Q_M1004_s
+ N_Q_M1023_s N_Q_c_1759_n N_Q_c_1763_n N_Q_c_1769_n N_Q_c_1752_n N_Q_c_1753_n
+ N_Q_c_1781_n N_Q_c_1785_n N_Q_c_1787_n N_Q_c_1754_n N_Q_c_1757_n N_Q_c_1755_n
+ N_Q_c_1797_n Q PM_SKY130_FD_SC_HDLL__SDFXTP_4%Q
x_PM_SKY130_FD_SC_HDLL__SDFXTP_4%VGND N_VGND_M1035_d N_VGND_M1016_d
+ N_VGND_M1029_d N_VGND_M1007_d N_VGND_M1005_d N_VGND_M1019_d N_VGND_M1011_d
+ N_VGND_M1017_d N_VGND_c_1838_n N_VGND_c_1839_n N_VGND_c_1840_n N_VGND_c_1841_n
+ N_VGND_c_1842_n N_VGND_c_1843_n N_VGND_c_1844_n N_VGND_c_1845_n
+ N_VGND_c_1846_n N_VGND_c_1847_n N_VGND_c_1848_n N_VGND_c_1849_n
+ N_VGND_c_1850_n N_VGND_c_1851_n N_VGND_c_1852_n N_VGND_c_1853_n
+ N_VGND_c_1854_n N_VGND_c_1855_n VGND N_VGND_c_1856_n N_VGND_c_1857_n
+ N_VGND_c_1858_n N_VGND_c_1859_n N_VGND_c_1860_n N_VGND_c_1861_n
+ PM_SKY130_FD_SC_HDLL__SDFXTP_4%VGND
cc_1 VNB N_CLK_c_218_n 0.0583772f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.325
cc_2 VNB N_CLK_c_219_n 0.0176355f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB CLK 0.0188196f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_4 VNB N_A_27_47#_M1009_g 0.0375848f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_5 VNB N_A_27_47#_M1034_g 0.0536074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_258_n 0.0165741f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_259_n 0.00252324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_260_n 0.0211715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1027_g 0.0463832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_262_n 0.00363705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_263_n 0.00651432f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_264_n 0.0026153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_265_n 0.0271693f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_266_n 0.0106206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_267_n 0.00181115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_SCE_M1016_g 0.0523637f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.74
cc_17 VNB N_SCE_M1036_g 0.0173106f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_18 VNB N_SCE_c_496_n 0.00782765f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_19 VNB N_SCE_c_497_n 0.00118673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_SCE_c_498_n 0.0313943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB SCE 0.00459496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_319_47#_M1020_g 0.0222638f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.665
cc_23 VNB N_A_319_47#_c_595_n 0.0138845f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_24 VNB N_A_319_47#_c_596_n 0.00234349f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_319_47#_c_597_n 0.0025595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_319_47#_c_598_n 0.00168005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_319_47#_c_599_n 0.0389429f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_D_M1002_g 0.0460082f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.74
cc_29 VNB N_SCD_M1029_g 0.0452314f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_30 VNB SCD 0.0074008f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_SCD_c_753_n 0.0152332f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_32 VNB N_A_203_47#_c_804_n 0.0187963f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_203_47#_c_805_n 0.0190457f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_34 VNB N_A_203_47#_c_806_n 0.00349774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_203_47#_c_807_n 0.00443734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_203_47#_c_808_n 0.00617897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_203_47#_c_809_n 0.00523362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_203_47#_c_810_n 0.0515315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_203_47#_c_811_n 0.00195192f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_203_47#_c_812_n 0.00133536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_203_47#_c_813_n 0.0100115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_203_47#_c_814_n 0.00514406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_203_47#_c_815_n 0.0322705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_203_47#_c_816_n 0.0341862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_203_47#_c_817_n 0.0158897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_1189_183#_c_1009_n 0.0156207f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=2.135
cc_47 VNB N_A_1189_183#_M1007_g 0.0217505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1189_183#_c_1011_n 0.00519749f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_49 VNB N_A_1189_183#_c_1012_n 0.00138644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1189_183#_c_1013_n 0.00316561f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1189_183#_c_1014_n 0.0360704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1011_47#_c_1107_n 0.0127956f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=2.135
cc_53 VNB N_A_1011_47#_c_1108_n 0.0160928f $X=-0.19 $Y=-0.24 $X2=0.33 $Y2=1.16
cc_54 VNB N_A_1011_47#_c_1109_n 0.017448f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_55 VNB N_A_1011_47#_c_1110_n 0.00885927f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_56 VNB N_A_1011_47#_c_1111_n 0.00101096f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1011_47#_c_1112_n 0.0110107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1011_47#_c_1113_n 0.00197131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1011_47#_c_1114_n 0.00260443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1667_315#_M1005_g 0.051678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1667_315#_c_1225_n 0.0166231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1667_315#_c_1226_n 0.0168542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1667_315#_c_1227_n 0.017288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1667_315#_c_1228_n 0.0200606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1667_315#_c_1229_n 0.00380558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1667_315#_c_1230_n 0.0058217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1667_315#_c_1231_n 0.00722612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1667_315#_c_1232_n 0.0766906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1474_413#_c_1363_n 0.0201833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1474_413#_c_1364_n 0.0399158f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.105
cc_71 VNB N_A_1474_413#_c_1365_n 0.0125491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_A_1474_413#_c_1366_n 0.0106267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_A_1474_413#_c_1367_n 0.00584041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1474_413#_c_1368_n 0.00355647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VPWR_c_1452_n 0.497461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_608_369#_c_1629_n 2.48589e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_608_369#_c_1630_n 0.0157766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_608_369#_c_1631_n 0.00126846f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_608_369#_c_1632_n 0.00359021f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_608_369#_c_1633_n 0.0101757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_608_369#_c_1634_n 0.00249978f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_608_369#_c_1635_n 0.00173494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_Q_c_1752_n 0.00252865f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_Q_c_1753_n 0.00251972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_Q_c_1754_n 0.00859613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_Q_c_1755_n 0.00262045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB Q 0.0209508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1838_n 0.00287347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1839_n 0.00491179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1840_n 0.0058544f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1841_n 0.0026572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1842_n 0.0046831f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1843_n 0.00469613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1844_n 0.0117774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1845_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1846_n 0.0318988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1847_n 0.00512961f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1848_n 0.0405598f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1849_n 0.00381885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1850_n 0.0504733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1851_n 0.00709041f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1852_n 0.0229461f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1853_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1854_n 0.0206863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1855_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1856_n 0.0154125f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1857_n 0.0481245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1858_n 0.0197764f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1859_n 0.0055668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1860_n 0.00610106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1861_n 0.561116f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VPB N_CLK_c_218_n 0.00482568f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_113 VPB N_CLK_c_222_n 0.0166215f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.59
cc_114 VPB N_CLK_c_223_n 0.0478608f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_115 VPB CLK 0.018034f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_116 VPB N_A_27_47#_c_268_n 0.0165313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_A_27_47#_c_269_n 0.0251878f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_118 VPB N_A_27_47#_c_258_n 0.0157764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_27_47#_c_259_n 0.0052974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_27_47#_c_272_n 0.0117186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_27_47#_c_273_n 0.0502981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_27_47#_c_274_n 0.015896f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_27_47#_c_275_n 0.0228905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_27_47#_c_260_n 0.0243073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_47#_c_277_n 0.00135894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_27_47#_c_264_n 0.00368748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_27_47#_c_279_n 0.00358354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_27_47#_c_280_n 0.00307948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_27_47#_c_281_n 0.00819854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_27_47#_c_282_n 0.0599261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_27_47#_c_283_n 9.26987e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_27_47#_c_284_n 0.0050591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_27_47#_c_285_n 0.00111253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_27_47#_c_265_n 0.0120872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_266_n 0.0223882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_27_47#_c_267_n 0.00457659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_SCE_c_500_n 0.0190803f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_138 VPB N_SCE_M1016_g 0.00528153f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_139 VPB N_SCE_c_502_n 0.0160063f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_140 VPB N_SCE_c_503_n 0.0654792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB SCE 0.00295547f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_319_47#_c_600_n 0.0519631f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.665
cc_143 VPB N_A_319_47#_c_595_n 0.0110225f $X=-0.19 $Y=1.305 $X2=0.33 $Y2=1.16
cc_144 VPB N_A_319_47#_c_602_n 0.00408285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_319_47#_c_596_n 0.00570519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_319_47#_c_604_n 0.00286307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_319_47#_c_605_n 0.00183048f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_D_c_713_n 0.0518998f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.325
cc_149 VPB N_D_M1002_g 0.00356251f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_150 VPB D 0.00796807f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_151 VPB N_SCD_c_754_n 0.0089876f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.74
cc_152 VPB N_SCD_c_755_n 0.0275418f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_153 VPB SCD 0.00585825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_SCD_c_753_n 0.0198457f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_155 VPB N_A_203_47#_c_818_n 0.0628983f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_156 VPB N_A_203_47#_c_819_n 0.0548605f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_157 VPB N_A_203_47#_c_806_n 0.00468188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_203_47#_c_807_n 0.00338744f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_203_47#_c_822_n 0.00620308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_203_47#_c_817_n 0.0177176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_1189_183#_c_1009_n 0.0311863f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_162 VPB N_A_1189_183#_c_1016_n 0.0245924f $X=-0.19 $Y=1.305 $X2=0.31
+ $Y2=1.665
cc_163 VPB N_A_1189_183#_c_1013_n 0.00253199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_1011_47#_c_1115_n 0.018063f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.665
cc_165 VPB N_A_1011_47#_c_1110_n 0.0189295f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_166 VPB N_A_1011_47#_c_1111_n 0.0158723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_1011_47#_c_1118_n 0.00162511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_1011_47#_c_1113_n 0.00398233f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_1011_47#_c_1114_n 0.00381428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_1667_315#_c_1233_n 0.0731764f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_171 VPB N_A_1667_315#_M1005_g 0.021917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_1667_315#_c_1235_n 0.0164389f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_173 VPB N_A_1667_315#_c_1236_n 0.016346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_1667_315#_c_1237_n 0.0163429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_1667_315#_c_1238_n 0.0191351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_1667_315#_c_1239_n 0.0129293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_1667_315#_c_1240_n 0.00551938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1667_315#_c_1230_n 0.00560408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1667_315#_c_1232_n 0.0465479f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1474_413#_c_1369_n 0.0198033f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=2.135
cc_181 VPB N_A_1474_413#_c_1364_n 0.0146935f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=1.105
cc_182 VPB N_A_1474_413#_c_1365_n 0.00732599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_1474_413#_c_1372_n 0.0143523f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1474_413#_c_1366_n 0.00422709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_1474_413#_c_1367_n 0.00709413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1453_n 0.00126291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1454_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1455_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1456_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1457_n 0.00548992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1458_n 0.00471485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1459_n 0.00471485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1460_n 0.0121437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1461_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1462_n 0.0429455f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1463_n 0.00324297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1464_n 0.0560185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1465_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1466_n 0.0513405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1467_n 0.00584025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1468_n 0.0234195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1469_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1470_n 0.0216564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_VPWR_c_1471_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_VPWR_c_1472_n 0.0156572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_VPWR_c_1473_n 0.0270443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_VPWR_c_1474_n 0.0213382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_VPWR_c_1475_n 0.0054556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_VPWR_c_1476_n 0.00502699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_VPWR_c_1452_n 0.0634477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_A_608_369#_c_1636_n 0.0113352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_608_369#_c_1637_n 5.59096e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_608_369#_c_1633_n 0.0122437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_608_369#_c_1639_n 0.00885905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_Q_c_1757_n 0.0082934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB Q 0.0101015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 N_CLK_c_218_n N_A_27_47#_M1009_g 0.00437311f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_218 N_CLK_c_219_n N_A_27_47#_M1009_g 0.0161772f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_219 CLK N_A_27_47#_M1009_g 3.44553e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_220 N_CLK_c_222_n N_A_27_47#_c_268_n 0.004446f $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_221 N_CLK_c_223_n N_A_27_47#_c_268_n 0.00668506f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_222 CLK N_A_27_47#_c_268_n 6.27642e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_223 N_CLK_c_223_n N_A_27_47#_c_269_n 0.0192752f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_224 N_CLK_c_218_n N_A_27_47#_c_262_n 0.00788454f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_225 N_CLK_c_219_n N_A_27_47#_c_262_n 0.00700547f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_226 CLK N_A_27_47#_c_262_n 0.00774265f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_227 N_CLK_c_218_n N_A_27_47#_c_263_n 0.00622672f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_228 CLK N_A_27_47#_c_263_n 0.0144574f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_229 N_CLK_c_223_n N_A_27_47#_c_277_n 0.0171149f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_230 CLK N_A_27_47#_c_277_n 0.00731943f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_231 N_CLK_c_218_n N_A_27_47#_c_264_n 0.0045363f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_232 N_CLK_c_222_n N_A_27_47#_c_264_n 7.61846e-19 $X=0.31 $Y=1.59 $X2=0 $Y2=0
cc_233 N_CLK_c_223_n N_A_27_47#_c_264_n 0.0042845f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_234 CLK N_A_27_47#_c_264_n 0.0429434f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_235 N_CLK_c_218_n N_A_27_47#_c_279_n 2.26313e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_236 N_CLK_c_223_n N_A_27_47#_c_279_n 0.007998f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_237 CLK N_A_27_47#_c_279_n 0.0153364f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_238 N_CLK_c_223_n N_A_27_47#_c_280_n 0.00150514f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_239 N_CLK_c_218_n N_A_27_47#_c_265_n 0.0130887f $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_240 CLK N_A_27_47#_c_265_n 0.00184424f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_241 N_CLK_c_223_n N_VPWR_c_1453_n 0.0125197f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_242 N_CLK_c_223_n N_VPWR_c_1472_n 0.00304525f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_243 N_CLK_c_223_n N_VPWR_c_1452_n 0.00455272f $X=0.5 $Y=1.74 $X2=0 $Y2=0
cc_244 N_CLK_c_218_n N_VGND_c_1856_n 4.61451e-19 $X=0.31 $Y=1.325 $X2=0 $Y2=0
cc_245 N_CLK_c_219_n N_VGND_c_1856_n 0.00340075f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_246 N_CLK_c_219_n N_VGND_c_1859_n 0.0115525f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_247 N_CLK_c_219_n N_VGND_c_1861_n 0.00497799f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_282_n N_SCE_c_500_n 0.00317255f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_249 N_A_27_47#_c_282_n N_SCE_c_502_n 0.00121046f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_282_n N_SCE_c_503_n 0.00470527f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_282_n SCE 0.00858979f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_282_n N_A_319_47#_c_600_n 0.00355626f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_253 N_A_27_47#_c_282_n N_A_319_47#_c_595_n 0.012706f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_282_n N_A_319_47#_c_608_n 0.0211859f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_282_n N_A_319_47#_c_596_n 0.00964382f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_256 N_A_27_47#_c_282_n N_A_319_47#_c_610_n 0.0357899f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_282_n N_A_319_47#_c_604_n 0.0130171f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_M1009_g N_A_319_47#_c_597_n 9.20042e-19 $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_c_282_n N_A_319_47#_c_605_n 0.0130533f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_282_n N_A_319_47#_c_599_n 0.00321182f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_282_n N_A_319_47#_c_615_n 0.00491135f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_262 N_A_27_47#_c_282_n N_D_c_713_n 0.00665992f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_263 N_A_27_47#_c_282_n D 0.0102357f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_282_n N_SCD_c_755_n 0.00274884f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_282_n SCD 0.00910253f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_282_n N_SCD_c_753_n 0.0013799f $X=5.555 $Y=1.825 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_282_n N_A_203_47#_M1026_d 7.52281e-19 $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_268 N_A_27_47#_c_259_n N_A_203_47#_c_818_n 0.0194945f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_273_n N_A_203_47#_c_818_n 0.0316637f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_281_n N_A_203_47#_c_818_n 0.00224123f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_271 N_A_27_47#_c_282_n N_A_203_47#_c_818_n 0.0095879f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_M1034_g N_A_203_47#_c_804_n 0.0121859f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_M1027_g N_A_203_47#_c_805_n 0.013629f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_274_n N_A_203_47#_c_819_n 0.0184424f $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_275_n N_A_203_47#_c_819_n 0.0117705f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_260_n N_A_203_47#_c_819_n 0.0237682f $X=7.975 $Y=1.32 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_284_n N_A_203_47#_c_819_n 6.9418e-19 $X=7.31 $Y=1.825 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_267_n N_A_203_47#_c_819_n 0.00177751f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_27_47#_M1034_g N_A_203_47#_c_806_n 0.00796706f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_280 N_A_27_47#_c_258_n N_A_203_47#_c_806_n 0.00910826f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_281 N_A_27_47#_c_259_n N_A_203_47#_c_806_n 0.00418731f $X=5.055 $Y=1.32 $X2=0
+ $Y2=0
cc_282 N_A_27_47#_c_272_n N_A_203_47#_c_806_n 0.00639348f $X=5.515 $Y=1.575
+ $X2=0 $Y2=0
cc_283 N_A_27_47#_c_273_n N_A_203_47#_c_806_n 7.35344e-19 $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_c_281_n N_A_203_47#_c_806_n 0.0169317f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_285 N_A_27_47#_c_282_n N_A_203_47#_c_806_n 0.0161657f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_286 N_A_27_47#_c_283_n N_A_203_47#_c_806_n 4.35179e-19 $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_287 N_A_27_47#_c_260_n N_A_203_47#_c_807_n 0.0120753f $X=7.975 $Y=1.32 $X2=0
+ $Y2=0
cc_288 N_A_27_47#_M1027_g N_A_203_47#_c_807_n 0.00393345f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_266_n N_A_203_47#_c_807_n 0.00416507f $X=7.275 $Y=1.32 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_267_n N_A_203_47#_c_807_n 0.023853f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_M1027_g N_A_203_47#_c_808_n 0.0022503f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_266_n N_A_203_47#_c_808_n 0.00228363f $X=7.275 $Y=1.32 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_c_267_n N_A_203_47#_c_808_n 0.0151119f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_c_274_n N_A_203_47#_c_822_n 0.0011999f $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_c_260_n N_A_203_47#_c_822_n 0.00449357f $X=7.975 $Y=1.32 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_284_n N_A_203_47#_c_822_n 0.00656065f $X=7.31 $Y=1.825 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_267_n N_A_203_47#_c_822_n 0.024565f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_M1009_g N_A_203_47#_c_809_n 0.00640849f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_262_n N_A_203_47#_c_809_n 0.00344258f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_c_264_n N_A_203_47#_c_809_n 0.00374014f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1034_g N_A_203_47#_c_810_n 0.00225641f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1034_g N_A_203_47#_c_811_n 3.57691e-19 $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_303 N_A_27_47#_c_266_n N_A_203_47#_c_812_n 0.00119328f $X=7.275 $Y=1.32 $X2=0
+ $Y2=0
cc_304 N_A_27_47#_c_267_n N_A_203_47#_c_812_n 0.00143873f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_305 N_A_27_47#_c_258_n N_A_203_47#_c_813_n 4.20893e-19 $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_306 N_A_27_47#_M1034_g N_A_203_47#_c_814_n 0.0122484f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_307 N_A_27_47#_c_258_n N_A_203_47#_c_814_n 0.00609027f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_308 N_A_27_47#_c_281_n N_A_203_47#_c_814_n 0.00398178f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_M1034_g N_A_203_47#_c_815_n 0.0163838f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_258_n N_A_203_47#_c_815_n 0.0211553f $X=5.415 $Y=1.32 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_273_n N_A_203_47#_c_815_n 5.43883e-19 $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_281_n N_A_203_47#_c_815_n 6.38247e-19 $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_313 N_A_27_47#_M1027_g N_A_203_47#_c_816_n 0.0118259f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_266_n N_A_203_47#_c_816_n 0.0234243f $X=7.275 $Y=1.32 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_267_n N_A_203_47#_c_816_n 3.7895e-19 $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_316 N_A_27_47#_M1009_g N_A_203_47#_c_817_n 0.0133504f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_269_n N_A_203_47#_c_817_n 0.00212706f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_262_n N_A_203_47#_c_817_n 0.00981189f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_384_p N_A_203_47#_c_817_n 0.006717f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_320 N_A_27_47#_c_264_n N_A_203_47#_c_817_n 0.0584555f $X=0.81 $Y=1.235 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_280_n N_A_203_47#_c_817_n 0.00207039f $X=0.895 $Y=1.825
+ $X2=0 $Y2=0
cc_322 N_A_27_47#_c_282_n N_A_203_47#_c_817_n 0.0255099f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_265_n N_A_203_47#_c_817_n 0.0167016f $X=0.97 $Y=1.235 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_285_n N_A_1189_183#_M1022_d 0.00523078f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_258_n N_A_1189_183#_c_1009_n 0.0118986f $X=5.415 $Y=1.32
+ $X2=0 $Y2=0
cc_326 N_A_27_47#_c_273_n N_A_1189_183#_c_1009_n 0.0209627f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_327 N_A_27_47#_c_281_n N_A_1189_183#_c_1009_n 0.00212256f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_328 N_A_27_47#_c_283_n N_A_1189_183#_c_1009_n 0.00152496f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_329 N_A_27_47#_c_285_n N_A_1189_183#_c_1009_n 0.00150072f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_330 N_A_27_47#_c_273_n N_A_1189_183#_c_1016_n 0.0264165f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_331 N_A_27_47#_c_285_n N_A_1189_183#_c_1016_n 0.00126931f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_275_n N_A_1189_183#_c_1026_n 0.00554009f $X=7.28 $Y=1.99
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_285_n N_A_1189_183#_c_1026_n 0.00261642f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_334 N_A_27_47#_c_274_n N_A_1189_183#_c_1013_n 0.00121845f $X=7.28 $Y=1.89
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_275_n N_A_1189_183#_c_1013_n 0.00370799f $X=7.28 $Y=1.99
+ $X2=0 $Y2=0
cc_336 N_A_27_47#_c_284_n N_A_1189_183#_c_1013_n 0.00281477f $X=7.31 $Y=1.825
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_285_n N_A_1189_183#_c_1013_n 0.0240109f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_338 N_A_27_47#_c_266_n N_A_1189_183#_c_1013_n 0.00232864f $X=7.275 $Y=1.32
+ $X2=0 $Y2=0
cc_339 N_A_27_47#_c_267_n N_A_1189_183#_c_1013_n 0.0530513f $X=7.25 $Y=1.41
+ $X2=0 $Y2=0
cc_340 N_A_27_47#_c_266_n N_A_1011_47#_c_1107_n 0.0159377f $X=7.275 $Y=1.32
+ $X2=0 $Y2=0
cc_341 N_A_27_47#_c_267_n N_A_1011_47#_c_1107_n 3.02222e-19 $X=7.25 $Y=1.41
+ $X2=0 $Y2=0
cc_342 N_A_27_47#_c_274_n N_A_1011_47#_c_1115_n 0.0116663f $X=7.28 $Y=1.89 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_c_275_n N_A_1011_47#_c_1115_n 0.0139731f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_c_285_n N_A_1011_47#_c_1115_n 0.00642704f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_345 N_A_27_47#_c_267_n N_A_1011_47#_c_1115_n 6.1879e-19 $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_346 N_A_27_47#_c_285_n N_A_1011_47#_c_1110_n 0.00109659f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_347 N_A_27_47#_c_274_n N_A_1011_47#_c_1111_n 0.00314415f $X=7.28 $Y=1.89
+ $X2=0 $Y2=0
cc_348 N_A_27_47#_c_285_n N_A_1011_47#_c_1111_n 2.82791e-19 $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_349 N_A_27_47#_c_267_n N_A_1011_47#_c_1111_n 2.11637e-19 $X=7.25 $Y=1.41
+ $X2=0 $Y2=0
cc_350 N_A_27_47#_c_273_n N_A_1011_47#_c_1131_n 0.0105456f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_351 N_A_27_47#_c_281_n N_A_1011_47#_c_1131_n 0.0282373f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_352 N_A_27_47#_c_282_n N_A_1011_47#_c_1131_n 0.00865498f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_353 N_A_27_47#_c_283_n N_A_1011_47#_c_1131_n 0.00430757f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_354 N_A_27_47#_M1034_g N_A_1011_47#_c_1135_n 0.0017473f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_355 N_A_27_47#_M1034_g N_A_1011_47#_c_1112_n 8.9875e-19 $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_356 N_A_27_47#_c_273_n N_A_1011_47#_c_1118_n 0.00172804f $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_357 N_A_27_47#_c_281_n N_A_1011_47#_c_1118_n 0.0253723f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_358 N_A_27_47#_c_283_n N_A_1011_47#_c_1118_n 0.00267624f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_359 N_A_27_47#_c_285_n N_A_1011_47#_c_1118_n 0.0230281f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_360 N_A_27_47#_c_258_n N_A_1011_47#_c_1113_n 0.00356727f $X=5.415 $Y=1.32
+ $X2=0 $Y2=0
cc_361 N_A_27_47#_c_272_n N_A_1011_47#_c_1113_n 4.58809e-19 $X=5.515 $Y=1.575
+ $X2=0 $Y2=0
cc_362 N_A_27_47#_c_273_n N_A_1011_47#_c_1113_n 2.56759e-19 $X=5.515 $Y=1.99
+ $X2=0 $Y2=0
cc_363 N_A_27_47#_c_281_n N_A_1011_47#_c_1113_n 0.012133f $X=5.75 $Y=1.825 $X2=0
+ $Y2=0
cc_364 N_A_27_47#_c_283_n N_A_1011_47#_c_1113_n 0.00215015f $X=5.895 $Y=1.825
+ $X2=0 $Y2=0
cc_365 N_A_27_47#_c_285_n N_A_1011_47#_c_1113_n 0.0053751f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_366 N_A_27_47#_c_285_n N_A_1011_47#_c_1114_n 0.0121788f $X=7.115 $Y=1.825
+ $X2=0 $Y2=0
cc_367 N_A_27_47#_M1027_g N_A_1667_315#_M1005_g 0.0463022f $X=8.05 $Y=0.415
+ $X2=0 $Y2=0
cc_368 N_A_27_47#_c_275_n N_A_1474_413#_c_1375_n 0.00455494f $X=7.28 $Y=1.99
+ $X2=0 $Y2=0
cc_369 N_A_27_47#_c_284_n N_A_1474_413#_c_1375_n 0.00192009f $X=7.31 $Y=1.825
+ $X2=0 $Y2=0
cc_370 N_A_27_47#_c_266_n N_A_1474_413#_c_1375_n 4.94934e-19 $X=7.275 $Y=1.32
+ $X2=0 $Y2=0
cc_371 N_A_27_47#_c_267_n N_A_1474_413#_c_1375_n 0.00520742f $X=7.25 $Y=1.41
+ $X2=0 $Y2=0
cc_372 N_A_27_47#_M1027_g N_A_1474_413#_c_1379_n 0.00860822f $X=8.05 $Y=0.415
+ $X2=0 $Y2=0
cc_373 N_A_27_47#_M1027_g N_A_1474_413#_c_1366_n 3.1587e-19 $X=8.05 $Y=0.415
+ $X2=0 $Y2=0
cc_374 N_A_27_47#_c_260_n N_A_1474_413#_c_1367_n 0.00730991f $X=7.975 $Y=1.32
+ $X2=0 $Y2=0
cc_375 N_A_27_47#_M1027_g N_A_1474_413#_c_1367_n 0.00725207f $X=8.05 $Y=0.415
+ $X2=0 $Y2=0
cc_376 N_A_27_47#_M1027_g N_A_1474_413#_c_1368_n 0.0132802f $X=8.05 $Y=0.415
+ $X2=0 $Y2=0
cc_377 N_A_27_47#_c_384_p N_VPWR_M1001_d 0.00171205f $X=0.78 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_378 N_A_27_47#_c_285_n N_VPWR_M1000_d 0.00711711f $X=7.115 $Y=1.825 $X2=0
+ $Y2=0
cc_379 N_A_27_47#_c_269_n N_VPWR_c_1453_n 0.00955536f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_380 N_A_27_47#_c_277_n N_VPWR_c_1453_n 0.00629408f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_381 N_A_27_47#_c_384_p N_VPWR_c_1453_n 0.0135522f $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_382 N_A_27_47#_c_279_n N_VPWR_c_1453_n 0.0246493f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_383 N_A_27_47#_c_280_n N_VPWR_c_1453_n 0.00146287f $X=0.895 $Y=1.825 $X2=0
+ $Y2=0
cc_384 N_A_27_47#_c_282_n N_VPWR_c_1454_n 0.00142595f $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_385 N_A_27_47#_c_282_n N_VPWR_c_1455_n 8.00522e-19 $X=5.555 $Y=1.825 $X2=0
+ $Y2=0
cc_386 N_A_27_47#_c_285_n N_VPWR_c_1456_n 0.00945054f $X=7.115 $Y=1.825 $X2=0
+ $Y2=0
cc_387 N_A_27_47#_c_273_n N_VPWR_c_1464_n 0.00454633f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_388 N_A_27_47#_c_275_n N_VPWR_c_1466_n 0.00519523f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_389 N_A_27_47#_c_267_n N_VPWR_c_1466_n 0.00189776f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_390 N_A_27_47#_c_277_n N_VPWR_c_1472_n 0.00180073f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_391 N_A_27_47#_c_279_n N_VPWR_c_1472_n 0.0120313f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_392 N_A_27_47#_c_269_n N_VPWR_c_1473_n 0.00590576f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_393 N_A_27_47#_c_269_n N_VPWR_c_1452_n 0.00667006f $X=0.97 $Y=1.74 $X2=0
+ $Y2=0
cc_394 N_A_27_47#_c_273_n N_VPWR_c_1452_n 0.00640619f $X=5.515 $Y=1.99 $X2=0
+ $Y2=0
cc_395 N_A_27_47#_c_275_n N_VPWR_c_1452_n 0.00684001f $X=7.28 $Y=1.99 $X2=0
+ $Y2=0
cc_396 N_A_27_47#_c_277_n N_VPWR_c_1452_n 0.00425497f $X=0.665 $Y=1.88 $X2=0
+ $Y2=0
cc_397 N_A_27_47#_c_384_p N_VPWR_c_1452_n 5.98513e-19 $X=0.78 $Y=1.795 $X2=0
+ $Y2=0
cc_398 N_A_27_47#_c_279_n N_VPWR_c_1452_n 0.00646745f $X=0.265 $Y=1.96 $X2=0
+ $Y2=0
cc_399 N_A_27_47#_c_280_n N_VPWR_c_1452_n 0.319583f $X=0.895 $Y=1.825 $X2=0
+ $Y2=0
cc_400 N_A_27_47#_c_267_n N_VPWR_c_1452_n 0.00165953f $X=7.25 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A_27_47#_c_282_n N_A_608_369#_c_1640_n 0.00705026f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_402 N_A_27_47#_c_282_n N_A_608_369#_c_1636_n 0.0293627f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_403 N_A_27_47#_c_282_n N_A_608_369#_c_1637_n 0.00852023f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_404 N_A_27_47#_M1034_g N_A_608_369#_c_1632_n 0.0044467f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_405 N_A_27_47#_M1034_g N_A_608_369#_c_1633_n 0.00914943f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_406 N_A_27_47#_c_282_n N_A_608_369#_c_1633_n 0.0104876f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_407 N_A_27_47#_M1034_g N_A_608_369#_c_1634_n 0.0020076f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_408 N_A_27_47#_M1034_g N_A_608_369#_c_1635_n 0.00164257f $X=4.98 $Y=0.415
+ $X2=0 $Y2=0
cc_409 N_A_27_47#_c_281_n N_A_608_369#_c_1639_n 0.00293569f $X=5.75 $Y=1.825
+ $X2=0 $Y2=0
cc_410 N_A_27_47#_c_282_n N_A_608_369#_c_1639_n 0.011045f $X=5.555 $Y=1.825
+ $X2=0 $Y2=0
cc_411 N_A_27_47#_c_282_n A_702_369# 0.00154833f $X=5.555 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_412 N_A_27_47#_c_262_n N_VGND_M1035_d 0.00215637f $X=0.665 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_413 N_A_27_47#_M1034_g N_VGND_c_1839_n 0.00339332f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_414 N_A_27_47#_M1027_g N_VGND_c_1841_n 0.00231736f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_415 N_A_27_47#_M1009_g N_VGND_c_1846_n 0.00468308f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_416 N_A_27_47#_M1034_g N_VGND_c_1850_n 0.00431421f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_417 N_A_27_47#_c_482_p N_VGND_c_1856_n 0.00713694f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_418 N_A_27_47#_c_262_n N_VGND_c_1856_n 0.00244629f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_419 N_A_27_47#_M1027_g N_VGND_c_1857_n 0.00379633f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_420 N_A_27_47#_M1009_g N_VGND_c_1859_n 0.0101565f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_421 N_A_27_47#_c_262_n N_VGND_c_1859_n 0.0211078f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_422 N_A_27_47#_c_265_n N_VGND_c_1859_n 5.78916e-19 $X=0.97 $Y=1.235 $X2=0
+ $Y2=0
cc_423 N_A_27_47#_M1035_s N_VGND_c_1861_n 0.003754f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_424 N_A_27_47#_M1009_g N_VGND_c_1861_n 0.00934478f $X=0.94 $Y=0.445 $X2=0
+ $Y2=0
cc_425 N_A_27_47#_M1034_g N_VGND_c_1861_n 0.00742063f $X=4.98 $Y=0.415 $X2=0
+ $Y2=0
cc_426 N_A_27_47#_M1027_g N_VGND_c_1861_n 0.00604059f $X=8.05 $Y=0.415 $X2=0
+ $Y2=0
cc_427 N_A_27_47#_c_482_p N_VGND_c_1861_n 0.00608739f $X=0.26 $Y=0.51 $X2=0
+ $Y2=0
cc_428 N_A_27_47#_c_262_n N_VGND_c_1861_n 0.00602661f $X=0.665 $Y=0.72 $X2=0
+ $Y2=0
cc_429 N_SCE_M1016_g N_A_319_47#_M1020_g 0.0172933f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_430 N_SCE_c_496_n N_A_319_47#_M1020_g 0.0115622f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_431 SCE N_A_319_47#_M1020_g 0.00149975f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_432 N_SCE_c_497_n N_A_319_47#_c_600_n 2.11997e-19 $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_433 N_SCE_c_498_n N_A_319_47#_c_600_n 0.0178626f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_434 N_SCE_c_500_n N_A_319_47#_c_595_n 0.00268171f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_435 N_SCE_M1016_g N_A_319_47#_c_595_n 0.0181395f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_436 N_SCE_c_503_n N_A_319_47#_c_595_n 0.0110375f $X=1.965 $Y=1.52 $X2=0 $Y2=0
cc_437 N_SCE_c_517_p N_A_319_47#_c_595_n 0.0128929f $X=2.047 $Y=0.785 $X2=0
+ $Y2=0
cc_438 SCE N_A_319_47#_c_595_n 0.065136f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_439 N_SCE_c_500_n N_A_319_47#_c_602_n 0.00579439f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_440 N_SCE_c_500_n N_A_319_47#_c_608_n 0.0137121f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_441 N_SCE_c_502_n N_A_319_47#_c_608_n 0.00528858f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_442 N_SCE_c_503_n N_A_319_47#_c_608_n 0.00610816f $X=1.965 $Y=1.52 $X2=0
+ $Y2=0
cc_443 SCE N_A_319_47#_c_608_n 0.0212535f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_444 N_SCE_c_500_n N_A_319_47#_c_596_n 6.74057e-19 $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_445 N_SCE_M1016_g N_A_319_47#_c_596_n 9.99138e-19 $X=1.95 $Y=0.445 $X2=0
+ $Y2=0
cc_446 N_SCE_c_502_n N_A_319_47#_c_596_n 0.00301815f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_447 N_SCE_c_503_n N_A_319_47#_c_596_n 0.0108547f $X=1.965 $Y=1.52 $X2=0 $Y2=0
cc_448 SCE N_A_319_47#_c_596_n 0.0429658f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_449 N_SCE_c_497_n N_A_319_47#_c_604_n 0.00960462f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_450 N_SCE_c_498_n N_A_319_47#_c_604_n 3.97341e-19 $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_451 N_SCE_M1016_g N_A_319_47#_c_597_n 0.0026078f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_452 N_SCE_c_517_p N_A_319_47#_c_597_n 0.00168685f $X=2.047 $Y=0.785 $X2=0
+ $Y2=0
cc_453 N_SCE_c_503_n N_A_319_47#_c_605_n 3.36465e-19 $X=1.965 $Y=1.52 $X2=0
+ $Y2=0
cc_454 N_SCE_c_496_n N_A_319_47#_c_598_n 0.0198926f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_455 N_SCE_c_497_n N_A_319_47#_c_598_n 0.00387695f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_456 SCE N_A_319_47#_c_598_n 0.0133755f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_457 N_SCE_M1016_g N_A_319_47#_c_599_n 0.0114642f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_458 N_SCE_c_496_n N_A_319_47#_c_599_n 0.0050517f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_459 N_SCE_c_503_n N_A_319_47#_c_599_n 0.00762323f $X=1.965 $Y=1.52 $X2=0
+ $Y2=0
cc_460 SCE N_A_319_47#_c_599_n 0.00357615f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_461 N_SCE_c_502_n N_A_319_47#_c_615_n 0.0087726f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_462 N_SCE_c_502_n N_D_c_713_n 0.0317564f $X=2.43 $Y=1.77 $X2=-0.19 $Y2=-0.24
cc_463 N_SCE_c_496_n N_D_c_713_n 9.61584e-19 $X=3.335 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_464 N_SCE_c_503_n N_D_c_713_n 0.0162646f $X=1.965 $Y=1.52 $X2=-0.19 $Y2=-0.24
cc_465 N_SCE_M1036_g N_D_M1002_g 0.0117556f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_466 N_SCE_c_496_n N_D_M1002_g 0.0132698f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_467 N_SCE_c_497_n N_D_M1002_g 0.00203037f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_468 N_SCE_c_498_n N_D_M1002_g 0.0215793f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_469 N_SCE_c_496_n D 0.00666421f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_470 N_SCE_c_503_n D 2.13149e-19 $X=1.965 $Y=1.52 $X2=0 $Y2=0
cc_471 N_SCE_M1036_g N_SCD_M1029_g 0.0574661f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_472 N_SCE_c_497_n N_SCD_M1029_g 0.00124626f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_473 N_SCE_c_497_n SCD 0.00503288f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_474 N_SCE_c_498_n SCD 5.8751e-19 $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_475 N_SCE_M1016_g N_A_203_47#_c_810_n 0.00255572f $X=1.95 $Y=0.445 $X2=0
+ $Y2=0
cc_476 N_SCE_M1036_g N_A_203_47#_c_810_n 0.00105565f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_477 N_SCE_c_496_n N_A_203_47#_c_810_n 0.0427685f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_478 N_SCE_c_497_n N_A_203_47#_c_810_n 0.0110804f $X=3.42 $Y=0.95 $X2=0 $Y2=0
cc_479 N_SCE_c_503_n N_A_203_47#_c_810_n 0.00375664f $X=1.965 $Y=1.52 $X2=0
+ $Y2=0
cc_480 N_SCE_c_498_n N_A_203_47#_c_810_n 0.00457721f $X=3.53 $Y=0.95 $X2=0 $Y2=0
cc_481 N_SCE_c_517_p N_A_203_47#_c_810_n 0.00679413f $X=2.047 $Y=0.785 $X2=0
+ $Y2=0
cc_482 SCE N_A_203_47#_c_810_n 0.0239947f $X=2.07 $Y=0.84 $X2=0 $Y2=0
cc_483 N_SCE_c_500_n N_A_203_47#_c_817_n 0.00143269f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_484 N_SCE_c_500_n N_VPWR_c_1454_n 0.0113766f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_485 N_SCE_c_502_n N_VPWR_c_1454_n 0.00947361f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_486 N_SCE_c_502_n N_VPWR_c_1462_n 0.00454152f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_487 N_SCE_c_500_n N_VPWR_c_1473_n 0.00312096f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_488 N_SCE_c_500_n N_VPWR_c_1452_n 0.00489637f $X=1.96 $Y=1.77 $X2=0 $Y2=0
cc_489 N_SCE_c_502_n N_VPWR_c_1452_n 0.00504866f $X=2.43 $Y=1.77 $X2=0 $Y2=0
cc_490 N_SCE_c_496_n N_A_608_369#_M1002_d 0.00271541f $X=3.335 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_491 N_SCE_c_502_n N_A_608_369#_c_1640_n 6.17318e-19 $X=2.43 $Y=1.77 $X2=0
+ $Y2=0
cc_492 N_SCE_M1036_g N_A_608_369#_c_1652_n 0.00787009f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_493 N_SCE_c_496_n N_A_608_369#_c_1652_n 0.0209567f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_494 N_SCE_c_498_n N_A_608_369#_c_1652_n 4.66881e-19 $X=3.53 $Y=0.95 $X2=0
+ $Y2=0
cc_495 N_SCE_M1036_g N_A_608_369#_c_1629_n 0.00410769f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_496 N_SCE_c_496_n N_A_608_369#_c_1629_n 0.00517226f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_497 N_SCE_M1036_g N_A_608_369#_c_1631_n 0.00111248f $X=3.53 $Y=0.445 $X2=0
+ $Y2=0
cc_498 N_SCE_c_496_n N_A_608_369#_c_1631_n 0.00650856f $X=3.335 $Y=0.7 $X2=0
+ $Y2=0
cc_499 N_SCE_c_497_n N_A_608_369#_c_1631_n 0.00423271f $X=3.42 $Y=0.95 $X2=0
+ $Y2=0
cc_500 N_SCE_c_496_n N_VGND_M1016_d 0.00173449f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_501 N_SCE_c_517_p N_VGND_M1016_d 0.00173341f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_502 N_SCE_M1016_g N_VGND_c_1838_n 0.0053869f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_503 N_SCE_c_496_n N_VGND_c_1838_n 0.0126787f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_504 N_SCE_c_517_p N_VGND_c_1838_n 0.0069839f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_505 N_SCE_M1016_g N_VGND_c_1846_n 0.00409976f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_506 N_SCE_c_517_p N_VGND_c_1846_n 0.00370519f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_507 N_SCE_M1036_g N_VGND_c_1848_n 0.00362032f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_508 N_SCE_c_496_n N_VGND_c_1848_n 0.0100187f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_509 N_SCE_M1016_g N_VGND_c_1861_n 0.00710252f $X=1.95 $Y=0.445 $X2=0 $Y2=0
cc_510 N_SCE_M1036_g N_VGND_c_1861_n 0.00537207f $X=3.53 $Y=0.445 $X2=0 $Y2=0
cc_511 N_SCE_c_496_n N_VGND_c_1861_n 0.00827087f $X=3.335 $Y=0.7 $X2=0 $Y2=0
cc_512 N_SCE_c_517_p N_VGND_c_1861_n 0.0032373f $X=2.047 $Y=0.785 $X2=0 $Y2=0
cc_513 N_SCE_c_496_n A_517_47# 0.00384984f $X=3.335 $Y=0.7 $X2=-0.19 $Y2=-0.24
cc_514 N_A_319_47#_c_600_n N_D_c_713_n 0.0473103f $X=3.42 $Y=1.77 $X2=-0.19
+ $Y2=-0.24
cc_515 N_A_319_47#_c_596_n N_D_c_713_n 0.00393982f $X=2.47 $Y=1.86 $X2=-0.19
+ $Y2=-0.24
cc_516 N_A_319_47#_c_610_n N_D_c_713_n 0.0170557f $X=3.33 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_517 N_A_319_47#_c_604_n N_D_c_713_n 0.00164299f $X=3.44 $Y=1.52 $X2=-0.19
+ $Y2=-0.24
cc_518 N_A_319_47#_M1020_g N_D_M1002_g 0.0291087f $X=2.51 $Y=0.445 $X2=0 $Y2=0
cc_519 N_A_319_47#_c_596_n N_D_M1002_g 0.00523437f $X=2.47 $Y=1.86 $X2=0 $Y2=0
cc_520 N_A_319_47#_c_598_n N_D_M1002_g 6.95674e-19 $X=2.55 $Y=1.04 $X2=0 $Y2=0
cc_521 N_A_319_47#_c_599_n N_D_M1002_g 0.0190245f $X=2.55 $Y=1.04 $X2=0 $Y2=0
cc_522 N_A_319_47#_c_600_n D 0.0019877f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_523 N_A_319_47#_c_596_n D 0.0232562f $X=2.47 $Y=1.86 $X2=0 $Y2=0
cc_524 N_A_319_47#_c_610_n D 0.0231586f $X=3.33 $Y=1.967 $X2=0 $Y2=0
cc_525 N_A_319_47#_c_604_n D 0.0244785f $X=3.44 $Y=1.52 $X2=0 $Y2=0
cc_526 N_A_319_47#_c_600_n N_SCD_c_755_n 0.0337486f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_527 N_A_319_47#_c_610_n N_SCD_c_755_n 2.1101e-19 $X=3.33 $Y=1.967 $X2=0 $Y2=0
cc_528 N_A_319_47#_c_604_n N_SCD_c_755_n 0.0024954f $X=3.44 $Y=1.52 $X2=0 $Y2=0
cc_529 N_A_319_47#_c_600_n SCD 0.00210871f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_530 N_A_319_47#_c_604_n SCD 0.0204455f $X=3.44 $Y=1.52 $X2=0 $Y2=0
cc_531 N_A_319_47#_c_600_n N_SCD_c_753_n 0.020449f $X=3.42 $Y=1.77 $X2=0 $Y2=0
cc_532 N_A_319_47#_c_604_n N_SCD_c_753_n 2.66358e-19 $X=3.44 $Y=1.52 $X2=0 $Y2=0
cc_533 N_A_319_47#_c_595_n N_A_203_47#_c_809_n 0.00266292f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_534 N_A_319_47#_M1020_g N_A_203_47#_c_810_n 0.00141103f $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_535 N_A_319_47#_c_600_n N_A_203_47#_c_810_n 8.89048e-19 $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_536 N_A_319_47#_c_595_n N_A_203_47#_c_810_n 0.0181694f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_537 N_A_319_47#_c_604_n N_A_203_47#_c_810_n 0.00172689f $X=3.44 $Y=1.52 $X2=0
+ $Y2=0
cc_538 N_A_319_47#_c_597_n N_A_203_47#_c_810_n 0.00465031f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_539 N_A_319_47#_c_598_n N_A_203_47#_c_810_n 0.00829416f $X=2.55 $Y=1.04 $X2=0
+ $Y2=0
cc_540 N_A_319_47#_c_599_n N_A_203_47#_c_810_n 0.00662895f $X=2.55 $Y=1.04 $X2=0
+ $Y2=0
cc_541 N_A_319_47#_c_595_n N_A_203_47#_c_817_n 0.0981154f $X=1.62 $Y=1.86 $X2=0
+ $Y2=0
cc_542 N_A_319_47#_c_602_n N_A_203_47#_c_817_n 0.0273077f $X=1.725 $Y=2.175
+ $X2=0 $Y2=0
cc_543 N_A_319_47#_c_597_n N_A_203_47#_c_817_n 0.00751789f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_544 N_A_319_47#_c_605_n N_A_203_47#_c_817_n 0.0159784f $X=1.672 $Y=1.967
+ $X2=0 $Y2=0
cc_545 N_A_319_47#_c_608_n N_VPWR_M1012_d 0.00351251f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_546 N_A_319_47#_c_602_n N_VPWR_c_1454_n 0.0154733f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_547 N_A_319_47#_c_608_n N_VPWR_c_1454_n 0.0184987f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_548 N_A_319_47#_c_600_n N_VPWR_c_1462_n 0.00441747f $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_549 N_A_319_47#_c_608_n N_VPWR_c_1462_n 3.89445e-19 $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_550 N_A_319_47#_c_610_n N_VPWR_c_1462_n 0.00525224f $X=3.33 $Y=1.967 $X2=0
+ $Y2=0
cc_551 N_A_319_47#_c_615_n N_VPWR_c_1462_n 0.00269709f $X=2.47 $Y=1.967 $X2=0
+ $Y2=0
cc_552 N_A_319_47#_c_602_n N_VPWR_c_1473_n 0.0170259f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_553 N_A_319_47#_c_608_n N_VPWR_c_1473_n 0.00234063f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_554 N_A_319_47#_M1012_s N_VPWR_c_1452_n 0.0019314f $X=1.6 $Y=1.845 $X2=0
+ $Y2=0
cc_555 N_A_319_47#_c_600_n N_VPWR_c_1452_n 0.00617905f $X=3.42 $Y=1.77 $X2=0
+ $Y2=0
cc_556 N_A_319_47#_c_602_n N_VPWR_c_1452_n 0.00494372f $X=1.725 $Y=2.175 $X2=0
+ $Y2=0
cc_557 N_A_319_47#_c_608_n N_VPWR_c_1452_n 0.00311756f $X=2.385 $Y=1.967 $X2=0
+ $Y2=0
cc_558 N_A_319_47#_c_610_n N_VPWR_c_1452_n 0.00494869f $X=3.33 $Y=1.967 $X2=0
+ $Y2=0
cc_559 N_A_319_47#_c_615_n N_VPWR_c_1452_n 0.0020288f $X=2.47 $Y=1.967 $X2=0
+ $Y2=0
cc_560 N_A_319_47#_c_610_n A_504_369# 0.00716796f $X=3.33 $Y=1.967 $X2=-0.19
+ $Y2=-0.24
cc_561 N_A_319_47#_c_610_n N_A_608_369#_M1037_d 0.00417681f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_562 N_A_319_47#_c_600_n N_A_608_369#_c_1640_n 0.0114679f $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_563 N_A_319_47#_c_610_n N_A_608_369#_c_1640_n 0.0324509f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_564 N_A_319_47#_M1020_g N_A_608_369#_c_1652_n 4.9735e-19 $X=2.51 $Y=0.445
+ $X2=0 $Y2=0
cc_565 N_A_319_47#_c_600_n N_A_608_369#_c_1664_n 0.00370813f $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_566 N_A_319_47#_c_600_n N_A_608_369#_c_1637_n 5.85164e-19 $X=3.42 $Y=1.77
+ $X2=0 $Y2=0
cc_567 N_A_319_47#_c_610_n N_A_608_369#_c_1637_n 0.00601338f $X=3.33 $Y=1.967
+ $X2=0 $Y2=0
cc_568 N_A_319_47#_c_604_n N_A_608_369#_c_1637_n 0.0019322f $X=3.44 $Y=1.52
+ $X2=0 $Y2=0
cc_569 N_A_319_47#_M1020_g N_VGND_c_1838_n 0.00899047f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_570 N_A_319_47#_c_597_n N_VGND_c_1838_n 0.0108298f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_571 N_A_319_47#_c_597_n N_VGND_c_1846_n 0.0193961f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_572 N_A_319_47#_M1020_g N_VGND_c_1848_n 0.00365142f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_573 N_A_319_47#_c_597_n N_VGND_c_1859_n 0.00203921f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_574 N_A_319_47#_M1016_s N_VGND_c_1861_n 0.00186585f $X=1.595 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_A_319_47#_M1020_g N_VGND_c_1861_n 0.00420825f $X=2.51 $Y=0.445 $X2=0
+ $Y2=0
cc_576 N_A_319_47#_c_597_n N_VGND_c_1861_n 0.00613328f $X=1.74 $Y=0.36 $X2=0
+ $Y2=0
cc_577 N_D_M1002_g SCD 0.00549163f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_578 N_D_c_713_n N_A_203_47#_c_810_n 4.1316e-19 $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_579 N_D_M1002_g N_A_203_47#_c_810_n 0.00364714f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_580 D N_A_203_47#_c_810_n 0.00875808f $X=2.905 $Y=1.445 $X2=0 $Y2=0
cc_581 N_D_c_713_n N_VPWR_c_1454_n 0.00170479f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_582 N_D_c_713_n N_VPWR_c_1462_n 0.00455384f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_583 N_D_c_713_n N_VPWR_c_1452_n 0.00628186f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_584 N_D_c_713_n N_A_608_369#_c_1640_n 0.00796293f $X=2.95 $Y=1.77 $X2=0 $Y2=0
cc_585 N_D_M1002_g N_A_608_369#_c_1652_n 0.00299076f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_586 N_D_M1002_g N_VGND_c_1838_n 0.00163883f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_587 N_D_M1002_g N_VGND_c_1848_n 0.0042011f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_588 N_D_M1002_g N_VGND_c_1861_n 0.00596315f $X=3 $Y=0.445 $X2=0 $Y2=0
cc_589 N_SCD_M1029_g N_A_203_47#_c_810_n 0.00245337f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_590 SCD N_A_203_47#_c_810_n 0.00958434f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_591 N_SCD_c_753_n N_A_203_47#_c_810_n 0.00138804f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_592 N_SCD_c_755_n N_VPWR_c_1455_n 0.00627598f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_593 N_SCD_c_755_n N_VPWR_c_1462_n 0.00504444f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_594 N_SCD_c_755_n N_VPWR_c_1452_n 0.00784388f $X=3.935 $Y=1.77 $X2=0 $Y2=0
cc_595 N_SCD_c_755_n N_A_608_369#_c_1640_n 0.00520197f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_596 N_SCD_M1029_g N_A_608_369#_c_1652_n 0.00468836f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_597 N_SCD_c_755_n N_A_608_369#_c_1664_n 0.0072605f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_598 N_SCD_M1029_g N_A_608_369#_c_1629_n 0.00659485f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_599 N_SCD_c_755_n N_A_608_369#_c_1636_n 0.0108115f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_600 SCD N_A_608_369#_c_1636_n 0.0138435f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_601 N_SCD_c_753_n N_A_608_369#_c_1636_n 0.00199327f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_602 N_SCD_c_755_n N_A_608_369#_c_1637_n 0.00271587f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_603 SCD N_A_608_369#_c_1637_n 0.0118154f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_604 N_SCD_M1029_g N_A_608_369#_c_1630_n 0.00830957f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_605 SCD N_A_608_369#_c_1630_n 0.0137228f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_606 N_SCD_c_753_n N_A_608_369#_c_1630_n 0.00215057f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_607 N_SCD_M1029_g N_A_608_369#_c_1631_n 0.00228168f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_608 SCD N_A_608_369#_c_1631_n 0.0120393f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_609 N_SCD_M1029_g N_A_608_369#_c_1632_n 0.00233059f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_610 N_SCD_M1029_g N_A_608_369#_c_1633_n 0.00400866f $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_611 N_SCD_c_754_n N_A_608_369#_c_1633_n 0.00345986f $X=3.935 $Y=1.67 $X2=0
+ $Y2=0
cc_612 N_SCD_c_755_n N_A_608_369#_c_1633_n 0.00105043f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_613 SCD N_A_608_369#_c_1633_n 0.0231455f $X=3.82 $Y=1.105 $X2=0 $Y2=0
cc_614 N_SCD_c_753_n N_A_608_369#_c_1633_n 0.00629503f $X=3.97 $Y=1.355 $X2=0
+ $Y2=0
cc_615 N_SCD_M1029_g N_A_608_369#_c_1634_n 4.17422e-19 $X=3.91 $Y=0.445 $X2=0
+ $Y2=0
cc_616 N_SCD_c_755_n N_A_608_369#_c_1639_n 0.00289044f $X=3.935 $Y=1.77 $X2=0
+ $Y2=0
cc_617 N_SCD_M1029_g N_VGND_c_1839_n 0.0104318f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_618 N_SCD_M1029_g N_VGND_c_1848_n 0.00404961f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_619 N_SCD_M1029_g N_VGND_c_1861_n 0.00679524f $X=3.91 $Y=0.445 $X2=0 $Y2=0
cc_620 N_A_203_47#_c_808_n N_A_1189_183#_M1032_d 9.85811e-19 $X=7.575 $Y=0.87
+ $X2=-0.19 $Y2=-0.24
cc_621 N_A_203_47#_c_812_n N_A_1189_183#_M1032_d 0.00132248f $X=7.31 $Y=0.805
+ $X2=-0.19 $Y2=-0.24
cc_622 N_A_203_47#_c_813_n N_A_1189_183#_M1032_d 8.90023e-19 $X=7.115 $Y=0.805
+ $X2=-0.19 $Y2=-0.24
cc_623 N_A_203_47#_c_804_n N_A_1189_183#_M1007_g 0.0116191f $X=5.56 $Y=0.705
+ $X2=0 $Y2=0
cc_624 N_A_203_47#_c_813_n N_A_1189_183#_M1007_g 7.75003e-19 $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_625 N_A_203_47#_c_813_n N_A_1189_183#_c_1011_n 0.0340036f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_626 N_A_203_47#_c_812_n N_A_1189_183#_c_1040_n 0.00269614f $X=7.31 $Y=0.805
+ $X2=0 $Y2=0
cc_627 N_A_203_47#_c_808_n N_A_1189_183#_c_1041_n 0.00684931f $X=7.575 $Y=0.87
+ $X2=0 $Y2=0
cc_628 N_A_203_47#_c_812_n N_A_1189_183#_c_1041_n 0.00281358f $X=7.31 $Y=0.805
+ $X2=0 $Y2=0
cc_629 N_A_203_47#_c_813_n N_A_1189_183#_c_1041_n 0.00335015f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_630 N_A_203_47#_c_807_n N_A_1189_183#_c_1012_n 0.00106902f $X=7.67 $Y=1.575
+ $X2=0 $Y2=0
cc_631 N_A_203_47#_c_808_n N_A_1189_183#_c_1012_n 0.0196063f $X=7.575 $Y=0.87
+ $X2=0 $Y2=0
cc_632 N_A_203_47#_c_812_n N_A_1189_183#_c_1012_n 4.81588e-19 $X=7.31 $Y=0.805
+ $X2=0 $Y2=0
cc_633 N_A_203_47#_c_813_n N_A_1189_183#_c_1012_n 0.0215929f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_634 N_A_203_47#_c_816_n N_A_1189_183#_c_1012_n 5.8166e-19 $X=7.53 $Y=0.87
+ $X2=0 $Y2=0
cc_635 N_A_203_47#_c_807_n N_A_1189_183#_c_1013_n 0.00592824f $X=7.67 $Y=1.575
+ $X2=0 $Y2=0
cc_636 N_A_203_47#_c_813_n N_A_1189_183#_c_1014_n 0.00314354f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_637 N_A_203_47#_c_815_n N_A_1189_183#_c_1014_n 0.0158555f $X=5.56 $Y=0.87
+ $X2=0 $Y2=0
cc_638 N_A_203_47#_c_805_n N_A_1011_47#_c_1108_n 0.00964531f $X=7.385 $Y=0.705
+ $X2=0 $Y2=0
cc_639 N_A_203_47#_c_808_n N_A_1011_47#_c_1108_n 0.00103154f $X=7.575 $Y=0.87
+ $X2=0 $Y2=0
cc_640 N_A_203_47#_c_807_n N_A_1011_47#_c_1109_n 3.2664e-19 $X=7.67 $Y=1.575
+ $X2=0 $Y2=0
cc_641 N_A_203_47#_c_816_n N_A_1011_47#_c_1109_n 0.00964531f $X=7.53 $Y=0.87
+ $X2=0 $Y2=0
cc_642 N_A_203_47#_c_818_n N_A_1011_47#_c_1131_n 0.00454283f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_643 N_A_203_47#_c_806_n N_A_1011_47#_c_1131_n 0.00454699f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_644 N_A_203_47#_c_804_n N_A_1011_47#_c_1135_n 0.00861823f $X=5.56 $Y=0.705
+ $X2=0 $Y2=0
cc_645 N_A_203_47#_c_811_n N_A_1011_47#_c_1135_n 0.0026338f $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_646 N_A_203_47#_c_813_n N_A_1011_47#_c_1135_n 0.00539305f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_647 N_A_203_47#_c_814_n N_A_1011_47#_c_1135_n 0.0239627f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_648 N_A_203_47#_c_815_n N_A_1011_47#_c_1135_n 0.00330834f $X=5.56 $Y=0.87
+ $X2=0 $Y2=0
cc_649 N_A_203_47#_c_804_n N_A_1011_47#_c_1112_n 0.00670209f $X=5.56 $Y=0.705
+ $X2=0 $Y2=0
cc_650 N_A_203_47#_c_806_n N_A_1011_47#_c_1112_n 0.00747938f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_651 N_A_203_47#_c_811_n N_A_1011_47#_c_1112_n 0.00103647f $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_652 N_A_203_47#_c_813_n N_A_1011_47#_c_1112_n 0.0189576f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_653 N_A_203_47#_c_814_n N_A_1011_47#_c_1112_n 0.0218614f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_654 N_A_203_47#_c_806_n N_A_1011_47#_c_1113_n 0.00886537f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_655 N_A_203_47#_c_813_n N_A_1011_47#_c_1113_n 0.00729071f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_656 N_A_203_47#_c_813_n N_A_1011_47#_c_1114_n 0.00196802f $X=7.115 $Y=0.805
+ $X2=0 $Y2=0
cc_657 N_A_203_47#_c_819_n N_A_1667_315#_c_1233_n 0.0249256f $X=7.75 $Y=1.99
+ $X2=0 $Y2=0
cc_658 N_A_203_47#_c_819_n N_A_1474_413#_c_1375_n 0.0143397f $X=7.75 $Y=1.99
+ $X2=0 $Y2=0
cc_659 N_A_203_47#_c_822_n N_A_1474_413#_c_1375_n 0.0153945f $X=7.81 $Y=1.74
+ $X2=0 $Y2=0
cc_660 N_A_203_47#_c_805_n N_A_1474_413#_c_1379_n 0.00196231f $X=7.385 $Y=0.705
+ $X2=0 $Y2=0
cc_661 N_A_203_47#_c_808_n N_A_1474_413#_c_1379_n 0.0153898f $X=7.575 $Y=0.87
+ $X2=0 $Y2=0
cc_662 N_A_203_47#_c_816_n N_A_1474_413#_c_1379_n 8.58658e-19 $X=7.53 $Y=0.87
+ $X2=0 $Y2=0
cc_663 N_A_203_47#_c_819_n N_A_1474_413#_c_1372_n 0.00714563f $X=7.75 $Y=1.99
+ $X2=0 $Y2=0
cc_664 N_A_203_47#_c_807_n N_A_1474_413#_c_1372_n 0.00712777f $X=7.67 $Y=1.575
+ $X2=0 $Y2=0
cc_665 N_A_203_47#_c_822_n N_A_1474_413#_c_1372_n 0.0208221f $X=7.81 $Y=1.74
+ $X2=0 $Y2=0
cc_666 N_A_203_47#_c_819_n N_A_1474_413#_c_1367_n 0.00102186f $X=7.75 $Y=1.99
+ $X2=0 $Y2=0
cc_667 N_A_203_47#_c_807_n N_A_1474_413#_c_1367_n 0.0226171f $X=7.67 $Y=1.575
+ $X2=0 $Y2=0
cc_668 N_A_203_47#_c_805_n N_A_1474_413#_c_1368_n 8.84292e-19 $X=7.385 $Y=0.705
+ $X2=0 $Y2=0
cc_669 N_A_203_47#_c_808_n N_A_1474_413#_c_1368_n 0.0214311f $X=7.575 $Y=0.87
+ $X2=0 $Y2=0
cc_670 N_A_203_47#_c_812_n N_A_1474_413#_c_1368_n 0.00119523f $X=7.31 $Y=0.805
+ $X2=0 $Y2=0
cc_671 N_A_203_47#_c_816_n N_A_1474_413#_c_1368_n 3.55894e-19 $X=7.53 $Y=0.87
+ $X2=0 $Y2=0
cc_672 N_A_203_47#_c_817_n N_VPWR_c_1453_n 0.0107869f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_673 N_A_203_47#_c_817_n N_VPWR_c_1454_n 5.70469e-19 $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_674 N_A_203_47#_c_818_n N_VPWR_c_1455_n 0.00261116f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_675 N_A_203_47#_c_818_n N_VPWR_c_1464_n 0.00659238f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_676 N_A_203_47#_c_819_n N_VPWR_c_1466_n 0.00460277f $X=7.75 $Y=1.99 $X2=0
+ $Y2=0
cc_677 N_A_203_47#_c_817_n N_VPWR_c_1473_n 0.0163465f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_678 N_A_203_47#_c_818_n N_VPWR_c_1452_n 0.00864761f $X=5 $Y=1.99 $X2=0 $Y2=0
cc_679 N_A_203_47#_c_819_n N_VPWR_c_1452_n 0.00672622f $X=7.75 $Y=1.99 $X2=0
+ $Y2=0
cc_680 N_A_203_47#_c_806_n N_VPWR_c_1452_n 0.00196481f $X=4.99 $Y=1.74 $X2=0
+ $Y2=0
cc_681 N_A_203_47#_c_817_n N_VPWR_c_1452_n 0.00418267f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_682 N_A_203_47#_c_810_n N_A_608_369#_c_1652_n 0.00642978f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_683 N_A_203_47#_c_810_n N_A_608_369#_c_1630_n 0.0286775f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_684 N_A_203_47#_c_810_n N_A_608_369#_c_1631_n 0.00791492f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_685 N_A_203_47#_c_818_n N_A_608_369#_c_1633_n 0.00543259f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_686 N_A_203_47#_c_806_n N_A_608_369#_c_1633_n 0.0594075f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_687 N_A_203_47#_c_810_n N_A_608_369#_c_1633_n 0.0123751f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_688 N_A_203_47#_c_814_n N_A_608_369#_c_1633_n 0.0127869f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_689 N_A_203_47#_c_810_n N_A_608_369#_c_1634_n 0.00506513f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_690 N_A_203_47#_c_814_n N_A_608_369#_c_1634_n 6.01474e-19 $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_691 N_A_203_47#_c_810_n N_A_608_369#_c_1635_n 0.00562077f $X=5.045 $Y=0.805
+ $X2=0 $Y2=0
cc_692 N_A_203_47#_c_811_n N_A_608_369#_c_1635_n 9.47294e-19 $X=5.385 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_A_203_47#_c_814_n N_A_608_369#_c_1635_n 0.0121034f $X=5.45 $Y=0.87
+ $X2=0 $Y2=0
cc_694 N_A_203_47#_c_818_n N_A_608_369#_c_1639_n 0.0110623f $X=5 $Y=1.99 $X2=0
+ $Y2=0
cc_695 N_A_203_47#_c_806_n N_A_608_369#_c_1639_n 0.00558961f $X=4.99 $Y=1.74
+ $X2=0 $Y2=0
cc_696 N_A_203_47#_c_810_n N_VGND_c_1838_n 0.00117832f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_697 N_A_203_47#_c_810_n N_VGND_c_1839_n 8.73533e-19 $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_698 N_A_203_47#_c_813_n N_VGND_c_1840_n 0.00197442f $X=7.115 $Y=0.805 $X2=0
+ $Y2=0
cc_699 N_A_203_47#_c_809_n N_VGND_c_1846_n 4.93882e-19 $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_700 N_A_203_47#_c_817_n N_VGND_c_1846_n 0.0101403f $X=1.2 $Y=0.51 $X2=0 $Y2=0
cc_701 N_A_203_47#_c_804_n N_VGND_c_1850_n 0.0037981f $X=5.56 $Y=0.705 $X2=0
+ $Y2=0
cc_702 N_A_203_47#_c_811_n N_VGND_c_1850_n 4.34458e-19 $X=5.385 $Y=0.805 $X2=0
+ $Y2=0
cc_703 N_A_203_47#_c_814_n N_VGND_c_1850_n 0.00334975f $X=5.45 $Y=0.87 $X2=0
+ $Y2=0
cc_704 N_A_203_47#_c_805_n N_VGND_c_1857_n 0.00435108f $X=7.385 $Y=0.705 $X2=0
+ $Y2=0
cc_705 N_A_203_47#_c_808_n N_VGND_c_1857_n 0.00392786f $X=7.575 $Y=0.87 $X2=0
+ $Y2=0
cc_706 N_A_203_47#_c_812_n N_VGND_c_1857_n 6.4045e-19 $X=7.31 $Y=0.805 $X2=0
+ $Y2=0
cc_707 N_A_203_47#_c_816_n N_VGND_c_1857_n 0.00152809f $X=7.53 $Y=0.87 $X2=0
+ $Y2=0
cc_708 N_A_203_47#_c_817_n N_VGND_c_1859_n 0.00751197f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_709 N_A_203_47#_M1009_d N_VGND_c_1861_n 0.00503858f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_710 N_A_203_47#_c_804_n N_VGND_c_1861_n 0.00595796f $X=5.56 $Y=0.705 $X2=0
+ $Y2=0
cc_711 N_A_203_47#_c_805_n N_VGND_c_1861_n 0.00633417f $X=7.385 $Y=0.705 $X2=0
+ $Y2=0
cc_712 N_A_203_47#_c_808_n N_VGND_c_1861_n 0.00410232f $X=7.575 $Y=0.87 $X2=0
+ $Y2=0
cc_713 N_A_203_47#_c_809_n N_VGND_c_1861_n 0.0161544f $X=1.385 $Y=0.805 $X2=0
+ $Y2=0
cc_714 N_A_203_47#_c_810_n N_VGND_c_1861_n 0.169172f $X=5.045 $Y=0.805 $X2=0
+ $Y2=0
cc_715 N_A_203_47#_c_811_n N_VGND_c_1861_n 0.0202259f $X=5.385 $Y=0.805 $X2=0
+ $Y2=0
cc_716 N_A_203_47#_c_812_n N_VGND_c_1861_n 0.0199172f $X=7.31 $Y=0.805 $X2=0
+ $Y2=0
cc_717 N_A_203_47#_c_813_n N_VGND_c_1861_n 0.079659f $X=7.115 $Y=0.805 $X2=0
+ $Y2=0
cc_718 N_A_203_47#_c_814_n N_VGND_c_1861_n 0.00195657f $X=5.45 $Y=0.87 $X2=0
+ $Y2=0
cc_719 N_A_203_47#_c_816_n N_VGND_c_1861_n 0.00255999f $X=7.53 $Y=0.87 $X2=0
+ $Y2=0
cc_720 N_A_203_47#_c_817_n N_VGND_c_1861_n 0.00363393f $X=1.2 $Y=0.51 $X2=0
+ $Y2=0
cc_721 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1107_n 0.00684338f $X=6.925
+ $Y=2.135 $X2=0 $Y2=0
cc_722 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1115_n 0.00419555f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_723 N_A_1189_183#_c_1016_n N_A_1011_47#_c_1115_n 0.00719967f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_724 N_A_1189_183#_c_1026_n N_A_1011_47#_c_1115_n 0.00529276f $X=6.99 $Y=2.3
+ $X2=0 $Y2=0
cc_725 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1115_n 0.0113977f $X=6.925 $Y=2.135
+ $X2=0 $Y2=0
cc_726 N_A_1189_183#_M1007_g N_A_1011_47#_c_1108_n 0.0088205f $X=6.1 $Y=0.445
+ $X2=0 $Y2=0
cc_727 N_A_1189_183#_c_1040_n N_A_1011_47#_c_1108_n 0.00613927f $X=6.885
+ $Y=0.765 $X2=0 $Y2=0
cc_728 N_A_1189_183#_c_1059_p N_A_1011_47#_c_1108_n 0.006045f $X=6.995 $Y=0.45
+ $X2=0 $Y2=0
cc_729 N_A_1189_183#_c_1012_n N_A_1011_47#_c_1108_n 0.006666f $X=6.885 $Y=0.915
+ $X2=0 $Y2=0
cc_730 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1108_n 0.00413625f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_731 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1109_n 0.00513715f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_732 N_A_1189_183#_c_1011_n N_A_1011_47#_c_1109_n 0.0102886f $X=6.775 $Y=0.915
+ $X2=0 $Y2=0
cc_733 N_A_1189_183#_c_1012_n N_A_1011_47#_c_1109_n 0.00358011f $X=6.885
+ $Y=0.915 $X2=0 $Y2=0
cc_734 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1109_n 0.00421879f $X=6.925
+ $Y=2.135 $X2=0 $Y2=0
cc_735 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1109_n 0.00574663f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_736 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1110_n 0.0175118f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_737 N_A_1189_183#_c_1011_n N_A_1011_47#_c_1110_n 0.0033172f $X=6.775 $Y=0.915
+ $X2=0 $Y2=0
cc_738 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1110_n 0.00246562f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_739 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1111_n 0.00204756f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_740 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1111_n 0.0109999f $X=6.925 $Y=2.135
+ $X2=0 $Y2=0
cc_741 N_A_1189_183#_c_1016_n N_A_1011_47#_c_1131_n 0.0109992f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_742 N_A_1189_183#_M1007_g N_A_1011_47#_c_1135_n 0.00184156f $X=6.1 $Y=0.445
+ $X2=0 $Y2=0
cc_743 N_A_1189_183#_M1007_g N_A_1011_47#_c_1112_n 0.00554565f $X=6.1 $Y=0.445
+ $X2=0 $Y2=0
cc_744 N_A_1189_183#_c_1011_n N_A_1011_47#_c_1112_n 0.0222221f $X=6.775 $Y=0.915
+ $X2=0 $Y2=0
cc_745 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1112_n 0.00910555f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_746 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1118_n 0.00883472f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_747 N_A_1189_183#_c_1016_n N_A_1011_47#_c_1118_n 0.00968806f $X=6.045 $Y=1.99
+ $X2=0 $Y2=0
cc_748 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1118_n 0.00780656f $X=6.925
+ $Y=2.135 $X2=0 $Y2=0
cc_749 N_A_1189_183#_c_1009_n N_A_1011_47#_c_1113_n 0.0180066f $X=6.045 $Y=1.89
+ $X2=0 $Y2=0
cc_750 N_A_1189_183#_c_1011_n N_A_1011_47#_c_1113_n 0.0144711f $X=6.775 $Y=0.915
+ $X2=0 $Y2=0
cc_751 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1113_n 0.00281809f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_752 N_A_1189_183#_c_1011_n N_A_1011_47#_c_1114_n 0.0244869f $X=6.775 $Y=0.915
+ $X2=0 $Y2=0
cc_753 N_A_1189_183#_c_1013_n N_A_1011_47#_c_1114_n 0.02555f $X=6.925 $Y=2.135
+ $X2=0 $Y2=0
cc_754 N_A_1189_183#_c_1014_n N_A_1011_47#_c_1114_n 0.00217631f $X=6.1 $Y=0.93
+ $X2=0 $Y2=0
cc_755 N_A_1189_183#_c_1026_n N_A_1474_413#_c_1375_n 0.0110665f $X=6.99 $Y=2.3
+ $X2=0 $Y2=0
cc_756 N_A_1189_183#_c_1009_n N_VPWR_c_1456_n 3.85242e-19 $X=6.045 $Y=1.89 $X2=0
+ $Y2=0
cc_757 N_A_1189_183#_c_1016_n N_VPWR_c_1456_n 0.00532796f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_758 N_A_1189_183#_c_1013_n N_VPWR_c_1456_n 0.0451396f $X=6.925 $Y=2.135 $X2=0
+ $Y2=0
cc_759 N_A_1189_183#_c_1016_n N_VPWR_c_1464_n 0.00457093f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_760 N_A_1189_183#_c_1026_n N_VPWR_c_1466_n 0.0185094f $X=6.99 $Y=2.3 $X2=0
+ $Y2=0
cc_761 N_A_1189_183#_M1022_d N_VPWR_c_1452_n 0.00306139f $X=6.845 $Y=1.735 $X2=0
+ $Y2=0
cc_762 N_A_1189_183#_c_1016_n N_VPWR_c_1452_n 0.00678138f $X=6.045 $Y=1.99 $X2=0
+ $Y2=0
cc_763 N_A_1189_183#_c_1026_n N_VPWR_c_1452_n 0.00522915f $X=6.99 $Y=2.3 $X2=0
+ $Y2=0
cc_764 N_A_1189_183#_c_1011_n N_VGND_M1007_d 0.00408144f $X=6.775 $Y=0.915 $X2=0
+ $Y2=0
cc_765 N_A_1189_183#_M1007_g N_VGND_c_1840_n 0.00626852f $X=6.1 $Y=0.445 $X2=0
+ $Y2=0
cc_766 N_A_1189_183#_c_1011_n N_VGND_c_1840_n 0.0258458f $X=6.775 $Y=0.915 $X2=0
+ $Y2=0
cc_767 N_A_1189_183#_c_1014_n N_VGND_c_1840_n 0.00120654f $X=6.1 $Y=0.93 $X2=0
+ $Y2=0
cc_768 N_A_1189_183#_M1007_g N_VGND_c_1850_n 0.00585385f $X=6.1 $Y=0.445 $X2=0
+ $Y2=0
cc_769 N_A_1189_183#_c_1059_p N_VGND_c_1857_n 0.00738334f $X=6.995 $Y=0.45 $X2=0
+ $Y2=0
cc_770 N_A_1189_183#_c_1041_n N_VGND_c_1857_n 0.0100275f $X=7.12 $Y=0.45 $X2=0
+ $Y2=0
cc_771 N_A_1189_183#_M1032_d N_VGND_c_1861_n 0.00241064f $X=6.955 $Y=0.235 $X2=0
+ $Y2=0
cc_772 N_A_1189_183#_M1007_g N_VGND_c_1861_n 0.00683784f $X=6.1 $Y=0.445 $X2=0
+ $Y2=0
cc_773 N_A_1189_183#_c_1011_n N_VGND_c_1861_n 0.0085019f $X=6.775 $Y=0.915 $X2=0
+ $Y2=0
cc_774 N_A_1189_183#_c_1059_p N_VGND_c_1861_n 0.00343551f $X=6.995 $Y=0.45 $X2=0
+ $Y2=0
cc_775 N_A_1189_183#_c_1041_n N_VGND_c_1861_n 0.00428466f $X=7.12 $Y=0.45 $X2=0
+ $Y2=0
cc_776 N_A_1011_47#_c_1131_n N_VPWR_M1000_d 0.00249014f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_777 N_A_1011_47#_c_1118_n N_VPWR_M1000_d 0.00416039f $X=6.155 $Y=2.19 $X2=0
+ $Y2=0
cc_778 N_A_1011_47#_c_1115_n N_VPWR_c_1456_n 0.00502749f $X=6.755 $Y=1.66 $X2=0
+ $Y2=0
cc_779 N_A_1011_47#_c_1110_n N_VPWR_c_1456_n 9.61279e-19 $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_780 N_A_1011_47#_c_1131_n N_VPWR_c_1456_n 0.0138309f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_781 N_A_1011_47#_c_1118_n N_VPWR_c_1456_n 0.0257292f $X=6.155 $Y=2.19 $X2=0
+ $Y2=0
cc_782 N_A_1011_47#_c_1114_n N_VPWR_c_1456_n 0.00744785f $X=6.52 $Y=1.41 $X2=0
+ $Y2=0
cc_783 N_A_1011_47#_c_1131_n N_VPWR_c_1464_n 0.0416565f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_784 N_A_1011_47#_c_1115_n N_VPWR_c_1466_n 0.00597712f $X=6.755 $Y=1.66 $X2=0
+ $Y2=0
cc_785 N_A_1011_47#_M1024_d N_VPWR_c_1452_n 0.00230779f $X=5.09 $Y=2.065 $X2=0
+ $Y2=0
cc_786 N_A_1011_47#_c_1115_n N_VPWR_c_1452_n 0.00740372f $X=6.755 $Y=1.66 $X2=0
+ $Y2=0
cc_787 N_A_1011_47#_c_1131_n N_VPWR_c_1452_n 0.0185811f $X=6.045 $Y=2.275 $X2=0
+ $Y2=0
cc_788 N_A_1011_47#_c_1135_n N_A_608_369#_c_1634_n 0.0114634f $X=5.725 $Y=0.45
+ $X2=0 $Y2=0
cc_789 N_A_1011_47#_c_1131_n N_A_608_369#_c_1639_n 0.0102205f $X=6.045 $Y=2.275
+ $X2=0 $Y2=0
cc_790 N_A_1011_47#_c_1131_n A_1121_413# 0.00508444f $X=6.045 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_791 N_A_1011_47#_c_1108_n N_VGND_c_1840_n 0.00671184f $X=6.805 $Y=0.95 $X2=0
+ $Y2=0
cc_792 N_A_1011_47#_c_1135_n N_VGND_c_1850_n 0.0268875f $X=5.725 $Y=0.45 $X2=0
+ $Y2=0
cc_793 N_A_1011_47#_c_1108_n N_VGND_c_1857_n 0.0037962f $X=6.805 $Y=0.95 $X2=0
+ $Y2=0
cc_794 N_A_1011_47#_M1034_d N_VGND_c_1861_n 0.00299383f $X=5.055 $Y=0.235 $X2=0
+ $Y2=0
cc_795 N_A_1011_47#_c_1108_n N_VGND_c_1861_n 0.0062043f $X=6.805 $Y=0.95 $X2=0
+ $Y2=0
cc_796 N_A_1011_47#_c_1135_n N_VGND_c_1861_n 0.011449f $X=5.725 $Y=0.45 $X2=0
+ $Y2=0
cc_797 N_A_1011_47#_c_1135_n A_1127_47# 0.0055768f $X=5.725 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_798 N_A_1011_47#_c_1112_n A_1127_47# 0.00313175f $X=5.81 $Y=1.245 $X2=-0.19
+ $Y2=-0.24
cc_799 N_A_1667_315#_c_1233_n N_A_1474_413#_c_1369_n 0.00271108f $X=8.435
+ $Y=1.99 $X2=0 $Y2=0
cc_800 N_A_1667_315#_c_1235_n N_A_1474_413#_c_1369_n 0.0179885f $X=10.01 $Y=1.41
+ $X2=0 $Y2=0
cc_801 N_A_1667_315#_c_1247_p N_A_1474_413#_c_1369_n 0.00777604f $X=9.305
+ $Y=1.95 $X2=0 $Y2=0
cc_802 N_A_1667_315#_c_1240_n N_A_1474_413#_c_1369_n 0.00606276f $X=9.412
+ $Y=1.575 $X2=0 $Y2=0
cc_803 N_A_1667_315#_c_1249_p N_A_1474_413#_c_1369_n 0.00844052f $X=9.362
+ $Y=1.74 $X2=0 $Y2=0
cc_804 N_A_1667_315#_c_1225_n N_A_1474_413#_c_1363_n 0.0217187f $X=9.985
+ $Y=0.995 $X2=0 $Y2=0
cc_805 N_A_1667_315#_c_1229_n N_A_1474_413#_c_1363_n 0.00463572f $X=9.41
+ $Y=1.075 $X2=0 $Y2=0
cc_806 N_A_1667_315#_c_1231_n N_A_1474_413#_c_1363_n 0.00596988f $X=9.305
+ $Y=0.385 $X2=0 $Y2=0
cc_807 N_A_1667_315#_M1005_g N_A_1474_413#_c_1364_n 0.0121169f $X=8.525 $Y=0.445
+ $X2=0 $Y2=0
cc_808 N_A_1667_315#_c_1239_n N_A_1474_413#_c_1364_n 0.00734699f $X=9.22 $Y=1.74
+ $X2=0 $Y2=0
cc_809 N_A_1667_315#_c_1229_n N_A_1474_413#_c_1364_n 0.00475015f $X=9.41
+ $Y=1.075 $X2=0 $Y2=0
cc_810 N_A_1667_315#_c_1231_n N_A_1474_413#_c_1364_n 0.00747686f $X=9.305
+ $Y=0.385 $X2=0 $Y2=0
cc_811 N_A_1667_315#_c_1249_p N_A_1474_413#_c_1364_n 0.00407845f $X=9.362
+ $Y=1.74 $X2=0 $Y2=0
cc_812 N_A_1667_315#_c_1258_p N_A_1474_413#_c_1364_n 0.00932867f $X=9.412 $Y=1.2
+ $X2=0 $Y2=0
cc_813 N_A_1667_315#_c_1229_n N_A_1474_413#_c_1365_n 0.00282378f $X=9.41
+ $Y=1.075 $X2=0 $Y2=0
cc_814 N_A_1667_315#_c_1240_n N_A_1474_413#_c_1365_n 0.00342329f $X=9.412
+ $Y=1.575 $X2=0 $Y2=0
cc_815 N_A_1667_315#_c_1230_n N_A_1474_413#_c_1365_n 0.0183287f $X=11.215
+ $Y=1.16 $X2=0 $Y2=0
cc_816 N_A_1667_315#_c_1258_p N_A_1474_413#_c_1365_n 0.00178975f $X=9.412 $Y=1.2
+ $X2=0 $Y2=0
cc_817 N_A_1667_315#_c_1232_n N_A_1474_413#_c_1365_n 0.0217187f $X=11.43
+ $Y=1.202 $X2=0 $Y2=0
cc_818 N_A_1667_315#_M1005_g N_A_1474_413#_c_1379_n 0.0011727f $X=8.525 $Y=0.445
+ $X2=0 $Y2=0
cc_819 N_A_1667_315#_c_1233_n N_A_1474_413#_c_1372_n 0.00953255f $X=8.435
+ $Y=1.99 $X2=0 $Y2=0
cc_820 N_A_1667_315#_c_1239_n N_A_1474_413#_c_1372_n 0.0215608f $X=9.22 $Y=1.74
+ $X2=0 $Y2=0
cc_821 N_A_1667_315#_c_1233_n N_A_1474_413#_c_1366_n 0.00844924f $X=8.435
+ $Y=1.99 $X2=0 $Y2=0
cc_822 N_A_1667_315#_M1005_g N_A_1474_413#_c_1366_n 0.0204137f $X=8.525 $Y=0.445
+ $X2=0 $Y2=0
cc_823 N_A_1667_315#_c_1239_n N_A_1474_413#_c_1366_n 0.0358014f $X=9.22 $Y=1.74
+ $X2=0 $Y2=0
cc_824 N_A_1667_315#_c_1229_n N_A_1474_413#_c_1366_n 0.00600727f $X=9.41
+ $Y=1.075 $X2=0 $Y2=0
cc_825 N_A_1667_315#_c_1231_n N_A_1474_413#_c_1366_n 7.42989e-19 $X=9.305
+ $Y=0.385 $X2=0 $Y2=0
cc_826 N_A_1667_315#_c_1258_p N_A_1474_413#_c_1366_n 0.0210781f $X=9.412 $Y=1.2
+ $X2=0 $Y2=0
cc_827 N_A_1667_315#_M1005_g N_A_1474_413#_c_1367_n 0.00886819f $X=8.525
+ $Y=0.445 $X2=0 $Y2=0
cc_828 N_A_1667_315#_M1005_g N_A_1474_413#_c_1368_n 0.00817634f $X=8.525
+ $Y=0.445 $X2=0 $Y2=0
cc_829 N_A_1667_315#_c_1233_n N_VPWR_c_1457_n 0.0165478f $X=8.435 $Y=1.99 $X2=0
+ $Y2=0
cc_830 N_A_1667_315#_c_1239_n N_VPWR_c_1457_n 0.018568f $X=9.22 $Y=1.74 $X2=0
+ $Y2=0
cc_831 N_A_1667_315#_c_1247_p N_VPWR_c_1457_n 0.0148444f $X=9.305 $Y=1.95 $X2=0
+ $Y2=0
cc_832 N_A_1667_315#_c_1235_n N_VPWR_c_1458_n 0.00699265f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_833 N_A_1667_315#_c_1247_p N_VPWR_c_1458_n 0.0375787f $X=9.305 $Y=1.95 $X2=0
+ $Y2=0
cc_834 N_A_1667_315#_c_1230_n N_VPWR_c_1458_n 0.00949052f $X=11.215 $Y=1.16
+ $X2=0 $Y2=0
cc_835 N_A_1667_315#_c_1249_p N_VPWR_c_1458_n 0.0206045f $X=9.362 $Y=1.74 $X2=0
+ $Y2=0
cc_836 N_A_1667_315#_c_1236_n N_VPWR_c_1459_n 0.00627841f $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_837 N_A_1667_315#_c_1237_n N_VPWR_c_1459_n 0.00591423f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_838 N_A_1667_315#_c_1238_n N_VPWR_c_1461_n 0.00797955f $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_839 N_A_1667_315#_c_1233_n N_VPWR_c_1466_n 0.00742119f $X=8.435 $Y=1.99 $X2=0
+ $Y2=0
cc_840 N_A_1667_315#_c_1247_p N_VPWR_c_1468_n 0.0166993f $X=9.305 $Y=1.95 $X2=0
+ $Y2=0
cc_841 N_A_1667_315#_c_1235_n N_VPWR_c_1470_n 0.00604256f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_842 N_A_1667_315#_c_1236_n N_VPWR_c_1470_n 0.00675419f $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_843 N_A_1667_315#_c_1237_n N_VPWR_c_1474_n 0.00604256f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_844 N_A_1667_315#_c_1238_n N_VPWR_c_1474_n 0.00675419f $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_845 N_A_1667_315#_M1030_s N_VPWR_c_1452_n 0.00242267f $X=9.18 $Y=1.485 $X2=0
+ $Y2=0
cc_846 N_A_1667_315#_c_1233_n N_VPWR_c_1452_n 0.0157102f $X=8.435 $Y=1.99 $X2=0
+ $Y2=0
cc_847 N_A_1667_315#_c_1235_n N_VPWR_c_1452_n 0.0101148f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_848 N_A_1667_315#_c_1236_n N_VPWR_c_1452_n 0.0118986f $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_849 N_A_1667_315#_c_1237_n N_VPWR_c_1452_n 0.0100363f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_850 N_A_1667_315#_c_1238_n N_VPWR_c_1452_n 0.0127906f $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_851 N_A_1667_315#_c_1239_n N_VPWR_c_1452_n 0.0145324f $X=9.22 $Y=1.74 $X2=0
+ $Y2=0
cc_852 N_A_1667_315#_c_1247_p N_VPWR_c_1452_n 0.0105267f $X=9.305 $Y=1.95 $X2=0
+ $Y2=0
cc_853 N_A_1667_315#_c_1225_n N_Q_c_1759_n 0.00506154f $X=9.985 $Y=0.995 $X2=0
+ $Y2=0
cc_854 N_A_1667_315#_c_1226_n N_Q_c_1759_n 0.00656316f $X=10.455 $Y=0.995 $X2=0
+ $Y2=0
cc_855 N_A_1667_315#_c_1227_n N_Q_c_1759_n 5.47459e-19 $X=10.935 $Y=0.995 $X2=0
+ $Y2=0
cc_856 N_A_1667_315#_c_1231_n N_Q_c_1759_n 0.00118849f $X=9.305 $Y=0.385 $X2=0
+ $Y2=0
cc_857 N_A_1667_315#_c_1235_n N_Q_c_1763_n 0.00428632f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_858 N_A_1667_315#_c_1236_n N_Q_c_1763_n 5.87864e-19 $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_859 N_A_1667_315#_c_1240_n N_Q_c_1763_n 0.00211109f $X=9.412 $Y=1.575 $X2=0
+ $Y2=0
cc_860 N_A_1667_315#_c_1230_n N_Q_c_1763_n 0.0242189f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_861 N_A_1667_315#_c_1249_p N_Q_c_1763_n 0.00167158f $X=9.362 $Y=1.74 $X2=0
+ $Y2=0
cc_862 N_A_1667_315#_c_1232_n N_Q_c_1763_n 0.00646999f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_863 N_A_1667_315#_c_1235_n N_Q_c_1769_n 0.0108367f $X=10.01 $Y=1.41 $X2=0
+ $Y2=0
cc_864 N_A_1667_315#_c_1236_n N_Q_c_1769_n 0.00992124f $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_865 N_A_1667_315#_c_1237_n N_Q_c_1769_n 6.04888e-19 $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_866 N_A_1667_315#_c_1226_n N_Q_c_1752_n 0.00885266f $X=10.455 $Y=0.995 $X2=0
+ $Y2=0
cc_867 N_A_1667_315#_c_1227_n N_Q_c_1752_n 0.00885266f $X=10.935 $Y=0.995 $X2=0
+ $Y2=0
cc_868 N_A_1667_315#_c_1230_n N_Q_c_1752_n 0.0409838f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_869 N_A_1667_315#_c_1232_n N_Q_c_1752_n 0.00369708f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_870 N_A_1667_315#_c_1225_n N_Q_c_1753_n 0.00369706f $X=9.985 $Y=0.995 $X2=0
+ $Y2=0
cc_871 N_A_1667_315#_c_1226_n N_Q_c_1753_n 0.0011376f $X=10.455 $Y=0.995 $X2=0
+ $Y2=0
cc_872 N_A_1667_315#_c_1230_n N_Q_c_1753_n 0.0308573f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_873 N_A_1667_315#_c_1231_n N_Q_c_1753_n 0.0052297f $X=9.305 $Y=0.385 $X2=0
+ $Y2=0
cc_874 N_A_1667_315#_c_1232_n N_Q_c_1753_n 0.00357417f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_875 N_A_1667_315#_c_1236_n N_Q_c_1781_n 0.0139158f $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_876 N_A_1667_315#_c_1237_n N_Q_c_1781_n 0.0102085f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_877 N_A_1667_315#_c_1230_n N_Q_c_1781_n 0.0347278f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_878 N_A_1667_315#_c_1232_n N_Q_c_1781_n 0.00653102f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_879 N_A_1667_315#_c_1226_n N_Q_c_1785_n 5.26331e-19 $X=10.455 $Y=0.995 $X2=0
+ $Y2=0
cc_880 N_A_1667_315#_c_1227_n N_Q_c_1785_n 0.00619901f $X=10.935 $Y=0.995 $X2=0
+ $Y2=0
cc_881 N_A_1667_315#_c_1236_n N_Q_c_1787_n 6.24109e-19 $X=10.48 $Y=1.41 $X2=0
+ $Y2=0
cc_882 N_A_1667_315#_c_1237_n N_Q_c_1787_n 0.0122088f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_883 N_A_1667_315#_c_1238_n N_Q_c_1787_n 0.0144343f $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_884 N_A_1667_315#_c_1228_n N_Q_c_1754_n 0.0138585f $X=11.455 $Y=0.995 $X2=0
+ $Y2=0
cc_885 N_A_1667_315#_c_1230_n N_Q_c_1754_n 0.00143455f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_886 N_A_1667_315#_c_1238_n N_Q_c_1757_n 0.0170109f $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_887 N_A_1667_315#_c_1230_n N_Q_c_1757_n 0.00130203f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_888 N_A_1667_315#_c_1227_n N_Q_c_1755_n 0.00116689f $X=10.935 $Y=0.995 $X2=0
+ $Y2=0
cc_889 N_A_1667_315#_c_1230_n N_Q_c_1755_n 0.0309896f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_890 N_A_1667_315#_c_1232_n N_Q_c_1755_n 0.00485066f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_891 N_A_1667_315#_c_1237_n N_Q_c_1797_n 0.00213487f $X=10.96 $Y=1.41 $X2=0
+ $Y2=0
cc_892 N_A_1667_315#_c_1238_n N_Q_c_1797_n 5.87864e-19 $X=11.43 $Y=1.41 $X2=0
+ $Y2=0
cc_893 N_A_1667_315#_c_1230_n N_Q_c_1797_n 0.0242189f $X=11.215 $Y=1.16 $X2=0
+ $Y2=0
cc_894 N_A_1667_315#_c_1232_n N_Q_c_1797_n 0.00627489f $X=11.43 $Y=1.202 $X2=0
+ $Y2=0
cc_895 N_A_1667_315#_c_1238_n Q 0.0036336f $X=11.43 $Y=1.41 $X2=0 $Y2=0
cc_896 N_A_1667_315#_c_1228_n Q 0.0197784f $X=11.455 $Y=0.995 $X2=0 $Y2=0
cc_897 N_A_1667_315#_c_1230_n Q 0.0206595f $X=11.215 $Y=1.16 $X2=0 $Y2=0
cc_898 N_A_1667_315#_M1005_g N_VGND_c_1841_n 0.0217281f $X=8.525 $Y=0.445 $X2=0
+ $Y2=0
cc_899 N_A_1667_315#_c_1231_n N_VGND_c_1841_n 0.0189502f $X=9.305 $Y=0.385 $X2=0
+ $Y2=0
cc_900 N_A_1667_315#_c_1225_n N_VGND_c_1842_n 0.00309623f $X=9.985 $Y=0.995
+ $X2=0 $Y2=0
cc_901 N_A_1667_315#_c_1230_n N_VGND_c_1842_n 0.00771963f $X=11.215 $Y=1.16
+ $X2=0 $Y2=0
cc_902 N_A_1667_315#_c_1226_n N_VGND_c_1843_n 0.00456672f $X=10.455 $Y=0.995
+ $X2=0 $Y2=0
cc_903 N_A_1667_315#_c_1227_n N_VGND_c_1843_n 0.00277568f $X=10.935 $Y=0.995
+ $X2=0 $Y2=0
cc_904 N_A_1667_315#_c_1228_n N_VGND_c_1845_n 0.00438629f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_905 N_A_1667_315#_c_1231_n N_VGND_c_1852_n 0.0178335f $X=9.305 $Y=0.385 $X2=0
+ $Y2=0
cc_906 N_A_1667_315#_c_1225_n N_VGND_c_1854_n 0.00543342f $X=9.985 $Y=0.995
+ $X2=0 $Y2=0
cc_907 N_A_1667_315#_c_1226_n N_VGND_c_1854_n 0.00426399f $X=10.455 $Y=0.995
+ $X2=0 $Y2=0
cc_908 N_A_1667_315#_c_1227_n N_VGND_c_1858_n 0.00426399f $X=10.935 $Y=0.995
+ $X2=0 $Y2=0
cc_909 N_A_1667_315#_c_1228_n N_VGND_c_1858_n 0.00439206f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_910 N_A_1667_315#_M1019_s N_VGND_c_1861_n 0.00253533f $X=9.18 $Y=0.235 $X2=0
+ $Y2=0
cc_911 N_A_1667_315#_M1005_g N_VGND_c_1861_n 9.61436e-19 $X=8.525 $Y=0.445 $X2=0
+ $Y2=0
cc_912 N_A_1667_315#_c_1225_n N_VGND_c_1861_n 0.00973629f $X=9.985 $Y=0.995
+ $X2=0 $Y2=0
cc_913 N_A_1667_315#_c_1226_n N_VGND_c_1861_n 0.00614062f $X=10.455 $Y=0.995
+ $X2=0 $Y2=0
cc_914 N_A_1667_315#_c_1227_n N_VGND_c_1861_n 0.0061332f $X=10.935 $Y=0.995
+ $X2=0 $Y2=0
cc_915 N_A_1667_315#_c_1228_n N_VGND_c_1861_n 0.00713978f $X=11.455 $Y=0.995
+ $X2=0 $Y2=0
cc_916 N_A_1667_315#_c_1231_n N_VGND_c_1861_n 0.013314f $X=9.305 $Y=0.385 $X2=0
+ $Y2=0
cc_917 N_A_1474_413#_c_1369_n N_VPWR_c_1457_n 0.00215411f $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_918 N_A_1474_413#_c_1369_n N_VPWR_c_1458_n 0.00616442f $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_919 N_A_1474_413#_c_1375_n N_VPWR_c_1466_n 0.0326463f $X=8.165 $Y=2.25 $X2=0
+ $Y2=0
cc_920 N_A_1474_413#_c_1369_n N_VPWR_c_1468_n 0.00621235f $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_921 N_A_1474_413#_M1003_d N_VPWR_c_1452_n 0.00237013f $X=7.37 $Y=2.065 $X2=0
+ $Y2=0
cc_922 N_A_1474_413#_c_1369_n N_VPWR_c_1452_n 0.0119363f $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_923 N_A_1474_413#_c_1375_n N_VPWR_c_1452_n 0.0316874f $X=8.165 $Y=2.25 $X2=0
+ $Y2=0
cc_924 N_A_1474_413#_c_1375_n A_1568_413# 0.0141044f $X=8.165 $Y=2.25 $X2=-0.19
+ $Y2=-0.24
cc_925 N_A_1474_413#_c_1372_n A_1568_413# 0.00197037f $X=8.25 $Y=2.165 $X2=-0.19
+ $Y2=-0.24
cc_926 N_A_1474_413#_c_1369_n N_Q_c_1763_n 3.18216e-19 $X=9.54 $Y=1.41 $X2=0
+ $Y2=0
cc_927 N_A_1474_413#_c_1363_n N_Q_c_1753_n 5.01468e-19 $X=9.565 $Y=0.995 $X2=0
+ $Y2=0
cc_928 N_A_1474_413#_c_1363_n N_VGND_c_1841_n 0.00252764f $X=9.565 $Y=0.995
+ $X2=0 $Y2=0
cc_929 N_A_1474_413#_c_1379_n N_VGND_c_1841_n 0.0107262f $X=7.985 $Y=0.45 $X2=0
+ $Y2=0
cc_930 N_A_1474_413#_c_1366_n N_VGND_c_1841_n 0.0179173f $X=9.065 $Y=1.16 $X2=0
+ $Y2=0
cc_931 N_A_1474_413#_c_1368_n N_VGND_c_1841_n 0.00460335f $X=8.16 $Y=0.995 $X2=0
+ $Y2=0
cc_932 N_A_1474_413#_c_1363_n N_VGND_c_1842_n 0.00309623f $X=9.565 $Y=0.995
+ $X2=0 $Y2=0
cc_933 N_A_1474_413#_c_1363_n N_VGND_c_1852_n 0.00572277f $X=9.565 $Y=0.995
+ $X2=0 $Y2=0
cc_934 N_A_1474_413#_c_1379_n N_VGND_c_1857_n 0.0223802f $X=7.985 $Y=0.45 $X2=0
+ $Y2=0
cc_935 N_A_1474_413#_M1014_d N_VGND_c_1861_n 0.00484466f $X=7.46 $Y=0.235 $X2=0
+ $Y2=0
cc_936 N_A_1474_413#_c_1363_n N_VGND_c_1861_n 0.0116721f $X=9.565 $Y=0.995 $X2=0
+ $Y2=0
cc_937 N_A_1474_413#_c_1379_n N_VGND_c_1861_n 0.0218104f $X=7.985 $Y=0.45 $X2=0
+ $Y2=0
cc_938 N_A_1474_413#_c_1379_n A_1625_47# 0.00202155f $X=7.985 $Y=0.45 $X2=-0.19
+ $Y2=-0.24
cc_939 N_A_1474_413#_c_1368_n A_1625_47# 0.00129936f $X=8.16 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_940 N_VPWR_c_1452_n A_504_369# 0.00301127f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_941 N_VPWR_c_1452_n N_A_608_369#_M1037_d 0.00192656f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_942 N_VPWR_c_1452_n N_A_608_369#_M1024_s 0.002768f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_943 N_VPWR_c_1454_n N_A_608_369#_c_1640_n 0.00527813f $X=2.195 $Y=2.33 $X2=0
+ $Y2=0
cc_944 N_VPWR_c_1455_n N_A_608_369#_c_1640_n 0.0109395f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_945 N_VPWR_c_1462_n N_A_608_369#_c_1640_n 0.0429697f $X=4.11 $Y=2.72 $X2=0
+ $Y2=0
cc_946 N_VPWR_c_1452_n N_A_608_369#_c_1640_n 0.0157065f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_947 N_VPWR_c_1455_n N_A_608_369#_c_1664_n 0.00457937f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_948 N_VPWR_M1028_d N_A_608_369#_c_1636_n 0.00399644f $X=4.025 $Y=1.845 $X2=0
+ $Y2=0
cc_949 N_VPWR_c_1455_n N_A_608_369#_c_1636_n 0.0119067f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_950 N_VPWR_c_1462_n N_A_608_369#_c_1636_n 0.00264158f $X=4.11 $Y=2.72 $X2=0
+ $Y2=0
cc_951 N_VPWR_c_1464_n N_A_608_369#_c_1636_n 0.00429797f $X=6.435 $Y=2.72 $X2=0
+ $Y2=0
cc_952 N_VPWR_c_1452_n N_A_608_369#_c_1636_n 0.00580702f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_953 N_VPWR_c_1455_n N_A_608_369#_c_1639_n 0.0144725f $X=4.195 $Y=2.33 $X2=0
+ $Y2=0
cc_954 N_VPWR_c_1464_n N_A_608_369#_c_1639_n 0.0140749f $X=6.435 $Y=2.72 $X2=0
+ $Y2=0
cc_955 N_VPWR_c_1452_n N_A_608_369#_c_1639_n 0.00421345f $X=11.73 $Y=2.72 $X2=0
+ $Y2=0
cc_956 N_VPWR_c_1452_n A_702_369# 0.00224063f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_957 N_VPWR_c_1452_n A_1121_413# 0.00241113f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_958 N_VPWR_c_1452_n A_1568_413# 0.00450219f $X=11.73 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_959 N_VPWR_c_1452_n N_Q_M1004_s 0.00237436f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_960 N_VPWR_c_1452_n N_Q_M1023_s 0.00237436f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_961 N_VPWR_c_1458_n N_Q_c_1763_n 0.0039299f $X=9.775 $Y=1.79 $X2=0 $Y2=0
cc_962 N_VPWR_c_1458_n N_Q_c_1769_n 0.0537133f $X=9.775 $Y=1.79 $X2=0 $Y2=0
cc_963 N_VPWR_c_1459_n N_Q_c_1769_n 0.0325368f $X=10.725 $Y=2.01 $X2=0 $Y2=0
cc_964 N_VPWR_c_1470_n N_Q_c_1769_n 0.0154447f $X=10.64 $Y=2.72 $X2=0 $Y2=0
cc_965 N_VPWR_c_1452_n N_Q_c_1769_n 0.0134778f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_966 N_VPWR_M1018_d N_Q_c_1781_n 0.00391612f $X=10.57 $Y=1.485 $X2=0 $Y2=0
cc_967 N_VPWR_c_1459_n N_Q_c_1781_n 0.0136682f $X=10.725 $Y=2.01 $X2=0 $Y2=0
cc_968 N_VPWR_c_1459_n N_Q_c_1787_n 0.0410603f $X=10.725 $Y=2.01 $X2=0 $Y2=0
cc_969 N_VPWR_c_1461_n N_Q_c_1787_n 0.0336646f $X=11.665 $Y=2.01 $X2=0 $Y2=0
cc_970 N_VPWR_c_1474_n N_Q_c_1787_n 0.0154447f $X=11.58 $Y=2.72 $X2=0 $Y2=0
cc_971 N_VPWR_c_1452_n N_Q_c_1787_n 0.0134778f $X=11.73 $Y=2.72 $X2=0 $Y2=0
cc_972 N_VPWR_M1025_d N_Q_c_1757_n 0.00619112f $X=11.52 $Y=1.485 $X2=0 $Y2=0
cc_973 N_VPWR_c_1461_n N_Q_c_1757_n 0.0151472f $X=11.665 $Y=2.01 $X2=0 $Y2=0
cc_974 N_A_608_369#_c_1640_n A_702_369# 0.0041021f $X=3.72 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_975 N_A_608_369#_c_1664_n A_702_369# 0.0027134f $X=3.805 $Y=2.245 $X2=-0.19
+ $Y2=-0.24
cc_976 N_A_608_369#_c_1637_n A_702_369# 0.00101879f $X=3.89 $Y=1.91 $X2=-0.19
+ $Y2=-0.24
cc_977 N_A_608_369#_c_1652_n N_VGND_c_1838_n 0.00460192f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_978 N_A_608_369#_c_1652_n N_VGND_c_1839_n 0.0110659f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_979 N_A_608_369#_c_1629_n N_VGND_c_1839_n 0.00463869f $X=3.81 $Y=0.695 $X2=0
+ $Y2=0
cc_980 N_A_608_369#_c_1630_n N_VGND_c_1839_n 0.0142693f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_981 N_A_608_369#_c_1634_n N_VGND_c_1839_n 0.00958988f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_982 N_A_608_369#_c_1652_n N_VGND_c_1848_n 0.0409414f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_983 N_A_608_369#_c_1630_n N_VGND_c_1848_n 0.00337254f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_984 N_A_608_369#_c_1630_n N_VGND_c_1850_n 0.00402378f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_985 N_A_608_369#_c_1634_n N_VGND_c_1850_n 0.012161f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_986 N_A_608_369#_M1002_d N_VGND_c_1861_n 0.00250516f $X=3.075 $Y=0.235 $X2=0
+ $Y2=0
cc_987 N_A_608_369#_M1034_s N_VGND_c_1861_n 0.00195217f $X=4.625 $Y=0.235 $X2=0
+ $Y2=0
cc_988 N_A_608_369#_c_1652_n N_VGND_c_1861_n 0.0135588f $X=3.725 $Y=0.36 $X2=0
+ $Y2=0
cc_989 N_A_608_369#_c_1630_n N_VGND_c_1861_n 0.00576196f $X=4.565 $Y=0.78 $X2=0
+ $Y2=0
cc_990 N_A_608_369#_c_1634_n N_VGND_c_1861_n 0.00544577f $X=4.75 $Y=0.45 $X2=0
+ $Y2=0
cc_991 N_A_608_369#_c_1652_n A_721_47# 0.00210886f $X=3.725 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_992 N_A_608_369#_c_1629_n A_721_47# 0.00225806f $X=3.81 $Y=0.695 $X2=-0.19
+ $Y2=-0.24
cc_993 N_Q_c_1752_n N_VGND_M1011_d 0.00270984f $X=10.98 $Y=0.82 $X2=0 $Y2=0
cc_994 N_Q_c_1754_n N_VGND_M1017_d 0.00337227f $X=11.55 $Y=0.82 $X2=0 $Y2=0
cc_995 N_Q_c_1759_n N_VGND_c_1843_n 0.0153813f $X=10.245 $Y=0.395 $X2=0 $Y2=0
cc_996 N_Q_c_1752_n N_VGND_c_1843_n 0.0127122f $X=10.98 $Y=0.82 $X2=0 $Y2=0
cc_997 N_Q_c_1754_n N_VGND_c_1844_n 0.00163214f $X=11.55 $Y=0.82 $X2=0 $Y2=0
cc_998 N_Q_c_1754_n N_VGND_c_1845_n 0.0140453f $X=11.55 $Y=0.82 $X2=0 $Y2=0
cc_999 N_Q_c_1759_n N_VGND_c_1854_n 0.0168847f $X=10.245 $Y=0.395 $X2=0 $Y2=0
cc_1000 N_Q_c_1752_n N_VGND_c_1854_n 0.00274274f $X=10.98 $Y=0.82 $X2=0 $Y2=0
cc_1001 N_Q_c_1752_n N_VGND_c_1858_n 0.00193763f $X=10.98 $Y=0.82 $X2=0 $Y2=0
cc_1002 N_Q_c_1785_n N_VGND_c_1858_n 0.0174926f $X=11.195 $Y=0.395 $X2=0 $Y2=0
cc_1003 N_Q_c_1754_n N_VGND_c_1858_n 0.00226277f $X=11.55 $Y=0.82 $X2=0 $Y2=0
cc_1004 N_Q_M1006_s N_VGND_c_1861_n 0.00259276f $X=10.06 $Y=0.235 $X2=0 $Y2=0
cc_1005 N_Q_M1015_s N_VGND_c_1861_n 0.00308722f $X=11.01 $Y=0.235 $X2=0 $Y2=0
cc_1006 N_Q_c_1759_n N_VGND_c_1861_n 0.0137257f $X=10.245 $Y=0.395 $X2=0 $Y2=0
cc_1007 N_Q_c_1752_n N_VGND_c_1861_n 0.00987236f $X=10.98 $Y=0.82 $X2=0 $Y2=0
cc_1008 N_Q_c_1785_n N_VGND_c_1861_n 0.0139324f $X=11.195 $Y=0.395 $X2=0 $Y2=0
cc_1009 N_Q_c_1754_n N_VGND_c_1861_n 0.00853011f $X=11.55 $Y=0.82 $X2=0 $Y2=0
cc_1010 N_VGND_c_1861_n A_517_47# 0.00293312f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1011 N_VGND_c_1861_n A_721_47# 0.00152414f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1012 N_VGND_c_1861_n A_1127_47# 0.00366632f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1013 N_VGND_c_1861_n A_1625_47# 0.0111093f $X=11.73 $Y=0 $X2=-0.19 $Y2=-0.24
