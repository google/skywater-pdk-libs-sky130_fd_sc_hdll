* NGSPICE file created from sky130_fd_sc_hdll__o21ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 VPWR B1 Y VPB phighvt w=700000u l=180000u
+  ad=6.515e+11p pd=5.03e+06u as=3.72e+11p ps=2.84e+06u
M1001 Y A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.3e+11p ps=2.46e+06u
M1002 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=3.8025e+11p pd=2.47e+06u as=3.77e+11p ps=3.76e+06u
M1004 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.535e+11p ps=2.08e+06u
M1005 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

