* File: sky130_fd_sc_hdll__and2_1.pxi.spice
* Created: Wed Sep  2 08:21:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2_1%A N_A_c_48_n N_A_c_49_n N_A_M1000_g N_A_M1005_g
+ N_A_c_50_n A N_A_c_47_n A A PM_SKY130_FD_SC_HDLL__AND2_1%A
x_PM_SKY130_FD_SC_HDLL__AND2_1%B N_B_M1003_g N_B_c_81_n N_B_c_82_n N_B_M1004_g B
+ N_B_c_80_n PM_SKY130_FD_SC_HDLL__AND2_1%B
x_PM_SKY130_FD_SC_HDLL__AND2_1%A_27_75# N_A_27_75#_M1005_s N_A_27_75#_M1000_d
+ N_A_27_75#_c_119_n N_A_27_75#_M1001_g N_A_27_75#_c_120_n N_A_27_75#_M1002_g
+ N_A_27_75#_c_121_n N_A_27_75#_c_122_n N_A_27_75#_c_123_n N_A_27_75#_c_126_n
+ N_A_27_75#_c_127_n N_A_27_75#_c_128_n N_A_27_75#_c_124_n N_A_27_75#_c_130_n
+ PM_SKY130_FD_SC_HDLL__AND2_1%A_27_75#
x_PM_SKY130_FD_SC_HDLL__AND2_1%VPWR N_VPWR_M1000_s N_VPWR_M1004_d N_VPWR_c_194_n
+ N_VPWR_c_195_n N_VPWR_c_196_n N_VPWR_c_197_n VPWR N_VPWR_c_198_n
+ N_VPWR_c_193_n N_VPWR_c_200_n PM_SKY130_FD_SC_HDLL__AND2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2_1%X N_X_M1001_d N_X_M1002_d N_X_c_225_n X X X X X X
+ N_X_c_222_n X PM_SKY130_FD_SC_HDLL__AND2_1%X
x_PM_SKY130_FD_SC_HDLL__AND2_1%VGND N_VGND_M1003_d N_VGND_c_244_n VGND
+ N_VGND_c_245_n N_VGND_c_246_n N_VGND_c_247_n N_VGND_c_248_n
+ PM_SKY130_FD_SC_HDLL__AND2_1%VGND
cc_1 VNB N_A_M1005_g 0.0275837f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_2 VNB A 0.0120843f $X=-0.19 $Y=-0.24 $X2=0.445 $Y2=1.105
cc_3 VNB N_A_c_47_n 0.0392204f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.16
cc_4 VNB N_B_M1003_g 0.0216209f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.78
cc_5 VNB B 0.00327428f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=1.325
cc_6 VNB N_B_c_80_n 0.0231255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_75#_c_119_n 0.0221896f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.585
cc_8 VNB N_A_27_75#_c_120_n 0.0231448f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=1.325
cc_9 VNB N_A_27_75#_c_121_n 0.0167456f $X=-0.19 $Y=-0.24 $X2=0.295 $Y2=1.16
cc_10 VNB N_A_27_75#_c_122_n 0.00771204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_75#_c_123_n 0.0102905f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_12 VNB N_A_27_75#_c_124_n 0.00423513f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=1.2
cc_13 VNB N_VPWR_c_193_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_14 VNB X 0.0377384f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=1.325
cc_15 VNB N_X_c_222_n 0.0152225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_244_n 0.00665189f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_17 VNB N_VGND_c_245_n 0.032298f $X=-0.19 $Y=-0.24 $X2=0.277 $Y2=1.325
cc_18 VNB N_VGND_c_246_n 0.0255308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_247_n 0.158319f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_20 VNB N_VGND_c_248_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_21 VPB N_A_c_48_n 0.0242463f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.68
cc_22 VPB N_A_c_49_n 0.0289472f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.78
cc_23 VPB N_A_c_50_n 0.0189912f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.325
cc_24 VPB A 0.001743f $X=-0.19 $Y=1.305 $X2=0.445 $Y2=1.105
cc_25 VPB N_A_c_47_n 0.00996509f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_26 VPB N_B_c_81_n 0.0207321f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_27 VPB N_B_c_82_n 0.0228578f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.585
cc_28 VPB B 5.68425e-19 $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.325
cc_29 VPB N_B_c_80_n 0.00419406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_27_75#_c_120_n 0.0321106f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.325
cc_31 VPB N_A_27_75#_c_126_n 0.00414045f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_32 VPB N_A_27_75#_c_127_n 0.0015776f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_75#_c_128_n 0.00550067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_75#_c_124_n 8.62065e-19 $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.2
cc_35 VPB N_A_27_75#_c_130_n 0.00171578f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.2
cc_36 VPB N_VPWR_c_194_n 0.0115481f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.585
cc_37 VPB N_VPWR_c_195_n 0.0305246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_196_n 0.0198843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_197_n 0.0101138f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_40 VPB N_VPWR_c_198_n 0.0260081f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_41 VPB N_VPWR_c_193_n 0.0575029f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_42 VPB N_VPWR_c_200_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.19
cc_43 VPB X 0.0257056f $X=-0.19 $Y=1.305 $X2=0.277 $Y2=1.325
cc_44 VPB X 0.0212237f $X=-0.19 $Y=1.305 $X2=0.295 $Y2=1.16
cc_45 N_A_M1005_g N_B_M1003_g 0.0183058f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_46 N_A_c_48_n N_B_c_81_n 0.0183058f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_47 N_A_c_50_n N_B_c_81_n 0.00124828f $X=0.277 $Y=1.325 $X2=0 $Y2=0
cc_48 N_A_c_49_n N_B_c_82_n 0.02956f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_49 A B 0.0171131f $X=0.445 $Y=1.105 $X2=0 $Y2=0
cc_50 N_A_c_47_n B 2.90198e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_51 A N_B_c_80_n 0.00100898f $X=0.445 $Y=1.105 $X2=0 $Y2=0
cc_52 N_A_c_47_n N_B_c_80_n 0.0183058f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_M1005_g N_A_27_75#_c_121_n 6.10868e-19 $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_54 N_A_M1005_g N_A_27_75#_c_122_n 0.0143388f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_55 A N_A_27_75#_c_122_n 0.0151799f $X=0.445 $Y=1.105 $X2=0 $Y2=0
cc_56 N_A_c_47_n N_A_27_75#_c_122_n 2.87475e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_57 A N_A_27_75#_c_123_n 0.0268484f $X=0.445 $Y=1.105 $X2=0 $Y2=0
cc_58 N_A_c_47_n N_A_27_75#_c_123_n 0.00844754f $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_c_49_n N_A_27_75#_c_126_n 0.00361973f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_60 N_A_c_48_n N_A_27_75#_c_128_n 0.00300726f $X=0.515 $Y=1.68 $X2=0 $Y2=0
cc_61 N_A_c_50_n N_A_27_75#_c_128_n 0.00928358f $X=0.277 $Y=1.325 $X2=0 $Y2=0
cc_62 A N_A_27_75#_c_128_n 0.00266042f $X=0.445 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_c_49_n N_VPWR_c_195_n 0.0052997f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_64 N_A_c_50_n N_VPWR_c_195_n 0.0158886f $X=0.277 $Y=1.325 $X2=0 $Y2=0
cc_65 N_A_c_47_n N_VPWR_c_195_n 9.93035e-19 $X=0.54 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A_c_49_n N_VPWR_c_196_n 0.00628791f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_67 N_A_c_49_n N_VPWR_c_193_n 0.00622823f $X=0.515 $Y=1.78 $X2=0 $Y2=0
cc_68 N_A_M1005_g N_VGND_c_245_n 0.0044865f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_69 N_A_M1005_g N_VGND_c_247_n 0.00541051f $X=0.54 $Y=0.585 $X2=0 $Y2=0
cc_70 N_B_M1003_g N_A_27_75#_c_119_n 0.0160918f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_71 N_B_c_81_n N_A_27_75#_c_120_n 0.0141895f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_72 N_B_c_82_n N_A_27_75#_c_120_n 0.00429099f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_73 B N_A_27_75#_c_120_n 7.73095e-19 $X=0.955 $Y=1.105 $X2=0 $Y2=0
cc_74 N_B_c_80_n N_A_27_75#_c_120_n 0.0184381f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_75 N_B_M1003_g N_A_27_75#_c_122_n 0.0133448f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_76 B N_A_27_75#_c_122_n 0.0255303f $X=0.955 $Y=1.105 $X2=0 $Y2=0
cc_77 N_B_c_80_n N_A_27_75#_c_122_n 0.00441634f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_78 N_B_c_82_n N_A_27_75#_c_126_n 0.0104432f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_79 N_B_c_81_n N_A_27_75#_c_127_n 0.00570157f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_80 N_B_c_82_n N_A_27_75#_c_127_n 0.00863235f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_81 B N_A_27_75#_c_127_n 0.0164878f $X=0.955 $Y=1.105 $X2=0 $Y2=0
cc_82 N_B_c_80_n N_A_27_75#_c_127_n 0.00254816f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_83 N_B_c_81_n N_A_27_75#_c_128_n 0.00207597f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_84 N_B_c_82_n N_A_27_75#_c_128_n 8.61603e-19 $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_85 B N_A_27_75#_c_128_n 0.00230715f $X=0.955 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B_M1003_g N_A_27_75#_c_124_n 0.00155172f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_87 B N_A_27_75#_c_124_n 0.0205328f $X=0.955 $Y=1.105 $X2=0 $Y2=0
cc_88 N_B_c_80_n N_A_27_75#_c_124_n 0.00249646f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_81_n N_A_27_75#_c_130_n 0.00317568f $X=0.985 $Y=1.68 $X2=0 $Y2=0
cc_90 N_B_c_82_n N_VPWR_c_196_n 0.00601158f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_91 N_B_c_82_n N_VPWR_c_197_n 0.00395776f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_92 N_B_c_82_n N_VPWR_c_193_n 0.00622823f $X=0.985 $Y=1.78 $X2=0 $Y2=0
cc_93 N_B_M1003_g N_VGND_c_244_n 0.00574637f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_94 N_B_M1003_g N_VGND_c_245_n 0.0044865f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_95 N_B_M1003_g N_VGND_c_247_n 0.00541051f $X=0.96 $Y=0.585 $X2=0 $Y2=0
cc_96 N_A_27_75#_c_127_n N_VPWR_M1004_d 0.00641453f $X=1.405 $Y=1.66 $X2=0 $Y2=0
cc_97 N_A_27_75#_c_126_n N_VPWR_c_195_n 0.00129362f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_98 N_A_27_75#_c_126_n N_VPWR_c_196_n 0.0101858f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_99 N_A_27_75#_c_120_n N_VPWR_c_197_n 0.00483431f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_27_75#_c_126_n N_VPWR_c_197_n 0.0148424f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_101 N_A_27_75#_c_127_n N_VPWR_c_197_n 0.0226396f $X=1.405 $Y=1.66 $X2=0 $Y2=0
cc_102 N_A_27_75#_c_120_n N_VPWR_c_198_n 0.00702461f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_27_75#_c_120_n N_VPWR_c_193_n 0.0149049f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_27_75#_c_126_n N_VPWR_c_193_n 0.0103957f $X=0.75 $Y=2.13 $X2=0 $Y2=0
cc_105 N_A_27_75#_c_119_n N_X_c_225_n 0.0120308f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_27_75#_c_120_n N_X_c_225_n 0.00170145f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_27_75#_c_124_n N_X_c_225_n 0.00574749f $X=1.49 $Y=1.325 $X2=0 $Y2=0
cc_108 N_A_27_75#_c_119_n X 0.0107224f $X=1.515 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_27_75#_c_120_n X 0.0218921f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_27_75#_c_127_n X 0.00932492f $X=1.405 $Y=1.66 $X2=0 $Y2=0
cc_111 N_A_27_75#_c_124_n X 0.0376283f $X=1.49 $Y=1.325 $X2=0 $Y2=0
cc_112 N_A_27_75#_c_130_n X 0.0125358f $X=1.49 $Y=1.575 $X2=0 $Y2=0
cc_113 N_A_27_75#_c_120_n X 0.0133542f $X=1.54 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_27_75#_c_122_n A_123_75# 0.00297727f $X=1.405 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_27_75#_c_122_n N_VGND_M1003_d 0.00373958f $X=1.405 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_27_75#_c_119_n N_VGND_c_244_n 0.00544651f $X=1.515 $Y=0.995 $X2=0
+ $Y2=0
cc_117 N_A_27_75#_c_121_n N_VGND_c_244_n 0.00297161f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_118 N_A_27_75#_c_122_n N_VGND_c_244_n 0.0195021f $X=1.405 $Y=0.81 $X2=0 $Y2=0
cc_119 N_A_27_75#_c_121_n N_VGND_c_245_n 0.0141462f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_120 N_A_27_75#_c_122_n N_VGND_c_245_n 0.00808217f $X=1.405 $Y=0.81 $X2=0
+ $Y2=0
cc_121 N_A_27_75#_c_119_n N_VGND_c_246_n 0.00402345f $X=1.515 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_27_75#_c_122_n N_VGND_c_246_n 5.84002e-19 $X=1.405 $Y=0.81 $X2=0
+ $Y2=0
cc_123 N_A_27_75#_c_124_n N_VGND_c_246_n 0.00156003f $X=1.49 $Y=1.325 $X2=0
+ $Y2=0
cc_124 N_A_27_75#_c_119_n N_VGND_c_247_n 0.00816168f $X=1.515 $Y=0.995 $X2=0
+ $Y2=0
cc_125 N_A_27_75#_c_121_n N_VGND_c_247_n 0.0118806f $X=0.28 $Y=0.52 $X2=0 $Y2=0
cc_126 N_A_27_75#_c_122_n N_VGND_c_247_n 0.0194226f $X=1.405 $Y=0.81 $X2=0 $Y2=0
cc_127 N_A_27_75#_c_124_n N_VGND_c_247_n 0.00301995f $X=1.49 $Y=1.325 $X2=0
+ $Y2=0
cc_128 N_VPWR_c_193_n N_X_M1002_d 0.00773898f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_129 N_VPWR_c_198_n X 0.0296119f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_c_193_n X 0.0162632f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_131 N_X_c_225_n N_VGND_c_244_n 0.0231208f $X=1.86 $Y=0.4 $X2=0 $Y2=0
cc_132 N_X_c_225_n N_VGND_c_246_n 0.0201254f $X=1.86 $Y=0.4 $X2=0 $Y2=0
cc_133 N_X_c_222_n N_VGND_c_246_n 0.0210195f $X=2.007 $Y=0.545 $X2=0 $Y2=0
cc_134 N_X_M1001_d N_VGND_c_247_n 0.00296227f $X=1.59 $Y=0.235 $X2=0 $Y2=0
cc_135 N_X_c_225_n N_VGND_c_247_n 0.0123242f $X=1.86 $Y=0.4 $X2=0 $Y2=0
cc_136 N_X_c_222_n N_VGND_c_247_n 0.011361f $X=2.007 $Y=0.545 $X2=0 $Y2=0
