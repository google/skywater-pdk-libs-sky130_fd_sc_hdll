# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__inv_16
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__inv_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  4.440000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 6.125000 1.315000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.984000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.580000 0.255000 0.960000 0.715000 ;
        RECT 0.580000 0.715000 7.540000 0.905000 ;
        RECT 0.580000 1.495000 7.540000 1.665000 ;
        RECT 0.580000 1.665000 0.960000 2.465000 ;
        RECT 1.520000 0.255000 1.900000 0.715000 ;
        RECT 1.520000 1.665000 1.900000 2.465000 ;
        RECT 2.460000 0.255000 2.840000 0.715000 ;
        RECT 2.460000 1.665000 2.840000 2.465000 ;
        RECT 3.400000 0.255000 3.780000 0.715000 ;
        RECT 3.400000 1.665000 3.780000 2.465000 ;
        RECT 4.340000 0.255000 4.720000 0.715000 ;
        RECT 4.340000 1.665000 4.720000 2.465000 ;
        RECT 5.280000 0.255000 5.660000 0.715000 ;
        RECT 5.280000 1.665000 5.660000 2.465000 ;
        RECT 6.220000 0.255000 6.600000 0.715000 ;
        RECT 6.220000 1.665000 6.600000 2.465000 ;
        RECT 7.015000 0.905000 7.540000 1.495000 ;
        RECT 7.160000 0.255000 7.540000 0.715000 ;
        RECT 7.160000 1.665000 7.540000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.180000  0.085000 0.410000 0.885000 ;
        RECT 1.180000  0.085000 1.350000 0.545000 ;
        RECT 2.120000  0.085000 2.290000 0.545000 ;
        RECT 3.060000  0.085000 3.230000 0.545000 ;
        RECT 4.000000  0.085000 4.170000 0.545000 ;
        RECT 4.940000  0.085000 5.110000 0.545000 ;
        RECT 5.880000  0.085000 6.050000 0.545000 ;
        RECT 6.820000  0.085000 6.990000 0.545000 ;
        RECT 7.760000  0.085000 7.970000 0.885000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.200000 1.485000 0.410000 2.635000 ;
        RECT 1.180000 1.835000 1.350000 2.635000 ;
        RECT 2.120000 1.835000 2.290000 2.635000 ;
        RECT 3.060000 1.835000 3.230000 2.635000 ;
        RECT 4.000000 1.835000 4.170000 2.635000 ;
        RECT 4.940000 1.835000 5.110000 2.635000 ;
        RECT 5.880000 1.835000 6.050000 2.635000 ;
        RECT 6.820000 1.835000 6.990000 2.635000 ;
        RECT 7.760000 1.835000 7.970000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__inv_16
