* File: sky130_fd_sc_hdll__or2_2.pxi.spice
* Created: Thu Aug 27 19:23:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR2_2%B N_B_M1006_g N_B_c_49_n N_B_M1002_g B B
+ N_B_c_48_n PM_SKY130_FD_SC_HDLL__OR2_2%B
x_PM_SKY130_FD_SC_HDLL__OR2_2%A N_A_M1003_g N_A_c_74_n N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__OR2_2%A
x_PM_SKY130_FD_SC_HDLL__OR2_2%A_39_297# N_A_39_297#_M1006_d N_A_39_297#_M1002_s
+ N_A_39_297#_c_106_n N_A_39_297#_M1004_g N_A_39_297#_c_111_n
+ N_A_39_297#_M1001_g N_A_39_297#_c_112_n N_A_39_297#_M1007_g
+ N_A_39_297#_c_107_n N_A_39_297#_M1005_g N_A_39_297#_c_108_n
+ N_A_39_297#_c_131_n N_A_39_297#_c_114_n N_A_39_297#_c_109_n
+ N_A_39_297#_c_124_n N_A_39_297#_c_110_n PM_SKY130_FD_SC_HDLL__OR2_2%A_39_297#
x_PM_SKY130_FD_SC_HDLL__OR2_2%VPWR N_VPWR_M1000_d N_VPWR_M1007_s N_VPWR_c_181_n
+ N_VPWR_c_182_n N_VPWR_c_183_n N_VPWR_c_184_n N_VPWR_c_185_n N_VPWR_c_186_n
+ VPWR N_VPWR_c_187_n N_VPWR_c_180_n PM_SKY130_FD_SC_HDLL__OR2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR2_2%X N_X_M1004_s N_X_M1001_d N_X_c_220_n N_X_c_214_n
+ X N_X_c_217_n PM_SKY130_FD_SC_HDLL__OR2_2%X
x_PM_SKY130_FD_SC_HDLL__OR2_2%VGND N_VGND_M1006_s N_VGND_M1003_d N_VGND_M1005_d
+ N_VGND_c_257_n N_VGND_c_258_n N_VGND_c_259_n N_VGND_c_260_n N_VGND_c_261_n
+ N_VGND_c_262_n VGND N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n
+ N_VGND_c_266_n PM_SKY130_FD_SC_HDLL__OR2_2%VGND
cc_1 VNB N_B_M1006_g 0.0331904f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB B 0.0118016f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B_c_48_n 0.0502927f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_4 VNB N_A_M1003_g 0.0296101f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_c_74_n 0.0240366f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.41
cc_6 VNB A 0.00507267f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_7 VNB N_A_39_297#_c_106_n 0.0179469f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.695
cc_8 VNB N_A_39_297#_c_107_n 0.0191903f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=1.202
cc_9 VNB N_A_39_297#_c_108_n 0.00425992f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_10 VNB N_A_39_297#_c_109_n 0.00128728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_39_297#_c_110_n 0.0414866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_180_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_X_c_214_n 0.00800337f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB X 0.022222f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_15 VNB N_VGND_c_257_n 0.0101374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_258_n 0.0191448f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_17 VNB N_VGND_c_259_n 0.0217535f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_18 VNB N_VGND_c_260_n 0.00265022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_261_n 0.0137002f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.16
cc_20 VNB N_VGND_c_262_n 0.0128151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_263_n 0.0138147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_264_n 0.172101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_265_n 0.00479031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_266_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_B_c_49_n 0.0231061f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.41
cc_26 VPB B 0.00291893f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_27 VPB N_B_c_48_n 0.0186624f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_28 VPB N_A_c_74_n 0.0285387f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.41
cc_29 VPB A 0.00300962f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_30 VPB N_A_39_297#_c_111_n 0.0188865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_39_297#_c_112_n 0.0195909f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_32 VPB N_A_39_297#_c_108_n 0.00166906f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_33 VPB N_A_39_297#_c_114_n 0.0157579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_39_297#_c_109_n 9.4971e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_39_297#_c_110_n 0.0220249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_181_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_37 VPB N_VPWR_c_182_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_38 VPB N_VPWR_c_183_n 0.0403297f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.202
cc_39 VPB N_VPWR_c_184_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=0.85
cc_40 VPB N_VPWR_c_185_n 0.0197179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_186_n 0.0032427f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_42 VPB N_VPWR_c_187_n 0.0160602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_180_n 0.0891847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB X 0.0226489f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_45 VPB N_X_c_217_n 0.00833419f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=1.202
cc_46 N_B_M1006_g N_A_M1003_g 0.0223994f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_47 N_B_c_49_n N_A_c_74_n 0.0358317f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_48 N_B_c_48_n N_A_c_74_n 0.025578f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_49 N_B_M1006_g A 2.09936e-19 $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_50 N_B_c_48_n A 3.14894e-19 $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_51 N_B_M1006_g N_A_39_297#_c_108_n 0.013749f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_52 N_B_c_49_n N_A_39_297#_c_108_n 0.00460399f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_53 B N_A_39_297#_c_108_n 0.0404819f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_54 N_B_c_48_n N_A_39_297#_c_108_n 0.0166619f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_55 N_B_c_49_n N_A_39_297#_c_114_n 0.018652f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_56 B N_A_39_297#_c_114_n 0.0155318f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B_c_48_n N_A_39_297#_c_114_n 0.00500354f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_58 N_B_M1006_g N_A_39_297#_c_124_n 0.00554026f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_59 N_B_c_49_n N_VPWR_c_183_n 0.00393512f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B_c_49_n N_VPWR_c_180_n 0.00500987f $X=0.555 $Y=1.41 $X2=0 $Y2=0
cc_61 N_B_M1006_g N_VGND_c_258_n 0.00538861f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_62 B N_VGND_c_258_n 0.0191398f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_B_c_48_n N_VGND_c_258_n 0.00102125f $X=0.52 $Y=1.202 $X2=0 $Y2=0
cc_64 N_B_M1006_g N_VGND_c_259_n 0.00465454f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_65 N_B_M1006_g N_VGND_c_264_n 0.00880113f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_66 B N_VGND_c_264_n 8.66838e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_67 N_A_M1003_g N_A_39_297#_c_106_n 0.0173772f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_68 A N_A_39_297#_c_106_n 0.00531148f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_69 N_A_c_74_n N_A_39_297#_c_111_n 0.0165933f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_M1003_g N_A_39_297#_c_108_n 0.00913305f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_c_74_n N_A_39_297#_c_108_n 0.00189596f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_72 A N_A_39_297#_c_108_n 0.0441306f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_73 N_A_c_74_n N_A_39_297#_c_131_n 0.0187423f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 A N_A_39_297#_c_131_n 0.0338186f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_75 N_A_c_74_n N_A_39_297#_c_114_n 8.77357e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_74_n N_A_39_297#_c_109_n 0.0010723f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_77 A N_A_39_297#_c_109_n 0.0260726f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_78 N_A_c_74_n N_A_39_297#_c_110_n 0.021386f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_74_n N_VPWR_c_181_n 0.00450741f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_74_n N_VPWR_c_183_n 0.00393512f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_74_n N_VPWR_c_180_n 0.00500987f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 A X 0.00415068f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_83 A N_VGND_M1003_d 0.00280213f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_M1003_g N_VGND_c_259_n 0.00585385f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_M1003_g N_VGND_c_260_n 0.00634679f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_c_74_n N_VGND_c_260_n 2.29546e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 A N_VGND_c_260_n 0.0195582f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_M1003_g N_VGND_c_264_n 0.00805218f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_89 A N_VGND_c_264_n 0.00921658f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_90 N_A_39_297#_c_131_n A_129_297# 0.0054944f $X=1.545 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_39_297#_c_114_n A_129_297# 0.00189464f $X=0.745 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_39_297#_c_131_n N_VPWR_M1000_d 0.00792181f $X=1.545 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_39_297#_c_111_n N_VPWR_c_181_n 0.00646392f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_39_297#_c_131_n N_VPWR_c_181_n 0.0136682f $X=1.545 $Y=1.58 $X2=0 $Y2=0
cc_95 N_A_39_297#_c_112_n N_VPWR_c_182_n 0.00570803f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_39_297#_c_111_n N_VPWR_c_185_n 0.00596719f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_39_297#_c_112_n N_VPWR_c_185_n 0.005138f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_39_297#_c_111_n N_VPWR_c_180_n 0.0112309f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_39_297#_c_112_n N_VPWR_c_180_n 0.00787528f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_39_297#_c_131_n N_X_M1001_d 0.00254051f $X=1.545 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_39_297#_c_111_n N_X_c_220_n 0.00743906f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_39_297#_c_112_n N_X_c_220_n 0.0112706f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_39_297#_c_106_n N_X_c_214_n 0.00533562f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_39_297#_c_107_n N_X_c_214_n 0.00939304f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_39_297#_c_109_n N_X_c_214_n 0.00794212f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_39_297#_c_110_n N_X_c_214_n 0.00427241f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_107 N_A_39_297#_c_106_n X 0.00110823f $X=1.495 $Y=0.995 $X2=0 $Y2=0
cc_108 N_A_39_297#_c_111_n X 0.00115531f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_39_297#_c_112_n X 0.0189003f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_39_297#_c_107_n X 0.00663439f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_39_297#_c_131_n X 0.0144166f $X=1.545 $Y=1.58 $X2=0 $Y2=0
cc_112 N_A_39_297#_c_109_n X 0.0380652f $X=1.63 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_39_297#_c_110_n X 0.0200277f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_114 N_A_39_297#_c_111_n N_X_c_217_n 0.00369948f $X=1.52 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_39_297#_c_112_n N_X_c_217_n 0.0124462f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_39_297#_c_131_n N_X_c_217_n 0.0130929f $X=1.545 $Y=1.58 $X2=0 $Y2=0
cc_117 N_A_39_297#_c_110_n N_X_c_217_n 0.00327757f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_118 N_A_39_297#_c_124_n N_VGND_c_258_n 0.0258175f $X=0.73 $Y=0.43 $X2=0 $Y2=0
cc_119 N_A_39_297#_c_124_n N_VGND_c_259_n 0.0197637f $X=0.73 $Y=0.43 $X2=0 $Y2=0
cc_120 N_A_39_297#_c_106_n N_VGND_c_260_n 0.0106811f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_A_39_297#_c_107_n N_VGND_c_260_n 8.80969e-19 $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_39_297#_c_106_n N_VGND_c_261_n 0.0046653f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_123 N_A_39_297#_c_107_n N_VGND_c_261_n 0.00198948f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_124 N_A_39_297#_c_106_n N_VGND_c_262_n 9.42871e-19 $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_125 N_A_39_297#_c_107_n N_VGND_c_262_n 0.0120866f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_126 N_A_39_297#_M1006_d N_VGND_c_264_n 0.00249917f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_127 N_A_39_297#_c_106_n N_VGND_c_264_n 0.00821929f $X=1.495 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_39_297#_c_107_n N_VGND_c_264_n 0.00290681f $X=2.015 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_A_39_297#_c_124_n N_VGND_c_264_n 0.0125114f $X=0.73 $Y=0.43 $X2=0 $Y2=0
cc_130 N_VPWR_c_180_n N_X_M1001_d 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_131 N_VPWR_c_181_n N_X_c_220_n 0.0343413f $X=1.285 $Y=2.01 $X2=0 $Y2=0
cc_132 N_VPWR_c_182_n N_X_c_220_n 0.0177504f $X=2.225 $Y=2.34 $X2=0 $Y2=0
cc_133 N_VPWR_c_185_n N_X_c_220_n 0.021848f $X=2.14 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_180_n N_X_c_220_n 0.0138674f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_135 N_VPWR_M1007_s X 0.00230341f $X=2.08 $Y=1.485 $X2=0 $Y2=0
cc_136 N_VPWR_M1007_s N_X_c_217_n 0.00396732f $X=2.08 $Y=1.485 $X2=0 $Y2=0
cc_137 N_VPWR_c_181_n N_X_c_217_n 0.0132045f $X=1.285 $Y=2.01 $X2=0 $Y2=0
cc_138 N_VPWR_c_182_n N_X_c_217_n 0.0131159f $X=2.225 $Y=2.34 $X2=0 $Y2=0
cc_139 N_VPWR_c_185_n N_X_c_217_n 0.00270601f $X=2.14 $Y=2.72 $X2=0 $Y2=0
cc_140 N_VPWR_c_187_n N_X_c_217_n 0.00158548f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_141 N_VPWR_c_180_n N_X_c_217_n 0.0085867f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_142 N_X_c_214_n N_VGND_M1005_d 0.00292162f $X=1.755 $Y=0.565 $X2=0 $Y2=0
cc_143 X N_VGND_M1005_d 2.61253e-19 $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_144 N_X_c_214_n N_VGND_c_260_n 0.0127239f $X=1.755 $Y=0.565 $X2=0 $Y2=0
cc_145 N_X_c_214_n N_VGND_c_261_n 0.00871279f $X=1.755 $Y=0.565 $X2=0 $Y2=0
cc_146 N_X_c_214_n N_VGND_c_262_n 0.0344032f $X=1.755 $Y=0.565 $X2=0 $Y2=0
cc_147 N_X_c_214_n N_VGND_c_263_n 4.7797e-19 $X=1.755 $Y=0.565 $X2=0 $Y2=0
cc_148 N_X_M1004_s N_VGND_c_264_n 0.00696682f $X=1.57 $Y=0.235 $X2=0 $Y2=0
cc_149 N_X_c_214_n N_VGND_c_264_n 0.0131318f $X=1.755 $Y=0.565 $X2=0 $Y2=0
