* File: sky130_fd_sc_hdll__or3b_4.spice
* Created: Wed Sep  2 08:49:05 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3b_4.pex.spice"
.subckt sky130_fd_sc_hdll__or3b_4  VNB VPB C_N A B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A	A
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_C_N_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1302 PD=0.773271 PS=1.46 NRD=5.712 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75003.6 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_186_21#_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.121799 PD=0.97 PS=1.19673 NRD=8.304 NRS=6.456 M=1 R=4.33333
+ SA=75000.5 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1001_d N_A_186_21#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1012_d N_A_186_21#_M1012_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333 SA=75001.5
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1012_d N_A_186_21#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=17.532 NRS=0 M=1 R=4.33333 SA=75002
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1002 N_A_186_21#_M1002_d N_A_M1002_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_B_M1006_g N_A_186_21#_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.08775 PD=1.03 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.9
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1003 N_A_186_21#_M1003_d N_A_27_47#_M1003_g N_VGND_M1006_d VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.1235 PD=1.92 PS=1.03 NRD=8.304 NRS=10.152 M=1 R=4.33333
+ SA=75003.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1009 N_VPWR_M1009_d N_C_N_M1009_g N_A_27_47#_M1009_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=75.1752 NRS=0 M=1 R=2.33333
+ SA=90000.2 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1009_d N_A_186_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.145 PD=1.90845 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_186_21#_M1004_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1004_d N_A_186_21#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.3 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_186_21#_M1011_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.8 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 A_600_297# N_A_M1015_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=17.7103 NRS=0.9653 M=1 R=5.55556 SA=90002.3
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1014 A_694_297# N_B_M1014_g A_600_297# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.145 PD=1.35 PS=1.29 NRD=23.6203 NRS=17.7103 M=1 R=5.55556 SA=90002.8
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_A_186_21#_M1005_d N_A_27_47#_M1005_g A_694_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.175 PD=2.54 PS=1.35 NRD=0.9653 NRS=23.6203 M=1 R=5.55556
+ SA=90003.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hdll__or3b_4.pxi.spice"
*
.ends
*
*
