* File: sky130_fd_sc_hdll__clkmux2_1.pex.spice
* Created: Thu Aug 27 19:03:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_79_21# 1 2 9 11 13 16 19 20 22 23 27
+ 29
c75 29 0 1.9931e-19 $X=1.525 $Y=0.54
c76 27 0 1.80039e-19 $X=2.67 $Y=2.04
r77 29 31 9.72055 $w=4.33e-07 $l=3.45e-07 $layer=LI1_cond $X=1.525 $Y=0.54
+ $X2=1.87 $Y2=0.54
r78 25 27 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.955 $Y=2.04
+ $X2=2.67 $Y2=2.04
r79 23 25 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.61 $Y=2.04
+ $X2=1.955 $Y2=2.04
r80 22 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.525 $Y=1.955
+ $X2=1.61 $Y2=2.04
r81 21 29 6.26295 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=0.54
r82 21 22 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=1.525 $Y=0.825
+ $X2=1.525 $Y2=1.955
r83 19 29 7.20249 $w=4.33e-07 $l=2.40832e-07 $layer=LI1_cond $X=1.435 $Y=0.74
+ $X2=1.525 $Y2=0.54
r84 19 20 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=1.435 $Y=0.74
+ $X2=0.685 $Y2=0.74
r85 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r86 14 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.6 $Y=0.825
+ $X2=0.685 $Y2=0.74
r87 14 16 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.6 $Y=0.825
+ $X2=0.6 $Y2=1.16
r88 11 17 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.565 $Y2=1.16
r89 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r90 7 17 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.565 $Y2=1.16
r91 7 9 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.495
r92 2 27 400 $w=1.7e-07 $l=1.07949e-06 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=1.545 $X2=2.67 $Y2=2.04
r93 2 25 400 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=1.81
+ $Y=1.545 $X2=1.955 $Y2=2.04
r94 1 31 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=1.735
+ $Y=0.235 $X2=1.87 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%S 1 3 6 8 10 13 16 17 18 19 20 21 23 27
+ 31 32
c93 16 0 1.20839e-19 $X=1.17 $Y=2.295
r94 31 32 13.2166 $w=3.58e-07 $l=3.33e-07 $layer=LI1_cond $X=3.472 $Y=1.535
+ $X2=3.805 $Y2=1.535
r95 27 30 7.79239 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=1.132 $Y=1.16
+ $X2=1.132 $Y2=1.325
r96 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.08
+ $Y=1.16 $X2=1.08 $Y2=1.16
r97 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.22 $X2=3.89 $Y2=1.22
r98 21 32 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=3.9 $Y=1.44 $X2=3.9
+ $Y2=1.535
r99 21 23 12.8421 $w=1.88e-07 $l=2.2e-07 $layer=LI1_cond $X=3.9 $Y=1.44 $X2=3.9
+ $Y2=1.22
r100 19 31 3.61205 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.33 $Y=1.63
+ $X2=3.33 $Y2=1.535
r101 19 20 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=3.33 $Y=1.63
+ $X2=3.33 $Y2=2.295
r102 17 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=3.33 $Y2=2.295
r103 17 18 128.85 $w=1.68e-07 $l=1.975e-06 $layer=LI1_cond $X=3.245 $Y=2.38
+ $X2=1.27 $Y2=2.38
r104 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.17 $Y=2.295
+ $X2=1.27 $Y2=2.38
r105 16 30 53.7909 $w=1.98e-07 $l=9.7e-07 $layer=LI1_cond $X=1.17 $Y=2.295
+ $X2=1.17 $Y2=1.325
r106 11 24 39.2931 $w=2.55e-07 $l=1.88348e-07 $layer=POLY_cond $X=3.94 $Y=1.055
+ $X2=3.89 $Y2=1.22
r107 11 13 287.149 $w=1.5e-07 $l=5.6e-07 $layer=POLY_cond $X=3.94 $Y=1.055
+ $X2=3.94 $Y2=0.495
r108 8 24 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=3.915 $Y=1.47
+ $X2=3.89 $Y2=1.22
r109 8 10 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.915 $Y=1.47
+ $X2=3.915 $Y2=2.015
r110 4 28 39.2931 $w=2.55e-07 $l=1.94808e-07 $layer=POLY_cond $X=1.15 $Y=0.995
+ $X2=1.085 $Y2=1.16
r111 4 6 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.15 $Y=0.995
+ $X2=1.15 $Y2=0.445
r112 1 28 62.8272 $w=2.55e-07 $l=3.29393e-07 $layer=POLY_cond $X=1.125 $Y=1.47
+ $X2=1.085 $Y2=1.16
r113 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.125 $Y=1.47
+ $X2=1.125 $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A1 3 5 7 10 11 13 14 16 17
c68 5 0 1.3232e-19 $X=2.905 $Y=1.47
r69 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.22 $X2=2.87 $Y2=1.22
r70 17 26 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=2.93 $Y=1.19 $X2=2.93
+ $Y2=1.22
r71 16 17 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.93 $Y=0.85
+ $X2=2.93 $Y2=1.19
r72 15 26 15.6971 $w=2.88e-07 $l=3.95e-07 $layer=LI1_cond $X=2.93 $Y=1.615
+ $X2=2.93 $Y2=1.22
r73 13 15 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.785 $Y=1.7
+ $X2=2.93 $Y2=1.615
r74 13 14 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=2.785 $Y=1.7
+ $X2=1.95 $Y2=1.7
r75 11 20 45.5456 $w=2.7e-07 $l=2.05e-07 $layer=POLY_cond $X=1.865 $Y=0.975
+ $X2=1.66 $Y2=0.975
r76 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.865
+ $Y=0.975 $X2=1.865 $Y2=0.975
r77 8 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=1.615
+ $X2=1.95 $Y2=1.7
r78 8 10 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.865 $Y=1.615
+ $X2=1.865 $Y2=0.975
r79 5 25 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.905 $Y=1.47
+ $X2=2.87 $Y2=1.22
r80 5 7 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.905 $Y=1.47
+ $X2=2.905 $Y2=2.015
r81 1 20 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.66 $Y=0.84
+ $X2=1.66 $Y2=0.975
r82 1 3 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.66 $Y=0.84 $X2=1.66
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A0 1 3 4 5 8 11 12 15 16
c50 1 0 1.20839e-19 $X=1.72 $Y=1.47
r51 15 18 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=0.98
+ $X2=2.375 $Y2=1.145
r52 15 17 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.375 $Y=0.98
+ $X2=2.375 $Y2=0.815
r53 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.375
+ $Y=0.98 $X2=2.375 $Y2=0.98
r54 12 16 7.44655 $w=3.23e-07 $l=2.1e-07 $layer=LI1_cond $X=2.452 $Y=1.19
+ $X2=2.452 $Y2=0.98
r55 11 18 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=2.34 $Y=1.32 $X2=2.34
+ $Y2=1.145
r56 8 17 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=2.315 $Y=0.445
+ $X2=2.315 $Y2=0.815
r57 4 11 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=2.24 $Y=1.395
+ $X2=2.34 $Y2=1.32
r58 4 5 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.24 $Y=1.395 $X2=1.81
+ $Y2=1.395
r59 1 5 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.72 $Y=1.47
+ $X2=1.81 $Y2=1.395
r60 1 3 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.72 $Y=1.47 $X2=1.72
+ $Y2=2.015
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_649_21# 1 2 9 12 13 15 18 19 21 22 27
+ 32 33 34
c68 18 0 1.3232e-19 $X=3.41 $Y=1.02
c69 13 0 1.80039e-19 $X=3.345 $Y=1.47
c70 9 0 1.95128e-19 $X=3.32 $Y=0.445
r71 32 33 8.64761 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=2
+ $X2=4.185 $Y2=1.835
r72 29 34 4.36305 $w=2.07e-07 $l=1.25499e-07 $layer=LI1_cond $X=4.3 $Y=0.865
+ $X2=4.21 $Y2=0.78
r73 29 33 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.3 $Y=0.865 $X2=4.3
+ $Y2=1.835
r74 25 34 4.36305 $w=2.07e-07 $l=1.08305e-07 $layer=LI1_cond $X=4.157 $Y=0.695
+ $X2=4.21 $Y2=0.78
r75 25 27 11.2892 $w=2.43e-07 $l=2.4e-07 $layer=LI1_cond $X=4.157 $Y=0.695
+ $X2=4.157 $Y2=0.455
r76 21 34 2.06925 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=4.035 $Y=0.78
+ $X2=4.21 $Y2=0.78
r77 21 22 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=4.035 $Y=0.78
+ $X2=3.495 $Y2=0.78
r78 19 37 39.6736 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.02
+ $X2=3.395 $Y2=1.185
r79 19 36 47.9795 $w=3e-07 $l=1.65e-07 $layer=POLY_cond $X=3.395 $Y=1.02
+ $X2=3.395 $Y2=0.855
r80 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.41
+ $Y=1.02 $X2=3.41 $Y2=1.02
r81 16 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.41 $Y=0.865
+ $X2=3.495 $Y2=0.78
r82 16 18 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=3.41 $Y=0.865
+ $X2=3.41 $Y2=1.02
r83 13 15 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=3.345 $Y=1.47
+ $X2=3.345 $Y2=2.015
r84 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.345 $Y=1.37 $X2=3.345
+ $Y2=1.47
r85 12 37 61.3418 $w=2e-07 $l=1.85e-07 $layer=POLY_cond $X=3.345 $Y=1.37
+ $X2=3.345 $Y2=1.185
r86 9 36 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=3.32 $Y=0.445
+ $X2=3.32 $Y2=0.855
r87 2 32 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=4.005
+ $Y=1.545 $X2=4.15 $Y2=2
r88 1 27 182 $w=1.7e-07 $l=2.79464e-07 $layer=licon1_NDIFF $count=1 $X=4.015
+ $Y=0.235 $X2=4.15 $Y2=0.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%X 1 2 10 12 13 14
r17 14 27 4.47217 $w=3.33e-07 $l=1.3e-07 $layer=LI1_cond $X=0.257 $Y=2.21
+ $X2=0.257 $Y2=2.34
r18 13 14 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=1.87
+ $X2=0.257 $Y2=2.21
r19 11 12 46.0977 $w=2.53e-07 $l=1.02e-06 $layer=LI1_cond $X=0.217 $Y=1.495
+ $X2=0.217 $Y2=0.475
r20 10 11 6.36149 $w=3.33e-07 $l=1.65e-07 $layer=LI1_cond $X=0.257 $Y=1.66
+ $X2=0.257 $Y2=1.495
r21 8 13 7.15547 $w=3.33e-07 $l=2.08e-07 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.87
r22 8 10 0.0688026 $w=3.33e-07 $l=2e-09 $layer=LI1_cond $X=0.257 $Y=1.662
+ $X2=0.257 $Y2=1.66
r23 2 27 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r24 2 10 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r25 1 12 182 $w=1.7e-07 $l=2.95973e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VPWR 1 2 11 17 20 21 22 32 33 36
r46 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r48 30 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r49 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r50 27 30 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r51 27 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 26 29 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 26 27 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 24 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.73 $Y2=2.72
r55 24 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r56 22 37 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 20 29 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 20 21 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.585 $Y=2.72
+ $X2=3.7 $Y2=2.72
r59 19 32 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=4.37 $Y2=2.72
r60 19 21 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.815 $Y=2.72
+ $X2=3.7 $Y2=2.72
r61 15 21 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=2.635 $X2=3.7
+ $Y2=2.72
r62 15 17 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.7 $Y=2.635
+ $X2=3.7 $Y2=2
r63 11 14 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.73 $Y=1.66
+ $X2=0.73 $Y2=2.34
r64 9 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635 $X2=0.73
+ $Y2=2.72
r65 9 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.34
r66 2 17 300 $w=1.7e-07 $l=5.60312e-07 $layer=licon1_PDIFF $count=2 $X=3.435
+ $Y=1.545 $X2=3.67 $Y2=2
r67 1 14 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r68 1 11 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VGND 1 2 9 11 13 18 28 29 32
c55 18 0 1.95128e-19 $X=3.25 $Y=0
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r57 29 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.45
+ $Y2=0
r58 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r59 26 28 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=3.765 $Y=0 $X2=4.37
+ $Y2=0
r60 25 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r61 24 25 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r62 22 25 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r63 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r64 21 24 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r65 21 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r66 19 32 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r67 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r68 18 39 8.36094 $w=5.13e-07 $l=3.6e-07 $layer=LI1_cond $X=3.507 $Y=0 $X2=3.507
+ $Y2=0.36
r69 18 26 7.34265 $w=1.7e-07 $l=2.58e-07 $layer=LI1_cond $X=3.507 $Y=0 $X2=3.765
+ $Y2=0
r70 18 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r71 18 24 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=2.99
+ $Y2=0
r72 13 32 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r73 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r74 11 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 7 32 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r77 7 9 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.38
r78 2 39 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=3.395
+ $Y=0.235 $X2=3.63 $Y2=0.36
r79 1 9 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

