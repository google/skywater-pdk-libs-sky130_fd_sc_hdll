* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a21o_8 A1 A2 B1 VGND VNB VPB VPWR X
X0 a_27_297# B1 a_213_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR a_213_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_213_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_213_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND B1 a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_213_47# A1 a_297_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_27_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 X a_213_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 X a_213_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR A2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_131_47# A1 a_213_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 X a_213_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND A2 a_131_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_213_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_213_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 X a_213_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VPWR a_213_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND a_213_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 X a_213_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_297_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VGND a_213_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR A1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND a_213_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR a_213_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VGND a_213_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_213_47# B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 X a_213_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
