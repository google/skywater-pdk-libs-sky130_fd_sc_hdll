# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkmux2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkmux2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.290000 0.255000 2.615000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.780000 0.810000 1.950000 1.615000 ;
        RECT 1.780000 1.615000 3.075000 1.785000 ;
        RECT 2.785000 0.255000 3.075000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.479400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.995000 1.270000 1.325000 ;
        RECT 1.070000 1.325000 1.270000 2.295000 ;
        RECT 1.070000 2.295000 3.415000 2.465000 ;
        RECT 3.245000 1.440000 3.995000 1.630000 ;
        RECT 3.245000 1.630000 3.415000 2.295000 ;
        RECT 3.805000 1.055000 3.995000 1.440000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.405200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.255000 0.345000 1.495000 ;
        RECT 0.090000 1.495000 0.425000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.485000 ;
      RECT 0.515000  0.655000 1.610000 0.825000 ;
      RECT 0.515000  0.825000 0.685000 1.325000 ;
      RECT 0.645000  1.495000 0.815000 2.635000 ;
      RECT 1.435000  0.255000 1.955000 0.620000 ;
      RECT 1.435000  0.620000 1.610000 0.655000 ;
      RECT 1.440000  0.825000 1.610000 1.955000 ;
      RECT 1.440000  1.955000 2.885000 2.125000 ;
      RECT 3.250000  0.085000 3.765000 0.525000 ;
      RECT 3.325000  0.695000 4.385000 0.865000 ;
      RECT 3.325000  0.865000 3.495000 1.185000 ;
      RECT 3.585000  1.835000 3.815000 2.635000 ;
      RECT 3.985000  1.835000 4.385000 2.465000 ;
      RECT 4.035000  0.255000 4.280000 0.695000 ;
      RECT 4.215000  0.865000 4.385000 1.835000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_1
END LIBRARY
