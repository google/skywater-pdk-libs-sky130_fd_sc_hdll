* File: sky130_fd_sc_hdll__muxb16to1_4.pxi.spice
* Created: Thu Aug 27 19:11:38 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VNB VNB VNB VNB
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VNB
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPB VPB VPB VPB VPB VPB N_VPB_c_1128_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPB
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[0] N_D[0]_M1014_g N_D[0]_M1084_g
+ N_D[0]_M1219_g N_D[0]_M1146_g N_D[0]_M1208_g N_D[0]_M1300_g N_D[0]_M1317_g
+ N_D[0]_M1294_g D[0] N_D[0]_c_1877_n N_D[0]_c_1878_n N_D[0]_c_1879_n
+ N_D[0]_c_1880_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[8] N_D[8]_M1023_g N_D[8]_M1085_g
+ N_D[8]_M1090_g N_D[8]_M1155_g N_D[8]_M1221_g N_D[8]_M1235_g N_D[8]_M1240_g
+ N_D[8]_M1304_g D[8] N_D[8]_c_1967_n N_D[8]_c_1968_n N_D[8]_c_1969_n
+ N_D[8]_c_1970_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_265# N_A_559_265#_M1139_d
+ N_A_559_265#_M1018_s N_A_559_265#_c_2052_n N_A_559_265#_M1137_g
+ N_A_559_265#_c_2053_n N_A_559_265#_c_2054_n N_A_559_265#_c_2055_n
+ N_A_559_265#_M1207_g N_A_559_265#_c_2056_n N_A_559_265#_c_2057_n
+ N_A_559_265#_M1249_g N_A_559_265#_c_2058_n N_A_559_265#_c_2059_n
+ N_A_559_265#_M1299_g N_A_559_265#_c_2060_n N_A_559_265#_c_2061_n
+ N_A_559_265#_c_2045_n N_A_559_265#_c_2046_n N_A_559_265#_c_2047_n
+ N_A_559_265#_c_2048_n N_A_559_265#_c_2064_n N_A_559_265#_c_2049_n
+ N_A_559_265#_c_2050_n N_A_559_265#_c_2066_n N_A_559_265#_c_2051_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_793# N_A_559_793#_M1017_d
+ N_A_559_793#_M1123_s N_A_559_793#_c_2170_n N_A_559_793#_M1026_g
+ N_A_559_793#_c_2171_n N_A_559_793#_c_2172_n N_A_559_793#_c_2173_n
+ N_A_559_793#_M1079_g N_A_559_793#_c_2174_n N_A_559_793#_c_2175_n
+ N_A_559_793#_M1127_g N_A_559_793#_c_2176_n N_A_559_793#_c_2177_n
+ N_A_559_793#_M1269_g N_A_559_793#_c_2178_n N_A_559_793#_c_2179_n
+ N_A_559_793#_c_2163_n N_A_559_793#_c_2164_n N_A_559_793#_c_2182_n
+ N_A_559_793#_c_2183_n N_A_559_793#_c_2165_n N_A_559_793#_c_2166_n
+ N_A_559_793#_c_2184_n N_A_559_793#_c_2167_n N_A_559_793#_c_2168_n
+ N_A_559_793#_c_2169_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_559_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[0] N_S[0]_c_2287_n N_S[0]_M1053_g
+ N_S[0]_c_2288_n N_S[0]_c_2289_n N_S[0]_c_2290_n N_S[0]_M1074_g N_S[0]_c_2291_n
+ N_S[0]_c_2292_n N_S[0]_M1105_g N_S[0]_c_2293_n N_S[0]_c_2294_n N_S[0]_M1125_g
+ N_S[0]_c_2295_n N_S[0]_c_2296_n N_S[0]_c_2297_n N_S[0]_c_2298_n
+ N_S[0]_c_2299_n N_S[0]_c_2310_n N_S[0]_M1018_g N_S[0]_c_2300_n N_S[0]_M1139_g
+ N_S[0]_c_2301_n N_S[0]_c_2302_n N_S[0]_M1192_g N_S[0]_c_2303_n N_S[0]_M1061_g
+ N_S[0]_c_2304_n N_S[0]_c_2305_n N_S[0]_c_2306_n N_S[0]_c_2307_n S[0]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[8] N_S[8]_c_2404_n N_S[8]_M1070_g
+ N_S[8]_c_2405_n N_S[8]_c_2406_n N_S[8]_c_2407_n N_S[8]_M1159_g N_S[8]_c_2408_n
+ N_S[8]_c_2409_n N_S[8]_M1236_g N_S[8]_c_2410_n N_S[8]_c_2411_n N_S[8]_M1302_g
+ N_S[8]_c_2412_n N_S[8]_c_2413_n N_S[8]_c_2414_n N_S[8]_c_2415_n
+ N_S[8]_c_2425_n N_S[8]_c_2416_n N_S[8]_c_2427_n N_S[8]_M1123_g N_S[8]_c_2417_n
+ N_S[8]_M1017_g N_S[8]_c_2418_n N_S[8]_c_2419_n N_S[8]_M1078_g N_S[8]_c_2429_n
+ N_S[8]_M1172_g N_S[8]_c_2420_n N_S[8]_c_2421_n N_S[8]_c_2422_n N_S[8]_c_2423_n
+ S[8] PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[8]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[1] N_S[1]_c_2529_n N_S[1]_c_2530_n
+ N_S[1]_M1133_g N_S[1]_c_2531_n N_S[1]_M1241_g N_S[1]_c_2532_n N_S[1]_c_2533_n
+ N_S[1]_M1288_g N_S[1]_c_2534_n N_S[1]_c_2554_n N_S[1]_M1180_g N_S[1]_c_2535_n
+ N_S[1]_c_2536_n N_S[1]_c_2537_n N_S[1]_c_2538_n N_S[1]_c_2539_n N_S[1]_M1039_g
+ N_S[1]_c_2540_n N_S[1]_c_2541_n N_S[1]_M1045_g N_S[1]_c_2542_n N_S[1]_c_2543_n
+ N_S[1]_M1093_g N_S[1]_c_2544_n N_S[1]_c_2545_n N_S[1]_M1113_g N_S[1]_c_2546_n
+ N_S[1]_c_2547_n N_S[1]_c_2548_n N_S[1]_c_2549_n S[1] N_S[1]_c_2550_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[9] N_S[9]_c_2649_n N_S[9]_c_2671_n
+ N_S[9]_M1225_g N_S[9]_c_2650_n N_S[9]_M1008_g N_S[9]_c_2651_n N_S[9]_c_2673_n
+ N_S[9]_c_2652_n N_S[9]_c_2653_n N_S[9]_M1107_g N_S[9]_c_2675_n N_S[9]_M1266_g
+ N_S[9]_c_2654_n N_S[9]_c_2655_n N_S[9]_c_2656_n N_S[9]_c_2657_n
+ N_S[9]_c_2658_n N_S[9]_M1027_g N_S[9]_c_2659_n N_S[9]_c_2660_n N_S[9]_M1032_g
+ N_S[9]_c_2661_n N_S[9]_c_2662_n N_S[9]_M1096_g N_S[9]_c_2663_n N_S[9]_c_2664_n
+ N_S[9]_M1259_g N_S[9]_c_2665_n N_S[9]_c_2666_n N_S[9]_c_2667_n N_S[9]_c_2668_n
+ S[9] N_S[9]_c_2669_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_325# N_A_1430_325#_M1241_s
+ N_A_1430_325#_M1133_s N_A_1430_325#_c_2784_n N_A_1430_325#_M1007_g
+ N_A_1430_325#_c_2785_n N_A_1430_325#_c_2777_n N_A_1430_325#_c_2787_n
+ N_A_1430_325#_M1048_g N_A_1430_325#_c_2788_n N_A_1430_325#_c_2789_n
+ N_A_1430_325#_M1140_g N_A_1430_325#_c_2790_n N_A_1430_325#_c_2791_n
+ N_A_1430_325#_M1284_g N_A_1430_325#_c_2792_n N_A_1430_325#_c_2793_n
+ N_A_1430_325#_c_2794_n N_A_1430_325#_c_2778_n N_A_1430_325#_c_2779_n
+ N_A_1430_325#_c_2780_n N_A_1430_325#_c_2796_n N_A_1430_325#_c_2781_n
+ N_A_1430_325#_c_2782_n N_A_1430_325#_c_2783_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_325#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_599# N_A_1430_599#_M1008_d
+ N_A_1430_599#_M1225_s N_A_1430_599#_c_2900_n N_A_1430_599#_M1112_g
+ N_A_1430_599#_c_2901_n N_A_1430_599#_c_2893_n N_A_1430_599#_c_2903_n
+ N_A_1430_599#_M1161_g N_A_1430_599#_c_2904_n N_A_1430_599#_c_2905_n
+ N_A_1430_599#_M1199_g N_A_1430_599#_c_2906_n N_A_1430_599#_c_2907_n
+ N_A_1430_599#_M1273_g N_A_1430_599#_c_2908_n N_A_1430_599#_c_2909_n
+ N_A_1430_599#_c_2910_n N_A_1430_599#_c_2894_n N_A_1430_599#_c_2895_n
+ N_A_1430_599#_c_2911_n N_A_1430_599#_c_2896_n N_A_1430_599#_c_2913_n
+ N_A_1430_599#_c_2897_n N_A_1430_599#_c_2898_n N_A_1430_599#_c_2899_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1430_599#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[1] N_D[1]_M1002_g N_D[1]_M1049_g
+ N_D[1]_M1098_g N_D[1]_M1038_g N_D[1]_M1134_g N_D[1]_M1167_g N_D[1]_M1315_g
+ N_D[1]_M1271_g D[1] N_D[1]_c_3023_n N_D[1]_c_3024_n N_D[1]_c_3025_n
+ N_D[1]_c_3026_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[9] N_D[9]_M1011_g N_D[9]_M1019_g
+ N_D[9]_M1111_g N_D[9]_M1051_g N_D[9]_M1148_g N_D[9]_M1178_g N_D[9]_M1276_g
+ N_D[9]_M1285_g D[9] N_D[9]_c_3116_n N_D[9]_c_3117_n N_D[9]_c_3118_n
+ N_D[9]_c_3119_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[9]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[2] N_D[2]_M1020_g N_D[2]_M1001_g
+ N_D[2]_M1062_g N_D[2]_M1067_g N_D[2]_M1157_g N_D[2]_M1110_g N_D[2]_M1182_g
+ N_D[2]_M1301_g D[2] N_D[2]_c_3207_n N_D[2]_c_3208_n N_D[2]_c_3209_n
+ N_D[2]_c_3210_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[10] N_D[10]_M1024_g N_D[10]_M1033_g
+ N_D[10]_M1143_g N_D[10]_M1076_g N_D[10]_M1164_g N_D[10]_M1195_g
+ N_D[10]_M1307_g N_D[10]_M1309_g D[10] N_D[10]_c_3302_n N_D[10]_c_3303_n
+ N_D[10]_c_3304_n N_D[10]_c_3305_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_265# N_A_3135_265#_M1222_s
+ N_A_3135_265#_M1065_d N_A_3135_265#_c_3392_n N_A_3135_265#_M1082_g
+ N_A_3135_265#_c_3393_n N_A_3135_265#_c_3394_n N_A_3135_265#_c_3395_n
+ N_A_3135_265#_M1138_g N_A_3135_265#_c_3396_n N_A_3135_265#_c_3397_n
+ N_A_3135_265#_M1181_g N_A_3135_265#_c_3398_n N_A_3135_265#_c_3399_n
+ N_A_3135_265#_M1250_g N_A_3135_265#_c_3400_n N_A_3135_265#_c_3401_n
+ N_A_3135_265#_c_3385_n N_A_3135_265#_c_3386_n N_A_3135_265#_c_3387_n
+ N_A_3135_265#_c_3388_n N_A_3135_265#_c_3404_n N_A_3135_265#_c_3389_n
+ N_A_3135_265#_c_3390_n N_A_3135_265#_c_3406_n N_A_3135_265#_c_3391_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_793# N_A_3135_793#_M1043_d
+ N_A_3135_793#_M1083_s N_A_3135_793#_c_3511_n N_A_3135_793#_M1000_g
+ N_A_3135_793#_c_3512_n N_A_3135_793#_c_3513_n N_A_3135_793#_c_3514_n
+ N_A_3135_793#_M1080_g N_A_3135_793#_c_3515_n N_A_3135_793#_c_3516_n
+ N_A_3135_793#_M1229_g N_A_3135_793#_c_3517_n N_A_3135_793#_c_3518_n
+ N_A_3135_793#_M1270_g N_A_3135_793#_c_3519_n N_A_3135_793#_c_3520_n
+ N_A_3135_793#_c_3504_n N_A_3135_793#_c_3505_n N_A_3135_793#_c_3523_n
+ N_A_3135_793#_c_3524_n N_A_3135_793#_c_3506_n N_A_3135_793#_c_3507_n
+ N_A_3135_793#_c_3525_n N_A_3135_793#_c_3508_n N_A_3135_793#_c_3509_n
+ N_A_3135_793#_c_3510_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_3135_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[2] N_S[2]_c_3629_n N_S[2]_M1035_g
+ N_S[2]_c_3630_n N_S[2]_c_3631_n N_S[2]_c_3632_n N_S[2]_M1036_g N_S[2]_c_3633_n
+ N_S[2]_c_3634_n N_S[2]_M1108_g N_S[2]_c_3635_n N_S[2]_c_3636_n N_S[2]_M1306_g
+ N_S[2]_c_3637_n N_S[2]_c_3638_n N_S[2]_c_3639_n N_S[2]_c_3640_n
+ N_S[2]_c_3641_n N_S[2]_c_3652_n N_S[2]_M1065_g N_S[2]_c_3642_n N_S[2]_M1222_g
+ N_S[2]_c_3643_n N_S[2]_c_3644_n N_S[2]_M1239_g N_S[2]_c_3645_n N_S[2]_M1308_g
+ N_S[2]_c_3646_n N_S[2]_c_3647_n N_S[2]_c_3648_n N_S[2]_c_3649_n S[2]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[10] N_S[10]_c_3746_n N_S[10]_M1010_g
+ N_S[10]_c_3747_n N_S[10]_c_3748_n N_S[10]_c_3749_n N_S[10]_M1214_g
+ N_S[10]_c_3750_n N_S[10]_c_3751_n N_S[10]_M1263_g N_S[10]_c_3752_n
+ N_S[10]_c_3753_n N_S[10]_M1268_g N_S[10]_c_3754_n N_S[10]_c_3755_n
+ N_S[10]_c_3756_n N_S[10]_c_3757_n N_S[10]_c_3767_n N_S[10]_c_3758_n
+ N_S[10]_c_3769_n N_S[10]_M1083_g N_S[10]_c_3759_n N_S[10]_M1043_g
+ N_S[10]_c_3760_n N_S[10]_c_3761_n N_S[10]_M1215_g N_S[10]_c_3771_n
+ N_S[10]_M1173_g N_S[10]_c_3762_n N_S[10]_c_3763_n N_S[10]_c_3764_n
+ N_S[10]_c_3765_n S[10] PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[10]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[3] N_S[3]_c_3871_n N_S[3]_c_3872_n
+ N_S[3]_M1150_g N_S[3]_c_3873_n N_S[3]_M1234_g N_S[3]_c_3874_n N_S[3]_c_3875_n
+ N_S[3]_M1291_g N_S[3]_c_3876_n N_S[3]_c_3896_n N_S[3]_M1280_g N_S[3]_c_3877_n
+ N_S[3]_c_3878_n N_S[3]_c_3879_n N_S[3]_c_3880_n N_S[3]_c_3881_n N_S[3]_M1030_g
+ N_S[3]_c_3882_n N_S[3]_c_3883_n N_S[3]_M1031_g N_S[3]_c_3884_n N_S[3]_c_3885_n
+ N_S[3]_M1059_g N_S[3]_c_3886_n N_S[3]_c_3887_n N_S[3]_M1106_g N_S[3]_c_3888_n
+ N_S[3]_c_3889_n N_S[3]_c_3890_n N_S[3]_c_3891_n S[3] N_S[3]_c_3892_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[11] N_S[11]_c_3991_n N_S[11]_c_4013_n
+ N_S[11]_M1066_g N_S[11]_c_3992_n N_S[11]_M1054_g N_S[11]_c_3993_n
+ N_S[11]_c_4015_n N_S[11]_c_3994_n N_S[11]_c_3995_n N_S[11]_M1072_g
+ N_S[11]_c_4017_n N_S[11]_M1237_g N_S[11]_c_3996_n N_S[11]_c_3997_n
+ N_S[11]_c_3998_n N_S[11]_c_3999_n N_S[11]_c_4000_n N_S[11]_M1047_g
+ N_S[11]_c_4001_n N_S[11]_c_4002_n N_S[11]_M1160_g N_S[11]_c_4003_n
+ N_S[11]_c_4004_n N_S[11]_M1316_g N_S[11]_c_4005_n N_S[11]_c_4006_n
+ N_S[11]_M1318_g N_S[11]_c_4007_n N_S[11]_c_4008_n N_S[11]_c_4009_n
+ N_S[11]_c_4010_n S[11] N_S[11]_c_4011_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_325# N_A_4006_325#_M1234_s
+ N_A_4006_325#_M1150_d N_A_4006_325#_c_4126_n N_A_4006_325#_M1121_g
+ N_A_4006_325#_c_4127_n N_A_4006_325#_c_4119_n N_A_4006_325#_c_4129_n
+ N_A_4006_325#_M1171_g N_A_4006_325#_c_4130_n N_A_4006_325#_c_4131_n
+ N_A_4006_325#_M1243_g N_A_4006_325#_c_4132_n N_A_4006_325#_c_4133_n
+ N_A_4006_325#_M1287_g N_A_4006_325#_c_4134_n N_A_4006_325#_c_4135_n
+ N_A_4006_325#_c_4136_n N_A_4006_325#_c_4120_n N_A_4006_325#_c_4121_n
+ N_A_4006_325#_c_4122_n N_A_4006_325#_c_4138_n N_A_4006_325#_c_4123_n
+ N_A_4006_325#_c_4124_n N_A_4006_325#_c_4125_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_325#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_599# N_A_4006_599#_M1054_s
+ N_A_4006_599#_M1066_s N_A_4006_599#_c_4242_n N_A_4006_599#_M1071_g
+ N_A_4006_599#_c_4243_n N_A_4006_599#_c_4235_n N_A_4006_599#_c_4245_n
+ N_A_4006_599#_M1114_g N_A_4006_599#_c_4246_n N_A_4006_599#_c_4247_n
+ N_A_4006_599#_M1260_g N_A_4006_599#_c_4248_n N_A_4006_599#_c_4249_n
+ N_A_4006_599#_M1313_g N_A_4006_599#_c_4250_n N_A_4006_599#_c_4251_n
+ N_A_4006_599#_c_4252_n N_A_4006_599#_c_4236_n N_A_4006_599#_c_4237_n
+ N_A_4006_599#_c_4253_n N_A_4006_599#_c_4238_n N_A_4006_599#_c_4255_n
+ N_A_4006_599#_c_4239_n N_A_4006_599#_c_4240_n N_A_4006_599#_c_4241_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4006_599#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[3] N_D[3]_M1042_g N_D[3]_M1041_g
+ N_D[3]_M1100_g N_D[3]_M1089_g N_D[3]_M1116_g N_D[3]_M1135_g N_D[3]_M1193_g
+ N_D[3]_M1289_g D[3] N_D[3]_c_4365_n N_D[3]_c_4366_n N_D[3]_c_4367_n
+ N_D[3]_c_4368_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[11] N_D[11]_M1052_g N_D[11]_M1245_g
+ N_D[11]_M1296_g N_D[11]_M1101_g N_D[11]_M1129_g N_D[11]_M1310_g
+ N_D[11]_M1311_g N_D[11]_M1297_g D[11] N_D[11]_c_4459_n N_D[11]_c_4460_n
+ N_D[11]_c_4461_n N_D[11]_c_4462_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[11]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[4] N_D[4]_M1158_g N_D[4]_M1021_g
+ N_D[4]_M1177_g N_D[4]_M1194_g N_D[4]_M1265_g N_D[4]_M1232_g N_D[4]_M1275_g
+ N_D[4]_M1319_g D[4] N_D[4]_c_4551_n N_D[4]_c_4552_n N_D[4]_c_4553_n
+ N_D[4]_c_4554_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[12] N_D[12]_M1006_g N_D[12]_M1012_g
+ N_D[12]_M1128_g N_D[12]_M1165_g N_D[12]_M1203_g N_D[12]_M1187_g
+ N_D[12]_M1267_g N_D[12]_M1277_g D[12] N_D[12]_c_4647_n N_D[12]_c_4648_n
+ N_D[12]_c_4649_n N_D[12]_c_4650_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_265# N_A_5803_265#_M1037_s
+ N_A_5803_265#_M1016_s N_A_5803_265#_c_4738_n N_A_5803_265#_M1050_g
+ N_A_5803_265#_c_4739_n N_A_5803_265#_c_4740_n N_A_5803_265#_c_4741_n
+ N_A_5803_265#_M1118_g N_A_5803_265#_c_4742_n N_A_5803_265#_c_4743_n
+ N_A_5803_265#_M1231_g N_A_5803_265#_c_4744_n N_A_5803_265#_c_4745_n
+ N_A_5803_265#_M1295_g N_A_5803_265#_c_4746_n N_A_5803_265#_c_4747_n
+ N_A_5803_265#_c_4731_n N_A_5803_265#_c_4732_n N_A_5803_265#_c_4733_n
+ N_A_5803_265#_c_4734_n N_A_5803_265#_c_4750_n N_A_5803_265#_c_4735_n
+ N_A_5803_265#_c_4736_n N_A_5803_265#_c_4752_n N_A_5803_265#_c_4737_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_793# N_A_5803_793#_M1188_d
+ N_A_5803_793#_M1120_s N_A_5803_793#_c_4857_n N_A_5803_793#_M1055_g
+ N_A_5803_793#_c_4858_n N_A_5803_793#_c_4859_n N_A_5803_793#_c_4860_n
+ N_A_5803_793#_M1119_g N_A_5803_793#_c_4861_n N_A_5803_793#_c_4862_n
+ N_A_5803_793#_M1200_g N_A_5803_793#_c_4863_n N_A_5803_793#_c_4864_n
+ N_A_5803_793#_M1257_g N_A_5803_793#_c_4865_n N_A_5803_793#_c_4866_n
+ N_A_5803_793#_c_4850_n N_A_5803_793#_c_4851_n N_A_5803_793#_c_4869_n
+ N_A_5803_793#_c_4870_n N_A_5803_793#_c_4852_n N_A_5803_793#_c_4853_n
+ N_A_5803_793#_c_4871_n N_A_5803_793#_c_4854_n N_A_5803_793#_c_4855_n
+ N_A_5803_793#_c_4856_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5803_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[4] N_S[4]_c_4975_n N_S[4]_M1154_g
+ N_S[4]_c_4976_n N_S[4]_c_4977_n N_S[4]_c_4978_n N_S[4]_M1191_g N_S[4]_c_4979_n
+ N_S[4]_c_4980_n N_S[4]_M1205_g N_S[4]_c_4981_n N_S[4]_c_4982_n N_S[4]_M1213_g
+ N_S[4]_c_4983_n N_S[4]_c_4984_n N_S[4]_c_4985_n N_S[4]_c_4986_n
+ N_S[4]_c_4987_n N_S[4]_c_4998_n N_S[4]_M1016_g N_S[4]_c_4988_n N_S[4]_M1037_g
+ N_S[4]_c_4989_n N_S[4]_c_4990_n N_S[4]_M1086_g N_S[4]_c_4991_n N_S[4]_M1095_g
+ N_S[4]_c_4992_n N_S[4]_c_4993_n N_S[4]_c_4994_n N_S[4]_c_4995_n S[4]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[12] N_S[12]_c_5092_n N_S[12]_M1044_g
+ N_S[12]_c_5093_n N_S[12]_c_5094_n N_S[12]_c_5095_n N_S[12]_M1091_g
+ N_S[12]_c_5096_n N_S[12]_c_5097_n N_S[12]_M1218_g N_S[12]_c_5098_n
+ N_S[12]_c_5099_n N_S[12]_M1312_g N_S[12]_c_5100_n N_S[12]_c_5101_n
+ N_S[12]_c_5102_n N_S[12]_c_5103_n N_S[12]_c_5113_n N_S[12]_c_5104_n
+ N_S[12]_c_5115_n N_S[12]_M1120_g N_S[12]_c_5105_n N_S[12]_M1188_g
+ N_S[12]_c_5106_n N_S[12]_c_5107_n N_S[12]_M1283_g N_S[12]_c_5117_n
+ N_S[12]_M1201_g N_S[12]_c_5108_n N_S[12]_c_5109_n N_S[12]_c_5110_n
+ N_S[12]_c_5111_n S[12] PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[12]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[5] N_S[5]_c_5217_n N_S[5]_c_5218_n
+ N_S[5]_M1022_g N_S[5]_c_5219_n N_S[5]_M1126_g N_S[5]_c_5220_n N_S[5]_c_5221_n
+ N_S[5]_M1152_g N_S[5]_c_5222_n N_S[5]_c_5242_n N_S[5]_M1256_g N_S[5]_c_5223_n
+ N_S[5]_c_5224_n N_S[5]_c_5225_n N_S[5]_c_5226_n N_S[5]_c_5227_n N_S[5]_M1175_g
+ N_S[5]_c_5228_n N_S[5]_c_5229_n N_S[5]_M1210_g N_S[5]_c_5230_n N_S[5]_c_5231_n
+ N_S[5]_M1220_g N_S[5]_c_5232_n N_S[5]_c_5233_n N_S[5]_M1228_g N_S[5]_c_5234_n
+ N_S[5]_c_5235_n N_S[5]_c_5236_n N_S[5]_c_5237_n S[5] N_S[5]_c_5238_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[13] N_S[13]_c_5337_n N_S[13]_c_5359_n
+ N_S[13]_M1034_g N_S[13]_c_5338_n N_S[13]_M1060_g N_S[13]_c_5339_n
+ N_S[13]_c_5361_n N_S[13]_c_5340_n N_S[13]_c_5341_n N_S[13]_M1211_g
+ N_S[13]_c_5363_n N_S[13]_M1130_g N_S[13]_c_5342_n N_S[13]_c_5343_n
+ N_S[13]_c_5344_n N_S[13]_c_5345_n N_S[13]_c_5346_n N_S[13]_M1149_g
+ N_S[13]_c_5347_n N_S[13]_c_5348_n N_S[13]_M1226_g N_S[13]_c_5349_n
+ N_S[13]_c_5350_n N_S[13]_M1242_g N_S[13]_c_5351_n N_S[13]_c_5352_n
+ N_S[13]_M1290_g N_S[13]_c_5353_n N_S[13]_c_5354_n N_S[13]_c_5355_n
+ N_S[13]_c_5356_n S[13] N_S[13]_c_5357_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_325# N_A_6674_325#_M1126_s
+ N_A_6674_325#_M1022_d N_A_6674_325#_c_5472_n N_A_6674_325#_M1046_g
+ N_A_6674_325#_c_5473_n N_A_6674_325#_c_5465_n N_A_6674_325#_c_5475_n
+ N_A_6674_325#_M1094_g N_A_6674_325#_c_5476_n N_A_6674_325#_c_5477_n
+ N_A_6674_325#_M1261_g N_A_6674_325#_c_5478_n N_A_6674_325#_c_5479_n
+ N_A_6674_325#_M1292_g N_A_6674_325#_c_5480_n N_A_6674_325#_c_5481_n
+ N_A_6674_325#_c_5482_n N_A_6674_325#_c_5466_n N_A_6674_325#_c_5467_n
+ N_A_6674_325#_c_5468_n N_A_6674_325#_c_5484_n N_A_6674_325#_c_5469_n
+ N_A_6674_325#_c_5470_n N_A_6674_325#_c_5471_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_325#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_599# N_A_6674_599#_M1060_s
+ N_A_6674_599#_M1034_s N_A_6674_599#_c_5588_n N_A_6674_599#_M1092_g
+ N_A_6674_599#_c_5589_n N_A_6674_599#_c_5581_n N_A_6674_599#_c_5591_n
+ N_A_6674_599#_M1117_g N_A_6674_599#_c_5592_n N_A_6674_599#_c_5593_n
+ N_A_6674_599#_M1196_g N_A_6674_599#_c_5594_n N_A_6674_599#_c_5595_n
+ N_A_6674_599#_M1238_g N_A_6674_599#_c_5596_n N_A_6674_599#_c_5597_n
+ N_A_6674_599#_c_5598_n N_A_6674_599#_c_5582_n N_A_6674_599#_c_5583_n
+ N_A_6674_599#_c_5599_n N_A_6674_599#_c_5584_n N_A_6674_599#_c_5601_n
+ N_A_6674_599#_c_5585_n N_A_6674_599#_c_5586_n N_A_6674_599#_c_5587_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6674_599#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[5] N_D[5]_M1088_g N_D[5]_M1029_g
+ N_D[5]_M1057_g N_D[5]_M1183_g N_D[5]_M1217_g N_D[5]_M1247_g N_D[5]_M1262_g
+ N_D[5]_M1255_g D[5] N_D[5]_c_5711_n N_D[5]_c_5712_n N_D[5]_c_5713_n
+ N_D[5]_c_5714_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[13] N_D[13]_M1102_g N_D[13]_M1132_g
+ N_D[13]_M1136_g N_D[13]_M1186_g N_D[13]_M1224_g N_D[13]_M1274_g
+ N_D[13]_M1298_g N_D[13]_M1264_g D[13] N_D[13]_c_5804_n N_D[13]_c_5805_n
+ N_D[13]_c_5806_n N_D[13]_c_5807_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[13]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[6] N_D[6]_M1099_g N_D[6]_M1069_g
+ N_D[6]_M1122_g N_D[6]_M1176_g N_D[6]_M1246_g N_D[6]_M1147_g N_D[6]_M1258_g
+ N_D[6]_M1282_g D[6] N_D[6]_c_5895_n N_D[6]_c_5896_n N_D[6]_c_5897_n
+ N_D[6]_c_5898_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[14] N_D[14]_M1109_g N_D[14]_M1004_g
+ N_D[14]_M1179_g N_D[14]_M1184_g N_D[14]_M1251_g N_D[14]_M1189_g
+ N_D[14]_M1305_g N_D[14]_M1293_g D[14] N_D[14]_c_5990_n N_D[14]_c_5991_n
+ N_D[14]_c_5992_n N_D[14]_c_5993_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_265# N_A_8379_265#_M1009_d
+ N_A_8379_265#_M1015_s N_A_8379_265#_c_6080_n N_A_8379_265#_M1081_g
+ N_A_8379_265#_c_6081_n N_A_8379_265#_c_6082_n N_A_8379_265#_c_6083_n
+ N_A_8379_265#_M1168_g N_A_8379_265#_c_6084_n N_A_8379_265#_c_6085_n
+ N_A_8379_265#_M1206_g N_A_8379_265#_c_6086_n N_A_8379_265#_c_6087_n
+ N_A_8379_265#_M1248_g N_A_8379_265#_c_6088_n N_A_8379_265#_c_6089_n
+ N_A_8379_265#_c_6073_n N_A_8379_265#_c_6074_n N_A_8379_265#_c_6075_n
+ N_A_8379_265#_c_6076_n N_A_8379_265#_c_6092_n N_A_8379_265#_c_6077_n
+ N_A_8379_265#_c_6078_n N_A_8379_265#_c_6094_n N_A_8379_265#_c_6079_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_265#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_793# N_A_8379_793#_M1028_d
+ N_A_8379_793#_M1124_s N_A_8379_793#_c_6199_n N_A_8379_793#_M1025_g
+ N_A_8379_793#_c_6200_n N_A_8379_793#_c_6201_n N_A_8379_793#_c_6202_n
+ N_A_8379_793#_M1077_g N_A_8379_793#_c_6203_n N_A_8379_793#_c_6204_n
+ N_A_8379_793#_M1227_g N_A_8379_793#_c_6205_n N_A_8379_793#_c_6206_n
+ N_A_8379_793#_M1314_g N_A_8379_793#_c_6207_n N_A_8379_793#_c_6208_n
+ N_A_8379_793#_c_6192_n N_A_8379_793#_c_6193_n N_A_8379_793#_c_6211_n
+ N_A_8379_793#_c_6212_n N_A_8379_793#_c_6194_n N_A_8379_793#_c_6195_n
+ N_A_8379_793#_c_6213_n N_A_8379_793#_c_6196_n N_A_8379_793#_c_6197_n
+ N_A_8379_793#_c_6198_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_8379_793#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[6] N_S[6]_c_6317_n N_S[6]_M1202_g
+ N_S[6]_c_6318_n N_S[6]_c_6319_n N_S[6]_c_6320_n N_S[6]_M1212_g N_S[6]_c_6321_n
+ N_S[6]_c_6322_n N_S[6]_M1244_g N_S[6]_c_6323_n N_S[6]_c_6324_n N_S[6]_M1254_g
+ N_S[6]_c_6325_n N_S[6]_c_6326_n N_S[6]_c_6327_n N_S[6]_c_6328_n
+ N_S[6]_c_6329_n N_S[6]_c_6340_n N_S[6]_M1015_g N_S[6]_c_6330_n N_S[6]_M1009_g
+ N_S[6]_c_6331_n N_S[6]_c_6332_n N_S[6]_M1075_g N_S[6]_c_6333_n N_S[6]_M1063_g
+ N_S[6]_c_6334_n N_S[6]_c_6335_n N_S[6]_c_6336_n N_S[6]_c_6337_n S[6]
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[14] N_S[14]_c_6434_n N_S[14]_M1005_g
+ N_S[14]_c_6435_n N_S[14]_c_6436_n N_S[14]_c_6437_n N_S[14]_M1064_g
+ N_S[14]_c_6438_n N_S[14]_c_6439_n N_S[14]_M1162_g N_S[14]_c_6440_n
+ N_S[14]_c_6441_n N_S[14]_M1230_g N_S[14]_c_6442_n N_S[14]_c_6443_n
+ N_S[14]_c_6444_n N_S[14]_c_6445_n N_S[14]_c_6455_n N_S[14]_c_6446_n
+ N_S[14]_c_6457_n N_S[14]_M1124_g N_S[14]_c_6447_n N_S[14]_M1028_g
+ N_S[14]_c_6448_n N_S[14]_c_6449_n N_S[14]_M1097_g N_S[14]_c_6459_n
+ N_S[14]_M1170_g N_S[14]_c_6450_n N_S[14]_c_6451_n N_S[14]_c_6452_n
+ N_S[14]_c_6453_n S[14] PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[14]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[7] N_S[7]_c_6559_n N_S[7]_c_6560_n
+ N_S[7]_M1142_g N_S[7]_c_6561_n N_S[7]_M1141_g N_S[7]_c_6562_n N_S[7]_c_6563_n
+ N_S[7]_M1198_g N_S[7]_c_6564_n N_S[7]_c_6584_n N_S[7]_M1185_g N_S[7]_c_6565_n
+ N_S[7]_c_6566_n N_S[7]_c_6567_n N_S[7]_c_6568_n N_S[7]_c_6569_n N_S[7]_M1003_g
+ N_S[7]_c_6570_n N_S[7]_c_6571_n N_S[7]_M1209_g N_S[7]_c_6572_n N_S[7]_c_6573_n
+ N_S[7]_M1253_g N_S[7]_c_6574_n N_S[7]_c_6575_n N_S[7]_M1272_g N_S[7]_c_6576_n
+ N_S[7]_c_6577_n N_S[7]_c_6578_n N_S[7]_c_6579_n S[7] N_S[7]_c_6580_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[15] N_S[15]_c_6679_n N_S[15]_c_6701_n
+ N_S[15]_M1233_g N_S[15]_c_6680_n N_S[15]_M1174_g N_S[15]_c_6681_n
+ N_S[15]_c_6703_n N_S[15]_c_6682_n N_S[15]_c_6683_n N_S[15]_M1223_g
+ N_S[15]_c_6705_n N_S[15]_M1279_g N_S[15]_c_6684_n N_S[15]_c_6685_n
+ N_S[15]_c_6686_n N_S[15]_c_6687_n N_S[15]_c_6688_n N_S[15]_M1104_g
+ N_S[15]_c_6689_n N_S[15]_c_6690_n N_S[15]_M1169_g N_S[15]_c_6691_n
+ N_S[15]_c_6692_n N_S[15]_M1197_g N_S[15]_c_6693_n N_S[15]_c_6694_n
+ N_S[15]_M1252_g N_S[15]_c_6695_n N_S[15]_c_6696_n N_S[15]_c_6697_n
+ N_S[15]_c_6698_n S[15] N_S[15]_c_6699_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%S[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_325# N_A_9250_325#_M1141_d
+ N_A_9250_325#_M1142_s N_A_9250_325#_c_6814_n N_A_9250_325#_M1013_g
+ N_A_9250_325#_c_6815_n N_A_9250_325#_c_6807_n N_A_9250_325#_c_6817_n
+ N_A_9250_325#_M1058_g N_A_9250_325#_c_6818_n N_A_9250_325#_c_6819_n
+ N_A_9250_325#_M1153_g N_A_9250_325#_c_6820_n N_A_9250_325#_c_6821_n
+ N_A_9250_325#_M1163_g N_A_9250_325#_c_6822_n N_A_9250_325#_c_6823_n
+ N_A_9250_325#_c_6824_n N_A_9250_325#_c_6808_n N_A_9250_325#_c_6809_n
+ N_A_9250_325#_c_6810_n N_A_9250_325#_c_6826_n N_A_9250_325#_c_6811_n
+ N_A_9250_325#_c_6812_n N_A_9250_325#_c_6813_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_325#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_599# N_A_9250_599#_M1174_d
+ N_A_9250_599#_M1233_s N_A_9250_599#_c_6929_n N_A_9250_599#_M1166_g
+ N_A_9250_599#_c_6930_n N_A_9250_599#_c_6922_n N_A_9250_599#_c_6932_n
+ N_A_9250_599#_M1204_g N_A_9250_599#_c_6933_n N_A_9250_599#_c_6934_n
+ N_A_9250_599#_M1286_g N_A_9250_599#_c_6935_n N_A_9250_599#_c_6936_n
+ N_A_9250_599#_M1303_g N_A_9250_599#_c_6937_n N_A_9250_599#_c_6938_n
+ N_A_9250_599#_c_6939_n N_A_9250_599#_c_6923_n N_A_9250_599#_c_6924_n
+ N_A_9250_599#_c_6940_n N_A_9250_599#_c_6925_n N_A_9250_599#_c_6942_n
+ N_A_9250_599#_c_6926_n N_A_9250_599#_c_6927_n N_A_9250_599#_c_6928_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9250_599#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[7] N_D[7]_M1040_g N_D[7]_M1068_g
+ N_D[7]_M1115_g N_D[7]_M1087_g N_D[7]_M1131_g N_D[7]_M1216_g N_D[7]_M1281_g
+ N_D[7]_M1151_g D[7] N_D[7]_c_7051_n N_D[7]_c_7052_n N_D[7]_c_7053_n
+ N_D[7]_c_7054_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[15] N_D[15]_M1056_g N_D[15]_M1073_g
+ N_D[15]_M1144_g N_D[15]_M1103_g N_D[15]_M1145_g N_D[15]_M1190_g
+ N_D[15]_M1278_g N_D[15]_M1156_g D[15] N_D[15]_c_7139_n N_D[15]_c_7140_n
+ N_D[15]_c_7141_n N_D[15]_c_7142_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%D[15]
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPWR N_VPWR_M1014_d N_VPWR_M1023_d
+ N_VPWR_M1146_d N_VPWR_M1155_d N_VPWR_M1294_d N_VPWR_M1304_d N_VPWR_M1018_d
+ N_VPWR_M1123_d N_VPWR_M1061_d N_VPWR_M1172_d N_VPWR_M1133_d N_VPWR_M1225_d
+ N_VPWR_M1180_d N_VPWR_M1266_d N_VPWR_M1002_s N_VPWR_M1011_s N_VPWR_M1038_s
+ N_VPWR_M1051_s N_VPWR_M1271_s N_VPWR_M1285_s N_VPWR_M1020_s N_VPWR_M1024_s
+ N_VPWR_M1067_s N_VPWR_M1076_s N_VPWR_M1301_s N_VPWR_M1309_s N_VPWR_M1065_s
+ N_VPWR_M1083_d N_VPWR_M1308_s N_VPWR_M1173_d N_VPWR_M1150_s N_VPWR_M1066_d
+ N_VPWR_M1280_s N_VPWR_M1237_d N_VPWR_M1042_d N_VPWR_M1052_d N_VPWR_M1089_d
+ N_VPWR_M1101_d N_VPWR_M1289_d N_VPWR_M1297_d N_VPWR_M1158_d N_VPWR_M1006_s
+ N_VPWR_M1194_d N_VPWR_M1165_s N_VPWR_M1319_d N_VPWR_M1277_s N_VPWR_M1016_d
+ N_VPWR_M1120_d N_VPWR_M1095_d N_VPWR_M1201_d N_VPWR_M1022_s N_VPWR_M1034_d
+ N_VPWR_M1256_s N_VPWR_M1130_d N_VPWR_M1088_d N_VPWR_M1102_d N_VPWR_M1183_d
+ N_VPWR_M1186_d N_VPWR_M1255_d N_VPWR_M1264_d N_VPWR_M1099_d N_VPWR_M1109_d
+ N_VPWR_M1176_d N_VPWR_M1184_d N_VPWR_M1282_d N_VPWR_M1293_d N_VPWR_M1015_d
+ N_VPWR_M1124_d N_VPWR_M1063_d N_VPWR_M1170_d N_VPWR_M1142_d N_VPWR_M1233_d
+ N_VPWR_M1185_d N_VPWR_M1279_d N_VPWR_M1040_d N_VPWR_M1056_d N_VPWR_M1087_d
+ N_VPWR_M1103_d N_VPWR_M1151_d N_VPWR_M1156_d N_VPWR_c_7217_n N_VPWR_c_7218_n
+ N_VPWR_c_7219_n N_VPWR_c_7220_n N_VPWR_c_7221_n N_VPWR_c_7222_n
+ N_VPWR_c_7223_n N_VPWR_c_7224_n N_VPWR_c_7225_n N_VPWR_c_7226_n
+ N_VPWR_c_7227_n N_VPWR_c_7228_n N_VPWR_c_7229_n N_VPWR_c_7230_n
+ N_VPWR_c_7231_n N_VPWR_c_7232_n N_VPWR_c_7233_n N_VPWR_c_7234_n
+ N_VPWR_c_7235_n N_VPWR_c_7236_n N_VPWR_c_7237_n N_VPWR_c_7238_n
+ N_VPWR_c_7239_n N_VPWR_c_7240_n N_VPWR_c_7241_n N_VPWR_c_7242_n
+ N_VPWR_c_7243_n N_VPWR_c_7244_n N_VPWR_c_7245_n N_VPWR_c_7246_n
+ N_VPWR_c_7247_n N_VPWR_c_7248_n N_VPWR_c_7249_n N_VPWR_c_7250_n
+ N_VPWR_c_7251_n N_VPWR_c_7252_n N_VPWR_c_7253_n N_VPWR_c_7254_n
+ N_VPWR_c_7255_n N_VPWR_c_7256_n N_VPWR_c_7257_n N_VPWR_c_7258_n
+ N_VPWR_c_7259_n N_VPWR_c_7260_n N_VPWR_c_7262_n N_VPWR_c_7264_n
+ N_VPWR_c_7266_n N_VPWR_c_7268_n N_VPWR_c_7269_n N_VPWR_c_7270_n
+ N_VPWR_c_7271_n N_VPWR_c_7272_n N_VPWR_c_7273_n N_VPWR_c_7274_n
+ N_VPWR_c_7275_n N_VPWR_c_7276_n N_VPWR_c_7277_n N_VPWR_c_7278_n
+ N_VPWR_c_7279_n N_VPWR_c_7280_n N_VPWR_c_7281_n N_VPWR_c_7282_n
+ N_VPWR_c_7283_n N_VPWR_c_7284_n N_VPWR_c_7285_n N_VPWR_c_7286_n
+ N_VPWR_c_7287_n N_VPWR_c_7288_n N_VPWR_c_7289_n N_VPWR_c_7290_n
+ N_VPWR_c_7291_n N_VPWR_c_7292_n N_VPWR_c_7293_n N_VPWR_c_7294_n
+ N_VPWR_c_7295_n N_VPWR_c_7296_n N_VPWR_c_7297_n N_VPWR_c_7298_n
+ N_VPWR_c_7299_n N_VPWR_c_7300_n N_VPWR_c_7301_n N_VPWR_c_7302_n
+ N_VPWR_c_7303_n N_VPWR_c_7304_n N_VPWR_c_7305_n N_VPWR_c_7306_n
+ N_VPWR_c_7307_n N_VPWR_c_7308_n N_VPWR_c_7309_n N_VPWR_c_7310_n
+ N_VPWR_c_7311_n N_VPWR_c_7312_n N_VPWR_c_7313_n N_VPWR_c_7314_n
+ N_VPWR_c_7315_n N_VPWR_c_7316_n N_VPWR_c_7317_n N_VPWR_c_7318_n
+ N_VPWR_c_7319_n N_VPWR_c_7320_n N_VPWR_c_7321_n N_VPWR_c_7322_n
+ N_VPWR_c_7323_n N_VPWR_c_7324_n N_VPWR_c_7325_n N_VPWR_c_7326_n
+ N_VPWR_c_7327_n N_VPWR_c_7328_n N_VPWR_c_7329_n N_VPWR_c_7330_n
+ N_VPWR_c_7331_n N_VPWR_c_7332_n N_VPWR_c_7333_n N_VPWR_c_7334_n
+ N_VPWR_c_7335_n N_VPWR_c_7336_n N_VPWR_c_7337_n N_VPWR_c_7338_n
+ N_VPWR_c_7339_n N_VPWR_c_7340_n N_VPWR_c_7341_n N_VPWR_c_7342_n
+ N_VPWR_c_7343_n N_VPWR_c_7344_n N_VPWR_c_7345_n N_VPWR_c_7346_n VPWR VPWR VPWR
+ VPWR VPWR VPWR VPWR VPWR VPWR N_VPWR_c_7350_n N_VPWR_c_7351_n N_VPWR_c_7352_n
+ N_VPWR_c_7353_n N_VPWR_c_7354_n N_VPWR_c_7355_n N_VPWR_c_7356_n
+ N_VPWR_c_7357_n N_VPWR_c_7358_n N_VPWR_c_7361_n N_VPWR_c_7362_n
+ N_VPWR_c_7363_n N_VPWR_c_7364_n N_VPWR_c_7365_n N_VPWR_c_7366_n
+ N_VPWR_c_7367_n N_VPWR_c_7368_n N_VPWR_c_7369_n N_VPWR_c_7370_n
+ N_VPWR_c_7371_n N_VPWR_c_7372_n N_VPWR_c_7373_n N_VPWR_c_7374_n
+ N_VPWR_c_7375_n N_VPWR_c_7376_n N_VPWR_c_7377_n N_VPWR_c_7378_n
+ N_VPWR_c_7379_n N_VPWR_c_7380_n N_VPWR_c_7381_n N_VPWR_c_7382_n
+ N_VPWR_c_7383_n N_VPWR_c_7384_n N_VPWR_c_7385_n N_VPWR_c_7386_n
+ N_VPWR_c_7387_n N_VPWR_c_7388_n N_VPWR_c_7389_n N_VPWR_c_7390_n
+ N_VPWR_c_7391_n N_VPWR_c_7392_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_297# N_A_117_297#_M1014_s
+ N_A_117_297#_M1208_s N_A_117_297#_M1137_d N_A_117_297#_M1207_d
+ N_A_117_297#_M1299_d N_A_117_297#_c_8776_n N_A_117_297#_c_8771_n
+ N_A_117_297#_c_8781_n N_A_117_297#_c_8785_n N_A_117_297#_c_8789_n
+ N_A_117_297#_c_8825_n N_A_117_297#_c_8772_n N_A_117_297#_c_8832_n
+ N_A_117_297#_c_8800_n N_A_117_297#_c_8836_n N_A_117_297#_c_8802_n
+ N_A_117_297#_c_8839_n N_A_117_297#_c_8792_n N_A_117_297#_c_8795_n
+ N_A_117_297#_c_8847_n N_A_117_297#_c_8773_n N_A_117_297#_c_8774_n
+ N_A_117_297#_c_8775_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_591# N_A_117_591#_M1023_s
+ N_A_117_591#_M1221_s N_A_117_591#_M1026_s N_A_117_591#_M1079_s
+ N_A_117_591#_M1269_s N_A_117_591#_c_8892_n N_A_117_591#_c_8887_n
+ N_A_117_591#_c_8897_n N_A_117_591#_c_8901_n N_A_117_591#_c_8905_n
+ N_A_117_591#_c_8941_n N_A_117_591#_c_8888_n N_A_117_591#_c_8948_n
+ N_A_117_591#_c_8916_n N_A_117_591#_c_8952_n N_A_117_591#_c_8918_n
+ N_A_117_591#_c_8955_n N_A_117_591#_c_8956_n N_A_117_591#_c_8908_n
+ N_A_117_591#_c_8911_n N_A_117_591#_c_8889_n N_A_117_591#_c_8890_n
+ N_A_117_591#_c_8891_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_117_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%Z N_Z_M1053_s N_Z_M1070_d N_Z_M1105_s
+ N_Z_M1236_d N_Z_M1039_d N_Z_M1027_d N_Z_M1093_d N_Z_M1096_d N_Z_M1035_d
+ N_Z_M1010_s N_Z_M1108_d N_Z_M1263_s N_Z_M1030_s N_Z_M1047_s N_Z_M1059_s
+ N_Z_M1316_s N_Z_M1154_d N_Z_M1044_s N_Z_M1205_d N_Z_M1218_s N_Z_M1175_s
+ N_Z_M1149_s N_Z_M1220_s N_Z_M1242_s N_Z_M1202_s N_Z_M1005_s N_Z_M1244_s
+ N_Z_M1162_s N_Z_M1003_s N_Z_M1104_d N_Z_M1253_s N_Z_M1197_d N_Z_M1137_s
+ N_Z_M1026_d N_Z_M1249_s N_Z_M1127_d N_Z_M1007_d N_Z_M1112_s N_Z_M1140_d
+ N_Z_M1199_s N_Z_M1082_s N_Z_M1000_s N_Z_M1181_s N_Z_M1229_s N_Z_M1121_s
+ N_Z_M1071_s N_Z_M1243_s N_Z_M1260_s N_Z_M1050_s N_Z_M1055_d N_Z_M1231_s
+ N_Z_M1200_d N_Z_M1046_d N_Z_M1092_d N_Z_M1261_d N_Z_M1196_d N_Z_M1081_s
+ N_Z_M1025_s N_Z_M1206_s N_Z_M1227_s N_Z_M1013_d N_Z_M1166_d N_Z_M1153_d
+ N_Z_M1286_d N_Z_c_9003_n N_Z_c_9004_n N_Z_c_9005_n N_Z_c_9006_n N_Z_c_9007_n
+ N_Z_c_9008_n N_Z_c_9009_n N_Z_c_9010_n N_Z_c_9011_n N_Z_c_9012_n N_Z_c_9013_n
+ N_Z_c_9014_n N_Z_c_9015_n N_Z_c_9016_n N_Z_c_9017_n N_Z_c_9018_n N_Z_c_9019_n
+ N_Z_c_9020_n N_Z_c_9021_n N_Z_c_9022_n N_Z_c_9023_n N_Z_c_9024_n N_Z_c_9025_n
+ N_Z_c_9026_n N_Z_c_9027_n N_Z_c_9028_n N_Z_c_9029_n N_Z_c_9030_n N_Z_c_9031_n
+ N_Z_c_9032_n N_Z_c_9033_n N_Z_c_9034_n N_Z_c_9035_n N_Z_c_9036_n N_Z_c_9037_n
+ N_Z_c_9038_n N_Z_c_9039_n N_Z_c_9040_n N_Z_c_9041_n N_Z_c_9042_n N_Z_c_9043_n
+ N_Z_c_9044_n N_Z_c_9045_n N_Z_c_9046_n N_Z_c_9047_n N_Z_c_9048_n N_Z_c_9049_n
+ N_Z_c_9050_n N_Z_c_9051_n N_Z_c_9052_n N_Z_c_9053_n N_Z_c_9054_n N_Z_c_9055_n
+ N_Z_c_9056_n N_Z_c_9057_n N_Z_c_9058_n N_Z_c_9059_n N_Z_c_9060_n N_Z_c_9061_n
+ N_Z_c_9062_n N_Z_c_9063_n N_Z_c_9064_n N_Z_c_9065_n N_Z_c_9066_n N_Z_c_9067_n
+ N_Z_c_9068_n N_Z_c_9069_n N_Z_c_9070_n N_Z_c_9071_n N_Z_c_9072_n N_Z_c_9073_n
+ N_Z_c_9074_n N_Z_c_9075_n N_Z_c_9076_n N_Z_c_9077_n N_Z_c_9078_n N_Z_c_9079_n
+ N_Z_c_9080_n N_Z_c_9081_n N_Z_c_9082_n N_Z_c_9083_n N_Z_c_9084_n N_Z_c_9085_n
+ N_Z_c_9086_n N_Z_c_9087_n N_Z_c_9088_n N_Z_c_9089_n N_Z_c_9090_n N_Z_c_9091_n
+ N_Z_c_9092_n N_Z_c_9093_n N_Z_c_9094_n N_Z_c_9095_n N_Z_c_9096_n N_Z_c_9097_n
+ N_Z_c_9098_n N_Z_c_9115_n N_Z_c_10135_n N_Z_c_9116_n N_Z_c_10163_n
+ N_Z_c_9117_n N_Z_c_10198_p N_Z_c_9118_n N_Z_c_10238_p N_Z_c_9119_n
+ N_Z_c_10282_p N_Z_c_9120_n N_Z_c_10322_p N_Z_c_9121_n N_Z_c_10358_p
+ N_Z_c_9123_n N_Z_c_10398_p N_Z_c_9125_n N_Z_c_10442_p N_Z_c_9126_n
+ N_Z_c_10482_p N_Z_c_9127_n N_Z_c_10518_p N_Z_c_9128_n N_Z_c_10558_p
+ N_Z_c_9129_n N_Z_c_10602_p N_Z_c_9130_n N_Z_c_10642_p N_Z_c_9288_n
+ N_Z_c_9317_n N_Z_c_10276_p N_Z_c_10316_p N_Z_c_9494_n N_Z_c_9523_n
+ N_Z_c_10436_p N_Z_c_10476_p N_Z_c_9700_n N_Z_c_9729_n N_Z_c_10596_p
+ N_Z_c_10636_p N_Z_c_9905_n N_Z_c_10675_p N_Z_c_9933_n N_Z_c_10703_p Z Z Z Z Z
+ Z Z Z Z Z Z Z Z Z Z Z Z Z N_Z_c_9131_n N_Z_c_9132_n N_Z_c_9133_n N_Z_c_9134_n
+ N_Z_c_9135_n N_Z_c_9136_n N_Z_c_9137_n N_Z_c_9138_n N_Z_c_9139_n N_Z_c_9140_n
+ N_Z_c_9141_n N_Z_c_9142_n N_Z_c_9143_n N_Z_c_9144_n N_Z_c_9145_n N_Z_c_9146_n
+ N_Z_c_10154_n N_Z_c_10182_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%Z
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_311# N_A_1643_311#_M1007_s
+ N_A_1643_311#_M1048_s N_A_1643_311#_M1284_s N_A_1643_311#_M1002_d
+ N_A_1643_311#_M1134_d N_A_1643_311#_c_10897_n N_A_1643_311#_c_10898_n
+ N_A_1643_311#_c_10919_n N_A_1643_311#_c_10923_n N_A_1643_311#_c_10927_n
+ N_A_1643_311#_c_10906_n N_A_1643_311#_c_10948_n N_A_1643_311#_c_10908_n
+ N_A_1643_311#_c_10951_n N_A_1643_311#_c_10899_n N_A_1643_311#_c_10956_n
+ N_A_1643_311#_c_10932_n N_A_1643_311#_c_10962_n N_A_1643_311#_c_10934_n
+ N_A_1643_311#_c_10969_n N_A_1643_311#_c_10937_n N_A_1643_311#_c_10900_n
+ N_A_1643_311#_c_10901_n N_A_1643_311#_c_10902_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_311#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_613# N_A_1643_613#_M1112_d
+ N_A_1643_613#_M1161_d N_A_1643_613#_M1273_d N_A_1643_613#_M1011_d
+ N_A_1643_613#_M1148_d N_A_1643_613#_c_11028_n N_A_1643_613#_c_11029_n
+ N_A_1643_613#_c_11050_n N_A_1643_613#_c_11054_n N_A_1643_613#_c_11058_n
+ N_A_1643_613#_c_11037_n N_A_1643_613#_c_11079_n N_A_1643_613#_c_11039_n
+ N_A_1643_613#_c_11082_n N_A_1643_613#_c_11030_n N_A_1643_613#_c_11087_n
+ N_A_1643_613#_c_11063_n N_A_1643_613#_c_11093_n N_A_1643_613#_c_11096_n
+ N_A_1643_613#_c_11031_n N_A_1643_613#_c_11032_n N_A_1643_613#_c_11033_n
+ N_A_1643_613#_c_11066_n N_A_1643_613#_c_11069_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1643_613#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_297# N_A_2693_297#_M1020_d
+ N_A_2693_297#_M1157_d N_A_2693_297#_M1082_d N_A_2693_297#_M1138_d
+ N_A_2693_297#_M1250_d N_A_2693_297#_c_11164_n N_A_2693_297#_c_11159_n
+ N_A_2693_297#_c_11169_n N_A_2693_297#_c_11173_n N_A_2693_297#_c_11177_n
+ N_A_2693_297#_c_11212_n N_A_2693_297#_c_11160_n N_A_2693_297#_c_11219_n
+ N_A_2693_297#_c_11188_n N_A_2693_297#_c_11223_n N_A_2693_297#_c_11190_n
+ N_A_2693_297#_c_11226_n N_A_2693_297#_c_11180_n N_A_2693_297#_c_11183_n
+ N_A_2693_297#_c_11235_n N_A_2693_297#_c_11161_n N_A_2693_297#_c_11162_n
+ N_A_2693_297#_c_11163_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_591# N_A_2693_591#_M1024_d
+ N_A_2693_591#_M1164_d N_A_2693_591#_M1000_d N_A_2693_591#_M1080_d
+ N_A_2693_591#_M1270_d N_A_2693_591#_c_11292_n N_A_2693_591#_c_11287_n
+ N_A_2693_591#_c_11297_n N_A_2693_591#_c_11301_n N_A_2693_591#_c_11305_n
+ N_A_2693_591#_c_11340_n N_A_2693_591#_c_11288_n N_A_2693_591#_c_11347_n
+ N_A_2693_591#_c_11316_n N_A_2693_591#_c_11351_n N_A_2693_591#_c_11318_n
+ N_A_2693_591#_c_11354_n N_A_2693_591#_c_11355_n N_A_2693_591#_c_11308_n
+ N_A_2693_591#_c_11311_n N_A_2693_591#_c_11289_n N_A_2693_591#_c_11290_n
+ N_A_2693_591#_c_11291_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2693_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_311# N_A_4219_311#_M1121_d
+ N_A_4219_311#_M1171_d N_A_4219_311#_M1287_d N_A_4219_311#_M1042_s
+ N_A_4219_311#_M1116_s N_A_4219_311#_c_11415_n N_A_4219_311#_c_11416_n
+ N_A_4219_311#_c_11437_n N_A_4219_311#_c_11441_n N_A_4219_311#_c_11445_n
+ N_A_4219_311#_c_11424_n N_A_4219_311#_c_11466_n N_A_4219_311#_c_11426_n
+ N_A_4219_311#_c_11469_n N_A_4219_311#_c_11417_n N_A_4219_311#_c_11474_n
+ N_A_4219_311#_c_11450_n N_A_4219_311#_c_11480_n N_A_4219_311#_c_11452_n
+ N_A_4219_311#_c_11487_n N_A_4219_311#_c_11455_n N_A_4219_311#_c_11418_n
+ N_A_4219_311#_c_11419_n N_A_4219_311#_c_11420_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_311#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_613# N_A_4219_613#_M1071_d
+ N_A_4219_613#_M1114_d N_A_4219_613#_M1313_d N_A_4219_613#_M1052_s
+ N_A_4219_613#_M1129_s N_A_4219_613#_c_11546_n N_A_4219_613#_c_11547_n
+ N_A_4219_613#_c_11568_n N_A_4219_613#_c_11572_n N_A_4219_613#_c_11576_n
+ N_A_4219_613#_c_11555_n N_A_4219_613#_c_11597_n N_A_4219_613#_c_11557_n
+ N_A_4219_613#_c_11600_n N_A_4219_613#_c_11548_n N_A_4219_613#_c_11605_n
+ N_A_4219_613#_c_11581_n N_A_4219_613#_c_11611_n N_A_4219_613#_c_11614_n
+ N_A_4219_613#_c_11549_n N_A_4219_613#_c_11550_n N_A_4219_613#_c_11551_n
+ N_A_4219_613#_c_11584_n N_A_4219_613#_c_11587_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4219_613#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_297# N_A_5361_297#_M1158_s
+ N_A_5361_297#_M1265_s N_A_5361_297#_M1050_d N_A_5361_297#_M1118_d
+ N_A_5361_297#_M1295_d N_A_5361_297#_c_11682_n N_A_5361_297#_c_11677_n
+ N_A_5361_297#_c_11687_n N_A_5361_297#_c_11691_n N_A_5361_297#_c_11695_n
+ N_A_5361_297#_c_11730_n N_A_5361_297#_c_11678_n N_A_5361_297#_c_11737_n
+ N_A_5361_297#_c_11706_n N_A_5361_297#_c_11741_n N_A_5361_297#_c_11708_n
+ N_A_5361_297#_c_11744_n N_A_5361_297#_c_11698_n N_A_5361_297#_c_11701_n
+ N_A_5361_297#_c_11753_n N_A_5361_297#_c_11679_n N_A_5361_297#_c_11680_n
+ N_A_5361_297#_c_11681_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_591# N_A_5361_591#_M1006_d
+ N_A_5361_591#_M1203_d N_A_5361_591#_M1055_s N_A_5361_591#_M1119_s
+ N_A_5361_591#_M1257_s N_A_5361_591#_c_11810_n N_A_5361_591#_c_11805_n
+ N_A_5361_591#_c_11815_n N_A_5361_591#_c_11819_n N_A_5361_591#_c_11823_n
+ N_A_5361_591#_c_11858_n N_A_5361_591#_c_11806_n N_A_5361_591#_c_11865_n
+ N_A_5361_591#_c_11834_n N_A_5361_591#_c_11869_n N_A_5361_591#_c_11836_n
+ N_A_5361_591#_c_11872_n N_A_5361_591#_c_11873_n N_A_5361_591#_c_11826_n
+ N_A_5361_591#_c_11829_n N_A_5361_591#_c_11807_n N_A_5361_591#_c_11808_n
+ N_A_5361_591#_c_11809_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5361_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_311# N_A_6887_311#_M1046_s
+ N_A_6887_311#_M1094_s N_A_6887_311#_M1292_s N_A_6887_311#_M1088_s
+ N_A_6887_311#_M1217_s N_A_6887_311#_c_11933_n N_A_6887_311#_c_11934_n
+ N_A_6887_311#_c_11955_n N_A_6887_311#_c_11959_n N_A_6887_311#_c_11963_n
+ N_A_6887_311#_c_11942_n N_A_6887_311#_c_11984_n N_A_6887_311#_c_11944_n
+ N_A_6887_311#_c_11987_n N_A_6887_311#_c_11935_n N_A_6887_311#_c_11992_n
+ N_A_6887_311#_c_11968_n N_A_6887_311#_c_11998_n N_A_6887_311#_c_11970_n
+ N_A_6887_311#_c_12005_n N_A_6887_311#_c_11973_n N_A_6887_311#_c_11936_n
+ N_A_6887_311#_c_11937_n N_A_6887_311#_c_11938_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_311#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_613# N_A_6887_613#_M1092_s
+ N_A_6887_613#_M1117_s N_A_6887_613#_M1238_s N_A_6887_613#_M1102_s
+ N_A_6887_613#_M1224_s N_A_6887_613#_c_12064_n N_A_6887_613#_c_12065_n
+ N_A_6887_613#_c_12086_n N_A_6887_613#_c_12090_n N_A_6887_613#_c_12094_n
+ N_A_6887_613#_c_12073_n N_A_6887_613#_c_12115_n N_A_6887_613#_c_12075_n
+ N_A_6887_613#_c_12118_n N_A_6887_613#_c_12066_n N_A_6887_613#_c_12123_n
+ N_A_6887_613#_c_12099_n N_A_6887_613#_c_12129_n N_A_6887_613#_c_12132_n
+ N_A_6887_613#_c_12067_n N_A_6887_613#_c_12068_n N_A_6887_613#_c_12069_n
+ N_A_6887_613#_c_12102_n N_A_6887_613#_c_12105_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6887_613#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_297# N_A_7937_297#_M1099_s
+ N_A_7937_297#_M1246_s N_A_7937_297#_M1081_d N_A_7937_297#_M1168_d
+ N_A_7937_297#_M1248_d N_A_7937_297#_c_12200_n N_A_7937_297#_c_12195_n
+ N_A_7937_297#_c_12205_n N_A_7937_297#_c_12209_n N_A_7937_297#_c_12213_n
+ N_A_7937_297#_c_12248_n N_A_7937_297#_c_12196_n N_A_7937_297#_c_12255_n
+ N_A_7937_297#_c_12224_n N_A_7937_297#_c_12259_n N_A_7937_297#_c_12226_n
+ N_A_7937_297#_c_12262_n N_A_7937_297#_c_12216_n N_A_7937_297#_c_12219_n
+ N_A_7937_297#_c_12271_n N_A_7937_297#_c_12197_n N_A_7937_297#_c_12198_n
+ N_A_7937_297#_c_12199_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_297#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_591# N_A_7937_591#_M1109_s
+ N_A_7937_591#_M1251_s N_A_7937_591#_M1025_d N_A_7937_591#_M1077_d
+ N_A_7937_591#_M1314_d N_A_7937_591#_c_12328_n N_A_7937_591#_c_12323_n
+ N_A_7937_591#_c_12333_n N_A_7937_591#_c_12337_n N_A_7937_591#_c_12341_n
+ N_A_7937_591#_c_12376_n N_A_7937_591#_c_12324_n N_A_7937_591#_c_12383_n
+ N_A_7937_591#_c_12352_n N_A_7937_591#_c_12387_n N_A_7937_591#_c_12354_n
+ N_A_7937_591#_c_12390_n N_A_7937_591#_c_12391_n N_A_7937_591#_c_12344_n
+ N_A_7937_591#_c_12347_n N_A_7937_591#_c_12325_n N_A_7937_591#_c_12326_n
+ N_A_7937_591#_c_12327_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7937_591#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_311# N_A_9463_311#_M1013_s
+ N_A_9463_311#_M1058_s N_A_9463_311#_M1163_s N_A_9463_311#_M1040_s
+ N_A_9463_311#_M1131_s N_A_9463_311#_c_12451_n N_A_9463_311#_c_12452_n
+ N_A_9463_311#_c_12473_n N_A_9463_311#_c_12477_n N_A_9463_311#_c_12481_n
+ N_A_9463_311#_c_12460_n N_A_9463_311#_c_12502_n N_A_9463_311#_c_12462_n
+ N_A_9463_311#_c_12505_n N_A_9463_311#_c_12453_n N_A_9463_311#_c_12510_n
+ N_A_9463_311#_c_12486_n N_A_9463_311#_c_12517_n N_A_9463_311#_c_12488_n
+ N_A_9463_311#_c_12524_n N_A_9463_311#_c_12491_n N_A_9463_311#_c_12454_n
+ N_A_9463_311#_c_12455_n N_A_9463_311#_c_12456_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_311#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_613# N_A_9463_613#_M1166_s
+ N_A_9463_613#_M1204_s N_A_9463_613#_M1303_s N_A_9463_613#_M1056_s
+ N_A_9463_613#_M1145_s N_A_9463_613#_c_12570_n N_A_9463_613#_c_12571_n
+ N_A_9463_613#_c_12592_n N_A_9463_613#_c_12596_n N_A_9463_613#_c_12600_n
+ N_A_9463_613#_c_12579_n N_A_9463_613#_c_12621_n N_A_9463_613#_c_12581_n
+ N_A_9463_613#_c_12624_n N_A_9463_613#_c_12572_n N_A_9463_613#_c_12629_n
+ N_A_9463_613#_c_12605_n N_A_9463_613#_c_12636_n N_A_9463_613#_c_12639_n
+ N_A_9463_613#_c_12573_n N_A_9463_613#_c_12574_n N_A_9463_613#_c_12575_n
+ N_A_9463_613#_c_12608_n N_A_9463_613#_c_12611_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9463_613#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VGND N_VGND_M1084_d N_VGND_M1085_d
+ N_VGND_M1219_d N_VGND_M1090_d N_VGND_M1317_d N_VGND_M1240_d N_VGND_M1139_s
+ N_VGND_M1017_s N_VGND_M1192_s N_VGND_M1078_s N_VGND_M1241_d N_VGND_M1008_s
+ N_VGND_M1288_d N_VGND_M1107_s N_VGND_M1049_d N_VGND_M1019_d N_VGND_M1098_d
+ N_VGND_M1111_d N_VGND_M1315_d N_VGND_M1276_d N_VGND_M1001_s N_VGND_M1033_d
+ N_VGND_M1062_s N_VGND_M1143_d N_VGND_M1182_s N_VGND_M1307_d N_VGND_M1222_d
+ N_VGND_M1043_s N_VGND_M1239_d N_VGND_M1215_s N_VGND_M1234_d N_VGND_M1054_d
+ N_VGND_M1291_d N_VGND_M1072_d N_VGND_M1041_d N_VGND_M1245_s N_VGND_M1100_d
+ N_VGND_M1296_s N_VGND_M1193_d N_VGND_M1311_s N_VGND_M1021_d N_VGND_M1012_d
+ N_VGND_M1177_d N_VGND_M1128_d N_VGND_M1275_d N_VGND_M1267_d N_VGND_M1037_d
+ N_VGND_M1188_s N_VGND_M1086_d N_VGND_M1283_s N_VGND_M1126_d N_VGND_M1060_d
+ N_VGND_M1152_d N_VGND_M1211_d N_VGND_M1029_d N_VGND_M1132_d N_VGND_M1057_d
+ N_VGND_M1136_d N_VGND_M1262_d N_VGND_M1298_d N_VGND_M1069_s N_VGND_M1004_s
+ N_VGND_M1122_s N_VGND_M1179_s N_VGND_M1258_s N_VGND_M1305_s N_VGND_M1009_s
+ N_VGND_M1028_s N_VGND_M1075_s N_VGND_M1097_s N_VGND_M1141_s N_VGND_M1174_s
+ N_VGND_M1198_s N_VGND_M1223_s N_VGND_M1068_d N_VGND_M1073_s N_VGND_M1115_d
+ N_VGND_M1144_s N_VGND_M1281_d N_VGND_M1278_s N_VGND_c_12689_n N_VGND_c_12690_n
+ N_VGND_c_12691_n N_VGND_c_12692_n N_VGND_c_12693_n N_VGND_c_12694_n
+ N_VGND_c_12695_n N_VGND_c_12696_n N_VGND_c_12697_n N_VGND_c_12698_n
+ N_VGND_c_12699_n N_VGND_c_12700_n N_VGND_c_12701_n N_VGND_c_12702_n
+ N_VGND_c_12703_n N_VGND_c_12704_n N_VGND_c_12705_n N_VGND_c_12706_n
+ N_VGND_c_12707_n N_VGND_c_12708_n N_VGND_c_12709_n N_VGND_c_12710_n
+ N_VGND_c_12711_n N_VGND_c_12712_n N_VGND_c_12713_n N_VGND_c_12714_n
+ N_VGND_c_12715_n N_VGND_c_12716_n N_VGND_c_12717_n N_VGND_c_12718_n
+ N_VGND_c_12719_n N_VGND_c_12720_n N_VGND_c_12721_n N_VGND_c_12722_n
+ N_VGND_c_12723_n N_VGND_c_12724_n N_VGND_c_12725_n N_VGND_c_12726_n
+ N_VGND_c_12727_n N_VGND_c_12728_n N_VGND_c_12729_n N_VGND_c_12730_n
+ N_VGND_c_12731_n N_VGND_c_12732_n N_VGND_c_12733_n N_VGND_c_12734_n
+ N_VGND_c_12735_n N_VGND_c_12737_n N_VGND_c_12738_n N_VGND_c_12740_n
+ N_VGND_c_12741_n N_VGND_c_12742_n N_VGND_c_12743_n N_VGND_c_12744_n
+ N_VGND_c_12745_n N_VGND_c_12746_n N_VGND_c_12747_n N_VGND_c_12748_n
+ N_VGND_c_12749_n N_VGND_c_12750_n N_VGND_c_12751_n N_VGND_c_12752_n
+ N_VGND_c_12753_n N_VGND_c_12754_n N_VGND_c_12755_n N_VGND_c_12756_n
+ N_VGND_c_12757_n N_VGND_c_12758_n N_VGND_c_12759_n N_VGND_c_12760_n
+ N_VGND_c_12761_n N_VGND_c_12762_n N_VGND_c_12763_n N_VGND_c_12764_n
+ N_VGND_c_12765_n N_VGND_c_12766_n N_VGND_c_12767_n N_VGND_c_12768_n
+ N_VGND_c_12769_n N_VGND_c_12770_n N_VGND_c_12771_n N_VGND_c_12772_n
+ N_VGND_c_12773_n N_VGND_c_12774_n N_VGND_c_12775_n N_VGND_c_12776_n
+ N_VGND_c_12777_n N_VGND_c_12778_n N_VGND_c_12779_n N_VGND_c_12780_n
+ N_VGND_c_12781_n N_VGND_c_12782_n N_VGND_c_12783_n N_VGND_c_12784_n
+ N_VGND_c_12785_n N_VGND_c_12786_n N_VGND_c_12787_n N_VGND_c_12788_n
+ N_VGND_c_12789_n N_VGND_c_12790_n N_VGND_c_12791_n N_VGND_c_12792_n
+ N_VGND_c_12793_n N_VGND_c_12794_n N_VGND_c_12795_n N_VGND_c_12796_n
+ N_VGND_c_12797_n N_VGND_c_12798_n N_VGND_c_12799_n N_VGND_c_12800_n
+ N_VGND_c_12801_n N_VGND_c_12802_n N_VGND_c_12803_n N_VGND_c_12804_n
+ N_VGND_c_12805_n N_VGND_c_12806_n N_VGND_c_12807_n N_VGND_c_12808_n
+ N_VGND_c_12809_n N_VGND_c_12810_n N_VGND_c_12811_n N_VGND_c_12812_n
+ N_VGND_c_12813_n N_VGND_c_12814_n N_VGND_c_12815_n N_VGND_c_12816_n
+ N_VGND_c_12817_n N_VGND_c_12818_n N_VGND_c_12819_n N_VGND_c_12820_n
+ N_VGND_c_12821_n N_VGND_c_12822_n N_VGND_c_12823_n N_VGND_c_12824_n
+ N_VGND_c_12825_n N_VGND_c_12826_n N_VGND_c_12827_n N_VGND_c_12828_n
+ N_VGND_c_12829_n N_VGND_c_12830_n N_VGND_c_12831_n N_VGND_c_12832_n
+ N_VGND_c_12833_n N_VGND_c_12834_n N_VGND_c_12835_n N_VGND_c_12836_n
+ N_VGND_c_12837_n N_VGND_c_12838_n N_VGND_c_12839_n N_VGND_c_12840_n
+ N_VGND_c_12841_n N_VGND_c_12842_n N_VGND_c_12843_n N_VGND_c_12844_n
+ N_VGND_c_12845_n N_VGND_c_12846_n N_VGND_c_12847_n N_VGND_c_12848_n
+ N_VGND_c_12849_n N_VGND_c_12850_n N_VGND_c_12851_n N_VGND_c_12852_n
+ N_VGND_c_12853_n N_VGND_c_12854_n N_VGND_c_12855_n N_VGND_c_12856_n
+ N_VGND_c_12857_n N_VGND_c_12858_n N_VGND_c_12859_n N_VGND_c_12860_n
+ N_VGND_c_12861_n N_VGND_c_12862_n N_VGND_c_12863_n N_VGND_c_12864_n
+ N_VGND_c_12865_n N_VGND_c_12866_n VGND VGND VGND VGND VGND VGND VGND VGND VGND
+ VGND VGND VGND VGND VGND VGND VGND VGND VGND N_VGND_c_12870_n N_VGND_c_12871_n
+ N_VGND_c_12872_n N_VGND_c_12873_n N_VGND_c_12874_n N_VGND_c_12875_n
+ N_VGND_c_12876_n N_VGND_c_12877_n N_VGND_c_12878_n N_VGND_c_12879_n
+ N_VGND_c_12880_n N_VGND_c_12881_n N_VGND_c_12882_n N_VGND_c_12884_n
+ N_VGND_c_12885_n N_VGND_c_12886_n N_VGND_c_12887_n N_VGND_c_12888_n
+ N_VGND_c_12889_n N_VGND_c_12890_n N_VGND_c_12891_n N_VGND_c_12892_n
+ N_VGND_c_12893_n N_VGND_c_12894_n N_VGND_c_12895_n N_VGND_c_12896_n
+ N_VGND_c_12897_n N_VGND_c_12898_n N_VGND_c_12899_n N_VGND_c_12900_n
+ N_VGND_c_12901_n N_VGND_c_12902_n N_VGND_c_12903_n N_VGND_c_12904_n
+ N_VGND_c_12905_n N_VGND_c_12906_n N_VGND_c_12907_n N_VGND_c_12908_n
+ N_VGND_c_12909_n N_VGND_c_12910_n N_VGND_c_12911_n N_VGND_c_12912_n
+ N_VGND_c_12913_n N_VGND_c_12914_n N_VGND_c_12915_n N_VGND_c_12916_n
+ N_VGND_c_12917_n N_VGND_c_12918_n N_VGND_c_12919_n N_VGND_c_12920_n
+ N_VGND_c_12921_n N_VGND_c_12922_n N_VGND_c_12923_n N_VGND_c_12924_n
+ N_VGND_c_12925_n N_VGND_c_12926_n N_VGND_c_12927_n N_VGND_c_12928_n
+ N_VGND_c_12929_n N_VGND_c_12930_n N_VGND_c_12931_n N_VGND_c_12932_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%VGND
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_47# N_A_119_47#_M1084_s
+ N_A_119_47#_M1300_s N_A_119_47#_M1053_d N_A_119_47#_M1074_d
+ N_A_119_47#_M1125_d N_A_119_47#_c_14057_n N_A_119_47#_c_14060_n
+ N_A_119_47#_c_14049_n N_A_119_47#_c_14068_n N_A_119_47#_c_14050_n
+ N_A_119_47#_c_14051_n N_A_119_47#_c_14052_n N_A_119_47#_c_14053_n
+ N_A_119_47#_c_14077_n N_A_119_47#_c_14054_n N_A_119_47#_c_14055_n
+ N_A_119_47#_c_14056_n N_A_119_47#_c_14090_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_911# N_A_119_911#_M1085_s
+ N_A_119_911#_M1235_s N_A_119_911#_M1070_s N_A_119_911#_M1159_s
+ N_A_119_911#_M1302_s N_A_119_911#_c_14140_n N_A_119_911#_c_14132_n
+ N_A_119_911#_c_14133_n N_A_119_911#_c_14134_n N_A_119_911#_c_14135_n
+ N_A_119_911#_c_14156_n N_A_119_911#_c_14136_n N_A_119_911#_c_14137_n
+ N_A_119_911#_c_14138_n N_A_119_911#_c_14139_n N_A_119_911#_c_14169_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_119_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_66# N_A_1693_66#_M1039_s
+ N_A_1693_66#_M1045_s N_A_1693_66#_M1113_s N_A_1693_66#_M1049_s
+ N_A_1693_66#_M1167_s N_A_1693_66#_c_14211_n N_A_1693_66#_c_14212_n
+ N_A_1693_66#_c_14213_n N_A_1693_66#_c_14233_n N_A_1693_66#_c_14214_n
+ N_A_1693_66#_c_14215_n N_A_1693_66#_c_14216_n N_A_1693_66#_c_14217_n
+ N_A_1693_66#_c_14236_n N_A_1693_66#_c_14218_n N_A_1693_66#_c_14245_n
+ N_A_1693_66#_c_14230_n N_A_1693_66#_c_14219_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_66#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_918# N_A_1693_918#_M1027_s
+ N_A_1693_918#_M1032_s N_A_1693_918#_M1259_s N_A_1693_918#_M1019_s
+ N_A_1693_918#_M1178_s N_A_1693_918#_c_14295_n N_A_1693_918#_c_14296_n
+ N_A_1693_918#_c_14297_n N_A_1693_918#_c_14317_n N_A_1693_918#_c_14298_n
+ N_A_1693_918#_c_14299_n N_A_1693_918#_c_14300_n N_A_1693_918#_c_14301_n
+ N_A_1693_918#_c_14320_n N_A_1693_918#_c_14314_n N_A_1693_918#_c_14302_n
+ N_A_1693_918#_c_14303_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_1693_918#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_47# N_A_2695_47#_M1001_d
+ N_A_2695_47#_M1110_d N_A_2695_47#_M1035_s N_A_2695_47#_M1036_s
+ N_A_2695_47#_M1306_s N_A_2695_47#_c_14385_n N_A_2695_47#_c_14388_n
+ N_A_2695_47#_c_14377_n N_A_2695_47#_c_14396_n N_A_2695_47#_c_14378_n
+ N_A_2695_47#_c_14379_n N_A_2695_47#_c_14380_n N_A_2695_47#_c_14381_n
+ N_A_2695_47#_c_14405_n N_A_2695_47#_c_14382_n N_A_2695_47#_c_14383_n
+ N_A_2695_47#_c_14384_n N_A_2695_47#_c_14418_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_911# N_A_2695_911#_M1033_s
+ N_A_2695_911#_M1195_s N_A_2695_911#_M1010_d N_A_2695_911#_M1214_d
+ N_A_2695_911#_M1268_d N_A_2695_911#_c_14468_n N_A_2695_911#_c_14460_n
+ N_A_2695_911#_c_14461_n N_A_2695_911#_c_14462_n N_A_2695_911#_c_14463_n
+ N_A_2695_911#_c_14484_n N_A_2695_911#_c_14464_n N_A_2695_911#_c_14465_n
+ N_A_2695_911#_c_14466_n N_A_2695_911#_c_14467_n N_A_2695_911#_c_14497_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_2695_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_66# N_A_4269_66#_M1030_d
+ N_A_4269_66#_M1031_d N_A_4269_66#_M1106_d N_A_4269_66#_M1041_s
+ N_A_4269_66#_M1135_s N_A_4269_66#_c_14539_n N_A_4269_66#_c_14540_n
+ N_A_4269_66#_c_14541_n N_A_4269_66#_c_14561_n N_A_4269_66#_c_14542_n
+ N_A_4269_66#_c_14543_n N_A_4269_66#_c_14544_n N_A_4269_66#_c_14545_n
+ N_A_4269_66#_c_14564_n N_A_4269_66#_c_14546_n N_A_4269_66#_c_14573_n
+ N_A_4269_66#_c_14558_n N_A_4269_66#_c_14547_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_66#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_918# N_A_4269_918#_M1047_d
+ N_A_4269_918#_M1160_d N_A_4269_918#_M1318_d N_A_4269_918#_M1245_d
+ N_A_4269_918#_M1310_d N_A_4269_918#_c_14623_n N_A_4269_918#_c_14624_n
+ N_A_4269_918#_c_14625_n N_A_4269_918#_c_14645_n N_A_4269_918#_c_14626_n
+ N_A_4269_918#_c_14627_n N_A_4269_918#_c_14628_n N_A_4269_918#_c_14629_n
+ N_A_4269_918#_c_14648_n N_A_4269_918#_c_14642_n N_A_4269_918#_c_14630_n
+ N_A_4269_918#_c_14631_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_4269_918#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_47# N_A_5363_47#_M1021_s
+ N_A_5363_47#_M1232_s N_A_5363_47#_M1154_s N_A_5363_47#_M1191_s
+ N_A_5363_47#_M1213_s N_A_5363_47#_c_14713_n N_A_5363_47#_c_14716_n
+ N_A_5363_47#_c_14705_n N_A_5363_47#_c_14724_n N_A_5363_47#_c_14706_n
+ N_A_5363_47#_c_14707_n N_A_5363_47#_c_14708_n N_A_5363_47#_c_14709_n
+ N_A_5363_47#_c_14733_n N_A_5363_47#_c_14710_n N_A_5363_47#_c_14711_n
+ N_A_5363_47#_c_14712_n N_A_5363_47#_c_14746_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_911# N_A_5363_911#_M1012_s
+ N_A_5363_911#_M1187_s N_A_5363_911#_M1044_d N_A_5363_911#_M1091_d
+ N_A_5363_911#_M1312_d N_A_5363_911#_c_14796_n N_A_5363_911#_c_14788_n
+ N_A_5363_911#_c_14789_n N_A_5363_911#_c_14790_n N_A_5363_911#_c_14791_n
+ N_A_5363_911#_c_14812_n N_A_5363_911#_c_14792_n N_A_5363_911#_c_14793_n
+ N_A_5363_911#_c_14794_n N_A_5363_911#_c_14795_n N_A_5363_911#_c_14825_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_5363_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_66# N_A_6937_66#_M1175_d
+ N_A_6937_66#_M1210_d N_A_6937_66#_M1228_d N_A_6937_66#_M1029_s
+ N_A_6937_66#_M1247_s N_A_6937_66#_c_14867_n N_A_6937_66#_c_14868_n
+ N_A_6937_66#_c_14869_n N_A_6937_66#_c_14889_n N_A_6937_66#_c_14870_n
+ N_A_6937_66#_c_14871_n N_A_6937_66#_c_14872_n N_A_6937_66#_c_14873_n
+ N_A_6937_66#_c_14892_n N_A_6937_66#_c_14874_n N_A_6937_66#_c_14901_n
+ N_A_6937_66#_c_14886_n N_A_6937_66#_c_14875_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_66#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_918# N_A_6937_918#_M1149_d
+ N_A_6937_918#_M1226_d N_A_6937_918#_M1290_d N_A_6937_918#_M1132_s
+ N_A_6937_918#_M1274_s N_A_6937_918#_c_14951_n N_A_6937_918#_c_14952_n
+ N_A_6937_918#_c_14953_n N_A_6937_918#_c_14973_n N_A_6937_918#_c_14954_n
+ N_A_6937_918#_c_14955_n N_A_6937_918#_c_14956_n N_A_6937_918#_c_14957_n
+ N_A_6937_918#_c_14976_n N_A_6937_918#_c_14970_n N_A_6937_918#_c_14958_n
+ N_A_6937_918#_c_14959_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_6937_918#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_47# N_A_7939_47#_M1069_d
+ N_A_7939_47#_M1147_d N_A_7939_47#_M1202_d N_A_7939_47#_M1212_d
+ N_A_7939_47#_M1254_d N_A_7939_47#_c_15041_n N_A_7939_47#_c_15044_n
+ N_A_7939_47#_c_15033_n N_A_7939_47#_c_15052_n N_A_7939_47#_c_15034_n
+ N_A_7939_47#_c_15035_n N_A_7939_47#_c_15036_n N_A_7939_47#_c_15037_n
+ N_A_7939_47#_c_15061_n N_A_7939_47#_c_15038_n N_A_7939_47#_c_15039_n
+ N_A_7939_47#_c_15040_n N_A_7939_47#_c_15074_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_47#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_911# N_A_7939_911#_M1004_d
+ N_A_7939_911#_M1189_d N_A_7939_911#_M1005_d N_A_7939_911#_M1064_d
+ N_A_7939_911#_M1230_d N_A_7939_911#_c_15124_n N_A_7939_911#_c_15116_n
+ N_A_7939_911#_c_15117_n N_A_7939_911#_c_15118_n N_A_7939_911#_c_15119_n
+ N_A_7939_911#_c_15140_n N_A_7939_911#_c_15120_n N_A_7939_911#_c_15121_n
+ N_A_7939_911#_c_15122_n N_A_7939_911#_c_15123_n N_A_7939_911#_c_15153_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_7939_911#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_66# N_A_9513_66#_M1003_d
+ N_A_9513_66#_M1209_d N_A_9513_66#_M1272_d N_A_9513_66#_M1068_s
+ N_A_9513_66#_M1216_s N_A_9513_66#_c_15195_n N_A_9513_66#_c_15196_n
+ N_A_9513_66#_c_15197_n N_A_9513_66#_c_15217_n N_A_9513_66#_c_15198_n
+ N_A_9513_66#_c_15199_n N_A_9513_66#_c_15200_n N_A_9513_66#_c_15201_n
+ N_A_9513_66#_c_15220_n N_A_9513_66#_c_15202_n N_A_9513_66#_c_15229_n
+ N_A_9513_66#_c_15214_n N_A_9513_66#_c_15203_n
+ PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_66#
x_PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_918# N_A_9513_918#_M1104_s
+ N_A_9513_918#_M1169_s N_A_9513_918#_M1252_s N_A_9513_918#_M1073_d
+ N_A_9513_918#_M1190_d N_A_9513_918#_c_15279_n N_A_9513_918#_c_15280_n
+ N_A_9513_918#_c_15281_n N_A_9513_918#_c_15301_n N_A_9513_918#_c_15282_n
+ N_A_9513_918#_c_15283_n N_A_9513_918#_c_15284_n N_A_9513_918#_c_15285_n
+ N_A_9513_918#_c_15304_n N_A_9513_918#_c_15298_n N_A_9513_918#_c_15286_n
+ N_A_9513_918#_c_15287_n PM_SKY130_FD_SC_HDLL__MUXB16TO1_4%A_9513_918#
cc_1 VNB VPB 0.00992071f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.145
cc_2 VNB N_VPB_c_1128_n 0.00992071f $X=25.905 $Y=0.425 $X2=25.99 $Y2=1.73
cc_3 VNB N_D[0]_M1014_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_4 VNB N_D[0]_M1084_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_5 VNB N_D[0]_M1219_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_6 VNB N_D[0]_M1146_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_D[0]_M1208_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_D[0]_M1300_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_D[0]_M1317_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_D[0]_M1294_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D[0]_c_1877_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_D[0]_c_1878_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_13 VNB N_D[0]_c_1879_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_D[0]_c_1880_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_D[8]_M1023_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D[8]_M1085_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_17 VNB N_D[8]_M1090_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_18 VNB N_D[8]_M1155_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_D[8]_M1221_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_D[8]_M1235_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_D[8]_M1240_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_D[8]_M1304_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_D[8]_c_1967_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D[8]_c_1968_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_25 VNB N_D[8]_c_1969_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_D[8]_c_1970_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_559_265#_c_2045_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_559_265#_c_2046_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_559_265#_c_2047_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.57
cc_30 VNB N_A_559_265#_c_2048_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_559_265#_c_2049_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_559_265#_c_2050_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_559_265#_c_2051_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_559_793#_c_2163_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_559_793#_c_2164_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_559_793#_c_2165_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_559_793#_c_2166_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_559_793#_c_2167_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_559_793#_c_2168_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_559_793#_c_2169_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_S[0]_c_2287_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_42 VNB N_S[0]_c_2288_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_S[0]_c_2289_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_S[0]_c_2290_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_S[0]_c_2291_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_46 VNB N_S[0]_c_2292_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_47 VNB N_S[0]_c_2293_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_S[0]_c_2294_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_S[0]_c_2295_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_S[0]_c_2296_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_S[0]_c_2297_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_S[0]_c_2298_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_S[0]_c_2299_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_54 VNB N_S[0]_c_2300_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_55 VNB N_S[0]_c_2301_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_56 VNB N_S[0]_c_2302_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_S[0]_c_2303_n 0.065295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_S[0]_c_2304_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_S[0]_c_2305_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_S[0]_c_2306_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_S[0]_c_2307_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB S[0] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_S[8]_c_2404_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_64 VNB N_S[8]_c_2405_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_S[8]_c_2406_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_S[8]_c_2407_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_S[8]_c_2408_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_68 VNB N_S[8]_c_2409_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_69 VNB N_S[8]_c_2410_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_S[8]_c_2411_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_S[8]_c_2412_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_S[8]_c_2413_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_S[8]_c_2414_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_S[8]_c_2415_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_S[8]_c_2416_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_76 VNB N_S[8]_c_2417_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_77 VNB N_S[8]_c_2418_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_78 VNB N_S[8]_c_2419_n 0.0848512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_S[8]_c_2420_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_S[8]_c_2421_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_S[8]_c_2422_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_S[8]_c_2423_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB S[8] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_S[1]_c_2529_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_85 VNB N_S[1]_c_2530_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_S[1]_c_2531_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_S[1]_c_2532_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_88 VNB N_S[1]_c_2533_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_89 VNB N_S[1]_c_2534_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_S[1]_c_2535_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_S[1]_c_2536_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_S[1]_c_2537_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_S[1]_c_2538_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_S[1]_c_2539_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_95 VNB N_S[1]_c_2540_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_96 VNB N_S[1]_c_2541_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_97 VNB N_S[1]_c_2542_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_98 VNB N_S[1]_c_2543_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_S[1]_c_2544_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_S[1]_c_2545_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_S[1]_c_2546_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_S[1]_c_2547_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_S[1]_c_2548_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_S[1]_c_2549_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_S[1]_c_2550_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_S[9]_c_2649_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_107 VNB N_S[9]_c_2650_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_S[9]_c_2651_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_109 VNB N_S[9]_c_2652_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_S[9]_c_2653_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_S[9]_c_2654_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_S[9]_c_2655_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_S[9]_c_2656_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_S[9]_c_2657_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_S[9]_c_2658_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_116 VNB N_S[9]_c_2659_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_117 VNB N_S[9]_c_2660_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_118 VNB N_S[9]_c_2661_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_119 VNB N_S[9]_c_2662_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_S[9]_c_2663_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_S[9]_c_2664_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_S[9]_c_2665_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_S[9]_c_2666_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_S[9]_c_2667_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_S[9]_c_2668_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_S[9]_c_2669_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_A_1430_325#_c_2777_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_128 VNB N_A_1430_325#_c_2778_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_129 VNB N_A_1430_325#_c_2779_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.29
cc_130 VNB N_A_1430_325#_c_2780_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_A_1430_325#_c_2781_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_A_1430_325#_c_2782_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_A_1430_325#_c_2783_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_A_1430_599#_c_2893_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_135 VNB N_A_1430_599#_c_2894_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_A_1430_599#_c_2895_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_137 VNB N_A_1430_599#_c_2896_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_A_1430_599#_c_2897_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_A_1430_599#_c_2898_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_A_1430_599#_c_2899_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_D[1]_M1002_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_D[1]_M1049_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_143 VNB N_D[1]_M1098_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_144 VNB N_D[1]_M1038_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_D[1]_M1134_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_D[1]_M1167_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_D[1]_M1315_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_D[1]_M1271_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_D[1]_c_3023_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_D[1]_c_3024_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_151 VNB N_D[1]_c_3025_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_D[1]_c_3026_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB N_D[9]_M1011_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_D[9]_M1019_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_155 VNB N_D[9]_M1111_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_156 VNB N_D[9]_M1051_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_157 VNB N_D[9]_M1148_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_158 VNB N_D[9]_M1178_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_159 VNB N_D[9]_M1276_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_160 VNB N_D[9]_M1285_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_161 VNB N_D[9]_c_3116_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_162 VNB N_D[9]_c_3117_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_163 VNB N_D[9]_c_3118_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_164 VNB N_D[9]_c_3119_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_165 VNB N_D[2]_M1020_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_166 VNB N_D[2]_M1001_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_167 VNB N_D[2]_M1062_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_168 VNB N_D[2]_M1067_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_169 VNB N_D[2]_M1157_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_170 VNB N_D[2]_M1110_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_171 VNB N_D[2]_M1182_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_172 VNB N_D[2]_M1301_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_173 VNB N_D[2]_c_3207_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_174 VNB N_D[2]_c_3208_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_175 VNB N_D[2]_c_3209_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_176 VNB N_D[2]_c_3210_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_177 VNB N_D[10]_M1024_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_178 VNB N_D[10]_M1033_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_179 VNB N_D[10]_M1143_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_180 VNB N_D[10]_M1076_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_181 VNB N_D[10]_M1164_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_182 VNB N_D[10]_M1195_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_183 VNB N_D[10]_M1307_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_184 VNB N_D[10]_M1309_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_185 VNB N_D[10]_c_3302_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_186 VNB N_D[10]_c_3303_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_187 VNB N_D[10]_c_3304_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_188 VNB N_D[10]_c_3305_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_189 VNB N_A_3135_265#_c_3385_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_190 VNB N_A_3135_265#_c_3386_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_191 VNB N_A_3135_265#_c_3387_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.57
cc_192 VNB N_A_3135_265#_c_3388_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_193 VNB N_A_3135_265#_c_3389_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_194 VNB N_A_3135_265#_c_3390_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_195 VNB N_A_3135_265#_c_3391_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_196 VNB N_A_3135_793#_c_3504_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_197 VNB N_A_3135_793#_c_3505_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_198 VNB N_A_3135_793#_c_3506_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_199 VNB N_A_3135_793#_c_3507_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_200 VNB N_A_3135_793#_c_3508_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_201 VNB N_A_3135_793#_c_3509_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_202 VNB N_A_3135_793#_c_3510_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_203 VNB N_S[2]_c_3629_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_204 VNB N_S[2]_c_3630_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_205 VNB N_S[2]_c_3631_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_206 VNB N_S[2]_c_3632_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_207 VNB N_S[2]_c_3633_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_208 VNB N_S[2]_c_3634_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_209 VNB N_S[2]_c_3635_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_210 VNB N_S[2]_c_3636_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_211 VNB N_S[2]_c_3637_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_212 VNB N_S[2]_c_3638_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_213 VNB N_S[2]_c_3639_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_214 VNB N_S[2]_c_3640_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_215 VNB N_S[2]_c_3641_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_216 VNB N_S[2]_c_3642_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_217 VNB N_S[2]_c_3643_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_218 VNB N_S[2]_c_3644_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_219 VNB N_S[2]_c_3645_n 0.065295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_220 VNB N_S[2]_c_3646_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_221 VNB N_S[2]_c_3647_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_222 VNB N_S[2]_c_3648_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_223 VNB N_S[2]_c_3649_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_224 VNB S[2] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_225 VNB N_S[10]_c_3746_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_226 VNB N_S[10]_c_3747_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_227 VNB N_S[10]_c_3748_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_228 VNB N_S[10]_c_3749_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_229 VNB N_S[10]_c_3750_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_230 VNB N_S[10]_c_3751_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_231 VNB N_S[10]_c_3752_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_232 VNB N_S[10]_c_3753_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_233 VNB N_S[10]_c_3754_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_234 VNB N_S[10]_c_3755_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_235 VNB N_S[10]_c_3756_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_236 VNB N_S[10]_c_3757_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_237 VNB N_S[10]_c_3758_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_238 VNB N_S[10]_c_3759_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_239 VNB N_S[10]_c_3760_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_240 VNB N_S[10]_c_3761_n 0.0848512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_241 VNB N_S[10]_c_3762_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_242 VNB N_S[10]_c_3763_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_243 VNB N_S[10]_c_3764_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_244 VNB N_S[10]_c_3765_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_245 VNB S[10] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_246 VNB N_S[3]_c_3871_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_247 VNB N_S[3]_c_3872_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_248 VNB N_S[3]_c_3873_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_249 VNB N_S[3]_c_3874_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_250 VNB N_S[3]_c_3875_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_251 VNB N_S[3]_c_3876_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_252 VNB N_S[3]_c_3877_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_253 VNB N_S[3]_c_3878_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_254 VNB N_S[3]_c_3879_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_255 VNB N_S[3]_c_3880_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_256 VNB N_S[3]_c_3881_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_257 VNB N_S[3]_c_3882_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_258 VNB N_S[3]_c_3883_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_259 VNB N_S[3]_c_3884_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_260 VNB N_S[3]_c_3885_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_261 VNB N_S[3]_c_3886_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_262 VNB N_S[3]_c_3887_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_263 VNB N_S[3]_c_3888_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_264 VNB N_S[3]_c_3889_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_265 VNB N_S[3]_c_3890_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_266 VNB N_S[3]_c_3891_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_267 VNB N_S[3]_c_3892_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_268 VNB N_S[11]_c_3991_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_269 VNB N_S[11]_c_3992_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_270 VNB N_S[11]_c_3993_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_271 VNB N_S[11]_c_3994_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_272 VNB N_S[11]_c_3995_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_273 VNB N_S[11]_c_3996_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_274 VNB N_S[11]_c_3997_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_275 VNB N_S[11]_c_3998_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_276 VNB N_S[11]_c_3999_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_277 VNB N_S[11]_c_4000_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_278 VNB N_S[11]_c_4001_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_279 VNB N_S[11]_c_4002_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_280 VNB N_S[11]_c_4003_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_281 VNB N_S[11]_c_4004_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_282 VNB N_S[11]_c_4005_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_283 VNB N_S[11]_c_4006_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_284 VNB N_S[11]_c_4007_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_285 VNB N_S[11]_c_4008_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_286 VNB N_S[11]_c_4009_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_287 VNB N_S[11]_c_4010_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_288 VNB N_S[11]_c_4011_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_289 VNB N_A_4006_325#_c_4119_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_290 VNB N_A_4006_325#_c_4120_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_291 VNB N_A_4006_325#_c_4121_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.29
cc_292 VNB N_A_4006_325#_c_4122_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_293 VNB N_A_4006_325#_c_4123_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_294 VNB N_A_4006_325#_c_4124_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_295 VNB N_A_4006_325#_c_4125_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_296 VNB N_A_4006_599#_c_4235_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_297 VNB N_A_4006_599#_c_4236_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_298 VNB N_A_4006_599#_c_4237_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_299 VNB N_A_4006_599#_c_4238_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_300 VNB N_A_4006_599#_c_4239_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_301 VNB N_A_4006_599#_c_4240_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_302 VNB N_A_4006_599#_c_4241_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_303 VNB N_D[3]_M1042_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_304 VNB N_D[3]_M1041_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_305 VNB N_D[3]_M1100_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_306 VNB N_D[3]_M1089_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_307 VNB N_D[3]_M1116_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_308 VNB N_D[3]_M1135_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_309 VNB N_D[3]_M1193_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_310 VNB N_D[3]_M1289_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_311 VNB N_D[3]_c_4365_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_312 VNB N_D[3]_c_4366_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_313 VNB N_D[3]_c_4367_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_314 VNB N_D[3]_c_4368_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_315 VNB N_D[11]_M1052_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_316 VNB N_D[11]_M1245_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_317 VNB N_D[11]_M1296_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_318 VNB N_D[11]_M1101_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_319 VNB N_D[11]_M1129_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_320 VNB N_D[11]_M1310_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_321 VNB N_D[11]_M1311_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_322 VNB N_D[11]_M1297_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_323 VNB N_D[11]_c_4459_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_324 VNB N_D[11]_c_4460_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_325 VNB N_D[11]_c_4461_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_326 VNB N_D[11]_c_4462_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_327 VNB N_D[4]_M1158_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_328 VNB N_D[4]_M1021_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_329 VNB N_D[4]_M1177_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_330 VNB N_D[4]_M1194_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_331 VNB N_D[4]_M1265_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_332 VNB N_D[4]_M1232_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_333 VNB N_D[4]_M1275_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_334 VNB N_D[4]_M1319_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_335 VNB N_D[4]_c_4551_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_336 VNB N_D[4]_c_4552_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_337 VNB N_D[4]_c_4553_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_338 VNB N_D[4]_c_4554_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_339 VNB N_D[12]_M1006_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_340 VNB N_D[12]_M1012_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_341 VNB N_D[12]_M1128_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_342 VNB N_D[12]_M1165_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_343 VNB N_D[12]_M1203_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_344 VNB N_D[12]_M1187_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_345 VNB N_D[12]_M1267_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_346 VNB N_D[12]_M1277_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_347 VNB N_D[12]_c_4647_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_348 VNB N_D[12]_c_4648_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_349 VNB N_D[12]_c_4649_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_350 VNB N_D[12]_c_4650_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_351 VNB N_A_5803_265#_c_4731_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_352 VNB N_A_5803_265#_c_4732_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_353 VNB N_A_5803_265#_c_4733_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.57
cc_354 VNB N_A_5803_265#_c_4734_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_355 VNB N_A_5803_265#_c_4735_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_356 VNB N_A_5803_265#_c_4736_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_357 VNB N_A_5803_265#_c_4737_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_358 VNB N_A_5803_793#_c_4850_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_359 VNB N_A_5803_793#_c_4851_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_360 VNB N_A_5803_793#_c_4852_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_361 VNB N_A_5803_793#_c_4853_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_362 VNB N_A_5803_793#_c_4854_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_363 VNB N_A_5803_793#_c_4855_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_364 VNB N_A_5803_793#_c_4856_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_365 VNB N_S[4]_c_4975_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_366 VNB N_S[4]_c_4976_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_367 VNB N_S[4]_c_4977_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_368 VNB N_S[4]_c_4978_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_369 VNB N_S[4]_c_4979_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_370 VNB N_S[4]_c_4980_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_371 VNB N_S[4]_c_4981_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_372 VNB N_S[4]_c_4982_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_373 VNB N_S[4]_c_4983_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_374 VNB N_S[4]_c_4984_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_375 VNB N_S[4]_c_4985_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_376 VNB N_S[4]_c_4986_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_377 VNB N_S[4]_c_4987_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_378 VNB N_S[4]_c_4988_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_379 VNB N_S[4]_c_4989_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_380 VNB N_S[4]_c_4990_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_381 VNB N_S[4]_c_4991_n 0.065295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_382 VNB N_S[4]_c_4992_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_383 VNB N_S[4]_c_4993_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_384 VNB N_S[4]_c_4994_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_385 VNB N_S[4]_c_4995_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_386 VNB S[4] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_387 VNB N_S[12]_c_5092_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_388 VNB N_S[12]_c_5093_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_389 VNB N_S[12]_c_5094_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_390 VNB N_S[12]_c_5095_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_391 VNB N_S[12]_c_5096_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_392 VNB N_S[12]_c_5097_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_393 VNB N_S[12]_c_5098_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_394 VNB N_S[12]_c_5099_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_395 VNB N_S[12]_c_5100_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_396 VNB N_S[12]_c_5101_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_397 VNB N_S[12]_c_5102_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_398 VNB N_S[12]_c_5103_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_399 VNB N_S[12]_c_5104_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_400 VNB N_S[12]_c_5105_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_401 VNB N_S[12]_c_5106_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_402 VNB N_S[12]_c_5107_n 0.0848512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_403 VNB N_S[12]_c_5108_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_404 VNB N_S[12]_c_5109_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_405 VNB N_S[12]_c_5110_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_406 VNB N_S[12]_c_5111_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_407 VNB S[12] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_408 VNB N_S[5]_c_5217_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_409 VNB N_S[5]_c_5218_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_410 VNB N_S[5]_c_5219_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_411 VNB N_S[5]_c_5220_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_412 VNB N_S[5]_c_5221_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_413 VNB N_S[5]_c_5222_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_414 VNB N_S[5]_c_5223_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_415 VNB N_S[5]_c_5224_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_416 VNB N_S[5]_c_5225_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_417 VNB N_S[5]_c_5226_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_418 VNB N_S[5]_c_5227_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_419 VNB N_S[5]_c_5228_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_420 VNB N_S[5]_c_5229_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_421 VNB N_S[5]_c_5230_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_422 VNB N_S[5]_c_5231_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_423 VNB N_S[5]_c_5232_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_424 VNB N_S[5]_c_5233_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_425 VNB N_S[5]_c_5234_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_426 VNB N_S[5]_c_5235_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_427 VNB N_S[5]_c_5236_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_428 VNB N_S[5]_c_5237_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_429 VNB N_S[5]_c_5238_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_430 VNB N_S[13]_c_5337_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_431 VNB N_S[13]_c_5338_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_432 VNB N_S[13]_c_5339_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_433 VNB N_S[13]_c_5340_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_434 VNB N_S[13]_c_5341_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_435 VNB N_S[13]_c_5342_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_436 VNB N_S[13]_c_5343_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_437 VNB N_S[13]_c_5344_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_438 VNB N_S[13]_c_5345_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_439 VNB N_S[13]_c_5346_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_440 VNB N_S[13]_c_5347_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_441 VNB N_S[13]_c_5348_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_442 VNB N_S[13]_c_5349_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_443 VNB N_S[13]_c_5350_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_444 VNB N_S[13]_c_5351_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_445 VNB N_S[13]_c_5352_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_446 VNB N_S[13]_c_5353_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_447 VNB N_S[13]_c_5354_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_448 VNB N_S[13]_c_5355_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_449 VNB N_S[13]_c_5356_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_450 VNB N_S[13]_c_5357_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_451 VNB N_A_6674_325#_c_5465_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_452 VNB N_A_6674_325#_c_5466_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_453 VNB N_A_6674_325#_c_5467_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.29
cc_454 VNB N_A_6674_325#_c_5468_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_455 VNB N_A_6674_325#_c_5469_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_456 VNB N_A_6674_325#_c_5470_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_457 VNB N_A_6674_325#_c_5471_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_458 VNB N_A_6674_599#_c_5581_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_459 VNB N_A_6674_599#_c_5582_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_460 VNB N_A_6674_599#_c_5583_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_461 VNB N_A_6674_599#_c_5584_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_462 VNB N_A_6674_599#_c_5585_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_463 VNB N_A_6674_599#_c_5586_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_464 VNB N_A_6674_599#_c_5587_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_465 VNB N_D[5]_M1088_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_466 VNB N_D[5]_M1029_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_467 VNB N_D[5]_M1057_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_468 VNB N_D[5]_M1183_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_469 VNB N_D[5]_M1217_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_470 VNB N_D[5]_M1247_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_471 VNB N_D[5]_M1262_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_472 VNB N_D[5]_M1255_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_473 VNB N_D[5]_c_5711_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_474 VNB N_D[5]_c_5712_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_475 VNB N_D[5]_c_5713_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_476 VNB N_D[5]_c_5714_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_477 VNB N_D[13]_M1102_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_478 VNB N_D[13]_M1132_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_479 VNB N_D[13]_M1136_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_480 VNB N_D[13]_M1186_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_481 VNB N_D[13]_M1224_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_482 VNB N_D[13]_M1274_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_483 VNB N_D[13]_M1298_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_484 VNB N_D[13]_M1264_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_485 VNB N_D[13]_c_5804_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_486 VNB N_D[13]_c_5805_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_487 VNB N_D[13]_c_5806_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_488 VNB N_D[13]_c_5807_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_489 VNB N_D[6]_M1099_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_490 VNB N_D[6]_M1069_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_491 VNB N_D[6]_M1122_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_492 VNB N_D[6]_M1176_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_493 VNB N_D[6]_M1246_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_494 VNB N_D[6]_M1147_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_495 VNB N_D[6]_M1258_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_496 VNB N_D[6]_M1282_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_497 VNB N_D[6]_c_5895_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_498 VNB N_D[6]_c_5896_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_499 VNB N_D[6]_c_5897_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_500 VNB N_D[6]_c_5898_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_501 VNB N_D[14]_M1109_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_502 VNB N_D[14]_M1004_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_503 VNB N_D[14]_M1179_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_504 VNB N_D[14]_M1184_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_505 VNB N_D[14]_M1251_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_506 VNB N_D[14]_M1189_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_507 VNB N_D[14]_M1305_g 0.024303f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_508 VNB N_D[14]_M1293_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_509 VNB N_D[14]_c_5990_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_510 VNB N_D[14]_c_5991_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_511 VNB N_D[14]_c_5992_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_512 VNB N_D[14]_c_5993_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_513 VNB N_A_8379_265#_c_6073_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_514 VNB N_A_8379_265#_c_6074_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_515 VNB N_A_8379_265#_c_6075_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.57
cc_516 VNB N_A_8379_265#_c_6076_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_517 VNB N_A_8379_265#_c_6077_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_518 VNB N_A_8379_265#_c_6078_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_519 VNB N_A_8379_265#_c_6079_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_520 VNB N_A_8379_793#_c_6192_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_521 VNB N_A_8379_793#_c_6193_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_522 VNB N_A_8379_793#_c_6194_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_523 VNB N_A_8379_793#_c_6195_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_524 VNB N_A_8379_793#_c_6196_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_525 VNB N_A_8379_793#_c_6197_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_526 VNB N_A_8379_793#_c_6198_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_527 VNB N_S[6]_c_6317_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_528 VNB N_S[6]_c_6318_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_529 VNB N_S[6]_c_6319_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_530 VNB N_S[6]_c_6320_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_531 VNB N_S[6]_c_6321_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_532 VNB N_S[6]_c_6322_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_533 VNB N_S[6]_c_6323_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_534 VNB N_S[6]_c_6324_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_535 VNB N_S[6]_c_6325_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_536 VNB N_S[6]_c_6326_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_537 VNB N_S[6]_c_6327_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_538 VNB N_S[6]_c_6328_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_539 VNB N_S[6]_c_6329_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_540 VNB N_S[6]_c_6330_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_541 VNB N_S[6]_c_6331_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_542 VNB N_S[6]_c_6332_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_543 VNB N_S[6]_c_6333_n 0.065295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_544 VNB N_S[6]_c_6334_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_545 VNB N_S[6]_c_6335_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_546 VNB N_S[6]_c_6336_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_547 VNB N_S[6]_c_6337_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_548 VNB S[6] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_549 VNB N_S[14]_c_6434_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_550 VNB N_S[14]_c_6435_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_551 VNB N_S[14]_c_6436_n 0.0125768f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_552 VNB N_S[14]_c_6437_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_553 VNB N_S[14]_c_6438_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_554 VNB N_S[14]_c_6439_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_555 VNB N_S[14]_c_6440_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_556 VNB N_S[14]_c_6441_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_557 VNB N_S[14]_c_6442_n 0.0567558f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_558 VNB N_S[14]_c_6443_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_559 VNB N_S[14]_c_6444_n 0.0166808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_560 VNB N_S[14]_c_6445_n 0.00917895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_561 VNB N_S[14]_c_6446_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_562 VNB N_S[14]_c_6447_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_563 VNB N_S[14]_c_6448_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_564 VNB N_S[14]_c_6449_n 0.0848512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_565 VNB N_S[14]_c_6450_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_566 VNB N_S[14]_c_6451_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_567 VNB N_S[14]_c_6452_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_568 VNB N_S[14]_c_6453_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_569 VNB S[14] 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_570 VNB N_S[7]_c_6559_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_571 VNB N_S[7]_c_6560_n 0.0330319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_572 VNB N_S[7]_c_6561_n 0.0195563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_573 VNB N_S[7]_c_6562_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_574 VNB N_S[7]_c_6563_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_575 VNB N_S[7]_c_6564_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_576 VNB N_S[7]_c_6565_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_577 VNB N_S[7]_c_6566_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_578 VNB N_S[7]_c_6567_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_579 VNB N_S[7]_c_6568_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_580 VNB N_S[7]_c_6569_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_581 VNB N_S[7]_c_6570_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_582 VNB N_S[7]_c_6571_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_583 VNB N_S[7]_c_6572_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_584 VNB N_S[7]_c_6573_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_585 VNB N_S[7]_c_6574_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_586 VNB N_S[7]_c_6575_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_587 VNB N_S[7]_c_6576_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_588 VNB N_S[7]_c_6577_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_589 VNB N_S[7]_c_6578_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_590 VNB N_S[7]_c_6579_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_591 VNB N_S[7]_c_6580_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_592 VNB N_S[15]_c_6679_n 0.032202f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=1.525
cc_593 VNB N_S[15]_c_6680_n 0.0525882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_594 VNB N_S[15]_c_6681_n 0.0101778f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=2.125
cc_595 VNB N_S[15]_c_6682_n 0.0259684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_596 VNB N_S[15]_c_6683_n 0.0150643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_597 VNB N_S[15]_c_6684_n 0.0258597f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_598 VNB N_S[15]_c_6685_n 0.0308948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_599 VNB N_S[15]_c_6686_n 0.046608f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_600 VNB N_S[15]_c_6687_n 0.0101478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_601 VNB N_S[15]_c_6688_n 0.0160363f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_602 VNB N_S[15]_c_6689_n 0.0152656f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.87
cc_603 VNB N_S[15]_c_6690_n 0.0120586f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=2.21
cc_604 VNB N_S[15]_c_6691_n 0.0159402f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.23
cc_605 VNB N_S[15]_c_6692_n 0.0120614f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_606 VNB N_S[15]_c_6693_n 0.0278425f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_607 VNB N_S[15]_c_6694_n 0.0174346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_608 VNB N_S[15]_c_6695_n 0.00318387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_609 VNB N_S[15]_c_6696_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_610 VNB N_S[15]_c_6697_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_611 VNB N_S[15]_c_6698_n 0.00749069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_612 VNB N_S[15]_c_6699_n 0.00265247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_613 VNB N_A_9250_325#_c_6807_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_614 VNB N_A_9250_325#_c_6808_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_615 VNB N_A_9250_325#_c_6809_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.29
cc_616 VNB N_A_9250_325#_c_6810_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_617 VNB N_A_9250_325#_c_6811_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_618 VNB N_A_9250_325#_c_6812_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_619 VNB N_A_9250_325#_c_6813_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_620 VNB N_A_9250_599#_c_6922_n 0.0183242f $X=-0.19 $Y=-0.24 $X2=25.905
+ $Y2=3.51
cc_621 VNB N_A_9250_599#_c_6923_n 3.3289e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_622 VNB N_A_9250_599#_c_6924_n 4.0898e-19 $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_623 VNB N_A_9250_599#_c_6925_n 0.0169775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_624 VNB N_A_9250_599#_c_6926_n 0.00144063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_625 VNB N_A_9250_599#_c_6927_n 0.00144707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_626 VNB N_A_9250_599#_c_6928_n 0.0181344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_627 VNB N_D[7]_M1040_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_628 VNB N_D[7]_M1068_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_629 VNB N_D[7]_M1115_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_630 VNB N_D[7]_M1087_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_631 VNB N_D[7]_M1131_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_632 VNB N_D[7]_M1216_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_633 VNB N_D[7]_M1281_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_634 VNB N_D[7]_M1151_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_635 VNB N_D[7]_c_7051_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_636 VNB N_D[7]_c_7052_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_637 VNB N_D[7]_c_7053_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_638 VNB N_D[7]_c_7054_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_639 VNB N_D[15]_M1056_g 7.61465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_640 VNB N_D[15]_M1073_g 0.024303f $X=-0.19 $Y=-0.24 $X2=-0.19 $Y2=1.305
cc_641 VNB N_D[15]_M1144_g 0.0193326f $X=-0.19 $Y=-0.24 $X2=25.905 $Y2=3.51
cc_642 VNB N_D[15]_M1103_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_643 VNB N_D[15]_M1145_g 4.18552e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_644 VNB N_D[15]_M1190_g 0.0184976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_645 VNB N_D[15]_M1278_g 0.0251977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_646 VNB N_D[15]_M1156_g 5.52889e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_647 VNB N_D[15]_c_7139_n 0.0160223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_648 VNB N_D[15]_c_7140_n 0.0405808f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=3.29
cc_649 VNB N_D[15]_c_7141_n 0.0102483f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_650 VNB N_D[15]_c_7142_n 0.0356842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_651 VNB N_Z_c_9003_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_652 VNB N_Z_c_9004_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_653 VNB N_Z_c_9005_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_654 VNB N_Z_c_9006_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_655 VNB N_Z_c_9007_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_656 VNB N_Z_c_9008_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_657 VNB N_Z_c_9009_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_658 VNB N_Z_c_9010_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_659 VNB N_Z_c_9011_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_660 VNB N_Z_c_9012_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_661 VNB N_Z_c_9013_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_662 VNB N_Z_c_9014_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_663 VNB N_Z_c_9015_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_664 VNB N_Z_c_9016_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_665 VNB N_Z_c_9017_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_666 VNB N_Z_c_9018_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_667 VNB N_Z_c_9019_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_668 VNB N_Z_c_9020_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_669 VNB N_Z_c_9021_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_670 VNB N_Z_c_9022_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_671 VNB N_Z_c_9023_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_672 VNB N_Z_c_9024_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_673 VNB N_Z_c_9025_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_674 VNB N_Z_c_9026_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_675 VNB N_Z_c_9027_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_676 VNB N_Z_c_9028_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_677 VNB N_Z_c_9029_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_678 VNB N_Z_c_9030_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_679 VNB N_Z_c_9031_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_680 VNB N_Z_c_9032_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_681 VNB N_Z_c_9033_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_682 VNB N_Z_c_9034_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_683 VNB N_Z_c_9035_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_684 VNB N_Z_c_9036_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_685 VNB N_Z_c_9037_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_686 VNB N_Z_c_9038_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_687 VNB N_Z_c_9039_n 0.00420252f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_688 VNB N_Z_c_9040_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_689 VNB N_Z_c_9041_n 0.00534541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_690 VNB N_Z_c_9042_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_691 VNB N_Z_c_9043_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_692 VNB N_Z_c_9044_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_693 VNB N_Z_c_9045_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_694 VNB N_Z_c_9046_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_695 VNB N_Z_c_9047_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_696 VNB N_Z_c_9048_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_697 VNB N_Z_c_9049_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_698 VNB N_Z_c_9050_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_699 VNB N_Z_c_9051_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_700 VNB N_Z_c_9052_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_701 VNB N_Z_c_9053_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_702 VNB N_Z_c_9054_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_703 VNB N_Z_c_9055_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_704 VNB N_Z_c_9056_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_705 VNB N_Z_c_9057_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_706 VNB N_Z_c_9058_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_707 VNB N_Z_c_9059_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_708 VNB N_Z_c_9060_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_709 VNB N_Z_c_9061_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_710 VNB N_Z_c_9062_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_711 VNB N_Z_c_9063_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_712 VNB N_Z_c_9064_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_713 VNB N_Z_c_9065_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_714 VNB N_Z_c_9066_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_715 VNB N_Z_c_9067_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_716 VNB N_Z_c_9068_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_717 VNB N_Z_c_9069_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_718 VNB N_Z_c_9070_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_719 VNB N_Z_c_9071_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_720 VNB N_Z_c_9072_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_721 VNB N_Z_c_9073_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_722 VNB N_Z_c_9074_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_723 VNB N_Z_c_9075_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_724 VNB N_Z_c_9076_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_725 VNB N_Z_c_9077_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_726 VNB N_Z_c_9078_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_727 VNB N_Z_c_9079_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_728 VNB N_Z_c_9080_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_729 VNB N_Z_c_9081_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_730 VNB N_Z_c_9082_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_731 VNB N_Z_c_9083_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_732 VNB N_Z_c_9084_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_733 VNB N_Z_c_9085_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_734 VNB N_Z_c_9086_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_735 VNB N_Z_c_9087_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_736 VNB N_Z_c_9088_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_737 VNB N_Z_c_9089_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_738 VNB N_Z_c_9090_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_739 VNB N_Z_c_9091_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_740 VNB N_Z_c_9092_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_741 VNB N_Z_c_9093_n 0.00392171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_742 VNB N_Z_c_9094_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_743 VNB N_Z_c_9095_n 0.0108049f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_744 VNB N_Z_c_9096_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_745 VNB N_Z_c_9097_n 9.07588e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_746 VNB N_Z_c_9098_n 0.0049568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_747 VNB N_VGND_c_12689_n 0.0116316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_748 VNB N_VGND_c_12690_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_749 VNB N_VGND_c_12691_n 0.0116057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_750 VNB N_VGND_c_12692_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_751 VNB N_VGND_c_12693_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_752 VNB N_VGND_c_12694_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_753 VNB N_VGND_c_12695_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_754 VNB N_VGND_c_12696_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_755 VNB N_VGND_c_12697_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_756 VNB N_VGND_c_12698_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_757 VNB N_VGND_c_12699_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_758 VNB N_VGND_c_12700_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_759 VNB N_VGND_c_12701_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_760 VNB N_VGND_c_12702_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_761 VNB N_VGND_c_12703_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_762 VNB N_VGND_c_12704_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_763 VNB N_VGND_c_12705_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_764 VNB N_VGND_c_12706_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_765 VNB N_VGND_c_12707_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_766 VNB N_VGND_c_12708_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_767 VNB N_VGND_c_12709_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_768 VNB N_VGND_c_12710_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_769 VNB N_VGND_c_12711_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_770 VNB N_VGND_c_12712_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_771 VNB N_VGND_c_12713_n 0.00916474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_772 VNB N_VGND_c_12714_n 0.00916474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_773 VNB N_VGND_c_12715_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_774 VNB N_VGND_c_12716_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_775 VNB N_VGND_c_12717_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_776 VNB N_VGND_c_12718_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_777 VNB N_VGND_c_12719_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_778 VNB N_VGND_c_12720_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_779 VNB N_VGND_c_12721_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_780 VNB N_VGND_c_12722_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_781 VNB N_VGND_c_12723_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_782 VNB N_VGND_c_12724_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_783 VNB N_VGND_c_12725_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_784 VNB N_VGND_c_12726_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_785 VNB N_VGND_c_12727_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_786 VNB N_VGND_c_12728_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_787 VNB N_VGND_c_12729_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_788 VNB N_VGND_c_12730_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_789 VNB N_VGND_c_12731_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_790 VNB N_VGND_c_12732_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_791 VNB N_VGND_c_12733_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_792 VNB N_VGND_c_12734_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_793 VNB N_VGND_c_12735_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_794 VNB N_VGND_c_12735_n 0.0347908f $X=25.905 $Y=0.425 $X2=0 $Y2=0
cc_795 VNB N_VGND_c_12737_n 0.0433975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_796 VNB N_VGND_c_12738_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_797 VNB N_VGND_c_12738_n 0.0347908f $X=25.905 $Y=0.425 $X2=0 $Y2=0
cc_798 VNB N_VGND_c_12740_n 0.0433975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_799 VNB N_VGND_c_12741_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_800 VNB N_VGND_c_12742_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_801 VNB N_VGND_c_12743_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_802 VNB N_VGND_c_12744_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_803 VNB N_VGND_c_12745_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_804 VNB N_VGND_c_12746_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_805 VNB N_VGND_c_12747_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_806 VNB N_VGND_c_12748_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_807 VNB N_VGND_c_12749_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_808 VNB N_VGND_c_12750_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_809 VNB N_VGND_c_12751_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_810 VNB N_VGND_c_12752_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_811 VNB N_VGND_c_12753_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_812 VNB N_VGND_c_12754_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_813 VNB N_VGND_c_12755_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_814 VNB N_VGND_c_12756_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_815 VNB N_VGND_c_12757_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_816 VNB N_VGND_c_12758_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_817 VNB N_VGND_c_12759_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_818 VNB N_VGND_c_12760_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_819 VNB N_VGND_c_12761_n 0.00916474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_820 VNB N_VGND_c_12762_n 0.00916474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_821 VNB N_VGND_c_12763_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_822 VNB N_VGND_c_12764_n 0.00746944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_823 VNB N_VGND_c_12765_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_824 VNB N_VGND_c_12766_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_825 VNB N_VGND_c_12767_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_826 VNB N_VGND_c_12768_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_827 VNB N_VGND_c_12769_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_828 VNB N_VGND_c_12770_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_829 VNB N_VGND_c_12771_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_830 VNB N_VGND_c_12772_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_831 VNB N_VGND_c_12773_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_832 VNB N_VGND_c_12774_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_833 VNB N_VGND_c_12775_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_834 VNB N_VGND_c_12776_n 0.00998524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_835 VNB N_VGND_c_12777_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_836 VNB N_VGND_c_12778_n 0.00992042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_837 VNB N_VGND_c_12779_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_838 VNB N_VGND_c_12780_n 0.0077543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_839 VNB N_VGND_c_12781_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_840 VNB N_VGND_c_12782_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_841 VNB N_VGND_c_12783_n 0.0116316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_842 VNB N_VGND_c_12784_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_843 VNB N_VGND_c_12785_n 0.0116057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_844 VNB N_VGND_c_12786_n 0.0086067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_845 VNB N_VGND_c_12787_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_846 VNB N_VGND_c_12788_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_847 VNB N_VGND_c_12789_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_848 VNB N_VGND_c_12790_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_849 VNB N_VGND_c_12791_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_850 VNB N_VGND_c_12792_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_851 VNB N_VGND_c_12793_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_852 VNB N_VGND_c_12794_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_853 VNB N_VGND_c_12795_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_854 VNB N_VGND_c_12796_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_855 VNB N_VGND_c_12797_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_856 VNB N_VGND_c_12798_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_857 VNB N_VGND_c_12799_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_858 VNB N_VGND_c_12800_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_859 VNB N_VGND_c_12801_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_860 VNB N_VGND_c_12802_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_861 VNB N_VGND_c_12803_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_862 VNB N_VGND_c_12804_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_863 VNB N_VGND_c_12805_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_864 VNB N_VGND_c_12806_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_865 VNB N_VGND_c_12807_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_866 VNB N_VGND_c_12808_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_867 VNB N_VGND_c_12809_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_868 VNB N_VGND_c_12810_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_869 VNB N_VGND_c_12811_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_870 VNB N_VGND_c_12812_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_871 VNB N_VGND_c_12813_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_872 VNB N_VGND_c_12814_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_873 VNB N_VGND_c_12815_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_874 VNB N_VGND_c_12816_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_875 VNB N_VGND_c_12817_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_876 VNB N_VGND_c_12818_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_877 VNB N_VGND_c_12819_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_878 VNB N_VGND_c_12820_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_879 VNB N_VGND_c_12821_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_880 VNB N_VGND_c_12822_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_881 VNB N_VGND_c_12823_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_882 VNB N_VGND_c_12824_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_883 VNB N_VGND_c_12825_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_884 VNB N_VGND_c_12826_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_885 VNB N_VGND_c_12827_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_886 VNB N_VGND_c_12828_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_887 VNB N_VGND_c_12829_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_888 VNB N_VGND_c_12830_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_889 VNB N_VGND_c_12831_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_890 VNB N_VGND_c_12832_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_891 VNB N_VGND_c_12833_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_892 VNB N_VGND_c_12834_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_893 VNB N_VGND_c_12835_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_894 VNB N_VGND_c_12836_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_895 VNB N_VGND_c_12837_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_896 VNB N_VGND_c_12838_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_897 VNB N_VGND_c_12839_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_898 VNB N_VGND_c_12840_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_899 VNB N_VGND_c_12841_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_900 VNB N_VGND_c_12842_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_901 VNB N_VGND_c_12843_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_902 VNB N_VGND_c_12844_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_903 VNB N_VGND_c_12845_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_904 VNB N_VGND_c_12846_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_905 VNB N_VGND_c_12847_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_906 VNB N_VGND_c_12848_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_907 VNB N_VGND_c_12849_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_908 VNB N_VGND_c_12850_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_909 VNB N_VGND_c_12851_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_910 VNB N_VGND_c_12852_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_911 VNB N_VGND_c_12853_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_912 VNB N_VGND_c_12854_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_913 VNB N_VGND_c_12855_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_914 VNB N_VGND_c_12856_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_915 VNB N_VGND_c_12857_n 0.0171202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_916 VNB N_VGND_c_12858_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_917 VNB N_VGND_c_12859_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_918 VNB N_VGND_c_12860_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_919 VNB N_VGND_c_12861_n 0.0177624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_920 VNB N_VGND_c_12862_n 0.00555283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_921 VNB N_VGND_c_12863_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_922 VNB N_VGND_c_12864_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_923 VNB N_VGND_c_12865_n 0.065778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_924 VNB N_VGND_c_12866_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_925 VNB VGND 2.38318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_926 VNB VGND 0.0109735f $X=25.905 $Y=0.425 $X2=0 $Y2=0
cc_927 VNB VGND 2.39416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_928 VNB N_VGND_c_12870_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_929 VNB N_VGND_c_12871_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_930 VNB N_VGND_c_12872_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_931 VNB N_VGND_c_12873_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_932 VNB N_VGND_c_12874_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_933 VNB N_VGND_c_12875_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_934 VNB N_VGND_c_12876_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_935 VNB N_VGND_c_12877_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_936 VNB N_VGND_c_12878_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_937 VNB N_VGND_c_12879_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_938 VNB N_VGND_c_12880_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_939 VNB N_VGND_c_12881_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_940 VNB N_VGND_c_12882_n 0.0211459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_941 VNB N_VGND_c_12882_n 0.0191027f $X=25.905 $Y=0.425 $X2=0 $Y2=0
cc_942 VNB N_VGND_c_12884_n 0.0402485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_943 VNB N_VGND_c_12885_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_944 VNB N_VGND_c_12886_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_945 VNB N_VGND_c_12887_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_946 VNB N_VGND_c_12888_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_947 VNB N_VGND_c_12889_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_948 VNB N_VGND_c_12890_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_949 VNB N_VGND_c_12891_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_950 VNB N_VGND_c_12892_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_951 VNB N_VGND_c_12893_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_952 VNB N_VGND_c_12894_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_953 VNB N_VGND_c_12895_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_954 VNB N_VGND_c_12896_n 0.017296f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_955 VNB N_VGND_c_12897_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_956 VNB N_VGND_c_12898_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_957 VNB N_VGND_c_12899_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_958 VNB N_VGND_c_12900_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_959 VNB N_VGND_c_12901_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_960 VNB N_VGND_c_12902_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_961 VNB N_VGND_c_12903_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_962 VNB N_VGND_c_12904_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_963 VNB N_VGND_c_12905_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_964 VNB N_VGND_c_12906_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_965 VNB N_VGND_c_12907_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_966 VNB N_VGND_c_12908_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_967 VNB N_VGND_c_12909_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_968 VNB N_VGND_c_12910_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_969 VNB N_VGND_c_12911_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_970 VNB N_VGND_c_12912_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_971 VNB N_VGND_c_12913_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_972 VNB N_VGND_c_12914_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_973 VNB N_VGND_c_12915_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_974 VNB N_VGND_c_12916_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_975 VNB N_VGND_c_12917_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_976 VNB N_VGND_c_12918_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_977 VNB N_VGND_c_12919_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_978 VNB N_VGND_c_12920_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_979 VNB N_VGND_c_12921_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_980 VNB N_VGND_c_12922_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_981 VNB N_VGND_c_12923_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_982 VNB N_VGND_c_12924_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_983 VNB N_VGND_c_12925_n 0.00480536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_984 VNB N_VGND_c_12926_n 0.00477947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_985 VNB N_VGND_c_12927_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_986 VNB N_VGND_c_12928_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_987 VNB N_VGND_c_12929_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_988 VNB N_VGND_c_12930_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_989 VNB N_VGND_c_12931_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_990 VNB N_VGND_c_12932_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_991 VNB N_A_119_47#_c_14049_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_992 VNB N_A_119_47#_c_14050_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=25.99 $Y2=1.73
cc_993 VNB N_A_119_47#_c_14051_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_994 VNB N_A_119_47#_c_14052_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_995 VNB N_A_119_47#_c_14053_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_996 VNB N_A_119_47#_c_14054_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_997 VNB N_A_119_47#_c_14055_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_998 VNB N_A_119_47#_c_14056_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_999 VNB N_A_119_911#_c_14132_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1000 VNB N_A_119_911#_c_14133_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1001 VNB N_A_119_911#_c_14134_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.87
cc_1002 VNB N_A_119_911#_c_14135_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1003 VNB N_A_119_911#_c_14136_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1004 VNB N_A_119_911#_c_14137_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1005 VNB N_A_119_911#_c_14138_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1006 VNB N_A_119_911#_c_14139_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1007 VNB N_A_1693_66#_c_14211_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1008 VNB N_A_1693_66#_c_14212_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1009 VNB N_A_1693_66#_c_14213_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1010 VNB N_A_1693_66#_c_14214_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1011 VNB N_A_1693_66#_c_14215_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1012 VNB N_A_1693_66#_c_14216_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1013 VNB N_A_1693_66#_c_14217_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1014 VNB N_A_1693_66#_c_14218_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1015 VNB N_A_1693_66#_c_14219_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1016 VNB N_A_1693_918#_c_14295_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1017 VNB N_A_1693_918#_c_14296_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1018 VNB N_A_1693_918#_c_14297_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1019 VNB N_A_1693_918#_c_14298_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1020 VNB N_A_1693_918#_c_14299_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1021 VNB N_A_1693_918#_c_14300_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1022 VNB N_A_1693_918#_c_14301_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1023 VNB N_A_1693_918#_c_14302_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1024 VNB N_A_1693_918#_c_14303_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1025 VNB N_A_2695_47#_c_14377_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1026 VNB N_A_2695_47#_c_14378_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1027 VNB N_A_2695_47#_c_14379_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1028 VNB N_A_2695_47#_c_14380_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1029 VNB N_A_2695_47#_c_14381_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1030 VNB N_A_2695_47#_c_14382_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1031 VNB N_A_2695_47#_c_14383_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1032 VNB N_A_2695_47#_c_14384_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1033 VNB N_A_2695_911#_c_14460_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1034 VNB N_A_2695_911#_c_14461_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1035 VNB N_A_2695_911#_c_14462_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.87
cc_1036 VNB N_A_2695_911#_c_14463_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1037 VNB N_A_2695_911#_c_14464_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1038 VNB N_A_2695_911#_c_14465_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1039 VNB N_A_2695_911#_c_14466_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1040 VNB N_A_2695_911#_c_14467_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1041 VNB N_A_4269_66#_c_14539_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1042 VNB N_A_4269_66#_c_14540_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1043 VNB N_A_4269_66#_c_14541_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1044 VNB N_A_4269_66#_c_14542_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1045 VNB N_A_4269_66#_c_14543_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1046 VNB N_A_4269_66#_c_14544_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1047 VNB N_A_4269_66#_c_14545_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1048 VNB N_A_4269_66#_c_14546_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1049 VNB N_A_4269_66#_c_14547_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1050 VNB N_A_4269_918#_c_14623_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1051 VNB N_A_4269_918#_c_14624_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1052 VNB N_A_4269_918#_c_14625_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1053 VNB N_A_4269_918#_c_14626_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1054 VNB N_A_4269_918#_c_14627_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1055 VNB N_A_4269_918#_c_14628_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1056 VNB N_A_4269_918#_c_14629_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1057 VNB N_A_4269_918#_c_14630_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1058 VNB N_A_4269_918#_c_14631_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1059 VNB N_A_5363_47#_c_14705_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1060 VNB N_A_5363_47#_c_14706_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1061 VNB N_A_5363_47#_c_14707_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1062 VNB N_A_5363_47#_c_14708_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1063 VNB N_A_5363_47#_c_14709_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1064 VNB N_A_5363_47#_c_14710_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1065 VNB N_A_5363_47#_c_14711_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1066 VNB N_A_5363_47#_c_14712_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1067 VNB N_A_5363_911#_c_14788_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1068 VNB N_A_5363_911#_c_14789_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1069 VNB N_A_5363_911#_c_14790_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.87
cc_1070 VNB N_A_5363_911#_c_14791_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1071 VNB N_A_5363_911#_c_14792_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1072 VNB N_A_5363_911#_c_14793_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1073 VNB N_A_5363_911#_c_14794_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1074 VNB N_A_5363_911#_c_14795_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1075 VNB N_A_6937_66#_c_14867_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1076 VNB N_A_6937_66#_c_14868_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1077 VNB N_A_6937_66#_c_14869_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1078 VNB N_A_6937_66#_c_14870_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1079 VNB N_A_6937_66#_c_14871_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1080 VNB N_A_6937_66#_c_14872_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1081 VNB N_A_6937_66#_c_14873_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1082 VNB N_A_6937_66#_c_14874_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1083 VNB N_A_6937_66#_c_14875_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1084 VNB N_A_6937_918#_c_14951_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1085 VNB N_A_6937_918#_c_14952_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1086 VNB N_A_6937_918#_c_14953_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1087 VNB N_A_6937_918#_c_14954_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1088 VNB N_A_6937_918#_c_14955_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1089 VNB N_A_6937_918#_c_14956_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1090 VNB N_A_6937_918#_c_14957_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1091 VNB N_A_6937_918#_c_14958_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1092 VNB N_A_6937_918#_c_14959_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1093 VNB N_A_7939_47#_c_15033_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1094 VNB N_A_7939_47#_c_15034_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1095 VNB N_A_7939_47#_c_15035_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1096 VNB N_A_7939_47#_c_15036_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1097 VNB N_A_7939_47#_c_15037_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1098 VNB N_A_7939_47#_c_15038_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1099 VNB N_A_7939_47#_c_15039_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1100 VNB N_A_7939_47#_c_15040_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1101 VNB N_A_7939_911#_c_15116_n 0.0126549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1102 VNB N_A_7939_911#_c_15117_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1103 VNB N_A_7939_911#_c_15118_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.87
cc_1104 VNB N_A_7939_911#_c_15119_n 0.00378884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1105 VNB N_A_7939_911#_c_15120_n 0.00453652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1106 VNB N_A_7939_911#_c_15121_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1107 VNB N_A_7939_911#_c_15122_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1108 VNB N_A_7939_911#_c_15123_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1109 VNB N_A_9513_66#_c_15195_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1110 VNB N_A_9513_66#_c_15196_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1111 VNB N_A_9513_66#_c_15197_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1112 VNB N_A_9513_66#_c_15198_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1113 VNB N_A_9513_66#_c_15199_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1114 VNB N_A_9513_66#_c_15200_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1115 VNB N_A_9513_66#_c_15201_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1116 VNB N_A_9513_66#_c_15202_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1117 VNB N_A_9513_66#_c_15203_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1118 VNB N_A_9513_918#_c_15279_n 0.0043971f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1119 VNB N_A_9513_918#_c_15280_n 0.00238176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1120 VNB N_A_9513_918#_c_15281_n 0.00215476f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1121 VNB N_A_9513_918#_c_15282_n 0.0061706f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=1.73
cc_1122 VNB N_A_9513_918#_c_15283_n 0.00317182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1123 VNB N_A_9513_918#_c_15284_n 0.00736637f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1124 VNB N_A_9513_918#_c_15285_n 0.00528854f $X=-0.19 $Y=-0.24 $X2=25.99
+ $Y2=3.23
cc_1125 VNB N_A_9513_918#_c_15286_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1126 VNB N_A_9513_918#_c_15287_n 0.00116392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_1127 VPB N_D[0]_M1014_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1128 VPB N_D[0]_M1146_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1129 VPB N_D[0]_M1208_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1130 VPB N_D[0]_M1294_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1131 VPB N_D[0]_c_1879_n 0.00910964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1132 VPB N_D[8]_M1023_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1133 VPB N_D[8]_M1155_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1134 VPB N_D[8]_M1221_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1135 VPB N_D[8]_M1304_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1136 VPB N_D[8]_c_1969_n 0.00910964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1137 VPB N_A_559_265#_c_2052_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1138 VPB N_A_559_265#_c_2053_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1139 VPB N_A_559_265#_c_2054_n 0.0168203f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1140 VPB N_A_559_265#_c_2055_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1141 VPB N_A_559_265#_c_2056_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1142 VPB N_A_559_265#_c_2057_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1143 VPB N_A_559_265#_c_2058_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1144 VPB N_A_559_265#_c_2059_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1145 VPB N_A_559_265#_c_2060_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1146 VPB N_A_559_265#_c_2061_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1147 VPB N_A_559_265#_c_2045_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1148 VPB N_A_559_265#_c_2046_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1149 VPB N_A_559_265#_c_2064_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1150 VPB N_A_559_265#_c_2050_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1151 VPB N_A_559_265#_c_2066_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1152 VPB N_A_559_265#_c_2051_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1153 VPB N_A_559_793#_c_2170_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1154 VPB N_A_559_793#_c_2171_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1155 VPB N_A_559_793#_c_2172_n 0.0168203f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1156 VPB N_A_559_793#_c_2173_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1157 VPB N_A_559_793#_c_2174_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1158 VPB N_A_559_793#_c_2175_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1159 VPB N_A_559_793#_c_2176_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1160 VPB N_A_559_793#_c_2177_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1161 VPB N_A_559_793#_c_2178_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1162 VPB N_A_559_793#_c_2179_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1163 VPB N_A_559_793#_c_2163_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1164 VPB N_A_559_793#_c_2164_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1165 VPB N_A_559_793#_c_2182_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1166 VPB N_A_559_793#_c_2183_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1167 VPB N_A_559_793#_c_2184_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1168 VPB N_A_559_793#_c_2167_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1169 VPB N_A_559_793#_c_2169_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1170 VPB N_S[0]_c_2299_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1171 VPB N_S[0]_c_2310_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1172 VPB N_S[0]_c_2303_n 0.0526479f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1173 VPB S[0] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1174 VPB N_S[8]_c_2425_n 0.00847786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1175 VPB N_S[8]_c_2416_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1176 VPB N_S[8]_c_2427_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1177 VPB N_S[8]_c_2419_n 0.0340992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1178 VPB N_S[8]_c_2429_n 0.0185487f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1179 VPB S[8] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1180 VPB N_S[1]_c_2529_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1181 VPB N_S[1]_c_2530_n 0.0394096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1182 VPB N_S[1]_c_2534_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1183 VPB N_S[1]_c_2554_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1184 VPB N_S[1]_c_2550_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1185 VPB N_S[9]_c_2649_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1186 VPB N_S[9]_c_2671_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1187 VPB N_S[9]_c_2650_n 0.0208609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1188 VPB N_S[9]_c_2673_n 0.00847786f $X=-0.19 $Y=1.305 $X2=25.905 $Y2=4.845
cc_1189 VPB N_S[9]_c_2652_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1190 VPB N_S[9]_c_2675_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1191 VPB N_S[9]_c_2669_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1192 VPB N_A_1430_325#_c_2784_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1193 VPB N_A_1430_325#_c_2785_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1194 VPB N_A_1430_325#_c_2777_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1195 VPB N_A_1430_325#_c_2787_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1196 VPB N_A_1430_325#_c_2788_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1197 VPB N_A_1430_325#_c_2789_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1198 VPB N_A_1430_325#_c_2790_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1199 VPB N_A_1430_325#_c_2791_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1200 VPB N_A_1430_325#_c_2792_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1201 VPB N_A_1430_325#_c_2793_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1202 VPB N_A_1430_325#_c_2794_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1203 VPB N_A_1430_325#_c_2780_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1204 VPB N_A_1430_325#_c_2796_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1205 VPB N_A_1430_325#_c_2782_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1206 VPB N_A_1430_325#_c_2783_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1207 VPB N_A_1430_599#_c_2900_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1208 VPB N_A_1430_599#_c_2901_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1209 VPB N_A_1430_599#_c_2893_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1210 VPB N_A_1430_599#_c_2903_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1211 VPB N_A_1430_599#_c_2904_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1212 VPB N_A_1430_599#_c_2905_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1213 VPB N_A_1430_599#_c_2906_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1214 VPB N_A_1430_599#_c_2907_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1215 VPB N_A_1430_599#_c_2908_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1216 VPB N_A_1430_599#_c_2909_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1217 VPB N_A_1430_599#_c_2910_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1218 VPB N_A_1430_599#_c_2911_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1219 VPB N_A_1430_599#_c_2896_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1220 VPB N_A_1430_599#_c_2913_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1221 VPB N_A_1430_599#_c_2898_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1222 VPB N_A_1430_599#_c_2899_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1223 VPB N_D[1]_M1002_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1224 VPB N_D[1]_M1038_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1225 VPB N_D[1]_M1134_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1226 VPB N_D[1]_M1271_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1227 VPB N_D[1]_c_3025_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1228 VPB N_D[9]_M1011_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1229 VPB N_D[9]_M1051_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1230 VPB N_D[9]_M1148_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1231 VPB N_D[9]_M1285_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1232 VPB N_D[9]_c_3118_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1233 VPB N_D[2]_M1020_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1234 VPB N_D[2]_M1067_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1235 VPB N_D[2]_M1157_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1236 VPB N_D[2]_M1301_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1237 VPB N_D[2]_c_3209_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1238 VPB N_D[10]_M1024_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1239 VPB N_D[10]_M1076_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1240 VPB N_D[10]_M1164_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1241 VPB N_D[10]_M1309_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1242 VPB N_D[10]_c_3304_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1243 VPB N_A_3135_265#_c_3392_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1244 VPB N_A_3135_265#_c_3393_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1245 VPB N_A_3135_265#_c_3394_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1246 VPB N_A_3135_265#_c_3395_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1247 VPB N_A_3135_265#_c_3396_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1248 VPB N_A_3135_265#_c_3397_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1249 VPB N_A_3135_265#_c_3398_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1250 VPB N_A_3135_265#_c_3399_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1251 VPB N_A_3135_265#_c_3400_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1252 VPB N_A_3135_265#_c_3401_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1253 VPB N_A_3135_265#_c_3385_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1254 VPB N_A_3135_265#_c_3386_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1255 VPB N_A_3135_265#_c_3404_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1256 VPB N_A_3135_265#_c_3390_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1257 VPB N_A_3135_265#_c_3406_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1258 VPB N_A_3135_265#_c_3391_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1259 VPB N_A_3135_793#_c_3511_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1260 VPB N_A_3135_793#_c_3512_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1261 VPB N_A_3135_793#_c_3513_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1262 VPB N_A_3135_793#_c_3514_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1263 VPB N_A_3135_793#_c_3515_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1264 VPB N_A_3135_793#_c_3516_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1265 VPB N_A_3135_793#_c_3517_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1266 VPB N_A_3135_793#_c_3518_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1267 VPB N_A_3135_793#_c_3519_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1268 VPB N_A_3135_793#_c_3520_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1269 VPB N_A_3135_793#_c_3504_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1270 VPB N_A_3135_793#_c_3505_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1271 VPB N_A_3135_793#_c_3523_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1272 VPB N_A_3135_793#_c_3524_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1273 VPB N_A_3135_793#_c_3525_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1274 VPB N_A_3135_793#_c_3508_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1275 VPB N_A_3135_793#_c_3510_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1276 VPB N_S[2]_c_3641_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1277 VPB N_S[2]_c_3652_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1278 VPB N_S[2]_c_3645_n 0.0526479f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1279 VPB S[2] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1280 VPB N_S[10]_c_3767_n 0.00847786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1281 VPB N_S[10]_c_3758_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1282 VPB N_S[10]_c_3769_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1283 VPB N_S[10]_c_3761_n 0.0340992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1284 VPB N_S[10]_c_3771_n 0.0185487f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1285 VPB S[10] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1286 VPB N_S[3]_c_3871_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1287 VPB N_S[3]_c_3872_n 0.0394096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1288 VPB N_S[3]_c_3876_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1289 VPB N_S[3]_c_3896_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1290 VPB N_S[3]_c_3892_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1291 VPB N_S[11]_c_3991_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1292 VPB N_S[11]_c_4013_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1293 VPB N_S[11]_c_3992_n 0.0208609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1294 VPB N_S[11]_c_4015_n 0.00847786f $X=-0.19 $Y=1.305 $X2=25.905 $Y2=4.845
cc_1295 VPB N_S[11]_c_3994_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1296 VPB N_S[11]_c_4017_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1297 VPB N_S[11]_c_4011_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1298 VPB N_A_4006_325#_c_4126_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1299 VPB N_A_4006_325#_c_4127_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1300 VPB N_A_4006_325#_c_4119_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1301 VPB N_A_4006_325#_c_4129_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1302 VPB N_A_4006_325#_c_4130_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1303 VPB N_A_4006_325#_c_4131_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1304 VPB N_A_4006_325#_c_4132_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1305 VPB N_A_4006_325#_c_4133_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1306 VPB N_A_4006_325#_c_4134_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1307 VPB N_A_4006_325#_c_4135_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1308 VPB N_A_4006_325#_c_4136_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1309 VPB N_A_4006_325#_c_4122_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1310 VPB N_A_4006_325#_c_4138_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1311 VPB N_A_4006_325#_c_4124_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1312 VPB N_A_4006_325#_c_4125_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1313 VPB N_A_4006_599#_c_4242_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1314 VPB N_A_4006_599#_c_4243_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1315 VPB N_A_4006_599#_c_4235_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1316 VPB N_A_4006_599#_c_4245_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1317 VPB N_A_4006_599#_c_4246_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1318 VPB N_A_4006_599#_c_4247_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1319 VPB N_A_4006_599#_c_4248_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1320 VPB N_A_4006_599#_c_4249_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1321 VPB N_A_4006_599#_c_4250_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1322 VPB N_A_4006_599#_c_4251_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1323 VPB N_A_4006_599#_c_4252_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1324 VPB N_A_4006_599#_c_4253_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1325 VPB N_A_4006_599#_c_4238_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1326 VPB N_A_4006_599#_c_4255_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1327 VPB N_A_4006_599#_c_4240_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1328 VPB N_A_4006_599#_c_4241_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1329 VPB N_D[3]_M1042_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1330 VPB N_D[3]_M1089_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1331 VPB N_D[3]_M1116_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1332 VPB N_D[3]_M1289_g 0.025177f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1333 N_VPB_c_1128_n N_D[3]_M1289_g 0.00204846f $X=25.99 $Y=1.73 $X2=25.99
+ $Y2=0.51
cc_1334 VPB N_D[3]_c_4367_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1335 VPB N_D[11]_M1052_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1336 VPB N_D[11]_M1101_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1337 VPB N_D[11]_M1129_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1338 VPB N_D[11]_M1297_g 0.025177f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1339 VPB N_D[11]_M1297_g 0.00204846f $X=25.905 $Y=3.145 $X2=25.99 $Y2=0.51
cc_1340 VPB N_D[11]_c_4461_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1341 VPB N_D[4]_M1158_g 0.025177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1342 N_VPB_c_1128_n N_D[4]_M1158_g 0.00204846f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1343 VPB N_D[4]_M1194_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1344 VPB N_D[4]_M1265_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1345 VPB N_D[4]_M1319_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1346 VPB N_D[4]_c_4553_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1347 VPB N_D[12]_M1006_g 0.025177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1348 VPB N_D[12]_M1006_g 0.00204846f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1349 VPB N_D[12]_M1165_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1350 VPB N_D[12]_M1203_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1351 VPB N_D[12]_M1277_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1352 VPB N_D[12]_c_4649_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1353 VPB N_A_5803_265#_c_4738_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1354 VPB N_A_5803_265#_c_4739_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1355 VPB N_A_5803_265#_c_4740_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1356 VPB N_A_5803_265#_c_4741_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1357 VPB N_A_5803_265#_c_4742_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1358 VPB N_A_5803_265#_c_4743_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1359 VPB N_A_5803_265#_c_4744_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1360 VPB N_A_5803_265#_c_4745_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1361 VPB N_A_5803_265#_c_4746_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1362 VPB N_A_5803_265#_c_4747_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1363 VPB N_A_5803_265#_c_4731_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1364 VPB N_A_5803_265#_c_4732_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1365 VPB N_A_5803_265#_c_4750_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1366 VPB N_A_5803_265#_c_4736_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1367 VPB N_A_5803_265#_c_4752_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1368 VPB N_A_5803_265#_c_4737_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1369 VPB N_A_5803_793#_c_4857_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1370 VPB N_A_5803_793#_c_4858_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1371 VPB N_A_5803_793#_c_4859_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1372 VPB N_A_5803_793#_c_4860_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1373 VPB N_A_5803_793#_c_4861_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1374 VPB N_A_5803_793#_c_4862_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1375 VPB N_A_5803_793#_c_4863_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1376 VPB N_A_5803_793#_c_4864_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1377 VPB N_A_5803_793#_c_4865_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1378 VPB N_A_5803_793#_c_4866_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1379 VPB N_A_5803_793#_c_4850_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1380 VPB N_A_5803_793#_c_4851_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1381 VPB N_A_5803_793#_c_4869_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1382 VPB N_A_5803_793#_c_4870_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1383 VPB N_A_5803_793#_c_4871_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1384 VPB N_A_5803_793#_c_4854_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1385 VPB N_A_5803_793#_c_4856_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1386 VPB N_S[4]_c_4987_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1387 VPB N_S[4]_c_4998_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1388 VPB N_S[4]_c_4991_n 0.0526479f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1389 VPB S[4] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1390 VPB N_S[12]_c_5113_n 0.00847786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1391 VPB N_S[12]_c_5104_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1392 VPB N_S[12]_c_5115_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1393 VPB N_S[12]_c_5107_n 0.0340992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1394 VPB N_S[12]_c_5117_n 0.0185487f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1395 VPB S[12] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1396 VPB N_S[5]_c_5217_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1397 VPB N_S[5]_c_5218_n 0.0394096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1398 VPB N_S[5]_c_5222_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1399 VPB N_S[5]_c_5242_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1400 VPB N_S[5]_c_5238_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1401 VPB N_S[13]_c_5337_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1402 VPB N_S[13]_c_5359_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1403 VPB N_S[13]_c_5338_n 0.0208609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1404 VPB N_S[13]_c_5361_n 0.00847786f $X=-0.19 $Y=1.305 $X2=25.905 $Y2=4.845
cc_1405 VPB N_S[13]_c_5340_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1406 VPB N_S[13]_c_5363_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1407 VPB N_S[13]_c_5357_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1408 VPB N_A_6674_325#_c_5472_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1409 VPB N_A_6674_325#_c_5473_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1410 VPB N_A_6674_325#_c_5465_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1411 VPB N_A_6674_325#_c_5475_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1412 VPB N_A_6674_325#_c_5476_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1413 VPB N_A_6674_325#_c_5477_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1414 VPB N_A_6674_325#_c_5478_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1415 VPB N_A_6674_325#_c_5479_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1416 VPB N_A_6674_325#_c_5480_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1417 VPB N_A_6674_325#_c_5481_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1418 VPB N_A_6674_325#_c_5482_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1419 VPB N_A_6674_325#_c_5468_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1420 VPB N_A_6674_325#_c_5484_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1421 VPB N_A_6674_325#_c_5470_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1422 VPB N_A_6674_325#_c_5471_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1423 VPB N_A_6674_599#_c_5588_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1424 VPB N_A_6674_599#_c_5589_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1425 VPB N_A_6674_599#_c_5581_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1426 VPB N_A_6674_599#_c_5591_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1427 VPB N_A_6674_599#_c_5592_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1428 VPB N_A_6674_599#_c_5593_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1429 VPB N_A_6674_599#_c_5594_n 0.0312612f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1430 VPB N_A_6674_599#_c_5595_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1431 VPB N_A_6674_599#_c_5596_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1432 VPB N_A_6674_599#_c_5597_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1433 VPB N_A_6674_599#_c_5598_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1434 VPB N_A_6674_599#_c_5599_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1435 VPB N_A_6674_599#_c_5584_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1436 VPB N_A_6674_599#_c_5601_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1437 VPB N_A_6674_599#_c_5586_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1438 VPB N_A_6674_599#_c_5587_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1439 VPB N_D[5]_M1088_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1440 VPB N_D[5]_M1183_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1441 VPB N_D[5]_M1217_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1442 VPB N_D[5]_M1255_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1443 VPB N_D[5]_c_5713_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1444 VPB N_D[13]_M1102_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1445 VPB N_D[13]_M1186_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1446 VPB N_D[13]_M1224_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1447 VPB N_D[13]_M1264_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1448 VPB N_D[13]_c_5806_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1449 VPB N_D[6]_M1099_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1450 VPB N_D[6]_M1176_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1451 VPB N_D[6]_M1246_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1452 VPB N_D[6]_M1282_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1453 VPB N_D[6]_c_5897_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1454 VPB N_D[14]_M1109_g 0.0254682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1455 VPB N_D[14]_M1184_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1456 VPB N_D[14]_M1251_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1457 VPB N_D[14]_M1293_g 0.0259085f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1458 VPB N_D[14]_c_5992_n 0.0083121f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1459 VPB N_A_8379_265#_c_6080_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1460 VPB N_A_8379_265#_c_6081_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1461 VPB N_A_8379_265#_c_6082_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1462 VPB N_A_8379_265#_c_6083_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1463 VPB N_A_8379_265#_c_6084_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1464 VPB N_A_8379_265#_c_6085_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1465 VPB N_A_8379_265#_c_6086_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1466 VPB N_A_8379_265#_c_6087_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1467 VPB N_A_8379_265#_c_6088_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1468 VPB N_A_8379_265#_c_6089_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1469 VPB N_A_8379_265#_c_6073_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1470 VPB N_A_8379_265#_c_6074_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1471 VPB N_A_8379_265#_c_6092_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1472 VPB N_A_8379_265#_c_6078_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1473 VPB N_A_8379_265#_c_6094_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1474 VPB N_A_8379_265#_c_6079_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1475 VPB N_A_8379_793#_c_6199_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1476 VPB N_A_8379_793#_c_6200_n 0.0145708f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1477 VPB N_A_8379_793#_c_6201_n 0.0166904f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1478 VPB N_A_8379_793#_c_6202_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1479 VPB N_A_8379_793#_c_6203_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1480 VPB N_A_8379_793#_c_6204_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1481 VPB N_A_8379_793#_c_6205_n 0.0140434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1482 VPB N_A_8379_793#_c_6206_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1483 VPB N_A_8379_793#_c_6207_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1484 VPB N_A_8379_793#_c_6208_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1485 VPB N_A_8379_793#_c_6192_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1486 VPB N_A_8379_793#_c_6193_n 0.0150864f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.64
cc_1487 VPB N_A_8379_793#_c_6211_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1488 VPB N_A_8379_793#_c_6212_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1489 VPB N_A_8379_793#_c_6213_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1490 VPB N_A_8379_793#_c_6196_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1491 VPB N_A_8379_793#_c_6198_n 0.0215299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1492 VPB N_S[6]_c_6329_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1493 VPB N_S[6]_c_6340_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1494 VPB N_S[6]_c_6333_n 0.0526479f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1495 VPB S[6] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1496 VPB N_S[14]_c_6455_n 0.00847786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1497 VPB N_S[14]_c_6446_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1498 VPB N_S[14]_c_6457_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1499 VPB N_S[14]_c_6449_n 0.0340992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1500 VPB N_S[14]_c_6459_n 0.0185487f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=4.8
cc_1501 VPB S[14] 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1502 VPB N_S[7]_c_6559_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1503 VPB N_S[7]_c_6560_n 0.0394096f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1504 VPB N_S[7]_c_6564_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1505 VPB N_S[7]_c_6584_n 0.0260812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1506 VPB N_S[7]_c_6580_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1507 VPB N_S[15]_c_6679_n 0.0132361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1508 VPB N_S[15]_c_6701_n 0.0185487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1509 VPB N_S[15]_c_6680_n 0.0208609f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1510 VPB N_S[15]_c_6703_n 0.00847786f $X=-0.19 $Y=1.305 $X2=25.905 $Y2=4.845
cc_1511 VPB N_S[15]_c_6682_n 0.00781808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1512 VPB N_S[15]_c_6705_n 0.0176033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1513 VPB N_S[15]_c_6699_n 4.51032e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1514 VPB N_A_9250_325#_c_6814_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1515 VPB N_A_9250_325#_c_6815_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1516 VPB N_A_9250_325#_c_6807_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1517 VPB N_A_9250_325#_c_6817_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1518 VPB N_A_9250_325#_c_6818_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1519 VPB N_A_9250_325#_c_6819_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1520 VPB N_A_9250_325#_c_6820_n 0.0313911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1521 VPB N_A_9250_325#_c_6821_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1522 VPB N_A_9250_325#_c_6822_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1523 VPB N_A_9250_325#_c_6823_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1524 VPB N_A_9250_325#_c_6824_n 0.00751381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1525 VPB N_A_9250_325#_c_6810_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1526 VPB N_A_9250_325#_c_6826_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1527 VPB N_A_9250_325#_c_6812_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1528 VPB N_A_9250_325#_c_6813_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1529 VPB N_A_9250_599#_c_6929_n 0.0231078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1530 VPB N_A_9250_599#_c_6930_n 0.0140434f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=0.425
cc_1531 VPB N_A_9250_599#_c_6922_n 0.0215299f $X=-0.19 $Y=1.305 $X2=25.905
+ $Y2=4.845
cc_1532 VPB N_A_9250_599#_c_6932_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1533 VPB N_A_9250_599#_c_6933_n 0.013221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1534 VPB N_A_9250_599#_c_6934_n 0.0174802f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1535 VPB N_A_9250_599#_c_6935_n 0.0313911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1536 VPB N_A_9250_599#_c_6936_n 0.0215147f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1537 VPB N_A_9250_599#_c_6937_n 0.00800249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1538 VPB N_A_9250_599#_c_6938_n 0.00747525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1539 VPB N_A_9250_599#_c_6939_n 0.0021116f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1540 VPB N_A_9250_599#_c_6940_n 0.00195069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1541 VPB N_A_9250_599#_c_6925_n 0.00733901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1542 VPB N_A_9250_599#_c_6942_n 0.00540221f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1543 VPB N_A_9250_599#_c_6927_n 9.02366e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1544 VPB N_A_9250_599#_c_6928_n 0.0150864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1545 VPB N_D[7]_M1040_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1546 VPB N_D[7]_M1087_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1547 VPB N_D[7]_M1131_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1548 VPB N_D[7]_M1151_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1549 VPB N_D[7]_c_7053_n 0.00910964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1550 VPB N_D[15]_M1056_g 0.0259085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1551 VPB N_D[15]_M1103_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1552 VPB N_D[15]_M1145_g 0.0177422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1553 VPB N_D[15]_M1156_g 0.0254682f $X=-0.19 $Y=1.305 $X2=25.99 $Y2=0.51
cc_1554 VPB N_D[15]_c_7141_n 0.00910964f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1555 VPB N_VPWR_c_7217_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1556 VPB N_VPWR_c_7218_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1557 VPB N_VPWR_c_7219_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1558 VPB N_VPWR_c_7220_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1559 VPB N_VPWR_c_7221_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1560 VPB N_VPWR_c_7222_n 0.00967963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1561 VPB N_VPWR_c_7223_n 0.00967963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1562 VPB N_VPWR_c_7224_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1563 VPB N_VPWR_c_7225_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1564 VPB N_VPWR_c_7226_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1565 VPB N_VPWR_c_7227_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1566 VPB N_VPWR_c_7228_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1567 VPB N_VPWR_c_7229_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1568 VPB N_VPWR_c_7230_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1569 VPB N_VPWR_c_7231_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1570 VPB N_VPWR_c_7232_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1571 VPB N_VPWR_c_7233_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1572 VPB N_VPWR_c_7234_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1573 VPB N_VPWR_c_7235_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1574 VPB N_VPWR_c_7236_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1575 VPB N_VPWR_c_7237_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1576 VPB N_VPWR_c_7238_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1577 VPB N_VPWR_c_7239_n 0.00789186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1578 VPB N_VPWR_c_7240_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1579 VPB N_VPWR_c_7241_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1580 VPB N_VPWR_c_7242_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1581 VPB N_VPWR_c_7243_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1582 VPB N_VPWR_c_7244_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1583 VPB N_VPWR_c_7245_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1584 VPB N_VPWR_c_7246_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1585 VPB N_VPWR_c_7247_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1586 VPB N_VPWR_c_7248_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1587 VPB N_VPWR_c_7249_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1588 VPB N_VPWR_c_7250_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1589 VPB N_VPWR_c_7251_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1590 VPB N_VPWR_c_7252_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1591 VPB N_VPWR_c_7253_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1592 VPB N_VPWR_c_7254_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1593 VPB N_VPWR_c_7255_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1594 VPB N_VPWR_c_7256_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1595 VPB N_VPWR_c_7257_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1596 VPB N_VPWR_c_7258_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1597 VPB N_VPWR_c_7259_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1598 VPB N_VPWR_c_7260_n 0.0151504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1599 N_VPB_c_1128_n N_VPWR_c_7260_n 0.0655801f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1600 VPB N_VPWR_c_7262_n 0.0151504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1601 VPB N_VPWR_c_7262_n 0.0655801f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1602 VPB N_VPWR_c_7264_n 0.0151504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1603 N_VPB_c_1128_n N_VPWR_c_7264_n 0.0655801f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1604 VPB N_VPWR_c_7266_n 0.0151504f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1605 VPB N_VPWR_c_7266_n 0.0655801f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1606 VPB N_VPWR_c_7268_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1607 VPB N_VPWR_c_7269_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1608 VPB N_VPWR_c_7270_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1609 VPB N_VPWR_c_7271_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1610 VPB N_VPWR_c_7272_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1611 VPB N_VPWR_c_7273_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1612 VPB N_VPWR_c_7274_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1613 VPB N_VPWR_c_7275_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1614 VPB N_VPWR_c_7276_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1615 VPB N_VPWR_c_7277_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1616 VPB N_VPWR_c_7278_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1617 VPB N_VPWR_c_7279_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1618 VPB N_VPWR_c_7280_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1619 VPB N_VPWR_c_7281_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1620 VPB N_VPWR_c_7282_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1621 VPB N_VPWR_c_7283_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1622 VPB N_VPWR_c_7284_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1623 VPB N_VPWR_c_7285_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1624 VPB N_VPWR_c_7286_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1625 VPB N_VPWR_c_7287_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1626 VPB N_VPWR_c_7288_n 0.00789186f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1627 VPB N_VPWR_c_7289_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1628 VPB N_VPWR_c_7290_n 0.0102368f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1629 VPB N_VPWR_c_7291_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1630 VPB N_VPWR_c_7292_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1631 VPB N_VPWR_c_7293_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1632 VPB N_VPWR_c_7294_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1633 VPB N_VPWR_c_7295_n 0.00924019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1634 VPB N_VPWR_c_7296_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1635 VPB N_VPWR_c_7297_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1636 VPB N_VPWR_c_7298_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1637 VPB N_VPWR_c_7299_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1638 VPB N_VPWR_c_7300_n 0.013938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1639 VPB N_VPWR_c_7301_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1640 VPB N_VPWR_c_7302_n 0.0187058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1641 VPB N_VPWR_c_7303_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1642 VPB N_VPWR_c_7304_n 0.0166787f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1643 VPB N_VPWR_c_7305_n 0.00967963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1644 VPB N_VPWR_c_7306_n 0.00967963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1645 VPB N_VPWR_c_7307_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1646 VPB N_VPWR_c_7308_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1647 VPB N_VPWR_c_7309_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1648 VPB N_VPWR_c_7310_n 0.0413001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1649 VPB N_VPWR_c_7311_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1650 VPB N_VPWR_c_7312_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1651 VPB N_VPWR_c_7313_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1652 VPB N_VPWR_c_7314_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1653 VPB N_VPWR_c_7315_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1654 VPB N_VPWR_c_7316_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1655 VPB N_VPWR_c_7317_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1656 VPB N_VPWR_c_7318_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1657 VPB N_VPWR_c_7319_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1658 VPB N_VPWR_c_7320_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1659 VPB N_VPWR_c_7321_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1660 VPB N_VPWR_c_7322_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1661 VPB N_VPWR_c_7323_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1662 VPB N_VPWR_c_7324_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1663 VPB N_VPWR_c_7325_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1664 VPB N_VPWR_c_7326_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1665 VPB N_VPWR_c_7327_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1666 VPB N_VPWR_c_7328_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1667 VPB N_VPWR_c_7329_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1668 VPB N_VPWR_c_7330_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1669 VPB N_VPWR_c_7331_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1670 VPB N_VPWR_c_7332_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1671 VPB N_VPWR_c_7333_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1672 VPB N_VPWR_c_7334_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1673 VPB N_VPWR_c_7335_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1674 VPB N_VPWR_c_7336_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1675 VPB N_VPWR_c_7337_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1676 VPB N_VPWR_c_7338_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1677 VPB N_VPWR_c_7339_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1678 VPB N_VPWR_c_7340_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1679 VPB N_VPWR_c_7341_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1680 VPB N_VPWR_c_7342_n 0.0121967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1681 VPB N_VPWR_c_7343_n 0.0154298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1682 VPB N_VPWR_c_7344_n 0.00172912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1683 VPB N_VPWR_c_7345_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1684 VPB N_VPWR_c_7346_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1685 VPB VPWR 0.306981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1686 VPB VPWR 0.00525875f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1687 N_VPB_c_1128_n VPWR 0.00525875f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1688 VPB N_VPWR_c_7350_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1689 VPB N_VPWR_c_7351_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1690 VPB N_VPWR_c_7352_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1691 VPB N_VPWR_c_7353_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1692 VPB N_VPWR_c_7354_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1693 VPB N_VPWR_c_7355_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1694 VPB N_VPWR_c_7356_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1695 VPB N_VPWR_c_7357_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1696 VPB N_VPWR_c_7358_n 0.017216f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1697 VPB N_VPWR_c_7358_n 0.0194225f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1698 N_VPB_c_1128_n N_VPWR_c_7358_n 0.0194225f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1699 VPB N_VPWR_c_7361_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1700 VPB N_VPWR_c_7362_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1701 VPB N_VPWR_c_7363_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1702 VPB N_VPWR_c_7364_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1703 VPB N_VPWR_c_7365_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1704 VPB N_VPWR_c_7366_n 0.0114011f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1705 VPB N_VPWR_c_7367_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1706 VPB N_VPWR_c_7368_n 0.0146409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1707 VPB N_VPWR_c_7369_n 0.00787932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1708 VPB N_VPWR_c_7370_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1709 VPB N_VPWR_c_7371_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1710 VPB N_VPWR_c_7372_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1711 VPB N_VPWR_c_7373_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1712 VPB N_VPWR_c_7374_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1713 VPB N_VPWR_c_7375_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1714 VPB N_VPWR_c_7376_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1715 VPB N_VPWR_c_7377_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1716 VPB N_VPWR_c_7378_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1717 VPB N_VPWR_c_7379_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1718 VPB N_VPWR_c_7380_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1719 VPB N_VPWR_c_7381_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1720 VPB N_VPWR_c_7382_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1721 VPB N_VPWR_c_7383_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1722 VPB N_VPWR_c_7384_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1723 VPB N_VPWR_c_7385_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1724 VPB N_VPWR_c_7386_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1725 VPB N_VPWR_c_7387_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1726 VPB N_VPWR_c_7388_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1727 VPB N_VPWR_c_7389_n 0.00169103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1728 VPB N_VPWR_c_7390_n 0.00187966f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1729 VPB N_VPWR_c_7391_n 0.00168437f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1730 VPB N_VPWR_c_7392_n 0.00787932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1731 VPB N_A_117_297#_c_8771_n 0.0158623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1732 VPB N_A_117_297#_c_8772_n 0.00328881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1733 VPB N_A_117_297#_c_8773_n 0.0109659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1734 VPB N_A_117_297#_c_8774_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1735 VPB N_A_117_297#_c_8775_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1736 VPB N_A_117_591#_c_8887_n 0.0158623f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1737 VPB N_A_117_591#_c_8888_n 0.00328881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1738 VPB N_A_117_591#_c_8889_n 0.0109659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1739 VPB N_A_117_591#_c_8890_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1740 VPB N_A_117_591#_c_8891_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1741 VPB N_Z_c_9046_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1742 VPB N_Z_c_9047_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1743 VPB N_Z_c_9052_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1744 VPB N_Z_c_9053_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1745 VPB N_Z_c_9060_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1746 VPB N_Z_c_9061_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1747 VPB N_Z_c_9066_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1748 VPB N_Z_c_9067_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1749 VPB N_Z_c_9074_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1750 VPB N_Z_c_9075_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1751 VPB N_Z_c_9080_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1752 VPB N_Z_c_9081_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1753 VPB N_Z_c_9088_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1754 VPB N_Z_c_9089_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1755 VPB N_Z_c_9094_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1756 VPB N_Z_c_9095_n 8.14549e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1757 VPB N_Z_c_9115_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1758 VPB N_Z_c_9116_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1759 VPB N_Z_c_9117_n 0.0192835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1760 VPB N_Z_c_9118_n 0.0192835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1761 VPB N_Z_c_9119_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1762 VPB N_Z_c_9120_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1763 VPB N_Z_c_9121_n 0.0274318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1764 N_VPB_c_1128_n N_Z_c_9121_n 0.029613f $X=25.99 $Y=1.73 $X2=0 $Y2=0
cc_1765 VPB N_Z_c_9123_n 0.0274318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1766 VPB N_Z_c_9123_n 0.029613f $X=25.905 $Y=3.145 $X2=0 $Y2=0
cc_1767 VPB N_Z_c_9125_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1768 VPB N_Z_c_9126_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1769 VPB N_Z_c_9127_n 0.0192835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1770 VPB N_Z_c_9128_n 0.0192835f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1771 VPB N_Z_c_9129_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1772 VPB N_Z_c_9130_n 0.0261782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1773 VPB N_Z_c_9131_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1774 VPB N_Z_c_9132_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1775 VPB N_Z_c_9133_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1776 VPB N_Z_c_9134_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1777 VPB N_Z_c_9135_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1778 VPB N_Z_c_9136_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1779 VPB N_Z_c_9137_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1780 VPB N_Z_c_9138_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1781 VPB N_Z_c_9139_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1782 VPB N_Z_c_9140_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1783 VPB N_Z_c_9141_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1784 VPB N_Z_c_9142_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1785 VPB N_Z_c_9143_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1786 VPB N_Z_c_9144_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1787 VPB N_Z_c_9145_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1788 VPB N_Z_c_9146_n 0.00296863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1789 VPB N_A_1643_311#_c_10897_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1790 VPB N_A_1643_311#_c_10898_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1791 VPB N_A_1643_311#_c_10899_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1792 VPB N_A_1643_311#_c_10900_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1793 VPB N_A_1643_311#_c_10901_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1794 VPB N_A_1643_311#_c_10902_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1795 VPB N_A_1643_613#_c_11028_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1796 VPB N_A_1643_613#_c_11029_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1797 VPB N_A_1643_613#_c_11030_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1798 VPB N_A_1643_613#_c_11031_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1799 VPB N_A_1643_613#_c_11032_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1800 VPB N_A_1643_613#_c_11033_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1801 VPB N_A_2693_297#_c_11159_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1802 VPB N_A_2693_297#_c_11160_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1803 VPB N_A_2693_297#_c_11161_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1804 VPB N_A_2693_297#_c_11162_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1805 VPB N_A_2693_297#_c_11163_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1806 VPB N_A_2693_591#_c_11287_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1807 VPB N_A_2693_591#_c_11288_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1808 VPB N_A_2693_591#_c_11289_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1809 VPB N_A_2693_591#_c_11290_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1810 VPB N_A_2693_591#_c_11291_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1811 VPB N_A_4219_311#_c_11415_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1812 VPB N_A_4219_311#_c_11416_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1813 VPB N_A_4219_311#_c_11417_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1814 VPB N_A_4219_311#_c_11418_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1815 VPB N_A_4219_311#_c_11419_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1816 VPB N_A_4219_311#_c_11420_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1817 VPB N_A_4219_613#_c_11546_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1818 VPB N_A_4219_613#_c_11547_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1819 VPB N_A_4219_613#_c_11548_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1820 VPB N_A_4219_613#_c_11549_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1821 VPB N_A_4219_613#_c_11550_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1822 VPB N_A_4219_613#_c_11551_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1823 VPB N_A_5361_297#_c_11677_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1824 VPB N_A_5361_297#_c_11678_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1825 VPB N_A_5361_297#_c_11679_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1826 VPB N_A_5361_297#_c_11680_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1827 VPB N_A_5361_297#_c_11681_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1828 VPB N_A_5361_591#_c_11805_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1829 VPB N_A_5361_591#_c_11806_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1830 VPB N_A_5361_591#_c_11807_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1831 VPB N_A_5361_591#_c_11808_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1832 VPB N_A_5361_591#_c_11809_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1833 VPB N_A_6887_311#_c_11933_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1834 VPB N_A_6887_311#_c_11934_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1835 VPB N_A_6887_311#_c_11935_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1836 VPB N_A_6887_311#_c_11936_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1837 VPB N_A_6887_311#_c_11937_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1838 VPB N_A_6887_311#_c_11938_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1839 VPB N_A_6887_613#_c_12064_n 0.0075016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1840 VPB N_A_6887_613#_c_12065_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1841 VPB N_A_6887_613#_c_12066_n 0.00219932f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1842 VPB N_A_6887_613#_c_12067_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1843 VPB N_A_6887_613#_c_12068_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1844 VPB N_A_6887_613#_c_12069_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1845 VPB N_A_7937_297#_c_12195_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1846 VPB N_A_7937_297#_c_12196_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1847 VPB N_A_7937_297#_c_12197_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1848 VPB N_A_7937_297#_c_12198_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1849 VPB N_A_7937_297#_c_12199_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1850 VPB N_A_7937_591#_c_12323_n 0.0147622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1851 VPB N_A_7937_591#_c_12324_n 0.00219932f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1852 VPB N_A_7937_591#_c_12325_n 0.0105341f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1853 VPB N_A_7937_591#_c_12326_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1854 VPB N_A_7937_591#_c_12327_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1855 VPB N_A_9463_311#_c_12451_n 0.00860164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1856 VPB N_A_9463_311#_c_12452_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1857 VPB N_A_9463_311#_c_12453_n 0.00328881f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1858 VPB N_A_9463_311#_c_12454_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1859 VPB N_A_9463_311#_c_12455_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1860 VPB N_A_9463_311#_c_12456_n 0.0109659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1861 VPB N_A_9463_613#_c_12570_n 0.00860164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1862 VPB N_A_9463_613#_c_12571_n 0.00726062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1863 VPB N_A_9463_613#_c_12572_n 0.00328881f $X=-0.19 $Y=1.305 $X2=25.99
+ $Y2=0.51
cc_1864 VPB N_A_9463_613#_c_12573_n 0.0123309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1865 VPB N_A_9463_613#_c_12574_n 0.00704236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1866 VPB N_A_9463_613#_c_12575_n 0.0109659f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_1867 N_D[0]_M1014_g N_D[8]_M1023_g 0.0130744f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_1868 N_D[0]_M1146_g N_D[8]_M1155_g 0.0130744f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_1869 N_D[0]_M1208_g N_D[8]_M1221_g 0.0130744f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_1870 N_D[0]_M1294_g N_D[8]_M1304_g 0.0130744f $X=1.905 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_1871 N_D[0]_M1014_g N_VPWR_c_7217_n 0.00354866f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_1872 N_D[0]_M1146_g N_VPWR_c_7219_n 0.00193762f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_1873 N_D[0]_M1208_g N_VPWR_c_7219_n 0.00193762f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_1874 N_D[0]_M1208_g N_VPWR_c_7221_n 0.0035837f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_1875 N_D[0]_M1294_g N_VPWR_c_7221_n 0.0035837f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_1876 N_D[0]_M1294_g N_VPWR_c_7222_n 0.00374733f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_1877 N_D[0]_M1014_g VPWR 0.0112159f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_1878 N_D[0]_M1146_g VPWR 0.00445624f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_1879 N_D[0]_M1208_g VPWR 0.00445624f $X=1.435 $Y=1.985 $X2=0 $Y2=0
cc_1880 N_D[0]_M1294_g VPWR 0.00573859f $X=1.905 $Y=1.985 $X2=0 $Y2=0
cc_1881 N_D[0]_M1014_g N_VPWR_c_7350_n 0.0035837f $X=0.495 $Y=1.985 $X2=0 $Y2=0
cc_1882 N_D[0]_M1146_g N_VPWR_c_7350_n 0.0035837f $X=0.965 $Y=1.985 $X2=0 $Y2=0
cc_1883 N_D[0]_M1146_g N_A_117_297#_c_8776_n 0.0102411f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_1884 N_D[0]_M1208_g N_A_117_297#_c_8776_n 0.0102411f $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1885 N_D[0]_c_1877_n N_A_117_297#_c_8776_n 7.15862e-19 $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_1886 N_D[0]_c_1879_n N_A_117_297#_c_8776_n 0.0405252f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1887 N_D[0]_M1294_g N_A_117_297#_c_8771_n 0.0143215f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_1888 N_D[0]_M1014_g N_A_117_297#_c_8781_n 0.00215964f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_1889 N_D[0]_M1146_g N_A_117_297#_c_8781_n 5.79575e-19 $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_1890 N_D[0]_c_1878_n N_A_117_297#_c_8781_n 8.03631e-19 $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_1891 N_D[0]_c_1879_n N_A_117_297#_c_8781_n 0.022724f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1892 N_D[0]_M1208_g N_A_117_297#_c_8785_n 5.79575e-19 $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1893 N_D[0]_M1294_g N_A_117_297#_c_8785_n 8.61029e-19 $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_1894 N_D[0]_c_1879_n N_A_117_297#_c_8785_n 0.0199757f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1895 N_D[0]_c_1880_n N_A_117_297#_c_8785_n 8.03631e-19 $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_1896 N_D[0]_M1146_g N_A_117_297#_c_8789_n 0.00316234f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_1897 N_D[0]_M1208_g N_A_117_297#_c_8789_n 0.00316234f $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1898 N_D[0]_M1294_g N_A_117_297#_c_8772_n 0.00316234f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_1899 N_D[0]_M1014_g N_A_117_297#_c_8792_n 0.00896273f $X=0.495 $Y=1.985 $X2=0
+ $Y2=0
cc_1900 N_D[0]_M1146_g N_A_117_297#_c_8792_n 0.0095928f $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_1901 N_D[0]_M1208_g N_A_117_297#_c_8792_n 6.38147e-19 $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1902 N_D[0]_M1146_g N_A_117_297#_c_8795_n 6.38147e-19 $X=0.965 $Y=1.985 $X2=0
+ $Y2=0
cc_1903 N_D[0]_M1208_g N_A_117_297#_c_8795_n 0.0095928f $X=1.435 $Y=1.985 $X2=0
+ $Y2=0
cc_1904 N_D[0]_M1294_g N_A_117_297#_c_8795_n 0.0104026f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_1905 N_D[0]_M1294_g N_A_117_297#_c_8773_n 0.0035027f $X=1.905 $Y=1.985 $X2=0
+ $Y2=0
cc_1906 N_D[0]_M1084_g N_VGND_c_12690_n 0.00345859f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_1907 N_D[0]_M1084_g N_VGND_c_12693_n 2.64031e-19 $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_1908 N_D[0]_M1219_g N_VGND_c_12693_n 0.00166854f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_1909 N_D[0]_M1300_g N_VGND_c_12693_n 0.0019152f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_1910 N_D[0]_M1300_g N_VGND_c_12695_n 0.00430643f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_1911 N_D[0]_M1317_g N_VGND_c_12695_n 0.00422241f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_1912 N_D[0]_M1300_g N_VGND_c_12697_n 2.6376e-19 $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_1913 N_D[0]_M1317_g N_VGND_c_12697_n 0.00321269f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_1914 N_D[0]_M1084_g VGND 0.0107845f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_1915 N_D[0]_M1219_g VGND 0.00593887f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_1916 N_D[0]_M1300_g VGND 0.00624811f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_1917 N_D[0]_M1317_g VGND 0.00702263f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_1918 N_D[0]_M1084_g N_VGND_c_12870_n 0.00551064f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_1919 N_D[0]_M1219_g N_VGND_c_12870_n 0.00422241f $X=0.94 $Y=0.56 $X2=0 $Y2=0
cc_1920 N_D[0]_M1084_g N_A_119_47#_c_14057_n 0.00529286f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_1921 N_D[0]_M1219_g N_A_119_47#_c_14057_n 0.00661134f $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1922 N_D[0]_M1300_g N_A_119_47#_c_14057_n 5.22365e-19 $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_1923 N_D[0]_M1219_g N_A_119_47#_c_14060_n 0.00899636f $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1924 N_D[0]_M1300_g N_A_119_47#_c_14060_n 0.00900364f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_1925 N_D[0]_c_1877_n N_A_119_47#_c_14060_n 0.00463549f $X=1.345 $Y=1.16 $X2=0
+ $Y2=0
cc_1926 N_D[0]_c_1879_n N_A_119_47#_c_14060_n 0.0394855f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1927 N_D[0]_M1084_g N_A_119_47#_c_14049_n 0.00228093f $X=0.52 $Y=0.56 $X2=0
+ $Y2=0
cc_1928 N_D[0]_M1219_g N_A_119_47#_c_14049_n 8.68782e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1929 N_D[0]_c_1878_n N_A_119_47#_c_14049_n 0.00208088f $X=1.055 $Y=1.16 $X2=0
+ $Y2=0
cc_1930 N_D[0]_c_1879_n N_A_119_47#_c_14049_n 0.021403f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1931 N_D[0]_M1219_g N_A_119_47#_c_14068_n 5.22365e-19 $X=0.94 $Y=0.56 $X2=0
+ $Y2=0
cc_1932 N_D[0]_M1300_g N_A_119_47#_c_14068_n 0.00661764f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_1933 N_D[0]_M1317_g N_A_119_47#_c_14068_n 0.00699463f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1934 N_D[0]_M1317_g N_A_119_47#_c_14050_n 0.0121912f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1935 N_D[0]_M1317_g N_A_119_47#_c_14051_n 0.00261078f $X=1.88 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_1936 N_D[0]_M1300_g N_A_119_47#_c_14056_n 8.68782e-19 $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_1937 N_D[0]_M1317_g N_A_119_47#_c_14056_n 0.00128201f $X=1.88 $Y=0.56 $X2=0
+ $Y2=0
cc_1938 N_D[0]_c_1879_n N_A_119_47#_c_14056_n 0.018367f $X=1.62 $Y=1.16 $X2=0
+ $Y2=0
cc_1939 N_D[0]_c_1880_n N_A_119_47#_c_14056_n 0.00208088f $X=1.905 $Y=1.16 $X2=0
+ $Y2=0
cc_1940 N_D[8]_M1023_g N_VPWR_c_7218_n 0.00354866f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_1941 N_D[8]_M1155_g N_VPWR_c_7220_n 0.00193762f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_1942 N_D[8]_M1221_g N_VPWR_c_7220_n 0.00193762f $X=1.435 $Y=3.455 $X2=0 $Y2=0
cc_1943 N_D[8]_M1221_g N_VPWR_c_7221_n 0.0035837f $X=1.435 $Y=3.455 $X2=0 $Y2=0
cc_1944 N_D[8]_M1304_g N_VPWR_c_7221_n 0.0035837f $X=1.905 $Y=3.455 $X2=0 $Y2=0
cc_1945 N_D[8]_M1304_g N_VPWR_c_7223_n 0.00374733f $X=1.905 $Y=3.455 $X2=0 $Y2=0
cc_1946 N_D[8]_M1023_g VPWR 0.0112159f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_1947 N_D[8]_M1155_g VPWR 0.00445624f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_1948 N_D[8]_M1221_g VPWR 0.00445624f $X=1.435 $Y=3.455 $X2=0 $Y2=0
cc_1949 N_D[8]_M1304_g VPWR 0.00573859f $X=1.905 $Y=3.455 $X2=0 $Y2=0
cc_1950 N_D[8]_M1023_g N_VPWR_c_7350_n 0.0035837f $X=0.495 $Y=3.455 $X2=0 $Y2=0
cc_1951 N_D[8]_M1155_g N_VPWR_c_7350_n 0.0035837f $X=0.965 $Y=3.455 $X2=0 $Y2=0
cc_1952 N_D[8]_M1155_g N_A_117_591#_c_8892_n 0.0102411f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_1953 N_D[8]_M1221_g N_A_117_591#_c_8892_n 0.0102411f $X=1.435 $Y=3.455 $X2=0
+ $Y2=0
cc_1954 N_D[8]_c_1967_n N_A_117_591#_c_8892_n 7.15862e-19 $X=1.345 $Y=4.28 $X2=0
+ $Y2=0
cc_1955 N_D[8]_c_1969_n N_A_117_591#_c_8892_n 0.0405252f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_1956 N_D[8]_M1304_g N_A_117_591#_c_8887_n 0.0143215f $X=1.905 $Y=3.455 $X2=0
+ $Y2=0
cc_1957 N_D[8]_M1023_g N_A_117_591#_c_8897_n 0.00215964f $X=0.495 $Y=3.455 $X2=0
+ $Y2=0
cc_1958 N_D[8]_M1155_g N_A_117_591#_c_8897_n 5.79575e-19 $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_1959 N_D[8]_c_1968_n N_A_117_591#_c_8897_n 8.03631e-19 $X=1.055 $Y=4.28 $X2=0
+ $Y2=0
cc_1960 N_D[8]_c_1969_n N_A_117_591#_c_8897_n 0.022724f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_1961 N_D[8]_M1221_g N_A_117_591#_c_8901_n 5.79575e-19 $X=1.435 $Y=3.455 $X2=0
+ $Y2=0
cc_1962 N_D[8]_M1304_g N_A_117_591#_c_8901_n 8.61029e-19 $X=1.905 $Y=3.455 $X2=0
+ $Y2=0
cc_1963 N_D[8]_c_1969_n N_A_117_591#_c_8901_n 0.0199757f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_1964 N_D[8]_c_1970_n N_A_117_591#_c_8901_n 8.03631e-19 $X=1.905 $Y=4.28 $X2=0
+ $Y2=0
cc_1965 N_D[8]_M1155_g N_A_117_591#_c_8905_n 0.00316234f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_1966 N_D[8]_M1221_g N_A_117_591#_c_8905_n 0.00316234f $X=1.435 $Y=3.455 $X2=0
+ $Y2=0
cc_1967 N_D[8]_M1304_g N_A_117_591#_c_8888_n 0.00316234f $X=1.905 $Y=3.455 $X2=0
+ $Y2=0
cc_1968 N_D[8]_M1023_g N_A_117_591#_c_8908_n 0.00896273f $X=0.495 $Y=3.455 $X2=0
+ $Y2=0
cc_1969 N_D[8]_M1155_g N_A_117_591#_c_8908_n 0.0095928f $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_1970 N_D[8]_M1221_g N_A_117_591#_c_8908_n 6.38147e-19 $X=1.435 $Y=3.455 $X2=0
+ $Y2=0
cc_1971 N_D[8]_M1155_g N_A_117_591#_c_8911_n 6.38147e-19 $X=0.965 $Y=3.455 $X2=0
+ $Y2=0
cc_1972 N_D[8]_M1221_g N_A_117_591#_c_8911_n 0.0095928f $X=1.435 $Y=3.455 $X2=0
+ $Y2=0
cc_1973 N_D[8]_M1304_g N_A_117_591#_c_8911_n 0.0104026f $X=1.905 $Y=3.455 $X2=0
+ $Y2=0
cc_1974 N_D[8]_M1304_g N_A_117_591#_c_8889_n 0.0035027f $X=1.905 $Y=3.455 $X2=0
+ $Y2=0
cc_1975 N_D[8]_M1085_g N_VGND_c_12692_n 0.00345859f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_1976 N_D[8]_M1085_g N_VGND_c_12694_n 2.64031e-19 $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_1977 N_D[8]_M1090_g N_VGND_c_12694_n 0.00166854f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_1978 N_D[8]_M1235_g N_VGND_c_12694_n 0.0019152f $X=1.46 $Y=4.88 $X2=0 $Y2=0
cc_1979 N_D[8]_M1235_g N_VGND_c_12696_n 0.00430643f $X=1.46 $Y=4.88 $X2=0 $Y2=0
cc_1980 N_D[8]_M1240_g N_VGND_c_12696_n 0.00422241f $X=1.88 $Y=4.88 $X2=0 $Y2=0
cc_1981 N_D[8]_M1235_g N_VGND_c_12698_n 2.6376e-19 $X=1.46 $Y=4.88 $X2=0 $Y2=0
cc_1982 N_D[8]_M1240_g N_VGND_c_12698_n 0.00321269f $X=1.88 $Y=4.88 $X2=0 $Y2=0
cc_1983 N_D[8]_M1085_g VGND 0.0107845f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_1984 N_D[8]_M1090_g VGND 0.00593887f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_1985 N_D[8]_M1235_g VGND 0.00624811f $X=1.46 $Y=4.88 $X2=0 $Y2=0
cc_1986 N_D[8]_M1240_g VGND 0.00702263f $X=1.88 $Y=4.88 $X2=0 $Y2=0
cc_1987 N_D[8]_M1085_g N_VGND_c_12871_n 0.00551064f $X=0.52 $Y=4.88 $X2=0 $Y2=0
cc_1988 N_D[8]_M1090_g N_VGND_c_12871_n 0.00422241f $X=0.94 $Y=4.88 $X2=0 $Y2=0
cc_1989 N_D[8]_M1090_g N_A_119_911#_c_14140_n 0.00899636f $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_1990 N_D[8]_M1235_g N_A_119_911#_c_14140_n 0.00900364f $X=1.46 $Y=4.88 $X2=0
+ $Y2=0
cc_1991 N_D[8]_c_1967_n N_A_119_911#_c_14140_n 0.00463549f $X=1.345 $Y=4.28
+ $X2=0 $Y2=0
cc_1992 N_D[8]_c_1969_n N_A_119_911#_c_14140_n 0.0394855f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_1993 N_D[8]_M1240_g N_A_119_911#_c_14132_n 0.0121912f $X=1.88 $Y=4.88 $X2=0
+ $Y2=0
cc_1994 N_D[8]_M1240_g N_A_119_911#_c_14133_n 0.00261078f $X=1.88 $Y=4.88 $X2=0
+ $Y2=0
cc_1995 N_D[8]_M1085_g N_A_119_911#_c_14138_n 0.00757379f $X=0.52 $Y=4.88 $X2=0
+ $Y2=0
cc_1996 N_D[8]_M1090_g N_A_119_911#_c_14138_n 0.00748012f $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_1997 N_D[8]_M1235_g N_A_119_911#_c_14138_n 5.22365e-19 $X=1.46 $Y=4.88 $X2=0
+ $Y2=0
cc_1998 N_D[8]_c_1968_n N_A_119_911#_c_14138_n 0.00208088f $X=1.055 $Y=4.28
+ $X2=0 $Y2=0
cc_1999 N_D[8]_c_1969_n N_A_119_911#_c_14138_n 0.021403f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_2000 N_D[8]_M1090_g N_A_119_911#_c_14139_n 5.22365e-19 $X=0.94 $Y=4.88 $X2=0
+ $Y2=0
cc_2001 N_D[8]_M1235_g N_A_119_911#_c_14139_n 0.00748643f $X=1.46 $Y=4.88 $X2=0
+ $Y2=0
cc_2002 N_D[8]_M1240_g N_A_119_911#_c_14139_n 0.00827664f $X=1.88 $Y=4.88 $X2=0
+ $Y2=0
cc_2003 N_D[8]_c_1969_n N_A_119_911#_c_14139_n 0.018367f $X=1.62 $Y=4.28 $X2=0
+ $Y2=0
cc_2004 N_D[8]_c_1970_n N_A_119_911#_c_14139_n 0.00208088f $X=1.905 $Y=4.28
+ $X2=0 $Y2=0
cc_2005 N_A_559_265#_c_2052_n N_A_559_793#_c_2170_n 0.0129371f $X=2.895 $Y=1.475
+ $X2=0 $Y2=0
cc_2006 N_A_559_265#_c_2055_n N_A_559_793#_c_2173_n 0.0129371f $X=3.365 $Y=1.475
+ $X2=0 $Y2=0
cc_2007 N_A_559_265#_c_2057_n N_A_559_793#_c_2175_n 0.0129371f $X=3.835 $Y=1.475
+ $X2=0 $Y2=0
cc_2008 N_A_559_265#_c_2059_n N_A_559_793#_c_2177_n 0.0129371f $X=4.305 $Y=1.475
+ $X2=0 $Y2=0
cc_2009 N_A_559_265#_c_2054_n N_S[0]_c_2287_n 0.00507426f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_2010 N_A_559_265#_c_2053_n N_S[0]_c_2290_n 0.00509391f $X=3.275 $Y=1.4 $X2=0
+ $Y2=0
cc_2011 N_A_559_265#_c_2056_n N_S[0]_c_2292_n 0.00509204f $X=3.745 $Y=1.4
+ $X2=25.905 $Y2=4.845
cc_2012 N_A_559_265#_c_2058_n N_S[0]_c_2294_n 0.00507688f $X=4.215 $Y=1.4 $X2=0
+ $Y2=0
cc_2013 N_A_559_265#_c_2047_n N_S[0]_c_2296_n 6.53442e-19 $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_2014 N_A_559_265#_c_2045_n N_S[0]_c_2298_n 0.0103812f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2015 N_A_559_265#_c_2046_n N_S[0]_c_2298_n 0.0179529f $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_2016 N_A_559_265#_c_2045_n N_S[0]_c_2299_n 0.0206368f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2017 N_A_559_265#_c_2046_n N_S[0]_c_2299_n 0.0175393f $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_2018 N_A_559_265#_c_2048_n N_S[0]_c_2299_n 0.0085951f $X=5.505 $Y=1.065 $X2=0
+ $Y2=0
cc_2019 N_A_559_265#_c_2050_n N_S[0]_c_2299_n 0.00322131f $X=5.505 $Y=1.23 $X2=0
+ $Y2=0
cc_2020 N_A_559_265#_c_2066_n N_S[0]_c_2299_n 0.00255921f $X=5.585 $Y=1.605
+ $X2=0 $Y2=0
cc_2021 N_A_559_265#_c_2051_n N_S[0]_c_2299_n 0.00262132f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_2022 N_A_559_265#_c_2064_n N_S[0]_c_2310_n 0.0118698f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_2023 N_A_559_265#_c_2066_n N_S[0]_c_2310_n 0.00762115f $X=5.585 $Y=1.605
+ $X2=0 $Y2=0
cc_2024 N_A_559_265#_c_2047_n N_S[0]_c_2300_n 0.00603996f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_2025 N_A_559_265#_c_2049_n N_S[0]_c_2300_n 9.67113e-19 $X=5.545 $Y=0.825
+ $X2=0 $Y2=0
cc_2026 N_A_559_265#_c_2048_n N_S[0]_c_2301_n 0.00429801f $X=5.505 $Y=1.065
+ $X2=0 $Y2=0
cc_2027 N_A_559_265#_c_2049_n N_S[0]_c_2301_n 0.0111895f $X=5.545 $Y=0.825 $X2=0
+ $Y2=0
cc_2028 N_A_559_265#_c_2047_n N_S[0]_c_2302_n 0.00207203f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_2029 N_A_559_265#_c_2048_n N_S[0]_c_2303_n 0.00289358f $X=5.505 $Y=1.065
+ $X2=25.99 $Y2=4.8
cc_2030 N_A_559_265#_c_2064_n N_S[0]_c_2303_n 0.0128834f $X=5.585 $Y=1.77
+ $X2=25.99 $Y2=4.8
cc_2031 N_A_559_265#_c_2050_n N_S[0]_c_2303_n 0.00416423f $X=5.505 $Y=1.23
+ $X2=25.99 $Y2=4.8
cc_2032 N_A_559_265#_c_2066_n N_S[0]_c_2303_n 0.00454075f $X=5.585 $Y=1.605
+ $X2=25.99 $Y2=4.8
cc_2033 N_A_559_265#_c_2048_n N_S[0]_c_2307_n 0.00268644f $X=5.505 $Y=1.065
+ $X2=0 $Y2=0
cc_2034 N_A_559_265#_c_2049_n N_S[0]_c_2307_n 0.00426435f $X=5.545 $Y=0.825
+ $X2=0 $Y2=0
cc_2035 N_A_559_265#_c_2048_n S[0] 0.00541767f $X=5.505 $Y=1.065 $X2=0 $Y2=0
cc_2036 N_A_559_265#_c_2050_n S[0] 0.0228692f $X=5.505 $Y=1.23 $X2=0 $Y2=0
cc_2037 N_A_559_265#_c_2052_n N_VPWR_c_7222_n 0.00331565f $X=2.895 $Y=1.475
+ $X2=0 $Y2=0
cc_2038 N_A_559_265#_c_2059_n N_VPWR_c_7224_n 0.00367058f $X=4.305 $Y=1.475
+ $X2=0 $Y2=0
cc_2039 N_A_559_265#_c_2045_n N_VPWR_c_7224_n 0.0193185f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2040 N_A_559_265#_c_2046_n N_VPWR_c_7224_n 6.4101e-19 $X=4.875 $Y=1.23 $X2=0
+ $Y2=0
cc_2041 N_A_559_265#_c_2064_n N_VPWR_c_7224_n 0.0316788f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_2042 N_A_559_265#_c_2064_n N_VPWR_c_7226_n 0.0356181f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_2043 N_A_559_265#_c_2064_n N_VPWR_c_7313_n 0.0233824f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_2044 N_A_559_265#_c_2052_n VPWR 0.00473731f $X=2.895 $Y=1.475 $X2=0 $Y2=0
cc_2045 N_A_559_265#_c_2055_n VPWR 0.00362156f $X=3.365 $Y=1.475 $X2=0 $Y2=0
cc_2046 N_A_559_265#_c_2057_n VPWR 0.00362156f $X=3.835 $Y=1.475 $X2=0 $Y2=0
cc_2047 N_A_559_265#_c_2059_n VPWR 0.00473731f $X=4.305 $Y=1.475 $X2=0 $Y2=0
cc_2048 N_A_559_265#_c_2064_n VPWR 0.00593513f $X=5.585 $Y=1.77 $X2=0 $Y2=0
cc_2049 N_A_559_265#_c_2052_n N_A_117_297#_c_8771_n 0.00151141f $X=2.895
+ $Y=1.475 $X2=0 $Y2=0
cc_2050 N_A_559_265#_c_2052_n N_A_117_297#_c_8800_n 0.00799829f $X=2.895
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_2051 N_A_559_265#_c_2055_n N_A_117_297#_c_8800_n 0.00307958f $X=3.365
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_2052 N_A_559_265#_c_2057_n N_A_117_297#_c_8802_n 0.00307958f $X=3.835
+ $Y=1.475 $X2=0 $Y2=0
cc_2053 N_A_559_265#_c_2059_n N_A_117_297#_c_8802_n 0.00307958f $X=4.305
+ $Y=1.475 $X2=0 $Y2=0
cc_2054 N_A_559_265#_c_2052_n N_A_117_297#_c_8773_n 0.00546785f $X=2.895
+ $Y=1.475 $X2=0 $Y2=0
cc_2055 N_A_559_265#_c_2055_n N_A_117_297#_c_8774_n 0.00210632f $X=3.365
+ $Y=1.475 $X2=0 $Y2=0
cc_2056 N_A_559_265#_c_2056_n N_A_117_297#_c_8774_n 0.00251792f $X=3.745 $Y=1.4
+ $X2=0 $Y2=0
cc_2057 N_A_559_265#_c_2057_n N_A_117_297#_c_8774_n 0.00210632f $X=3.835
+ $Y=1.475 $X2=0 $Y2=0
cc_2058 N_A_559_265#_c_2059_n N_A_117_297#_c_8775_n 0.00499839f $X=4.305
+ $Y=1.475 $X2=0 $Y2=0
cc_2059 N_A_559_265#_c_2045_n N_A_117_297#_c_8775_n 0.0218124f $X=5.42 $Y=1.23
+ $X2=0 $Y2=0
cc_2060 N_A_559_265#_c_2046_n N_A_117_297#_c_8775_n 5.74251e-19 $X=4.875 $Y=1.23
+ $X2=0 $Y2=0
cc_2061 N_A_559_265#_c_2051_n N_A_117_297#_c_8775_n 0.00561627f $X=4.625 $Y=1.23
+ $X2=0 $Y2=0
cc_2062 N_A_559_265#_c_2056_n N_Z_c_9004_n 0.00762343f $X=3.745 $Y=1.4 $X2=0
+ $Y2=0
cc_2063 N_A_559_265#_c_2060_n N_Z_c_9004_n 0.00704092f $X=3.365 $Y=1.4 $X2=0
+ $Y2=0
cc_2064 N_A_559_265#_c_2054_n N_Z_c_9043_n 0.00248496f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_2065 N_A_559_265#_c_2053_n N_Z_c_9046_n 0.00678861f $X=3.275 $Y=1.4 $X2=0
+ $Y2=0
cc_2066 N_A_559_265#_c_2054_n N_Z_c_9046_n 0.00239476f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_2067 N_A_559_265#_c_2060_n N_Z_c_9046_n 2.98555e-19 $X=3.365 $Y=1.4 $X2=0
+ $Y2=0
cc_2068 N_A_559_265#_c_2056_n N_Z_c_9048_n 0.00145542f $X=3.745 $Y=1.4 $X2=0
+ $Y2=0
cc_2069 N_A_559_265#_c_2058_n N_Z_c_9048_n 0.00597584f $X=4.215 $Y=1.4 $X2=0
+ $Y2=0
cc_2070 N_A_559_265#_c_2061_n N_Z_c_9048_n 0.00909323f $X=3.835 $Y=1.4 $X2=0
+ $Y2=0
cc_2071 N_A_559_265#_c_2045_n N_Z_c_9048_n 0.0266078f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2072 N_A_559_265#_c_2051_n N_Z_c_9048_n 0.00747617f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_2073 N_A_559_265#_c_2059_n N_Z_c_9115_n 0.00795576f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_2074 N_A_559_265#_c_2045_n N_Z_c_9115_n 0.0186685f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2075 N_A_559_265#_c_2064_n N_Z_c_9115_n 0.0329704f $X=5.585 $Y=1.77 $X2=0
+ $Y2=0
cc_2076 N_A_559_265#_c_2051_n N_Z_c_9115_n 2.19754e-19 $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_2077 N_A_559_265#_c_2055_n Z 0.00372458f $X=3.365 $Y=1.475 $X2=0 $Y2=0
cc_2078 N_A_559_265#_c_2057_n Z 0.00372248f $X=3.835 $Y=1.475 $X2=0 $Y2=0
cc_2079 N_A_559_265#_c_2052_n N_Z_c_9131_n 0.020403f $X=2.895 $Y=1.475 $X2=0
+ $Y2=0
cc_2080 N_A_559_265#_c_2053_n N_Z_c_9131_n 0.00560592f $X=3.275 $Y=1.4 $X2=0
+ $Y2=0
cc_2081 N_A_559_265#_c_2054_n N_Z_c_9131_n 0.00474497f $X=2.985 $Y=1.4 $X2=0
+ $Y2=0
cc_2082 N_A_559_265#_c_2055_n N_Z_c_9131_n 0.0181262f $X=3.365 $Y=1.475 $X2=0
+ $Y2=0
cc_2083 N_A_559_265#_c_2057_n N_Z_c_9131_n 9.74366e-19 $X=3.835 $Y=1.475 $X2=0
+ $Y2=0
cc_2084 N_A_559_265#_c_2060_n N_Z_c_9131_n 0.00415268f $X=3.365 $Y=1.4 $X2=0
+ $Y2=0
cc_2085 N_A_559_265#_c_2055_n N_Z_c_9132_n 9.74366e-19 $X=3.365 $Y=1.475 $X2=0
+ $Y2=0
cc_2086 N_A_559_265#_c_2057_n N_Z_c_9132_n 0.0181262f $X=3.835 $Y=1.475 $X2=0
+ $Y2=0
cc_2087 N_A_559_265#_c_2058_n N_Z_c_9132_n 0.00560592f $X=4.215 $Y=1.4 $X2=0
+ $Y2=0
cc_2088 N_A_559_265#_c_2059_n N_Z_c_9132_n 0.0221748f $X=4.305 $Y=1.475 $X2=0
+ $Y2=0
cc_2089 N_A_559_265#_c_2061_n N_Z_c_9132_n 0.00181273f $X=3.835 $Y=1.4 $X2=0
+ $Y2=0
cc_2090 N_A_559_265#_c_2045_n N_Z_c_9132_n 0.00240108f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2091 N_A_559_265#_c_2051_n N_Z_c_9132_n 0.00425035f $X=4.625 $Y=1.23 $X2=0
+ $Y2=0
cc_2092 N_A_559_265#_c_2045_n N_VGND_c_12699_n 0.0123065f $X=5.42 $Y=1.23 $X2=0
+ $Y2=0
cc_2093 N_A_559_265#_c_2046_n N_VGND_c_12699_n 2.04129e-19 $X=4.875 $Y=1.23
+ $X2=0 $Y2=0
cc_2094 N_A_559_265#_c_2047_n N_VGND_c_12791_n 0.0129994f $X=5.585 $Y=0.445
+ $X2=0 $Y2=0
cc_2095 N_A_559_265#_M1139_d VGND 0.00394793f $X=5.45 $Y=0.235 $X2=0 $Y2=0
cc_2096 N_A_559_265#_c_2047_n VGND 0.00927134f $X=5.585 $Y=0.445 $X2=0 $Y2=0
cc_2097 N_A_559_265#_c_2060_n N_A_119_47#_c_14077_n 7.0477e-19 $X=3.365 $Y=1.4
+ $X2=0 $Y2=0
cc_2098 N_A_559_265#_c_2045_n N_A_119_47#_c_14055_n 0.0028695f $X=5.42 $Y=1.23
+ $X2=25.99 $Y2=4.93
cc_2099 N_A_559_265#_c_2051_n N_A_119_47#_c_14055_n 0.00589316f $X=4.625 $Y=1.23
+ $X2=25.99 $Y2=4.93
cc_2100 N_A_559_793#_c_2172_n N_S[8]_c_2404_n 0.00507426f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_2101 N_A_559_793#_c_2171_n N_S[8]_c_2407_n 0.00509391f $X=3.275 $Y=4.04 $X2=0
+ $Y2=0
cc_2102 N_A_559_793#_c_2174_n N_S[8]_c_2409_n 0.00509204f $X=3.745 $Y=4.04
+ $X2=25.905 $Y2=4.845
cc_2103 N_A_559_793#_c_2176_n N_S[8]_c_2411_n 0.00507688f $X=4.215 $Y=4.04 $X2=0
+ $Y2=0
cc_2104 N_A_559_793#_c_2165_n N_S[8]_c_2413_n 6.53442e-19 $X=5.545 $Y=4.74 $X2=0
+ $Y2=0
cc_2105 N_A_559_793#_c_2163_n N_S[8]_c_2415_n 0.0103812f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2106 N_A_559_793#_c_2164_n N_S[8]_c_2415_n 0.0179529f $X=4.875 $Y=4.21 $X2=0
+ $Y2=0
cc_2107 N_A_559_793#_c_2183_n N_S[8]_c_2425_n 0.00508008f $X=5.505 $Y=4.045
+ $X2=0 $Y2=0
cc_2108 N_A_559_793#_c_2169_n N_S[8]_c_2425_n 0.00262132f $X=4.625 $Y=4.21 $X2=0
+ $Y2=0
cc_2109 N_A_559_793#_c_2163_n N_S[8]_c_2416_n 0.0206368f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2110 N_A_559_793#_c_2164_n N_S[8]_c_2416_n 0.0175393f $X=4.875 $Y=4.21 $X2=0
+ $Y2=0
cc_2111 N_A_559_793#_c_2183_n N_S[8]_c_2416_n 0.00255921f $X=5.505 $Y=4.045
+ $X2=0 $Y2=0
cc_2112 N_A_559_793#_c_2167_n N_S[8]_c_2416_n 0.00322131f $X=5.505 $Y=4.21 $X2=0
+ $Y2=0
cc_2113 N_A_559_793#_c_2168_n N_S[8]_c_2416_n 0.0085951f $X=5.545 $Y=4.615 $X2=0
+ $Y2=0
cc_2114 N_A_559_793#_c_2182_n N_S[8]_c_2427_n 0.00970559f $X=5.585 $Y=3.14 $X2=0
+ $Y2=0
cc_2115 N_A_559_793#_c_2183_n N_S[8]_c_2427_n 0.00254107f $X=5.505 $Y=4.045
+ $X2=0 $Y2=0
cc_2116 N_A_559_793#_c_2184_n N_S[8]_c_2427_n 0.00216424f $X=5.585 $Y=3.835
+ $X2=0 $Y2=0
cc_2117 N_A_559_793#_c_2165_n N_S[8]_c_2417_n 9.67113e-19 $X=5.545 $Y=4.74 $X2=0
+ $Y2=0
cc_2118 N_A_559_793#_c_2166_n N_S[8]_c_2417_n 0.00603996f $X=5.585 $Y=4.995
+ $X2=0 $Y2=0
cc_2119 N_A_559_793#_c_2165_n N_S[8]_c_2418_n 0.0111895f $X=5.545 $Y=4.74 $X2=0
+ $Y2=0
cc_2120 N_A_559_793#_c_2168_n N_S[8]_c_2418_n 0.00429801f $X=5.545 $Y=4.615
+ $X2=0 $Y2=0
cc_2121 N_A_559_793#_c_2183_n N_S[8]_c_2419_n 0.00336772f $X=5.505 $Y=4.045
+ $X2=0 $Y2=0
cc_2122 N_A_559_793#_c_2165_n N_S[8]_c_2419_n 0.00207203f $X=5.545 $Y=4.74 $X2=0
+ $Y2=0
cc_2123 N_A_559_793#_c_2184_n N_S[8]_c_2419_n 5.48523e-19 $X=5.585 $Y=3.835
+ $X2=0 $Y2=0
cc_2124 N_A_559_793#_c_2167_n N_S[8]_c_2419_n 0.00416423f $X=5.505 $Y=4.21 $X2=0
+ $Y2=0
cc_2125 N_A_559_793#_c_2168_n N_S[8]_c_2419_n 0.00289358f $X=5.545 $Y=4.615
+ $X2=0 $Y2=0
cc_2126 N_A_559_793#_c_2182_n N_S[8]_c_2429_n 0.00929139f $X=5.585 $Y=3.14
+ $X2=25.99 $Y2=4.8
cc_2127 N_A_559_793#_c_2183_n N_S[8]_c_2429_n 0.00117303f $X=5.505 $Y=4.045
+ $X2=25.99 $Y2=4.8
cc_2128 N_A_559_793#_c_2184_n N_S[8]_c_2429_n 0.00304348f $X=5.585 $Y=3.835
+ $X2=25.99 $Y2=4.8
cc_2129 N_A_559_793#_c_2165_n N_S[8]_c_2423_n 0.00426435f $X=5.545 $Y=4.74 $X2=0
+ $Y2=0
cc_2130 N_A_559_793#_c_2168_n N_S[8]_c_2423_n 0.00268644f $X=5.545 $Y=4.615
+ $X2=0 $Y2=0
cc_2131 N_A_559_793#_c_2167_n S[8] 0.0228692f $X=5.505 $Y=4.21 $X2=0 $Y2=0
cc_2132 N_A_559_793#_c_2168_n S[8] 0.00541767f $X=5.545 $Y=4.615 $X2=0 $Y2=0
cc_2133 N_A_559_793#_c_2170_n N_VPWR_c_7223_n 0.00331565f $X=2.895 $Y=3.965
+ $X2=0 $Y2=0
cc_2134 N_A_559_793#_c_2177_n N_VPWR_c_7225_n 0.00367058f $X=4.305 $Y=3.965
+ $X2=0 $Y2=0
cc_2135 N_A_559_793#_c_2163_n N_VPWR_c_7225_n 0.0193185f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2136 N_A_559_793#_c_2164_n N_VPWR_c_7225_n 6.4101e-19 $X=4.875 $Y=4.21 $X2=0
+ $Y2=0
cc_2137 N_A_559_793#_c_2182_n N_VPWR_c_7225_n 0.0316788f $X=5.585 $Y=3.14 $X2=0
+ $Y2=0
cc_2138 N_A_559_793#_c_2182_n N_VPWR_c_7227_n 0.0356181f $X=5.585 $Y=3.14 $X2=0
+ $Y2=0
cc_2139 N_A_559_793#_c_2182_n N_VPWR_c_7313_n 0.0233824f $X=5.585 $Y=3.14 $X2=0
+ $Y2=0
cc_2140 N_A_559_793#_c_2170_n VPWR 0.00473731f $X=2.895 $Y=3.965 $X2=0 $Y2=0
cc_2141 N_A_559_793#_c_2173_n VPWR 0.00362156f $X=3.365 $Y=3.965 $X2=0 $Y2=0
cc_2142 N_A_559_793#_c_2175_n VPWR 0.00362156f $X=3.835 $Y=3.965 $X2=0 $Y2=0
cc_2143 N_A_559_793#_c_2177_n VPWR 0.00473731f $X=4.305 $Y=3.965 $X2=0 $Y2=0
cc_2144 N_A_559_793#_c_2182_n VPWR 0.00593513f $X=5.585 $Y=3.14 $X2=0 $Y2=0
cc_2145 N_A_559_793#_c_2170_n N_A_117_591#_c_8887_n 0.00151141f $X=2.895
+ $Y=3.965 $X2=0 $Y2=0
cc_2146 N_A_559_793#_c_2170_n N_A_117_591#_c_8916_n 0.00799829f $X=2.895
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_2147 N_A_559_793#_c_2173_n N_A_117_591#_c_8916_n 0.00307958f $X=3.365
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_2148 N_A_559_793#_c_2175_n N_A_117_591#_c_8918_n 0.00307958f $X=3.835
+ $Y=3.965 $X2=0 $Y2=0
cc_2149 N_A_559_793#_c_2177_n N_A_117_591#_c_8918_n 0.00307958f $X=4.305
+ $Y=3.965 $X2=0 $Y2=0
cc_2150 N_A_559_793#_c_2170_n N_A_117_591#_c_8889_n 0.00546785f $X=2.895
+ $Y=3.965 $X2=0 $Y2=0
cc_2151 N_A_559_793#_c_2173_n N_A_117_591#_c_8890_n 0.00210632f $X=3.365
+ $Y=3.965 $X2=0 $Y2=0
cc_2152 N_A_559_793#_c_2174_n N_A_117_591#_c_8890_n 0.00251792f $X=3.745 $Y=4.04
+ $X2=0 $Y2=0
cc_2153 N_A_559_793#_c_2175_n N_A_117_591#_c_8890_n 0.00210632f $X=3.835
+ $Y=3.965 $X2=0 $Y2=0
cc_2154 N_A_559_793#_c_2177_n N_A_117_591#_c_8891_n 0.00499839f $X=4.305
+ $Y=3.965 $X2=0 $Y2=0
cc_2155 N_A_559_793#_c_2163_n N_A_117_591#_c_8891_n 0.0218124f $X=5.42 $Y=4.21
+ $X2=0 $Y2=0
cc_2156 N_A_559_793#_c_2164_n N_A_117_591#_c_8891_n 5.74251e-19 $X=4.875 $Y=4.21
+ $X2=0 $Y2=0
cc_2157 N_A_559_793#_c_2169_n N_A_117_591#_c_8891_n 0.00561627f $X=4.625 $Y=4.21
+ $X2=0 $Y2=0
cc_2158 N_A_559_793#_c_2174_n N_Z_c_9005_n 0.00762343f $X=3.745 $Y=4.04 $X2=0
+ $Y2=0
cc_2159 N_A_559_793#_c_2178_n N_Z_c_9005_n 0.00704092f $X=3.365 $Y=4.04 $X2=0
+ $Y2=0
cc_2160 N_A_559_793#_c_2172_n N_Z_c_9044_n 0.00248496f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_2161 N_A_559_793#_c_2171_n N_Z_c_9047_n 0.00678861f $X=3.275 $Y=4.04 $X2=0
+ $Y2=0
cc_2162 N_A_559_793#_c_2172_n N_Z_c_9047_n 0.00239476f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_2163 N_A_559_793#_c_2178_n N_Z_c_9047_n 2.98555e-19 $X=3.365 $Y=4.04 $X2=0
+ $Y2=0
cc_2164 N_A_559_793#_c_2174_n N_Z_c_9049_n 0.00145542f $X=3.745 $Y=4.04 $X2=0
+ $Y2=0
cc_2165 N_A_559_793#_c_2176_n N_Z_c_9049_n 0.00597584f $X=4.215 $Y=4.04 $X2=0
+ $Y2=0
cc_2166 N_A_559_793#_c_2179_n N_Z_c_9049_n 0.00909323f $X=3.835 $Y=4.04 $X2=0
+ $Y2=0
cc_2167 N_A_559_793#_c_2163_n N_Z_c_9049_n 0.0266078f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2168 N_A_559_793#_c_2169_n N_Z_c_9049_n 0.00747617f $X=4.625 $Y=4.21 $X2=0
+ $Y2=0
cc_2169 N_A_559_793#_c_2177_n N_Z_c_9116_n 0.00795576f $X=4.305 $Y=3.965 $X2=0
+ $Y2=0
cc_2170 N_A_559_793#_c_2163_n N_Z_c_9116_n 0.0186685f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2171 N_A_559_793#_c_2182_n N_Z_c_9116_n 0.0329704f $X=5.585 $Y=3.14 $X2=0
+ $Y2=0
cc_2172 N_A_559_793#_c_2169_n N_Z_c_9116_n 2.19754e-19 $X=4.625 $Y=4.21 $X2=0
+ $Y2=0
cc_2173 N_A_559_793#_c_2173_n Z 0.00372458f $X=3.365 $Y=3.965 $X2=0 $Y2=0
cc_2174 N_A_559_793#_c_2175_n Z 0.00372248f $X=3.835 $Y=3.965 $X2=0 $Y2=0
cc_2175 N_A_559_793#_c_2170_n N_Z_c_9131_n 0.020403f $X=2.895 $Y=3.965 $X2=0
+ $Y2=0
cc_2176 N_A_559_793#_c_2171_n N_Z_c_9131_n 0.00560592f $X=3.275 $Y=4.04 $X2=0
+ $Y2=0
cc_2177 N_A_559_793#_c_2172_n N_Z_c_9131_n 0.00474497f $X=2.985 $Y=4.04 $X2=0
+ $Y2=0
cc_2178 N_A_559_793#_c_2173_n N_Z_c_9131_n 0.0181262f $X=3.365 $Y=3.965 $X2=0
+ $Y2=0
cc_2179 N_A_559_793#_c_2175_n N_Z_c_9131_n 9.74366e-19 $X=3.835 $Y=3.965 $X2=0
+ $Y2=0
cc_2180 N_A_559_793#_c_2178_n N_Z_c_9131_n 0.00415268f $X=3.365 $Y=4.04 $X2=0
+ $Y2=0
cc_2181 N_A_559_793#_c_2173_n N_Z_c_9132_n 9.74366e-19 $X=3.365 $Y=3.965 $X2=0
+ $Y2=0
cc_2182 N_A_559_793#_c_2175_n N_Z_c_9132_n 0.0181262f $X=3.835 $Y=3.965 $X2=0
+ $Y2=0
cc_2183 N_A_559_793#_c_2176_n N_Z_c_9132_n 0.00560592f $X=4.215 $Y=4.04 $X2=0
+ $Y2=0
cc_2184 N_A_559_793#_c_2177_n N_Z_c_9132_n 0.0221748f $X=4.305 $Y=3.965 $X2=0
+ $Y2=0
cc_2185 N_A_559_793#_c_2179_n N_Z_c_9132_n 0.00181273f $X=3.835 $Y=4.04 $X2=0
+ $Y2=0
cc_2186 N_A_559_793#_c_2163_n N_Z_c_9132_n 0.00240108f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2187 N_A_559_793#_c_2169_n N_Z_c_9132_n 0.00425035f $X=4.625 $Y=4.21 $X2=0
+ $Y2=0
cc_2188 N_A_559_793#_c_2163_n N_VGND_c_12700_n 0.0123065f $X=5.42 $Y=4.21 $X2=0
+ $Y2=0
cc_2189 N_A_559_793#_c_2164_n N_VGND_c_12700_n 2.04129e-19 $X=4.875 $Y=4.21
+ $X2=0 $Y2=0
cc_2190 N_A_559_793#_c_2166_n N_VGND_c_12793_n 0.0129994f $X=5.585 $Y=4.995
+ $X2=0 $Y2=0
cc_2191 N_A_559_793#_M1017_d VGND 0.00394793f $X=5.45 $Y=4.785 $X2=0 $Y2=0
cc_2192 N_A_559_793#_c_2166_n VGND 0.00927134f $X=5.585 $Y=4.995 $X2=0 $Y2=0
cc_2193 N_A_559_793#_c_2178_n N_A_119_911#_c_14156_n 7.0477e-19 $X=3.365 $Y=4.04
+ $X2=0 $Y2=0
cc_2194 N_A_559_793#_c_2163_n N_A_119_911#_c_14137_n 0.0028695f $X=5.42 $Y=4.21
+ $X2=25.99 $Y2=4.8
cc_2195 N_A_559_793#_c_2169_n N_A_119_911#_c_14137_n 0.00589316f $X=4.625
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_2196 N_S[0]_c_2310_n N_S[8]_c_2427_n 0.0130744f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_2197 N_S[0]_c_2303_n N_S[8]_c_2429_n 0.0130744f $X=5.82 $Y=1.55 $X2=25.99
+ $Y2=4.8
cc_2198 N_S[0]_c_2303_n N_S[1]_c_2529_n 0.0215827f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2199 S[0] N_S[1]_c_2529_n 0.00113563f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_2200 N_S[0]_c_2303_n N_S[1]_c_2550_n 0.00113563f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2201 S[0] N_S[1]_c_2550_n 0.0301108f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_2202 N_S[0]_c_2310_n N_VPWR_c_7224_n 0.00950399f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_2203 N_S[0]_c_2303_n N_VPWR_c_7226_n 0.016386f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2204 S[0] N_VPWR_c_7226_n 0.0157609f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_2205 N_S[0]_c_2310_n N_VPWR_c_7313_n 0.0035837f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_2206 N_S[0]_c_2303_n N_VPWR_c_7313_n 0.0035837f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2207 N_S[0]_c_2310_n VPWR 0.00711603f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_2208 N_S[0]_c_2303_n VPWR 0.0070533f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2209 N_S[0]_c_2287_n N_A_117_297#_c_8771_n 0.00168571f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_2210 N_S[0]_c_2310_n N_A_117_297#_c_8775_n 0.00239129f $X=5.35 $Y=1.55 $X2=0
+ $Y2=0
cc_2211 N_S[0]_c_2287_n N_Z_c_9003_n 0.002324f $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_2212 N_S[0]_c_2290_n N_Z_c_9003_n 0.00283489f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_2213 N_S[0]_c_2290_n N_Z_c_9004_n 3.10191e-19 $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_2214 N_S[0]_c_2292_n N_Z_c_9004_n 0.00190704f $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_2215 N_S[0]_c_2290_n N_Z_c_9006_n 6.35774e-19 $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_2216 N_S[0]_c_2292_n N_Z_c_9006_n 0.0077801f $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_2217 N_S[0]_c_2294_n N_Z_c_9006_n 0.0134253f $X=4.08 $Y=0.255 $X2=0 $Y2=0
cc_2218 N_S[0]_c_2287_n N_Z_c_9043_n 0.00443615f $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_2219 N_S[0]_c_2290_n N_Z_c_9043_n 0.00462308f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_2220 N_S[0]_c_2292_n N_Z_c_9043_n 6.35664e-19 $X=3.66 $Y=0.255 $X2=0 $Y2=0
cc_2221 N_S[0]_c_2290_n N_Z_c_9046_n 0.00180363f $X=3.24 $Y=0.255 $X2=0 $Y2=0
cc_2222 N_S[0]_c_2294_n N_Z_c_9048_n 0.00216436f $X=4.08 $Y=0.255 $X2=0 $Y2=0
cc_2223 N_S[0]_c_2310_n N_Z_c_9115_n 0.00478771f $X=5.35 $Y=1.55 $X2=0 $Y2=0
cc_2224 N_S[0]_c_2303_n N_Z_c_9115_n 0.00760321f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2225 S[0] N_Z_c_9115_n 0.010609f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_2226 N_S[0]_c_2287_n N_VGND_c_12697_n 5.5039e-19 $X=2.82 $Y=0.255 $X2=0 $Y2=0
cc_2227 N_S[0]_c_2289_n N_VGND_c_12697_n 0.0028166f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_2228 N_S[0]_c_2295_n N_VGND_c_12699_n 0.00862298f $X=4.765 $Y=0.18 $X2=0
+ $Y2=0
cc_2229 N_S[0]_c_2297_n N_VGND_c_12699_n 0.00525833f $X=5.25 $Y=0.81 $X2=0 $Y2=0
cc_2230 N_S[0]_c_2300_n N_VGND_c_12699_n 0.00173127f $X=5.375 $Y=0.735 $X2=0
+ $Y2=0
cc_2231 N_S[0]_c_2302_n N_VGND_c_12701_n 0.00374526f $X=5.795 $Y=0.735 $X2=0
+ $Y2=0
cc_2232 N_S[0]_c_2303_n N_VGND_c_12701_n 0.00578076f $X=5.82 $Y=1.55 $X2=0 $Y2=0
cc_2233 S[0] N_VGND_c_12701_n 0.0116413f $X=6.125 $Y=1.105 $X2=0 $Y2=0
cc_2234 N_S[0]_c_2289_n N_VGND_c_12787_n 0.0559651f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_2235 N_S[0]_c_2300_n N_VGND_c_12791_n 0.00542362f $X=5.375 $Y=0.735 $X2=0
+ $Y2=0
cc_2236 N_S[0]_c_2301_n N_VGND_c_12791_n 2.16067e-19 $X=5.72 $Y=0.81 $X2=0 $Y2=0
cc_2237 N_S[0]_c_2302_n N_VGND_c_12791_n 0.00585385f $X=5.795 $Y=0.735 $X2=0
+ $Y2=0
cc_2238 N_S[0]_c_2288_n VGND 0.00642387f $X=3.165 $Y=0.18 $X2=0 $Y2=0
cc_2239 N_S[0]_c_2289_n VGND 0.00591981f $X=2.895 $Y=0.18 $X2=0 $Y2=0
cc_2240 N_S[0]_c_2291_n VGND 0.0064237f $X=3.585 $Y=0.18 $X2=0 $Y2=0
cc_2241 N_S[0]_c_2293_n VGND 0.00642387f $X=4.005 $Y=0.18 $X2=0 $Y2=0
cc_2242 N_S[0]_c_2295_n VGND 0.0345801f $X=4.765 $Y=0.18 $X2=0 $Y2=0
cc_2243 N_S[0]_c_2300_n VGND 0.00990284f $X=5.375 $Y=0.735 $X2=0 $Y2=0
cc_2244 N_S[0]_c_2302_n VGND 0.0119653f $X=5.795 $Y=0.735 $X2=0 $Y2=0
cc_2245 N_S[0]_c_2304_n VGND 0.00366655f $X=3.24 $Y=0.18 $X2=0 $Y2=0
cc_2246 N_S[0]_c_2305_n VGND 0.00366655f $X=3.66 $Y=0.18 $X2=0 $Y2=0
cc_2247 N_S[0]_c_2306_n VGND 0.00366655f $X=4.08 $Y=0.18 $X2=0 $Y2=0
cc_2248 N_S[0]_c_2287_n N_A_119_47#_c_14050_n 0.00206084f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_2249 N_S[0]_c_2287_n N_A_119_47#_c_14052_n 0.0139014f $X=2.82 $Y=0.255 $X2=0
+ $Y2=0
cc_2250 N_S[0]_c_2288_n N_A_119_47#_c_14052_n 0.00211351f $X=3.165 $Y=0.18 $X2=0
+ $Y2=0
cc_2251 N_S[0]_c_2290_n N_A_119_47#_c_14052_n 0.0106826f $X=3.24 $Y=0.255 $X2=0
+ $Y2=0
cc_2252 N_S[0]_c_2292_n N_A_119_47#_c_14054_n 0.0106844f $X=3.66 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_2253 N_S[0]_c_2293_n N_A_119_47#_c_14054_n 0.00211351f $X=4.005 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_2254 N_S[0]_c_2294_n N_A_119_47#_c_14054_n 0.0112916f $X=4.08 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_2255 N_S[0]_c_2295_n N_A_119_47#_c_14054_n 0.00685838f $X=4.765 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_2256 N_S[0]_c_2296_n N_A_119_47#_c_14054_n 0.00189496f $X=4.84 $Y=0.735
+ $X2=25.99 $Y2=4.8
cc_2257 N_S[0]_c_2296_n N_A_119_47#_c_14055_n 0.00529837f $X=4.84 $Y=0.735
+ $X2=25.99 $Y2=4.93
cc_2258 N_S[0]_c_2291_n N_A_119_47#_c_14090_n 0.0034777f $X=3.585 $Y=0.18 $X2=0
+ $Y2=0
cc_2259 N_S[8]_c_2419_n N_S[9]_c_2649_n 0.0215827f $X=5.795 $Y=4.705 $X2=0 $Y2=0
cc_2260 S[8] N_S[9]_c_2649_n 0.00113563f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_2261 N_S[8]_c_2419_n N_S[9]_c_2669_n 0.00113563f $X=5.795 $Y=4.705 $X2=0
+ $Y2=0
cc_2262 S[8] N_S[9]_c_2669_n 0.0301108f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_2263 N_S[8]_c_2427_n N_VPWR_c_7225_n 0.00950399f $X=5.35 $Y=3.89 $X2=0 $Y2=0
cc_2264 N_S[8]_c_2419_n N_VPWR_c_7227_n 0.00652399f $X=5.795 $Y=4.705 $X2=0
+ $Y2=0
cc_2265 N_S[8]_c_2429_n N_VPWR_c_7227_n 0.00986205f $X=5.82 $Y=3.89 $X2=0 $Y2=0
cc_2266 S[8] N_VPWR_c_7227_n 0.0157609f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_2267 N_S[8]_c_2427_n N_VPWR_c_7313_n 0.0035837f $X=5.35 $Y=3.89 $X2=0 $Y2=0
cc_2268 N_S[8]_c_2429_n N_VPWR_c_7313_n 0.0035837f $X=5.82 $Y=3.89 $X2=0 $Y2=0
cc_2269 N_S[8]_c_2427_n VPWR 0.00711603f $X=5.35 $Y=3.89 $X2=0 $Y2=0
cc_2270 N_S[8]_c_2429_n VPWR 0.0070533f $X=5.82 $Y=3.89 $X2=0 $Y2=0
cc_2271 N_S[8]_c_2404_n N_A_117_591#_c_8887_n 0.00168571f $X=2.82 $Y=5.185 $X2=0
+ $Y2=0
cc_2272 N_S[8]_c_2427_n N_A_117_591#_c_8891_n 0.00239129f $X=5.35 $Y=3.89 $X2=0
+ $Y2=0
cc_2273 N_S[8]_c_2407_n N_Z_c_9005_n 3.10191e-19 $X=3.24 $Y=5.185 $X2=0 $Y2=0
cc_2274 N_S[8]_c_2409_n N_Z_c_9005_n 0.00190704f $X=3.66 $Y=5.185 $X2=0 $Y2=0
cc_2275 N_S[8]_c_2407_n N_Z_c_9007_n 6.35774e-19 $X=3.24 $Y=5.185 $X2=0 $Y2=0
cc_2276 N_S[8]_c_2409_n N_Z_c_9007_n 0.0077801f $X=3.66 $Y=5.185 $X2=0 $Y2=0
cc_2277 N_S[8]_c_2411_n N_Z_c_9007_n 0.0134253f $X=4.08 $Y=5.185 $X2=0 $Y2=0
cc_2278 N_S[8]_c_2404_n N_Z_c_9044_n 0.00443615f $X=2.82 $Y=5.185 $X2=0 $Y2=0
cc_2279 N_S[8]_c_2407_n N_Z_c_9044_n 0.00462308f $X=3.24 $Y=5.185 $X2=0 $Y2=0
cc_2280 N_S[8]_c_2404_n N_Z_c_9045_n 0.002324f $X=2.82 $Y=5.185 $X2=0 $Y2=0
cc_2281 N_S[8]_c_2407_n N_Z_c_9045_n 0.00283489f $X=3.24 $Y=5.185 $X2=0 $Y2=0
cc_2282 N_S[8]_c_2409_n N_Z_c_9045_n 6.35664e-19 $X=3.66 $Y=5.185 $X2=0 $Y2=0
cc_2283 N_S[8]_c_2407_n N_Z_c_9047_n 0.00180363f $X=3.24 $Y=5.185 $X2=0 $Y2=0
cc_2284 N_S[8]_c_2411_n N_Z_c_9049_n 0.00216436f $X=4.08 $Y=5.185 $X2=0 $Y2=0
cc_2285 N_S[8]_c_2425_n N_Z_c_9116_n 2.55735e-19 $X=5.35 $Y=3.99 $X2=0 $Y2=0
cc_2286 N_S[8]_c_2427_n N_Z_c_9116_n 0.00453198f $X=5.35 $Y=3.89 $X2=0 $Y2=0
cc_2287 N_S[8]_c_2419_n N_Z_c_9116_n 0.00258545f $X=5.795 $Y=4.705 $X2=0 $Y2=0
cc_2288 N_S[8]_c_2429_n N_Z_c_9116_n 0.00501777f $X=5.82 $Y=3.89 $X2=0 $Y2=0
cc_2289 S[8] N_Z_c_9116_n 0.010609f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_2290 N_S[8]_c_2404_n N_VGND_c_12698_n 5.5039e-19 $X=2.82 $Y=5.185 $X2=0 $Y2=0
cc_2291 N_S[8]_c_2406_n N_VGND_c_12698_n 0.0028166f $X=2.895 $Y=5.26 $X2=0 $Y2=0
cc_2292 N_S[8]_c_2413_n N_VGND_c_12700_n 0.00862298f $X=4.84 $Y=5.185 $X2=0
+ $Y2=0
cc_2293 N_S[8]_c_2414_n N_VGND_c_12700_n 0.00525833f $X=5.25 $Y=4.63 $X2=0 $Y2=0
cc_2294 N_S[8]_c_2417_n N_VGND_c_12700_n 0.00173127f $X=5.375 $Y=4.705 $X2=0
+ $Y2=0
cc_2295 N_S[8]_c_2419_n N_VGND_c_12702_n 0.00952602f $X=5.795 $Y=4.705 $X2=0
+ $Y2=0
cc_2296 S[8] N_VGND_c_12702_n 0.0116413f $X=6.125 $Y=4.165 $X2=0 $Y2=0
cc_2297 N_S[8]_c_2406_n N_VGND_c_12789_n 0.0559651f $X=2.895 $Y=5.26 $X2=0 $Y2=0
cc_2298 N_S[8]_c_2417_n N_VGND_c_12793_n 0.00542362f $X=5.375 $Y=4.705 $X2=0
+ $Y2=0
cc_2299 N_S[8]_c_2418_n N_VGND_c_12793_n 2.16067e-19 $X=5.72 $Y=4.63 $X2=0 $Y2=0
cc_2300 N_S[8]_c_2419_n N_VGND_c_12793_n 0.00585385f $X=5.795 $Y=4.705 $X2=0
+ $Y2=0
cc_2301 N_S[8]_c_2405_n VGND 0.00642387f $X=3.165 $Y=5.26 $X2=0 $Y2=0
cc_2302 N_S[8]_c_2406_n VGND 0.00591981f $X=2.895 $Y=5.26 $X2=0 $Y2=0
cc_2303 N_S[8]_c_2408_n VGND 0.0064237f $X=3.585 $Y=5.26 $X2=0 $Y2=0
cc_2304 N_S[8]_c_2410_n VGND 0.00642387f $X=4.005 $Y=5.26 $X2=0 $Y2=0
cc_2305 N_S[8]_c_2412_n VGND 0.0345801f $X=4.765 $Y=5.26 $X2=0 $Y2=0
cc_2306 N_S[8]_c_2417_n VGND 0.00990284f $X=5.375 $Y=4.705 $X2=0 $Y2=0
cc_2307 N_S[8]_c_2419_n VGND 0.0119653f $X=5.795 $Y=4.705 $X2=0 $Y2=0
cc_2308 N_S[8]_c_2420_n VGND 0.00366655f $X=3.24 $Y=5.26 $X2=0 $Y2=0
cc_2309 N_S[8]_c_2421_n VGND 0.00366655f $X=3.66 $Y=5.26 $X2=0 $Y2=0
cc_2310 N_S[8]_c_2422_n VGND 0.00366655f $X=4.08 $Y=5.26 $X2=0 $Y2=0
cc_2311 N_S[8]_c_2404_n N_A_119_911#_c_14132_n 0.00206084f $X=2.82 $Y=5.185
+ $X2=0 $Y2=0
cc_2312 N_S[8]_c_2404_n N_A_119_911#_c_14134_n 0.0139014f $X=2.82 $Y=5.185 $X2=0
+ $Y2=0
cc_2313 N_S[8]_c_2405_n N_A_119_911#_c_14134_n 0.00211351f $X=3.165 $Y=5.26
+ $X2=0 $Y2=0
cc_2314 N_S[8]_c_2407_n N_A_119_911#_c_14134_n 0.0106826f $X=3.24 $Y=5.185 $X2=0
+ $Y2=0
cc_2315 N_S[8]_c_2409_n N_A_119_911#_c_14136_n 0.0106844f $X=3.66 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_2316 N_S[8]_c_2410_n N_A_119_911#_c_14136_n 0.00211351f $X=4.005 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_2317 N_S[8]_c_2411_n N_A_119_911#_c_14136_n 0.0112916f $X=4.08 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_2318 N_S[8]_c_2412_n N_A_119_911#_c_14136_n 0.00685838f $X=4.765 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_2319 N_S[8]_c_2413_n N_A_119_911#_c_14136_n 0.00189496f $X=4.84 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_2320 N_S[8]_c_2415_n N_A_119_911#_c_14137_n 0.00529837f $X=4.915 $Y=4.63
+ $X2=25.99 $Y2=4.8
cc_2321 N_S[8]_c_2408_n N_A_119_911#_c_14169_n 0.0034777f $X=3.585 $Y=5.26 $X2=0
+ $Y2=0
cc_2322 N_S[1]_c_2530_n N_S[9]_c_2671_n 0.0130744f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_2323 N_S[1]_c_2554_n N_S[9]_c_2675_n 0.0130744f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_2324 N_S[1]_c_2539_n N_A_1430_325#_c_2785_n 0.00507688f $X=8.8 $Y=0.255
+ $X2=25.905 $Y2=0.425
cc_2325 N_S[1]_c_2534_n N_A_1430_325#_c_2777_n 0.00262132f $X=7.53 $Y=1.45
+ $X2=25.905 $Y2=4.845
cc_2326 N_S[1]_c_2541_n N_A_1430_325#_c_2788_n 0.00509204f $X=9.22 $Y=0.255
+ $X2=0 $Y2=0
cc_2327 N_S[1]_c_2545_n N_A_1430_325#_c_2790_n 0.00507426f $X=10.06 $Y=0.255
+ $X2=0 $Y2=0
cc_2328 N_S[1]_c_2543_n N_A_1430_325#_c_2793_n 0.00509391f $X=9.64 $Y=0.255
+ $X2=0 $Y2=0
cc_2329 N_S[1]_c_2530_n N_A_1430_325#_c_2794_n 0.0128834f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_2330 N_S[1]_c_2554_n N_A_1430_325#_c_2794_n 0.0118698f $X=7.53 $Y=1.55 $X2=0
+ $Y2=0
cc_2331 N_S[1]_c_2531_n N_A_1430_325#_c_2778_n 0.00207203f $X=7.085 $Y=0.735
+ $X2=0 $Y2=0
cc_2332 N_S[1]_c_2533_n N_A_1430_325#_c_2778_n 0.00603996f $X=7.505 $Y=0.735
+ $X2=0 $Y2=0
cc_2333 N_S[1]_c_2536_n N_A_1430_325#_c_2778_n 6.53442e-19 $X=8.04 $Y=0.735
+ $X2=0 $Y2=0
cc_2334 N_S[1]_c_2530_n N_A_1430_325#_c_2779_n 0.00289358f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_2335 N_S[1]_c_2532_n N_A_1430_325#_c_2779_n 0.00429801f $X=7.43 $Y=0.81 $X2=0
+ $Y2=0
cc_2336 N_S[1]_c_2534_n N_A_1430_325#_c_2779_n 0.0085951f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_2337 N_S[1]_c_2546_n N_A_1430_325#_c_2779_n 0.00268644f $X=7.53 $Y=0.81 $X2=0
+ $Y2=0
cc_2338 N_S[1]_c_2550_n N_A_1430_325#_c_2779_n 0.00541767f $X=7.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2339 N_S[1]_c_2534_n N_A_1430_325#_c_2780_n 0.0206368f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_2340 N_S[1]_c_2535_n N_A_1430_325#_c_2780_n 0.0103812f $X=7.965 $Y=0.81 $X2=0
+ $Y2=0
cc_2341 N_S[1]_c_2530_n N_A_1430_325#_c_2796_n 0.00454075f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_2342 N_S[1]_c_2534_n N_A_1430_325#_c_2796_n 0.00255921f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_2343 N_S[1]_c_2554_n N_A_1430_325#_c_2796_n 0.00762115f $X=7.53 $Y=1.55 $X2=0
+ $Y2=0
cc_2344 N_S[1]_c_2532_n N_A_1430_325#_c_2781_n 0.0111895f $X=7.43 $Y=0.81 $X2=0
+ $Y2=0
cc_2345 N_S[1]_c_2533_n N_A_1430_325#_c_2781_n 9.67113e-19 $X=7.505 $Y=0.735
+ $X2=0 $Y2=0
cc_2346 N_S[1]_c_2546_n N_A_1430_325#_c_2781_n 0.00426435f $X=7.53 $Y=0.81 $X2=0
+ $Y2=0
cc_2347 N_S[1]_c_2530_n N_A_1430_325#_c_2782_n 0.00416423f $X=7.06 $Y=1.55 $X2=0
+ $Y2=0
cc_2348 N_S[1]_c_2534_n N_A_1430_325#_c_2782_n 0.00322131f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_2349 N_S[1]_c_2550_n N_A_1430_325#_c_2782_n 0.0228692f $X=7.02 $Y=1.16 $X2=0
+ $Y2=0
cc_2350 N_S[1]_c_2534_n N_A_1430_325#_c_2783_n 0.0175393f $X=7.53 $Y=1.45 $X2=0
+ $Y2=0
cc_2351 N_S[1]_c_2535_n N_A_1430_325#_c_2783_n 0.0179529f $X=7.965 $Y=0.81 $X2=0
+ $Y2=0
cc_2352 N_S[1]_c_2529_n N_VPWR_c_7229_n 0.00652399f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_2353 N_S[1]_c_2530_n N_VPWR_c_7229_n 0.00986205f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_2354 N_S[1]_c_2550_n N_VPWR_c_7229_n 0.0157609f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_2355 N_S[1]_c_2554_n N_VPWR_c_7231_n 0.00950399f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_2356 N_S[1]_c_2530_n N_VPWR_c_7316_n 0.0035837f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_2357 N_S[1]_c_2554_n N_VPWR_c_7316_n 0.0035837f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_2358 N_S[1]_c_2530_n VPWR 0.0070533f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_2359 N_S[1]_c_2554_n VPWR 0.00711603f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_2360 N_S[1]_c_2539_n N_Z_c_9008_n 0.0134253f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_2361 N_S[1]_c_2541_n N_Z_c_9008_n 0.0077801f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_2362 N_S[1]_c_2543_n N_Z_c_9008_n 6.35774e-19 $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_2363 N_S[1]_c_2541_n N_Z_c_9010_n 0.00190704f $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_2364 N_S[1]_c_2543_n N_Z_c_9010_n 3.10191e-19 $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_2365 N_S[1]_c_2543_n N_Z_c_9012_n 0.00283489f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_2366 N_S[1]_c_2545_n N_Z_c_9012_n 0.002324f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_2367 N_S[1]_c_2539_n N_Z_c_9050_n 0.00216436f $X=8.8 $Y=0.255 $X2=0 $Y2=0
cc_2368 N_S[1]_c_2543_n N_Z_c_9052_n 0.00180363f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_2369 N_S[1]_c_2541_n N_Z_c_9054_n 6.35664e-19 $X=9.22 $Y=0.255 $X2=0 $Y2=0
cc_2370 N_S[1]_c_2543_n N_Z_c_9054_n 0.00462308f $X=9.64 $Y=0.255 $X2=0 $Y2=0
cc_2371 N_S[1]_c_2545_n N_Z_c_9054_n 0.00443615f $X=10.06 $Y=0.255 $X2=0 $Y2=0
cc_2372 N_S[1]_c_2529_n N_Z_c_9115_n 0.00234109f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_2373 N_S[1]_c_2530_n N_Z_c_9115_n 0.0052507f $X=7.06 $Y=1.55 $X2=0 $Y2=0
cc_2374 N_S[1]_c_2554_n N_Z_c_9115_n 0.00478771f $X=7.53 $Y=1.55 $X2=0 $Y2=0
cc_2375 N_S[1]_c_2550_n N_Z_c_9115_n 0.0105931f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_2376 N_S[1]_c_2545_n N_A_1643_311#_c_10898_n 0.00168571f $X=10.06 $Y=0.255
+ $X2=0 $Y2=0
cc_2377 N_S[1]_c_2554_n N_A_1643_311#_c_10900_n 0.00239129f $X=7.53 $Y=1.55
+ $X2=0 $Y2=0
cc_2378 N_S[1]_c_2529_n N_VGND_c_12703_n 0.00576464f $X=6.96 $Y=1.16 $X2=0 $Y2=0
cc_2379 N_S[1]_c_2531_n N_VGND_c_12703_n 0.00374526f $X=7.085 $Y=0.735 $X2=0
+ $Y2=0
cc_2380 N_S[1]_c_2550_n N_VGND_c_12703_n 0.0116218f $X=7.02 $Y=1.16 $X2=0 $Y2=0
cc_2381 N_S[1]_c_2533_n N_VGND_c_12705_n 0.00173127f $X=7.505 $Y=0.735 $X2=0
+ $Y2=0
cc_2382 N_S[1]_c_2535_n N_VGND_c_12705_n 0.00525833f $X=7.965 $Y=0.81 $X2=0
+ $Y2=0
cc_2383 N_S[1]_c_2538_n N_VGND_c_12705_n 0.00862298f $X=8.115 $Y=0.18 $X2=0
+ $Y2=0
cc_2384 N_S[1]_c_2544_n N_VGND_c_12707_n 0.0028166f $X=9.985 $Y=0.18 $X2=0 $Y2=0
cc_2385 N_S[1]_c_2545_n N_VGND_c_12707_n 5.5039e-19 $X=10.06 $Y=0.255 $X2=0
+ $Y2=0
cc_2386 N_S[1]_c_2531_n N_VGND_c_12799_n 0.00585385f $X=7.085 $Y=0.735 $X2=0
+ $Y2=0
cc_2387 N_S[1]_c_2532_n N_VGND_c_12799_n 2.16067e-19 $X=7.43 $Y=0.81 $X2=0 $Y2=0
cc_2388 N_S[1]_c_2533_n N_VGND_c_12799_n 0.00542362f $X=7.505 $Y=0.735 $X2=0
+ $Y2=0
cc_2389 N_S[1]_c_2538_n N_VGND_c_12803_n 0.0559651f $X=8.115 $Y=0.18 $X2=0 $Y2=0
cc_2390 N_S[1]_c_2531_n VGND 0.0119653f $X=7.085 $Y=0.735 $X2=0 $Y2=0
cc_2391 N_S[1]_c_2533_n VGND 0.00990284f $X=7.505 $Y=0.735 $X2=0 $Y2=0
cc_2392 N_S[1]_c_2537_n VGND 0.0244174f $X=8.725 $Y=0.18 $X2=0 $Y2=0
cc_2393 N_S[1]_c_2538_n VGND 0.0101627f $X=8.115 $Y=0.18 $X2=0 $Y2=0
cc_2394 N_S[1]_c_2540_n VGND 0.00642387f $X=9.145 $Y=0.18 $X2=0 $Y2=0
cc_2395 N_S[1]_c_2542_n VGND 0.0064237f $X=9.565 $Y=0.18 $X2=0 $Y2=0
cc_2396 N_S[1]_c_2544_n VGND 0.0123437f $X=9.985 $Y=0.18 $X2=0 $Y2=0
cc_2397 N_S[1]_c_2547_n VGND 0.00366655f $X=8.8 $Y=0.18 $X2=0 $Y2=0
cc_2398 N_S[1]_c_2548_n VGND 0.00366655f $X=9.22 $Y=0.18 $X2=0 $Y2=0
cc_2399 N_S[1]_c_2549_n VGND 0.00366655f $X=9.64 $Y=0.18 $X2=0 $Y2=0
cc_2400 N_S[1]_c_2536_n N_A_1693_66#_c_14211_n 0.00529837f $X=8.04 $Y=0.735
+ $X2=0 $Y2=0
cc_2401 N_S[1]_c_2539_n N_A_1693_66#_c_14212_n 0.0112916f $X=8.8 $Y=0.255 $X2=0
+ $Y2=0
cc_2402 N_S[1]_c_2540_n N_A_1693_66#_c_14212_n 0.00211351f $X=9.145 $Y=0.18
+ $X2=0 $Y2=0
cc_2403 N_S[1]_c_2541_n N_A_1693_66#_c_14212_n 0.0106844f $X=9.22 $Y=0.255 $X2=0
+ $Y2=0
cc_2404 N_S[1]_c_2536_n N_A_1693_66#_c_14213_n 0.00189496f $X=8.04 $Y=0.735
+ $X2=0 $Y2=0
cc_2405 N_S[1]_c_2537_n N_A_1693_66#_c_14213_n 0.00685838f $X=8.725 $Y=0.18
+ $X2=0 $Y2=0
cc_2406 N_S[1]_c_2543_n N_A_1693_66#_c_14214_n 0.0106826f $X=9.64 $Y=0.255 $X2=0
+ $Y2=0
cc_2407 N_S[1]_c_2544_n N_A_1693_66#_c_14214_n 0.00211351f $X=9.985 $Y=0.18
+ $X2=0 $Y2=0
cc_2408 N_S[1]_c_2545_n N_A_1693_66#_c_14214_n 0.0139014f $X=10.06 $Y=0.255
+ $X2=0 $Y2=0
cc_2409 N_S[1]_c_2545_n N_A_1693_66#_c_14217_n 0.00206084f $X=10.06 $Y=0.255
+ $X2=0 $Y2=0
cc_2410 N_S[1]_c_2542_n N_A_1693_66#_c_14230_n 0.0034777f $X=9.565 $Y=0.18 $X2=0
+ $Y2=0
cc_2411 N_S[9]_c_2658_n N_A_1430_599#_c_2901_n 0.00507688f $X=8.8 $Y=5.185
+ $X2=25.905 $Y2=0.425
cc_2412 N_S[9]_c_2673_n N_A_1430_599#_c_2893_n 0.00262132f $X=7.53 $Y=3.99
+ $X2=25.905 $Y2=4.845
cc_2413 N_S[9]_c_2660_n N_A_1430_599#_c_2904_n 0.00509204f $X=9.22 $Y=5.185
+ $X2=0 $Y2=0
cc_2414 N_S[9]_c_2664_n N_A_1430_599#_c_2906_n 0.00507426f $X=10.06 $Y=5.185
+ $X2=0 $Y2=0
cc_2415 N_S[9]_c_2662_n N_A_1430_599#_c_2909_n 0.00509391f $X=9.64 $Y=5.185
+ $X2=0 $Y2=0
cc_2416 N_S[9]_c_2671_n N_A_1430_599#_c_2910_n 0.00929139f $X=7.06 $Y=3.89 $X2=0
+ $Y2=0
cc_2417 N_S[9]_c_2675_n N_A_1430_599#_c_2910_n 0.00970559f $X=7.53 $Y=3.89 $X2=0
+ $Y2=0
cc_2418 N_S[9]_c_2650_n N_A_1430_599#_c_2894_n 0.00207203f $X=7.085 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_2419 N_S[9]_c_2651_n N_A_1430_599#_c_2894_n 0.0111895f $X=7.43 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_2420 N_S[9]_c_2653_n N_A_1430_599#_c_2894_n 9.67113e-19 $X=7.505 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_2421 N_S[9]_c_2655_n N_A_1430_599#_c_2894_n 6.53442e-19 $X=8.04 $Y=5.185
+ $X2=25.99 $Y2=0.51
cc_2422 N_S[9]_c_2665_n N_A_1430_599#_c_2894_n 0.00426435f $X=7.53 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_2423 N_S[9]_c_2653_n N_A_1430_599#_c_2895_n 0.00603996f $X=7.505 $Y=4.705
+ $X2=0 $Y2=0
cc_2424 N_S[9]_c_2671_n N_A_1430_599#_c_2911_n 0.00117303f $X=7.06 $Y=3.89 $X2=0
+ $Y2=0
cc_2425 N_S[9]_c_2650_n N_A_1430_599#_c_2911_n 0.00336772f $X=7.085 $Y=4.705
+ $X2=0 $Y2=0
cc_2426 N_S[9]_c_2673_n N_A_1430_599#_c_2911_n 0.00508008f $X=7.53 $Y=3.99 $X2=0
+ $Y2=0
cc_2427 N_S[9]_c_2652_n N_A_1430_599#_c_2911_n 0.00255921f $X=7.53 $Y=4.555
+ $X2=0 $Y2=0
cc_2428 N_S[9]_c_2675_n N_A_1430_599#_c_2911_n 0.00254107f $X=7.53 $Y=3.89 $X2=0
+ $Y2=0
cc_2429 N_S[9]_c_2652_n N_A_1430_599#_c_2896_n 0.0206368f $X=7.53 $Y=4.555 $X2=0
+ $Y2=0
cc_2430 N_S[9]_c_2654_n N_A_1430_599#_c_2896_n 0.0103812f $X=7.965 $Y=4.63 $X2=0
+ $Y2=0
cc_2431 N_S[9]_c_2671_n N_A_1430_599#_c_2913_n 0.00304348f $X=7.06 $Y=3.89 $X2=0
+ $Y2=0
cc_2432 N_S[9]_c_2650_n N_A_1430_599#_c_2913_n 5.48523e-19 $X=7.085 $Y=4.705
+ $X2=0 $Y2=0
cc_2433 N_S[9]_c_2675_n N_A_1430_599#_c_2913_n 0.00216424f $X=7.53 $Y=3.89 $X2=0
+ $Y2=0
cc_2434 N_S[9]_c_2650_n N_A_1430_599#_c_2897_n 0.00289358f $X=7.085 $Y=4.705
+ $X2=0 $Y2=0
cc_2435 N_S[9]_c_2651_n N_A_1430_599#_c_2897_n 0.00429801f $X=7.43 $Y=4.63 $X2=0
+ $Y2=0
cc_2436 N_S[9]_c_2652_n N_A_1430_599#_c_2897_n 0.0085951f $X=7.53 $Y=4.555 $X2=0
+ $Y2=0
cc_2437 N_S[9]_c_2665_n N_A_1430_599#_c_2897_n 0.00268644f $X=7.53 $Y=4.63 $X2=0
+ $Y2=0
cc_2438 N_S[9]_c_2669_n N_A_1430_599#_c_2897_n 0.00541767f $X=7.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2439 N_S[9]_c_2650_n N_A_1430_599#_c_2898_n 0.00416423f $X=7.085 $Y=4.705
+ $X2=0 $Y2=0
cc_2440 N_S[9]_c_2652_n N_A_1430_599#_c_2898_n 0.00322131f $X=7.53 $Y=4.555
+ $X2=0 $Y2=0
cc_2441 N_S[9]_c_2669_n N_A_1430_599#_c_2898_n 0.0228692f $X=7.02 $Y=4.28 $X2=0
+ $Y2=0
cc_2442 N_S[9]_c_2652_n N_A_1430_599#_c_2899_n 0.0175393f $X=7.53 $Y=4.555 $X2=0
+ $Y2=0
cc_2443 N_S[9]_c_2654_n N_A_1430_599#_c_2899_n 0.0179529f $X=7.965 $Y=4.63 $X2=0
+ $Y2=0
cc_2444 N_S[9]_c_2649_n N_VPWR_c_7230_n 0.00652399f $X=6.96 $Y=4.28 $X2=0 $Y2=0
cc_2445 N_S[9]_c_2671_n N_VPWR_c_7230_n 0.00986205f $X=7.06 $Y=3.89 $X2=0 $Y2=0
cc_2446 N_S[9]_c_2669_n N_VPWR_c_7230_n 0.0157609f $X=7.02 $Y=4.28 $X2=0 $Y2=0
cc_2447 N_S[9]_c_2675_n N_VPWR_c_7232_n 0.00950399f $X=7.53 $Y=3.89 $X2=0 $Y2=0
cc_2448 N_S[9]_c_2671_n N_VPWR_c_7316_n 0.0035837f $X=7.06 $Y=3.89 $X2=0 $Y2=0
cc_2449 N_S[9]_c_2675_n N_VPWR_c_7316_n 0.0035837f $X=7.53 $Y=3.89 $X2=0 $Y2=0
cc_2450 N_S[9]_c_2671_n VPWR 0.0070533f $X=7.06 $Y=3.89 $X2=0 $Y2=0
cc_2451 N_S[9]_c_2675_n VPWR 0.00711603f $X=7.53 $Y=3.89 $X2=0 $Y2=0
cc_2452 N_S[9]_c_2658_n N_Z_c_9009_n 0.0134253f $X=8.8 $Y=5.185 $X2=0 $Y2=0
cc_2453 N_S[9]_c_2660_n N_Z_c_9009_n 0.0077801f $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_2454 N_S[9]_c_2662_n N_Z_c_9009_n 6.35774e-19 $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_2455 N_S[9]_c_2660_n N_Z_c_9011_n 0.00190704f $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_2456 N_S[9]_c_2662_n N_Z_c_9011_n 3.10191e-19 $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_2457 N_S[9]_c_2658_n N_Z_c_9051_n 0.00216436f $X=8.8 $Y=5.185 $X2=0 $Y2=0
cc_2458 N_S[9]_c_2662_n N_Z_c_9053_n 0.00180363f $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_2459 N_S[9]_c_2662_n N_Z_c_9055_n 0.00462308f $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_2460 N_S[9]_c_2664_n N_Z_c_9055_n 0.00443615f $X=10.06 $Y=5.185 $X2=0 $Y2=0
cc_2461 N_S[9]_c_2660_n N_Z_c_9056_n 6.35664e-19 $X=9.22 $Y=5.185 $X2=0 $Y2=0
cc_2462 N_S[9]_c_2662_n N_Z_c_9056_n 0.00283489f $X=9.64 $Y=5.185 $X2=0 $Y2=0
cc_2463 N_S[9]_c_2664_n N_Z_c_9056_n 0.002324f $X=10.06 $Y=5.185 $X2=0 $Y2=0
cc_2464 N_S[9]_c_2649_n N_Z_c_9116_n 0.00234109f $X=6.96 $Y=4.28 $X2=0 $Y2=0
cc_2465 N_S[9]_c_2671_n N_Z_c_9116_n 0.00501777f $X=7.06 $Y=3.89 $X2=0 $Y2=0
cc_2466 N_S[9]_c_2650_n N_Z_c_9116_n 2.32936e-19 $X=7.085 $Y=4.705 $X2=0 $Y2=0
cc_2467 N_S[9]_c_2673_n N_Z_c_9116_n 2.55735e-19 $X=7.53 $Y=3.99 $X2=0 $Y2=0
cc_2468 N_S[9]_c_2675_n N_Z_c_9116_n 0.00453198f $X=7.53 $Y=3.89 $X2=0 $Y2=0
cc_2469 N_S[9]_c_2669_n N_Z_c_9116_n 0.0105931f $X=7.02 $Y=4.28 $X2=0 $Y2=0
cc_2470 N_S[9]_c_2664_n N_A_1643_613#_c_11029_n 0.00168571f $X=10.06 $Y=5.185
+ $X2=0 $Y2=0
cc_2471 N_S[9]_c_2675_n N_A_1643_613#_c_11031_n 0.00239129f $X=7.53 $Y=3.89
+ $X2=0 $Y2=0
cc_2472 N_S[9]_c_2649_n N_VGND_c_12704_n 0.00576464f $X=6.96 $Y=4.28 $X2=0 $Y2=0
cc_2473 N_S[9]_c_2650_n N_VGND_c_12704_n 0.00374526f $X=7.085 $Y=4.705 $X2=0
+ $Y2=0
cc_2474 N_S[9]_c_2669_n N_VGND_c_12704_n 0.0116218f $X=7.02 $Y=4.28 $X2=0 $Y2=0
cc_2475 N_S[9]_c_2653_n N_VGND_c_12706_n 0.00173127f $X=7.505 $Y=4.705 $X2=0
+ $Y2=0
cc_2476 N_S[9]_c_2654_n N_VGND_c_12706_n 0.00525833f $X=7.965 $Y=4.63 $X2=0
+ $Y2=0
cc_2477 N_S[9]_c_2655_n N_VGND_c_12706_n 0.00862298f $X=8.04 $Y=5.185 $X2=0
+ $Y2=0
cc_2478 N_S[9]_c_2663_n N_VGND_c_12708_n 0.0028166f $X=9.985 $Y=5.26 $X2=0 $Y2=0
cc_2479 N_S[9]_c_2664_n N_VGND_c_12708_n 5.5039e-19 $X=10.06 $Y=5.185 $X2=0
+ $Y2=0
cc_2480 N_S[9]_c_2650_n N_VGND_c_12801_n 0.00585385f $X=7.085 $Y=4.705 $X2=0
+ $Y2=0
cc_2481 N_S[9]_c_2651_n N_VGND_c_12801_n 2.16067e-19 $X=7.43 $Y=4.63 $X2=0 $Y2=0
cc_2482 N_S[9]_c_2653_n N_VGND_c_12801_n 0.00542362f $X=7.505 $Y=4.705 $X2=0
+ $Y2=0
cc_2483 N_S[9]_c_2657_n N_VGND_c_12805_n 0.0559651f $X=8.115 $Y=5.26 $X2=0 $Y2=0
cc_2484 N_S[9]_c_2650_n VGND 0.0119653f $X=7.085 $Y=4.705 $X2=0 $Y2=0
cc_2485 N_S[9]_c_2653_n VGND 0.00990284f $X=7.505 $Y=4.705 $X2=0 $Y2=0
cc_2486 N_S[9]_c_2656_n VGND 0.0244174f $X=8.725 $Y=5.26 $X2=0 $Y2=0
cc_2487 N_S[9]_c_2657_n VGND 0.0101627f $X=8.115 $Y=5.26 $X2=0 $Y2=0
cc_2488 N_S[9]_c_2659_n VGND 0.00642387f $X=9.145 $Y=5.26 $X2=0 $Y2=0
cc_2489 N_S[9]_c_2661_n VGND 0.0064237f $X=9.565 $Y=5.26 $X2=0 $Y2=0
cc_2490 N_S[9]_c_2663_n VGND 0.0123437f $X=9.985 $Y=5.26 $X2=0 $Y2=0
cc_2491 N_S[9]_c_2666_n VGND 0.00366655f $X=8.8 $Y=5.26 $X2=0 $Y2=0
cc_2492 N_S[9]_c_2667_n VGND 0.00366655f $X=9.22 $Y=5.26 $X2=0 $Y2=0
cc_2493 N_S[9]_c_2668_n VGND 0.00366655f $X=9.64 $Y=5.26 $X2=0 $Y2=0
cc_2494 N_S[9]_c_2654_n N_A_1693_918#_c_14295_n 0.00529837f $X=7.965 $Y=4.63
+ $X2=0 $Y2=0
cc_2495 N_S[9]_c_2658_n N_A_1693_918#_c_14296_n 0.0112916f $X=8.8 $Y=5.185 $X2=0
+ $Y2=0
cc_2496 N_S[9]_c_2659_n N_A_1693_918#_c_14296_n 0.00211351f $X=9.145 $Y=5.26
+ $X2=0 $Y2=0
cc_2497 N_S[9]_c_2660_n N_A_1693_918#_c_14296_n 0.0106844f $X=9.22 $Y=5.185
+ $X2=0 $Y2=0
cc_2498 N_S[9]_c_2655_n N_A_1693_918#_c_14297_n 0.00189496f $X=8.04 $Y=5.185
+ $X2=0 $Y2=0
cc_2499 N_S[9]_c_2656_n N_A_1693_918#_c_14297_n 0.00685838f $X=8.725 $Y=5.26
+ $X2=0 $Y2=0
cc_2500 N_S[9]_c_2662_n N_A_1693_918#_c_14298_n 0.0106826f $X=9.64 $Y=5.185
+ $X2=0 $Y2=0
cc_2501 N_S[9]_c_2663_n N_A_1693_918#_c_14298_n 0.00211351f $X=9.985 $Y=5.26
+ $X2=0 $Y2=0
cc_2502 N_S[9]_c_2664_n N_A_1693_918#_c_14298_n 0.0139014f $X=10.06 $Y=5.185
+ $X2=0 $Y2=0
cc_2503 N_S[9]_c_2664_n N_A_1693_918#_c_14301_n 0.00206084f $X=10.06 $Y=5.185
+ $X2=0 $Y2=0
cc_2504 N_S[9]_c_2661_n N_A_1693_918#_c_14314_n 0.0034777f $X=9.565 $Y=5.26
+ $X2=0 $Y2=0
cc_2505 N_A_1430_325#_c_2784_n N_A_1430_599#_c_2900_n 0.0129371f $X=8.575
+ $Y=1.475 $X2=0 $Y2=0
cc_2506 N_A_1430_325#_c_2787_n N_A_1430_599#_c_2903_n 0.0129371f $X=9.045
+ $Y=1.475 $X2=0 $Y2=0
cc_2507 N_A_1430_325#_c_2789_n N_A_1430_599#_c_2905_n 0.0129371f $X=9.515
+ $Y=1.475 $X2=0 $Y2=0
cc_2508 N_A_1430_325#_c_2791_n N_A_1430_599#_c_2907_n 0.0129371f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_2509 N_A_1430_325#_c_2794_n N_VPWR_c_7229_n 0.0356181f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_2510 N_A_1430_325#_c_2784_n N_VPWR_c_7231_n 0.00367058f $X=8.575 $Y=1.475
+ $X2=0 $Y2=0
cc_2511 N_A_1430_325#_c_2794_n N_VPWR_c_7231_n 0.0316788f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_2512 N_A_1430_325#_c_2780_n N_VPWR_c_7231_n 0.0193185f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_2513 N_A_1430_325#_c_2783_n N_VPWR_c_7231_n 6.4101e-19 $X=8.255 $Y=1.23 $X2=0
+ $Y2=0
cc_2514 N_A_1430_325#_c_2791_n N_VPWR_c_7233_n 0.00324472f $X=9.985 $Y=1.475
+ $X2=0 $Y2=0
cc_2515 N_A_1430_325#_c_2794_n N_VPWR_c_7316_n 0.0233824f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_2516 N_A_1430_325#_c_2784_n VPWR 0.00473731f $X=8.575 $Y=1.475 $X2=0 $Y2=0
cc_2517 N_A_1430_325#_c_2787_n VPWR 0.00362156f $X=9.045 $Y=1.475 $X2=0 $Y2=0
cc_2518 N_A_1430_325#_c_2789_n VPWR 0.00362156f $X=9.515 $Y=1.475 $X2=0 $Y2=0
cc_2519 N_A_1430_325#_c_2791_n VPWR 0.00473731f $X=9.985 $Y=1.475 $X2=0 $Y2=0
cc_2520 N_A_1430_325#_c_2794_n VPWR 0.00593513f $X=7.295 $Y=1.77 $X2=0 $Y2=0
cc_2521 N_A_1430_325#_c_2788_n N_Z_c_9010_n 0.00762343f $X=9.425 $Y=1.4 $X2=0
+ $Y2=0
cc_2522 N_A_1430_325#_c_2793_n N_Z_c_9010_n 0.00704092f $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_2523 N_A_1430_325#_c_2785_n N_Z_c_9050_n 0.00597584f $X=8.955 $Y=1.4 $X2=0
+ $Y2=0
cc_2524 N_A_1430_325#_c_2777_n N_Z_c_9050_n 0.00747617f $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_2525 N_A_1430_325#_c_2788_n N_Z_c_9050_n 0.00145542f $X=9.425 $Y=1.4 $X2=0
+ $Y2=0
cc_2526 N_A_1430_325#_c_2792_n N_Z_c_9050_n 0.00909323f $X=9.045 $Y=1.4 $X2=0
+ $Y2=0
cc_2527 N_A_1430_325#_c_2780_n N_Z_c_9050_n 0.0266078f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_2528 N_A_1430_325#_c_2790_n N_Z_c_9052_n 0.00918337f $X=9.895 $Y=1.4 $X2=0
+ $Y2=0
cc_2529 N_A_1430_325#_c_2793_n N_Z_c_9052_n 2.98555e-19 $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_2530 N_A_1430_325#_c_2790_n N_Z_c_9054_n 0.00248496f $X=9.895 $Y=1.4 $X2=0
+ $Y2=0
cc_2531 N_A_1430_325#_c_2784_n N_Z_c_9115_n 0.00795576f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_2532 N_A_1430_325#_c_2777_n N_Z_c_9115_n 2.19754e-19 $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_2533 N_A_1430_325#_c_2794_n N_Z_c_9115_n 0.0329704f $X=7.295 $Y=1.77 $X2=0
+ $Y2=0
cc_2534 N_A_1430_325#_c_2780_n N_Z_c_9115_n 0.0186685f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_2535 N_A_1430_325#_c_2791_n N_Z_c_9117_n 0.00834829f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_2536 N_A_1430_325#_c_2787_n N_Z_c_9288_n 0.00372248f $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_2537 N_A_1430_325#_c_2789_n N_Z_c_9288_n 0.00372458f $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_2538 N_A_1430_325#_c_2784_n N_Z_c_9133_n 0.0221748f $X=8.575 $Y=1.475 $X2=0
+ $Y2=0
cc_2539 N_A_1430_325#_c_2785_n N_Z_c_9133_n 0.00560592f $X=8.955 $Y=1.4 $X2=0
+ $Y2=0
cc_2540 N_A_1430_325#_c_2777_n N_Z_c_9133_n 0.00425035f $X=8.665 $Y=1.4 $X2=0
+ $Y2=0
cc_2541 N_A_1430_325#_c_2787_n N_Z_c_9133_n 0.0181262f $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_2542 N_A_1430_325#_c_2789_n N_Z_c_9133_n 9.74366e-19 $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_2543 N_A_1430_325#_c_2792_n N_Z_c_9133_n 0.00181273f $X=9.045 $Y=1.4 $X2=0
+ $Y2=0
cc_2544 N_A_1430_325#_c_2780_n N_Z_c_9133_n 0.00240108f $X=8.345 $Y=1.23 $X2=0
+ $Y2=0
cc_2545 N_A_1430_325#_c_2787_n N_Z_c_9134_n 9.74366e-19 $X=9.045 $Y=1.475 $X2=0
+ $Y2=0
cc_2546 N_A_1430_325#_c_2789_n N_Z_c_9134_n 0.0181262f $X=9.515 $Y=1.475 $X2=0
+ $Y2=0
cc_2547 N_A_1430_325#_c_2790_n N_Z_c_9134_n 0.0103509f $X=9.895 $Y=1.4 $X2=0
+ $Y2=0
cc_2548 N_A_1430_325#_c_2791_n N_Z_c_9134_n 0.0199111f $X=9.985 $Y=1.475 $X2=0
+ $Y2=0
cc_2549 N_A_1430_325#_c_2793_n N_Z_c_9134_n 0.00415268f $X=9.515 $Y=1.4 $X2=0
+ $Y2=0
cc_2550 N_A_1430_325#_c_2791_n N_A_1643_311#_c_10898_n 0.00151141f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_2551 N_A_1430_325#_c_2784_n N_A_1643_311#_c_10906_n 0.00307958f $X=8.575
+ $Y=1.475 $X2=0 $Y2=0
cc_2552 N_A_1430_325#_c_2787_n N_A_1643_311#_c_10906_n 0.00307958f $X=9.045
+ $Y=1.475 $X2=0 $Y2=0
cc_2553 N_A_1430_325#_c_2789_n N_A_1643_311#_c_10908_n 0.00307958f $X=9.515
+ $Y=1.475 $X2=0 $Y2=0
cc_2554 N_A_1430_325#_c_2791_n N_A_1643_311#_c_10908_n 0.00307958f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_2555 N_A_1430_325#_c_2784_n N_A_1643_311#_c_10900_n 0.00499839f $X=8.575
+ $Y=1.475 $X2=0 $Y2=0
cc_2556 N_A_1430_325#_c_2777_n N_A_1643_311#_c_10900_n 0.00561627f $X=8.665
+ $Y=1.4 $X2=0 $Y2=0
cc_2557 N_A_1430_325#_c_2780_n N_A_1643_311#_c_10900_n 0.0218124f $X=8.345
+ $Y=1.23 $X2=0 $Y2=0
cc_2558 N_A_1430_325#_c_2783_n N_A_1643_311#_c_10900_n 5.74251e-19 $X=8.255
+ $Y=1.23 $X2=0 $Y2=0
cc_2559 N_A_1430_325#_c_2787_n N_A_1643_311#_c_10901_n 0.00210632f $X=9.045
+ $Y=1.475 $X2=0 $Y2=0
cc_2560 N_A_1430_325#_c_2788_n N_A_1643_311#_c_10901_n 0.00251792f $X=9.425
+ $Y=1.4 $X2=0 $Y2=0
cc_2561 N_A_1430_325#_c_2789_n N_A_1643_311#_c_10901_n 0.00210632f $X=9.515
+ $Y=1.475 $X2=0 $Y2=0
cc_2562 N_A_1430_325#_c_2791_n N_A_1643_311#_c_10902_n 0.00554566f $X=9.985
+ $Y=1.475 $X2=0 $Y2=0
cc_2563 N_A_1430_325#_c_2780_n N_VGND_c_12705_n 0.0123065f $X=8.345 $Y=1.23
+ $X2=0 $Y2=0
cc_2564 N_A_1430_325#_c_2783_n N_VGND_c_12705_n 2.04129e-19 $X=8.255 $Y=1.23
+ $X2=0 $Y2=0
cc_2565 N_A_1430_325#_c_2778_n N_VGND_c_12799_n 0.0129994f $X=7.295 $Y=0.445
+ $X2=0 $Y2=0
cc_2566 N_A_1430_325#_M1241_s VGND 0.00394793f $X=7.16 $Y=0.235 $X2=0 $Y2=0
cc_2567 N_A_1430_325#_c_2778_n VGND 0.00927134f $X=7.295 $Y=0.445 $X2=0 $Y2=0
cc_2568 N_A_1430_325#_c_2777_n N_A_1693_66#_c_14211_n 0.00600378f $X=8.665
+ $Y=1.4 $X2=0 $Y2=0
cc_2569 N_A_1430_325#_c_2780_n N_A_1693_66#_c_14211_n 0.0028695f $X=8.345
+ $Y=1.23 $X2=0 $Y2=0
cc_2570 N_A_1430_325#_c_2788_n N_A_1693_66#_c_14233_n 7.0477e-19 $X=9.425 $Y=1.4
+ $X2=0 $Y2=0
cc_2571 N_A_1430_599#_c_2910_n N_VPWR_c_7230_n 0.0356181f $X=7.295 $Y=3.14 $X2=0
+ $Y2=0
cc_2572 N_A_1430_599#_c_2900_n N_VPWR_c_7232_n 0.00367058f $X=8.575 $Y=3.965
+ $X2=0 $Y2=0
cc_2573 N_A_1430_599#_c_2910_n N_VPWR_c_7232_n 0.0316788f $X=7.295 $Y=3.14 $X2=0
+ $Y2=0
cc_2574 N_A_1430_599#_c_2896_n N_VPWR_c_7232_n 0.0193185f $X=8.345 $Y=4.21 $X2=0
+ $Y2=0
cc_2575 N_A_1430_599#_c_2899_n N_VPWR_c_7232_n 6.4101e-19 $X=8.255 $Y=4.21 $X2=0
+ $Y2=0
cc_2576 N_A_1430_599#_c_2907_n N_VPWR_c_7234_n 0.00324472f $X=9.985 $Y=3.965
+ $X2=0 $Y2=0
cc_2577 N_A_1430_599#_c_2910_n N_VPWR_c_7316_n 0.0233824f $X=7.295 $Y=3.14 $X2=0
+ $Y2=0
cc_2578 N_A_1430_599#_c_2900_n VPWR 0.00473731f $X=8.575 $Y=3.965 $X2=0 $Y2=0
cc_2579 N_A_1430_599#_c_2903_n VPWR 0.00362156f $X=9.045 $Y=3.965 $X2=0 $Y2=0
cc_2580 N_A_1430_599#_c_2905_n VPWR 0.00362156f $X=9.515 $Y=3.965 $X2=0 $Y2=0
cc_2581 N_A_1430_599#_c_2907_n VPWR 0.00473731f $X=9.985 $Y=3.965 $X2=0 $Y2=0
cc_2582 N_A_1430_599#_c_2910_n VPWR 0.00593513f $X=7.295 $Y=3.14 $X2=0 $Y2=0
cc_2583 N_A_1430_599#_c_2904_n N_Z_c_9011_n 0.00762343f $X=9.425 $Y=4.04 $X2=0
+ $Y2=0
cc_2584 N_A_1430_599#_c_2909_n N_Z_c_9011_n 0.00704092f $X=9.515 $Y=4.04 $X2=0
+ $Y2=0
cc_2585 N_A_1430_599#_c_2901_n N_Z_c_9051_n 0.00597584f $X=8.955 $Y=4.04 $X2=0
+ $Y2=0
cc_2586 N_A_1430_599#_c_2893_n N_Z_c_9051_n 0.00747617f $X=8.665 $Y=4.04 $X2=0
+ $Y2=0
cc_2587 N_A_1430_599#_c_2904_n N_Z_c_9051_n 0.00145542f $X=9.425 $Y=4.04 $X2=0
+ $Y2=0
cc_2588 N_A_1430_599#_c_2908_n N_Z_c_9051_n 0.00909323f $X=9.045 $Y=4.04 $X2=0
+ $Y2=0
cc_2589 N_A_1430_599#_c_2896_n N_Z_c_9051_n 0.0266078f $X=8.345 $Y=4.21 $X2=0
+ $Y2=0
cc_2590 N_A_1430_599#_c_2906_n N_Z_c_9053_n 0.00918337f $X=9.895 $Y=4.04 $X2=0
+ $Y2=0
cc_2591 N_A_1430_599#_c_2909_n N_Z_c_9053_n 2.98555e-19 $X=9.515 $Y=4.04 $X2=0
+ $Y2=0
cc_2592 N_A_1430_599#_c_2906_n N_Z_c_9055_n 0.00248496f $X=9.895 $Y=4.04 $X2=0
+ $Y2=0
cc_2593 N_A_1430_599#_c_2900_n N_Z_c_9116_n 0.00795576f $X=8.575 $Y=3.965 $X2=0
+ $Y2=0
cc_2594 N_A_1430_599#_c_2893_n N_Z_c_9116_n 2.19754e-19 $X=8.665 $Y=4.04 $X2=0
+ $Y2=0
cc_2595 N_A_1430_599#_c_2910_n N_Z_c_9116_n 0.0329704f $X=7.295 $Y=3.14 $X2=0
+ $Y2=0
cc_2596 N_A_1430_599#_c_2896_n N_Z_c_9116_n 0.0186685f $X=8.345 $Y=4.21 $X2=0
+ $Y2=0
cc_2597 N_A_1430_599#_c_2907_n N_Z_c_9118_n 0.00834829f $X=9.985 $Y=3.965 $X2=0
+ $Y2=0
cc_2598 N_A_1430_599#_c_2903_n N_Z_c_9317_n 0.00372248f $X=9.045 $Y=3.965 $X2=0
+ $Y2=0
cc_2599 N_A_1430_599#_c_2905_n N_Z_c_9317_n 0.00372458f $X=9.515 $Y=3.965 $X2=0
+ $Y2=0
cc_2600 N_A_1430_599#_c_2900_n N_Z_c_9133_n 0.0221748f $X=8.575 $Y=3.965 $X2=0
+ $Y2=0
cc_2601 N_A_1430_599#_c_2901_n N_Z_c_9133_n 0.00560592f $X=8.955 $Y=4.04 $X2=0
+ $Y2=0
cc_2602 N_A_1430_599#_c_2893_n N_Z_c_9133_n 0.00425035f $X=8.665 $Y=4.04 $X2=0
+ $Y2=0
cc_2603 N_A_1430_599#_c_2903_n N_Z_c_9133_n 0.0181262f $X=9.045 $Y=3.965 $X2=0
+ $Y2=0
cc_2604 N_A_1430_599#_c_2905_n N_Z_c_9133_n 9.74366e-19 $X=9.515 $Y=3.965 $X2=0
+ $Y2=0
cc_2605 N_A_1430_599#_c_2908_n N_Z_c_9133_n 0.00181273f $X=9.045 $Y=4.04 $X2=0
+ $Y2=0
cc_2606 N_A_1430_599#_c_2896_n N_Z_c_9133_n 0.00240108f $X=8.345 $Y=4.21 $X2=0
+ $Y2=0
cc_2607 N_A_1430_599#_c_2903_n N_Z_c_9134_n 9.74366e-19 $X=9.045 $Y=3.965 $X2=0
+ $Y2=0
cc_2608 N_A_1430_599#_c_2905_n N_Z_c_9134_n 0.0181262f $X=9.515 $Y=3.965 $X2=0
+ $Y2=0
cc_2609 N_A_1430_599#_c_2906_n N_Z_c_9134_n 0.0103509f $X=9.895 $Y=4.04 $X2=0
+ $Y2=0
cc_2610 N_A_1430_599#_c_2907_n N_Z_c_9134_n 0.0199111f $X=9.985 $Y=3.965 $X2=0
+ $Y2=0
cc_2611 N_A_1430_599#_c_2909_n N_Z_c_9134_n 0.00415268f $X=9.515 $Y=4.04 $X2=0
+ $Y2=0
cc_2612 N_A_1430_599#_c_2907_n N_A_1643_613#_c_11029_n 0.00151141f $X=9.985
+ $Y=3.965 $X2=0 $Y2=0
cc_2613 N_A_1430_599#_c_2900_n N_A_1643_613#_c_11037_n 0.00307958f $X=8.575
+ $Y=3.965 $X2=0 $Y2=0
cc_2614 N_A_1430_599#_c_2903_n N_A_1643_613#_c_11037_n 0.00307958f $X=9.045
+ $Y=3.965 $X2=0 $Y2=0
cc_2615 N_A_1430_599#_c_2905_n N_A_1643_613#_c_11039_n 0.00307958f $X=9.515
+ $Y=3.965 $X2=0 $Y2=0
cc_2616 N_A_1430_599#_c_2907_n N_A_1643_613#_c_11039_n 0.00307958f $X=9.985
+ $Y=3.965 $X2=0 $Y2=0
cc_2617 N_A_1430_599#_c_2900_n N_A_1643_613#_c_11031_n 0.00499839f $X=8.575
+ $Y=3.965 $X2=0 $Y2=0
cc_2618 N_A_1430_599#_c_2893_n N_A_1643_613#_c_11031_n 0.00561627f $X=8.665
+ $Y=4.04 $X2=0 $Y2=0
cc_2619 N_A_1430_599#_c_2896_n N_A_1643_613#_c_11031_n 0.0218124f $X=8.345
+ $Y=4.21 $X2=0 $Y2=0
cc_2620 N_A_1430_599#_c_2899_n N_A_1643_613#_c_11031_n 5.74251e-19 $X=8.255
+ $Y=4.21 $X2=0 $Y2=0
cc_2621 N_A_1430_599#_c_2903_n N_A_1643_613#_c_11032_n 0.00210632f $X=9.045
+ $Y=3.965 $X2=0 $Y2=0
cc_2622 N_A_1430_599#_c_2904_n N_A_1643_613#_c_11032_n 0.00251792f $X=9.425
+ $Y=4.04 $X2=0 $Y2=0
cc_2623 N_A_1430_599#_c_2905_n N_A_1643_613#_c_11032_n 0.00210632f $X=9.515
+ $Y=3.965 $X2=0 $Y2=0
cc_2624 N_A_1430_599#_c_2907_n N_A_1643_613#_c_11033_n 0.00554566f $X=9.985
+ $Y=3.965 $X2=0 $Y2=0
cc_2625 N_A_1430_599#_c_2896_n N_VGND_c_12706_n 0.0123065f $X=8.345 $Y=4.21
+ $X2=0 $Y2=0
cc_2626 N_A_1430_599#_c_2899_n N_VGND_c_12706_n 2.04129e-19 $X=8.255 $Y=4.21
+ $X2=0 $Y2=0
cc_2627 N_A_1430_599#_c_2895_n N_VGND_c_12801_n 0.0129994f $X=7.295 $Y=4.995
+ $X2=0 $Y2=0
cc_2628 N_A_1430_599#_M1008_d VGND 0.00394793f $X=7.16 $Y=4.785 $X2=0 $Y2=0
cc_2629 N_A_1430_599#_c_2895_n VGND 0.00927134f $X=7.295 $Y=4.995 $X2=0 $Y2=0
cc_2630 N_A_1430_599#_c_2893_n N_A_1693_918#_c_14295_n 0.00600378f $X=8.665
+ $Y=4.04 $X2=0 $Y2=0
cc_2631 N_A_1430_599#_c_2896_n N_A_1693_918#_c_14295_n 0.0028695f $X=8.345
+ $Y=4.21 $X2=0 $Y2=0
cc_2632 N_A_1430_599#_c_2904_n N_A_1693_918#_c_14317_n 7.0477e-19 $X=9.425
+ $Y=4.04 $X2=0 $Y2=0
cc_2633 N_D[1]_M1002_g N_D[9]_M1011_g 0.0130744f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_2634 N_D[1]_M1038_g N_D[9]_M1051_g 0.0130744f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_2635 N_D[1]_M1134_g N_D[9]_M1148_g 0.0130744f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_2636 N_D[1]_M1271_g N_D[9]_M1285_g 0.0130744f $X=12.385 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_2637 N_D[1]_M1002_g N_VPWR_c_7233_n 0.00389633f $X=10.975 $Y=1.985 $X2=0
+ $Y2=0
cc_2638 N_D[1]_M1038_g N_VPWR_c_7235_n 0.00208662f $X=11.445 $Y=1.985 $X2=0
+ $Y2=0
cc_2639 N_D[1]_M1134_g N_VPWR_c_7235_n 0.00208662f $X=11.915 $Y=1.985 $X2=0
+ $Y2=0
cc_2640 N_D[1]_M1271_g N_VPWR_c_7237_n 0.00374733f $X=12.385 $Y=1.985 $X2=0
+ $Y2=0
cc_2641 N_D[1]_M1002_g VPWR 0.00573859f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_2642 N_D[1]_M1038_g VPWR 0.00445624f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_2643 N_D[1]_M1134_g VPWR 0.00445624f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_2644 N_D[1]_M1271_g VPWR 0.00691494f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_2645 N_D[1]_M1002_g N_VPWR_c_7352_n 0.0035837f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_2646 N_D[1]_M1038_g N_VPWR_c_7352_n 0.0035837f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_2647 N_D[1]_M1134_g N_VPWR_c_7353_n 0.0035837f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_2648 N_D[1]_M1271_g N_VPWR_c_7353_n 0.0035837f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_2649 N_D[1]_M1002_g N_Z_c_9117_n 0.00311896f $X=10.975 $Y=1.985 $X2=0 $Y2=0
cc_2650 N_D[1]_M1038_g N_Z_c_9117_n 0.00306964f $X=11.445 $Y=1.985 $X2=0 $Y2=0
cc_2651 N_D[1]_M1134_g N_Z_c_9117_n 0.00306964f $X=11.915 $Y=1.985 $X2=0 $Y2=0
cc_2652 N_D[1]_M1271_g N_Z_c_9117_n 0.00470782f $X=12.385 $Y=1.985 $X2=0 $Y2=0
cc_2653 N_D[1]_c_3025_n N_Z_c_9117_n 0.00846955f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_2654 N_D[1]_M1002_g N_A_1643_311#_c_10897_n 0.013247f $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_2655 N_D[1]_M1038_g N_A_1643_311#_c_10919_n 0.00916655f $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_2656 N_D[1]_M1134_g N_A_1643_311#_c_10919_n 0.00916655f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_2657 N_D[1]_c_3023_n N_A_1643_311#_c_10919_n 7.15862e-19 $X=11.825 $Y=1.16
+ $X2=0 $Y2=0
cc_2658 N_D[1]_c_3025_n N_A_1643_311#_c_10919_n 0.0387168f $X=12.28 $Y=1.16
+ $X2=0 $Y2=0
cc_2659 N_D[1]_M1002_g N_A_1643_311#_c_10923_n 8.61029e-19 $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_2660 N_D[1]_M1038_g N_A_1643_311#_c_10923_n 5.79575e-19 $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_2661 N_D[1]_c_3024_n N_A_1643_311#_c_10923_n 8.03631e-19 $X=11.535 $Y=1.16
+ $X2=0 $Y2=0
cc_2662 N_D[1]_c_3025_n N_A_1643_311#_c_10923_n 0.0191156f $X=12.28 $Y=1.16
+ $X2=0 $Y2=0
cc_2663 N_D[1]_M1134_g N_A_1643_311#_c_10927_n 5.79575e-19 $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_2664 N_D[1]_M1271_g N_A_1643_311#_c_10927_n 0.00215964f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_2665 N_D[1]_c_3025_n N_A_1643_311#_c_10927_n 0.0217153f $X=12.28 $Y=1.16
+ $X2=0 $Y2=0
cc_2666 N_D[1]_c_3026_n N_A_1643_311#_c_10927_n 8.03631e-19 $X=12.385 $Y=1.16
+ $X2=0 $Y2=0
cc_2667 N_D[1]_M1002_g N_A_1643_311#_c_10899_n 0.00232998f $X=10.975 $Y=1.985
+ $X2=25.99 $Y2=0.51
cc_2668 N_D[1]_M1038_g N_A_1643_311#_c_10932_n 0.00232998f $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_2669 N_D[1]_M1134_g N_A_1643_311#_c_10932_n 0.00232998f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_2670 N_D[1]_M1002_g N_A_1643_311#_c_10934_n 0.00977623f $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_2671 N_D[1]_M1038_g N_A_1643_311#_c_10934_n 0.00911325f $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_2672 N_D[1]_M1134_g N_A_1643_311#_c_10934_n 7.05028e-19 $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_2673 N_D[1]_M1038_g N_A_1643_311#_c_10937_n 7.05028e-19 $X=11.445 $Y=1.985
+ $X2=0 $Y2=0
cc_2674 N_D[1]_M1134_g N_A_1643_311#_c_10937_n 0.00911325f $X=11.915 $Y=1.985
+ $X2=0 $Y2=0
cc_2675 N_D[1]_M1271_g N_A_1643_311#_c_10937_n 0.00847082f $X=12.385 $Y=1.985
+ $X2=0 $Y2=0
cc_2676 N_D[1]_M1002_g N_A_1643_311#_c_10902_n 0.00333758f $X=10.975 $Y=1.985
+ $X2=0 $Y2=0
cc_2677 N_D[1]_M1049_g N_VGND_c_12707_n 0.00321269f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_2678 N_D[1]_M1098_g N_VGND_c_12707_n 2.6376e-19 $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_2679 N_D[1]_M1098_g N_VGND_c_12709_n 0.0019152f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_2680 N_D[1]_M1167_g N_VGND_c_12709_n 0.00166854f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_2681 N_D[1]_M1315_g N_VGND_c_12709_n 2.64031e-19 $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_2682 N_D[1]_M1315_g N_VGND_c_12711_n 0.00345859f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_2683 N_D[1]_M1049_g VGND 0.00702263f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_2684 N_D[1]_M1098_g VGND 0.00624811f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_2685 N_D[1]_M1167_g VGND 0.00593887f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_2686 N_D[1]_M1315_g VGND 0.0111368f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_2687 N_D[1]_M1049_g N_VGND_c_12872_n 0.00422241f $X=11 $Y=0.56 $X2=0 $Y2=0
cc_2688 N_D[1]_M1098_g N_VGND_c_12872_n 0.00430643f $X=11.42 $Y=0.56 $X2=0 $Y2=0
cc_2689 N_D[1]_M1167_g N_VGND_c_12874_n 0.00422241f $X=11.94 $Y=0.56 $X2=0 $Y2=0
cc_2690 N_D[1]_M1315_g N_VGND_c_12874_n 0.00551064f $X=12.36 $Y=0.56 $X2=0 $Y2=0
cc_2691 N_D[1]_M1049_g N_A_1693_66#_c_14215_n 0.00261078f $X=11 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_2692 N_D[1]_M1049_g N_A_1693_66#_c_14216_n 0.0121912f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_2693 N_D[1]_M1049_g N_A_1693_66#_c_14236_n 0.00699463f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_2694 N_D[1]_M1098_g N_A_1693_66#_c_14236_n 0.00661764f $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_2695 N_D[1]_M1167_g N_A_1693_66#_c_14236_n 5.22365e-19 $X=11.94 $Y=0.56 $X2=0
+ $Y2=0
cc_2696 N_D[1]_M1098_g N_A_1693_66#_c_14218_n 0.00900364f $X=11.42 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_2697 N_D[1]_M1167_g N_A_1693_66#_c_14218_n 0.00986515f $X=11.94 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_2698 N_D[1]_M1315_g N_A_1693_66#_c_14218_n 0.00228093f $X=12.36 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_2699 N_D[1]_c_3023_n N_A_1693_66#_c_14218_n 0.00463549f $X=11.825 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_2700 N_D[1]_c_3025_n N_A_1693_66#_c_14218_n 0.0608884f $X=12.28 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_2701 N_D[1]_c_3026_n N_A_1693_66#_c_14218_n 0.00208088f $X=12.385 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_2702 N_D[1]_M1098_g N_A_1693_66#_c_14245_n 5.22365e-19 $X=11.42 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_2703 N_D[1]_M1167_g N_A_1693_66#_c_14245_n 0.00661134f $X=11.94 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_2704 N_D[1]_M1315_g N_A_1693_66#_c_14245_n 0.00529286f $X=12.36 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_2705 N_D[1]_M1049_g N_A_1693_66#_c_14219_n 0.00128201f $X=11 $Y=0.56 $X2=0
+ $Y2=0
cc_2706 N_D[1]_M1098_g N_A_1693_66#_c_14219_n 8.68782e-19 $X=11.42 $Y=0.56 $X2=0
+ $Y2=0
cc_2707 N_D[1]_c_3024_n N_A_1693_66#_c_14219_n 0.00208088f $X=11.535 $Y=1.16
+ $X2=0 $Y2=0
cc_2708 N_D[1]_c_3025_n N_A_1693_66#_c_14219_n 0.018367f $X=12.28 $Y=1.16 $X2=0
+ $Y2=0
cc_2709 N_D[9]_M1011_g N_VPWR_c_7234_n 0.00389633f $X=10.975 $Y=3.455 $X2=0
+ $Y2=0
cc_2710 N_D[9]_M1051_g N_VPWR_c_7236_n 0.00208662f $X=11.445 $Y=3.455 $X2=0
+ $Y2=0
cc_2711 N_D[9]_M1148_g N_VPWR_c_7236_n 0.00208662f $X=11.915 $Y=3.455 $X2=0
+ $Y2=0
cc_2712 N_D[9]_M1285_g N_VPWR_c_7238_n 0.00374733f $X=12.385 $Y=3.455 $X2=0
+ $Y2=0
cc_2713 N_D[9]_M1011_g VPWR 0.00573859f $X=10.975 $Y=3.455 $X2=0 $Y2=0
cc_2714 N_D[9]_M1051_g VPWR 0.00445624f $X=11.445 $Y=3.455 $X2=0 $Y2=0
cc_2715 N_D[9]_M1148_g VPWR 0.00445624f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_2716 N_D[9]_M1285_g VPWR 0.00691494f $X=12.385 $Y=3.455 $X2=0 $Y2=0
cc_2717 N_D[9]_M1011_g N_VPWR_c_7352_n 0.0035837f $X=10.975 $Y=3.455 $X2=0 $Y2=0
cc_2718 N_D[9]_M1051_g N_VPWR_c_7352_n 0.0035837f $X=11.445 $Y=3.455 $X2=0 $Y2=0
cc_2719 N_D[9]_M1148_g N_VPWR_c_7353_n 0.0035837f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_2720 N_D[9]_M1285_g N_VPWR_c_7353_n 0.0035837f $X=12.385 $Y=3.455 $X2=0 $Y2=0
cc_2721 N_D[9]_M1011_g N_Z_c_9118_n 0.00311896f $X=10.975 $Y=3.455 $X2=0 $Y2=0
cc_2722 N_D[9]_M1051_g N_Z_c_9118_n 0.00306964f $X=11.445 $Y=3.455 $X2=0 $Y2=0
cc_2723 N_D[9]_M1148_g N_Z_c_9118_n 0.00306964f $X=11.915 $Y=3.455 $X2=0 $Y2=0
cc_2724 N_D[9]_M1285_g N_Z_c_9118_n 0.00470782f $X=12.385 $Y=3.455 $X2=0 $Y2=0
cc_2725 N_D[9]_c_3118_n N_Z_c_9118_n 0.00846955f $X=12.28 $Y=4.28 $X2=0 $Y2=0
cc_2726 N_D[9]_M1011_g N_A_1643_613#_c_11028_n 0.013247f $X=10.975 $Y=3.455
+ $X2=0 $Y2=0
cc_2727 N_D[9]_M1051_g N_A_1643_613#_c_11050_n 0.00916655f $X=11.445 $Y=3.455
+ $X2=0 $Y2=0
cc_2728 N_D[9]_M1148_g N_A_1643_613#_c_11050_n 0.00916655f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_2729 N_D[9]_c_3116_n N_A_1643_613#_c_11050_n 7.15862e-19 $X=11.825 $Y=4.28
+ $X2=0 $Y2=0
cc_2730 N_D[9]_c_3118_n N_A_1643_613#_c_11050_n 0.0387168f $X=12.28 $Y=4.28
+ $X2=0 $Y2=0
cc_2731 N_D[9]_M1011_g N_A_1643_613#_c_11054_n 8.61029e-19 $X=10.975 $Y=3.455
+ $X2=0 $Y2=0
cc_2732 N_D[9]_M1051_g N_A_1643_613#_c_11054_n 5.79575e-19 $X=11.445 $Y=3.455
+ $X2=0 $Y2=0
cc_2733 N_D[9]_c_3117_n N_A_1643_613#_c_11054_n 8.03631e-19 $X=11.535 $Y=4.28
+ $X2=0 $Y2=0
cc_2734 N_D[9]_c_3118_n N_A_1643_613#_c_11054_n 0.0191156f $X=12.28 $Y=4.28
+ $X2=0 $Y2=0
cc_2735 N_D[9]_M1148_g N_A_1643_613#_c_11058_n 5.79575e-19 $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_2736 N_D[9]_M1285_g N_A_1643_613#_c_11058_n 0.00215964f $X=12.385 $Y=3.455
+ $X2=0 $Y2=0
cc_2737 N_D[9]_c_3118_n N_A_1643_613#_c_11058_n 0.0217153f $X=12.28 $Y=4.28
+ $X2=0 $Y2=0
cc_2738 N_D[9]_c_3119_n N_A_1643_613#_c_11058_n 8.03631e-19 $X=12.385 $Y=4.28
+ $X2=0 $Y2=0
cc_2739 N_D[9]_M1011_g N_A_1643_613#_c_11030_n 0.00232998f $X=10.975 $Y=3.455
+ $X2=25.99 $Y2=0.51
cc_2740 N_D[9]_M1051_g N_A_1643_613#_c_11063_n 0.00232998f $X=11.445 $Y=3.455
+ $X2=0 $Y2=0
cc_2741 N_D[9]_M1148_g N_A_1643_613#_c_11063_n 0.00232998f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_2742 N_D[9]_M1011_g N_A_1643_613#_c_11033_n 0.00333758f $X=10.975 $Y=3.455
+ $X2=0 $Y2=0
cc_2743 N_D[9]_M1011_g N_A_1643_613#_c_11066_n 0.00977623f $X=10.975 $Y=3.455
+ $X2=0 $Y2=0
cc_2744 N_D[9]_M1051_g N_A_1643_613#_c_11066_n 0.00911325f $X=11.445 $Y=3.455
+ $X2=0 $Y2=0
cc_2745 N_D[9]_M1148_g N_A_1643_613#_c_11066_n 7.05028e-19 $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_2746 N_D[9]_M1051_g N_A_1643_613#_c_11069_n 7.05028e-19 $X=11.445 $Y=3.455
+ $X2=0 $Y2=0
cc_2747 N_D[9]_M1148_g N_A_1643_613#_c_11069_n 0.00911325f $X=11.915 $Y=3.455
+ $X2=0 $Y2=0
cc_2748 N_D[9]_M1285_g N_A_1643_613#_c_11069_n 0.00847082f $X=12.385 $Y=3.455
+ $X2=0 $Y2=0
cc_2749 N_D[9]_M1019_g N_VGND_c_12708_n 0.00321269f $X=11 $Y=4.88 $X2=0 $Y2=0
cc_2750 N_D[9]_M1111_g N_VGND_c_12708_n 2.6376e-19 $X=11.42 $Y=4.88 $X2=0 $Y2=0
cc_2751 N_D[9]_M1111_g N_VGND_c_12710_n 0.0019152f $X=11.42 $Y=4.88 $X2=0 $Y2=0
cc_2752 N_D[9]_M1178_g N_VGND_c_12710_n 0.00166854f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_2753 N_D[9]_M1276_g N_VGND_c_12710_n 2.64031e-19 $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_2754 N_D[9]_M1276_g N_VGND_c_12712_n 0.00345859f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_2755 N_D[9]_M1019_g VGND 0.00702263f $X=11 $Y=4.88 $X2=0 $Y2=0
cc_2756 N_D[9]_M1111_g VGND 0.00624811f $X=11.42 $Y=4.88 $X2=0 $Y2=0
cc_2757 N_D[9]_M1178_g VGND 0.00593887f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_2758 N_D[9]_M1276_g VGND 0.0111368f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_2759 N_D[9]_M1019_g N_VGND_c_12873_n 0.00422241f $X=11 $Y=4.88 $X2=0 $Y2=0
cc_2760 N_D[9]_M1111_g N_VGND_c_12873_n 0.00430643f $X=11.42 $Y=4.88 $X2=0 $Y2=0
cc_2761 N_D[9]_M1178_g N_VGND_c_12875_n 0.00422241f $X=11.94 $Y=4.88 $X2=0 $Y2=0
cc_2762 N_D[9]_M1276_g N_VGND_c_12875_n 0.00551064f $X=12.36 $Y=4.88 $X2=0 $Y2=0
cc_2763 N_D[9]_M1019_g N_A_1693_918#_c_14299_n 0.00261078f $X=11 $Y=4.88
+ $X2=25.99 $Y2=0.51
cc_2764 N_D[9]_M1019_g N_A_1693_918#_c_14300_n 0.0121912f $X=11 $Y=4.88 $X2=0
+ $Y2=0
cc_2765 N_D[9]_M1111_g N_A_1693_918#_c_14320_n 0.00900364f $X=11.42 $Y=4.88
+ $X2=0 $Y2=0
cc_2766 N_D[9]_M1178_g N_A_1693_918#_c_14320_n 0.00899636f $X=11.94 $Y=4.88
+ $X2=0 $Y2=0
cc_2767 N_D[9]_c_3116_n N_A_1693_918#_c_14320_n 0.00463549f $X=11.825 $Y=4.28
+ $X2=0 $Y2=0
cc_2768 N_D[9]_c_3118_n N_A_1693_918#_c_14320_n 0.0394855f $X=12.28 $Y=4.28
+ $X2=0 $Y2=0
cc_2769 N_D[9]_M1019_g N_A_1693_918#_c_14302_n 0.00827664f $X=11 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_2770 N_D[9]_M1111_g N_A_1693_918#_c_14302_n 0.00748643f $X=11.42 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_2771 N_D[9]_M1178_g N_A_1693_918#_c_14302_n 5.22365e-19 $X=11.94 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_2772 N_D[9]_c_3117_n N_A_1693_918#_c_14302_n 0.00208088f $X=11.535 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_2773 N_D[9]_c_3118_n N_A_1693_918#_c_14302_n 0.018367f $X=12.28 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_2774 N_D[9]_M1111_g N_A_1693_918#_c_14303_n 5.22365e-19 $X=11.42 $Y=4.88
+ $X2=0 $Y2=0
cc_2775 N_D[9]_M1178_g N_A_1693_918#_c_14303_n 0.00748012f $X=11.94 $Y=4.88
+ $X2=0 $Y2=0
cc_2776 N_D[9]_M1276_g N_A_1693_918#_c_14303_n 0.00757379f $X=12.36 $Y=4.88
+ $X2=0 $Y2=0
cc_2777 N_D[9]_c_3118_n N_A_1693_918#_c_14303_n 0.021403f $X=12.28 $Y=4.28 $X2=0
+ $Y2=0
cc_2778 N_D[9]_c_3119_n N_A_1693_918#_c_14303_n 0.00208088f $X=12.385 $Y=4.28
+ $X2=0 $Y2=0
cc_2779 N_D[2]_M1020_g N_D[10]_M1024_g 0.0130744f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2780 N_D[2]_M1067_g N_D[10]_M1076_g 0.0130744f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2781 N_D[2]_M1157_g N_D[10]_M1164_g 0.0130744f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_2782 N_D[2]_M1301_g N_D[10]_M1309_g 0.0130744f $X=14.785 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_2783 N_D[2]_M1020_g N_VPWR_c_7240_n 0.00374733f $X=13.375 $Y=1.985 $X2=0
+ $Y2=0
cc_2784 N_D[2]_M1067_g N_VPWR_c_7242_n 0.00208662f $X=13.845 $Y=1.985 $X2=0
+ $Y2=0
cc_2785 N_D[2]_M1157_g N_VPWR_c_7242_n 0.00208662f $X=14.315 $Y=1.985 $X2=0
+ $Y2=0
cc_2786 N_D[2]_M1157_g N_VPWR_c_7244_n 0.0035837f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_2787 N_D[2]_M1301_g N_VPWR_c_7244_n 0.0035837f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_2788 N_D[2]_M1301_g N_VPWR_c_7245_n 0.00389633f $X=14.785 $Y=1.985 $X2=0
+ $Y2=0
cc_2789 N_D[2]_M1020_g VPWR 0.00691494f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2790 N_D[2]_M1067_g VPWR 0.00445624f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2791 N_D[2]_M1157_g VPWR 0.00445624f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_2792 N_D[2]_M1301_g VPWR 0.00573859f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_2793 N_D[2]_M1020_g N_VPWR_c_7354_n 0.0035837f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2794 N_D[2]_M1067_g N_VPWR_c_7354_n 0.0035837f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2795 N_D[2]_M1020_g N_Z_c_9117_n 0.00470782f $X=13.375 $Y=1.985 $X2=0 $Y2=0
cc_2796 N_D[2]_M1067_g N_Z_c_9117_n 0.00306964f $X=13.845 $Y=1.985 $X2=0 $Y2=0
cc_2797 N_D[2]_M1157_g N_Z_c_9117_n 0.00306964f $X=14.315 $Y=1.985 $X2=0 $Y2=0
cc_2798 N_D[2]_M1301_g N_Z_c_9117_n 0.00311896f $X=14.785 $Y=1.985 $X2=0 $Y2=0
cc_2799 N_D[2]_c_3209_n N_Z_c_9117_n 0.00846955f $X=14.5 $Y=1.16 $X2=0 $Y2=0
cc_2800 N_D[2]_M1067_g N_A_2693_297#_c_11164_n 0.00916655f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2801 N_D[2]_M1157_g N_A_2693_297#_c_11164_n 0.00916655f $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_2802 N_D[2]_c_3207_n N_A_2693_297#_c_11164_n 7.15862e-19 $X=14.225 $Y=1.16
+ $X2=0 $Y2=0
cc_2803 N_D[2]_c_3209_n N_A_2693_297#_c_11164_n 0.0387168f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2804 N_D[2]_M1301_g N_A_2693_297#_c_11159_n 0.013247f $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_2805 N_D[2]_M1020_g N_A_2693_297#_c_11169_n 0.00215964f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_2806 N_D[2]_M1067_g N_A_2693_297#_c_11169_n 5.79575e-19 $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2807 N_D[2]_c_3208_n N_A_2693_297#_c_11169_n 8.03631e-19 $X=13.935 $Y=1.16
+ $X2=0 $Y2=0
cc_2808 N_D[2]_c_3209_n N_A_2693_297#_c_11169_n 0.0217153f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2809 N_D[2]_M1157_g N_A_2693_297#_c_11173_n 5.79575e-19 $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_2810 N_D[2]_M1301_g N_A_2693_297#_c_11173_n 8.61029e-19 $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_2811 N_D[2]_c_3209_n N_A_2693_297#_c_11173_n 0.0191156f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2812 N_D[2]_c_3210_n N_A_2693_297#_c_11173_n 8.03631e-19 $X=14.785 $Y=1.16
+ $X2=0 $Y2=0
cc_2813 N_D[2]_M1067_g N_A_2693_297#_c_11177_n 0.00232998f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2814 N_D[2]_M1157_g N_A_2693_297#_c_11177_n 0.00232998f $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_2815 N_D[2]_M1301_g N_A_2693_297#_c_11160_n 0.00232998f $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_2816 N_D[2]_M1020_g N_A_2693_297#_c_11180_n 0.00847082f $X=13.375 $Y=1.985
+ $X2=0 $Y2=0
cc_2817 N_D[2]_M1067_g N_A_2693_297#_c_11180_n 0.00911325f $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2818 N_D[2]_M1157_g N_A_2693_297#_c_11180_n 7.05028e-19 $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_2819 N_D[2]_M1067_g N_A_2693_297#_c_11183_n 7.05028e-19 $X=13.845 $Y=1.985
+ $X2=0 $Y2=0
cc_2820 N_D[2]_M1157_g N_A_2693_297#_c_11183_n 0.00911325f $X=14.315 $Y=1.985
+ $X2=0 $Y2=0
cc_2821 N_D[2]_M1301_g N_A_2693_297#_c_11183_n 0.00977623f $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_2822 N_D[2]_M1301_g N_A_2693_297#_c_11161_n 0.00333758f $X=14.785 $Y=1.985
+ $X2=0 $Y2=0
cc_2823 N_D[2]_M1001_g N_VGND_c_12715_n 0.00345859f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2824 N_D[2]_M1001_g N_VGND_c_12717_n 2.64031e-19 $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2825 N_D[2]_M1062_g N_VGND_c_12717_n 0.00166854f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2826 N_D[2]_M1110_g N_VGND_c_12717_n 0.0019152f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_2827 N_D[2]_M1110_g N_VGND_c_12719_n 0.00430643f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_2828 N_D[2]_M1182_g N_VGND_c_12719_n 0.00422241f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_2829 N_D[2]_M1110_g N_VGND_c_12721_n 2.6376e-19 $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_2830 N_D[2]_M1182_g N_VGND_c_12721_n 0.00321269f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_2831 N_D[2]_M1001_g VGND 0.0111368f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2832 N_D[2]_M1062_g VGND 0.00593887f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2833 N_D[2]_M1110_g VGND 0.00624811f $X=14.34 $Y=0.56 $X2=0 $Y2=0
cc_2834 N_D[2]_M1182_g VGND 0.00702263f $X=14.76 $Y=0.56 $X2=0 $Y2=0
cc_2835 N_D[2]_M1001_g N_VGND_c_12876_n 0.00551064f $X=13.4 $Y=0.56 $X2=0 $Y2=0
cc_2836 N_D[2]_M1062_g N_VGND_c_12876_n 0.00422241f $X=13.82 $Y=0.56 $X2=0 $Y2=0
cc_2837 N_D[2]_M1001_g N_A_2695_47#_c_14385_n 0.00529286f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2838 N_D[2]_M1062_g N_A_2695_47#_c_14385_n 0.00661134f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2839 N_D[2]_M1110_g N_A_2695_47#_c_14385_n 5.22365e-19 $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2840 N_D[2]_M1062_g N_A_2695_47#_c_14388_n 0.00899636f $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2841 N_D[2]_M1110_g N_A_2695_47#_c_14388_n 0.00900364f $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2842 N_D[2]_c_3207_n N_A_2695_47#_c_14388_n 0.00463549f $X=14.225 $Y=1.16
+ $X2=0 $Y2=0
cc_2843 N_D[2]_c_3209_n N_A_2695_47#_c_14388_n 0.0394855f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2844 N_D[2]_M1001_g N_A_2695_47#_c_14377_n 0.00228093f $X=13.4 $Y=0.56 $X2=0
+ $Y2=0
cc_2845 N_D[2]_M1062_g N_A_2695_47#_c_14377_n 8.68782e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2846 N_D[2]_c_3208_n N_A_2695_47#_c_14377_n 0.00208088f $X=13.935 $Y=1.16
+ $X2=0 $Y2=0
cc_2847 N_D[2]_c_3209_n N_A_2695_47#_c_14377_n 0.021403f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2848 N_D[2]_M1062_g N_A_2695_47#_c_14396_n 5.22365e-19 $X=13.82 $Y=0.56 $X2=0
+ $Y2=0
cc_2849 N_D[2]_M1110_g N_A_2695_47#_c_14396_n 0.00661764f $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2850 N_D[2]_M1182_g N_A_2695_47#_c_14396_n 0.00699463f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_2851 N_D[2]_M1182_g N_A_2695_47#_c_14378_n 0.0121912f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_2852 N_D[2]_M1182_g N_A_2695_47#_c_14379_n 0.00261078f $X=14.76 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_2853 N_D[2]_M1110_g N_A_2695_47#_c_14384_n 8.68782e-19 $X=14.34 $Y=0.56 $X2=0
+ $Y2=0
cc_2854 N_D[2]_M1182_g N_A_2695_47#_c_14384_n 0.00128201f $X=14.76 $Y=0.56 $X2=0
+ $Y2=0
cc_2855 N_D[2]_c_3209_n N_A_2695_47#_c_14384_n 0.018367f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_2856 N_D[2]_c_3210_n N_A_2695_47#_c_14384_n 0.00208088f $X=14.785 $Y=1.16
+ $X2=0 $Y2=0
cc_2857 N_D[10]_M1024_g N_VPWR_c_7241_n 0.00374733f $X=13.375 $Y=3.455 $X2=0
+ $Y2=0
cc_2858 N_D[10]_M1076_g N_VPWR_c_7243_n 0.00208662f $X=13.845 $Y=3.455 $X2=0
+ $Y2=0
cc_2859 N_D[10]_M1164_g N_VPWR_c_7243_n 0.00208662f $X=14.315 $Y=3.455 $X2=0
+ $Y2=0
cc_2860 N_D[10]_M1164_g N_VPWR_c_7244_n 0.0035837f $X=14.315 $Y=3.455 $X2=0
+ $Y2=0
cc_2861 N_D[10]_M1309_g N_VPWR_c_7244_n 0.0035837f $X=14.785 $Y=3.455 $X2=0
+ $Y2=0
cc_2862 N_D[10]_M1309_g N_VPWR_c_7246_n 0.00389633f $X=14.785 $Y=3.455 $X2=0
+ $Y2=0
cc_2863 N_D[10]_M1024_g VPWR 0.00691494f $X=13.375 $Y=3.455 $X2=0 $Y2=0
cc_2864 N_D[10]_M1076_g VPWR 0.00445624f $X=13.845 $Y=3.455 $X2=0 $Y2=0
cc_2865 N_D[10]_M1164_g VPWR 0.00445624f $X=14.315 $Y=3.455 $X2=0 $Y2=0
cc_2866 N_D[10]_M1309_g VPWR 0.00573859f $X=14.785 $Y=3.455 $X2=0 $Y2=0
cc_2867 N_D[10]_M1024_g N_VPWR_c_7354_n 0.0035837f $X=13.375 $Y=3.455 $X2=0
+ $Y2=0
cc_2868 N_D[10]_M1076_g N_VPWR_c_7354_n 0.0035837f $X=13.845 $Y=3.455 $X2=0
+ $Y2=0
cc_2869 N_D[10]_M1024_g N_Z_c_9118_n 0.00470782f $X=13.375 $Y=3.455 $X2=0 $Y2=0
cc_2870 N_D[10]_M1076_g N_Z_c_9118_n 0.00306964f $X=13.845 $Y=3.455 $X2=0 $Y2=0
cc_2871 N_D[10]_M1164_g N_Z_c_9118_n 0.00306964f $X=14.315 $Y=3.455 $X2=0 $Y2=0
cc_2872 N_D[10]_M1309_g N_Z_c_9118_n 0.00311896f $X=14.785 $Y=3.455 $X2=0 $Y2=0
cc_2873 N_D[10]_c_3304_n N_Z_c_9118_n 0.00846955f $X=14.5 $Y=4.28 $X2=0 $Y2=0
cc_2874 N_D[10]_M1076_g N_A_2693_591#_c_11292_n 0.00916655f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2875 N_D[10]_M1164_g N_A_2693_591#_c_11292_n 0.00916655f $X=14.315 $Y=3.455
+ $X2=0 $Y2=0
cc_2876 N_D[10]_c_3302_n N_A_2693_591#_c_11292_n 7.15862e-19 $X=14.225 $Y=4.28
+ $X2=0 $Y2=0
cc_2877 N_D[10]_c_3304_n N_A_2693_591#_c_11292_n 0.0387168f $X=14.5 $Y=4.28
+ $X2=0 $Y2=0
cc_2878 N_D[10]_M1309_g N_A_2693_591#_c_11287_n 0.013247f $X=14.785 $Y=3.455
+ $X2=0 $Y2=0
cc_2879 N_D[10]_M1024_g N_A_2693_591#_c_11297_n 0.00215964f $X=13.375 $Y=3.455
+ $X2=0 $Y2=0
cc_2880 N_D[10]_M1076_g N_A_2693_591#_c_11297_n 5.79575e-19 $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2881 N_D[10]_c_3303_n N_A_2693_591#_c_11297_n 8.03631e-19 $X=13.935 $Y=4.28
+ $X2=0 $Y2=0
cc_2882 N_D[10]_c_3304_n N_A_2693_591#_c_11297_n 0.0217153f $X=14.5 $Y=4.28
+ $X2=0 $Y2=0
cc_2883 N_D[10]_M1164_g N_A_2693_591#_c_11301_n 5.79575e-19 $X=14.315 $Y=3.455
+ $X2=0 $Y2=0
cc_2884 N_D[10]_M1309_g N_A_2693_591#_c_11301_n 8.61029e-19 $X=14.785 $Y=3.455
+ $X2=0 $Y2=0
cc_2885 N_D[10]_c_3304_n N_A_2693_591#_c_11301_n 0.0191156f $X=14.5 $Y=4.28
+ $X2=0 $Y2=0
cc_2886 N_D[10]_c_3305_n N_A_2693_591#_c_11301_n 8.03631e-19 $X=14.785 $Y=4.28
+ $X2=0 $Y2=0
cc_2887 N_D[10]_M1076_g N_A_2693_591#_c_11305_n 0.00232998f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2888 N_D[10]_M1164_g N_A_2693_591#_c_11305_n 0.00232998f $X=14.315 $Y=3.455
+ $X2=0 $Y2=0
cc_2889 N_D[10]_M1309_g N_A_2693_591#_c_11288_n 0.00232998f $X=14.785 $Y=3.455
+ $X2=0 $Y2=0
cc_2890 N_D[10]_M1024_g N_A_2693_591#_c_11308_n 0.00847082f $X=13.375 $Y=3.455
+ $X2=0 $Y2=0
cc_2891 N_D[10]_M1076_g N_A_2693_591#_c_11308_n 0.00911325f $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2892 N_D[10]_M1164_g N_A_2693_591#_c_11308_n 7.05028e-19 $X=14.315 $Y=3.455
+ $X2=0 $Y2=0
cc_2893 N_D[10]_M1076_g N_A_2693_591#_c_11311_n 7.05028e-19 $X=13.845 $Y=3.455
+ $X2=0 $Y2=0
cc_2894 N_D[10]_M1164_g N_A_2693_591#_c_11311_n 0.00911325f $X=14.315 $Y=3.455
+ $X2=0 $Y2=0
cc_2895 N_D[10]_M1309_g N_A_2693_591#_c_11311_n 0.00977623f $X=14.785 $Y=3.455
+ $X2=0 $Y2=0
cc_2896 N_D[10]_M1309_g N_A_2693_591#_c_11289_n 0.00333758f $X=14.785 $Y=3.455
+ $X2=0 $Y2=0
cc_2897 N_D[10]_M1033_g N_VGND_c_12716_n 0.00345859f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2898 N_D[10]_M1033_g N_VGND_c_12718_n 2.64031e-19 $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2899 N_D[10]_M1143_g N_VGND_c_12718_n 0.00166854f $X=13.82 $Y=4.88 $X2=0
+ $Y2=0
cc_2900 N_D[10]_M1195_g N_VGND_c_12718_n 0.0019152f $X=14.34 $Y=4.88 $X2=0 $Y2=0
cc_2901 N_D[10]_M1195_g N_VGND_c_12720_n 0.00430643f $X=14.34 $Y=4.88 $X2=0
+ $Y2=0
cc_2902 N_D[10]_M1307_g N_VGND_c_12720_n 0.00422241f $X=14.76 $Y=4.88 $X2=0
+ $Y2=0
cc_2903 N_D[10]_M1195_g N_VGND_c_12722_n 2.6376e-19 $X=14.34 $Y=4.88 $X2=0 $Y2=0
cc_2904 N_D[10]_M1307_g N_VGND_c_12722_n 0.00321269f $X=14.76 $Y=4.88 $X2=0
+ $Y2=0
cc_2905 N_D[10]_M1033_g VGND 0.0111368f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2906 N_D[10]_M1143_g VGND 0.00593887f $X=13.82 $Y=4.88 $X2=0 $Y2=0
cc_2907 N_D[10]_M1195_g VGND 0.00624811f $X=14.34 $Y=4.88 $X2=0 $Y2=0
cc_2908 N_D[10]_M1307_g VGND 0.00702263f $X=14.76 $Y=4.88 $X2=0 $Y2=0
cc_2909 N_D[10]_M1033_g N_VGND_c_12877_n 0.00551064f $X=13.4 $Y=4.88 $X2=0 $Y2=0
cc_2910 N_D[10]_M1143_g N_VGND_c_12877_n 0.00422241f $X=13.82 $Y=4.88 $X2=0
+ $Y2=0
cc_2911 N_D[10]_M1143_g N_A_2695_911#_c_14468_n 0.00899636f $X=13.82 $Y=4.88
+ $X2=0 $Y2=0
cc_2912 N_D[10]_M1195_g N_A_2695_911#_c_14468_n 0.00900364f $X=14.34 $Y=4.88
+ $X2=0 $Y2=0
cc_2913 N_D[10]_c_3302_n N_A_2695_911#_c_14468_n 0.00463549f $X=14.225 $Y=4.28
+ $X2=0 $Y2=0
cc_2914 N_D[10]_c_3304_n N_A_2695_911#_c_14468_n 0.0394855f $X=14.5 $Y=4.28
+ $X2=0 $Y2=0
cc_2915 N_D[10]_M1307_g N_A_2695_911#_c_14460_n 0.0121912f $X=14.76 $Y=4.88
+ $X2=0 $Y2=0
cc_2916 N_D[10]_M1307_g N_A_2695_911#_c_14461_n 0.00261078f $X=14.76 $Y=4.88
+ $X2=0 $Y2=0
cc_2917 N_D[10]_M1033_g N_A_2695_911#_c_14466_n 0.00757379f $X=13.4 $Y=4.88
+ $X2=0 $Y2=0
cc_2918 N_D[10]_M1143_g N_A_2695_911#_c_14466_n 0.00748012f $X=13.82 $Y=4.88
+ $X2=0 $Y2=0
cc_2919 N_D[10]_M1195_g N_A_2695_911#_c_14466_n 5.22365e-19 $X=14.34 $Y=4.88
+ $X2=0 $Y2=0
cc_2920 N_D[10]_c_3303_n N_A_2695_911#_c_14466_n 0.00208088f $X=13.935 $Y=4.28
+ $X2=0 $Y2=0
cc_2921 N_D[10]_c_3304_n N_A_2695_911#_c_14466_n 0.021403f $X=14.5 $Y=4.28 $X2=0
+ $Y2=0
cc_2922 N_D[10]_M1143_g N_A_2695_911#_c_14467_n 5.22365e-19 $X=13.82 $Y=4.88
+ $X2=0 $Y2=0
cc_2923 N_D[10]_M1195_g N_A_2695_911#_c_14467_n 0.00748643f $X=14.34 $Y=4.88
+ $X2=0 $Y2=0
cc_2924 N_D[10]_M1307_g N_A_2695_911#_c_14467_n 0.00827664f $X=14.76 $Y=4.88
+ $X2=0 $Y2=0
cc_2925 N_D[10]_c_3304_n N_A_2695_911#_c_14467_n 0.018367f $X=14.5 $Y=4.28 $X2=0
+ $Y2=0
cc_2926 N_D[10]_c_3305_n N_A_2695_911#_c_14467_n 0.00208088f $X=14.785 $Y=4.28
+ $X2=0 $Y2=0
cc_2927 N_A_3135_265#_c_3392_n N_A_3135_793#_c_3511_n 0.0129371f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_2928 N_A_3135_265#_c_3395_n N_A_3135_793#_c_3514_n 0.0129371f $X=16.245
+ $Y=1.475 $X2=0 $Y2=0
cc_2929 N_A_3135_265#_c_3397_n N_A_3135_793#_c_3516_n 0.0129371f $X=16.715
+ $Y=1.475 $X2=0 $Y2=0
cc_2930 N_A_3135_265#_c_3399_n N_A_3135_793#_c_3518_n 0.0129371f $X=17.185
+ $Y=1.475 $X2=0 $Y2=0
cc_2931 N_A_3135_265#_c_3394_n N_S[2]_c_3629_n 0.00507426f $X=15.865 $Y=1.4
+ $X2=0 $Y2=0
cc_2932 N_A_3135_265#_c_3393_n N_S[2]_c_3632_n 0.00509391f $X=16.155 $Y=1.4
+ $X2=0 $Y2=0
cc_2933 N_A_3135_265#_c_3396_n N_S[2]_c_3634_n 0.00509204f $X=16.625 $Y=1.4
+ $X2=25.905 $Y2=4.845
cc_2934 N_A_3135_265#_c_3398_n N_S[2]_c_3636_n 0.00507688f $X=17.095 $Y=1.4
+ $X2=0 $Y2=0
cc_2935 N_A_3135_265#_c_3387_n N_S[2]_c_3638_n 6.53442e-19 $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_2936 N_A_3135_265#_c_3385_n N_S[2]_c_3640_n 0.0103812f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_2937 N_A_3135_265#_c_3386_n N_S[2]_c_3640_n 0.0179529f $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_2938 N_A_3135_265#_c_3385_n N_S[2]_c_3641_n 0.0206368f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_2939 N_A_3135_265#_c_3386_n N_S[2]_c_3641_n 0.0175393f $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_2940 N_A_3135_265#_c_3388_n N_S[2]_c_3641_n 0.0085951f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_2941 N_A_3135_265#_c_3390_n N_S[2]_c_3641_n 0.00322131f $X=18.385 $Y=1.23
+ $X2=0 $Y2=0
cc_2942 N_A_3135_265#_c_3406_n N_S[2]_c_3641_n 0.00255921f $X=18.465 $Y=1.605
+ $X2=0 $Y2=0
cc_2943 N_A_3135_265#_c_3391_n N_S[2]_c_3641_n 0.00262132f $X=17.505 $Y=1.23
+ $X2=0 $Y2=0
cc_2944 N_A_3135_265#_c_3404_n N_S[2]_c_3652_n 0.0118698f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_2945 N_A_3135_265#_c_3406_n N_S[2]_c_3652_n 0.00762115f $X=18.465 $Y=1.605
+ $X2=0 $Y2=0
cc_2946 N_A_3135_265#_c_3387_n N_S[2]_c_3642_n 0.00603996f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_2947 N_A_3135_265#_c_3389_n N_S[2]_c_3642_n 9.67113e-19 $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_2948 N_A_3135_265#_c_3388_n N_S[2]_c_3643_n 0.00429801f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_2949 N_A_3135_265#_c_3389_n N_S[2]_c_3643_n 0.0111895f $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_2950 N_A_3135_265#_c_3387_n N_S[2]_c_3644_n 0.00207203f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_2951 N_A_3135_265#_c_3388_n N_S[2]_c_3645_n 0.00289358f $X=18.385 $Y=1.065
+ $X2=25.99 $Y2=4.8
cc_2952 N_A_3135_265#_c_3404_n N_S[2]_c_3645_n 0.0128834f $X=18.465 $Y=1.77
+ $X2=25.99 $Y2=4.8
cc_2953 N_A_3135_265#_c_3390_n N_S[2]_c_3645_n 0.00416423f $X=18.385 $Y=1.23
+ $X2=25.99 $Y2=4.8
cc_2954 N_A_3135_265#_c_3406_n N_S[2]_c_3645_n 0.00454075f $X=18.465 $Y=1.605
+ $X2=25.99 $Y2=4.8
cc_2955 N_A_3135_265#_c_3388_n N_S[2]_c_3649_n 0.00268644f $X=18.385 $Y=1.065
+ $X2=0 $Y2=0
cc_2956 N_A_3135_265#_c_3389_n N_S[2]_c_3649_n 0.00426435f $X=18.425 $Y=0.825
+ $X2=0 $Y2=0
cc_2957 N_A_3135_265#_c_3388_n S[2] 0.00541767f $X=18.385 $Y=1.065 $X2=0 $Y2=0
cc_2958 N_A_3135_265#_c_3390_n S[2] 0.0228692f $X=18.385 $Y=1.23 $X2=0 $Y2=0
cc_2959 N_A_3135_265#_c_3392_n N_VPWR_c_7245_n 0.00324472f $X=15.775 $Y=1.475
+ $X2=0 $Y2=0
cc_2960 N_A_3135_265#_c_3399_n N_VPWR_c_7247_n 0.00367058f $X=17.185 $Y=1.475
+ $X2=0 $Y2=0
cc_2961 N_A_3135_265#_c_3385_n N_VPWR_c_7247_n 0.0193185f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_2962 N_A_3135_265#_c_3386_n N_VPWR_c_7247_n 6.4101e-19 $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_2963 N_A_3135_265#_c_3404_n N_VPWR_c_7247_n 0.0316788f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_2964 N_A_3135_265#_c_3404_n N_VPWR_c_7249_n 0.0356181f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_2965 N_A_3135_265#_c_3404_n N_VPWR_c_7322_n 0.0233824f $X=18.465 $Y=1.77
+ $X2=0 $Y2=0
cc_2966 N_A_3135_265#_c_3392_n VPWR 0.00473731f $X=15.775 $Y=1.475 $X2=0 $Y2=0
cc_2967 N_A_3135_265#_c_3395_n VPWR 0.00362156f $X=16.245 $Y=1.475 $X2=0 $Y2=0
cc_2968 N_A_3135_265#_c_3397_n VPWR 0.00362156f $X=16.715 $Y=1.475 $X2=0 $Y2=0
cc_2969 N_A_3135_265#_c_3399_n VPWR 0.00473731f $X=17.185 $Y=1.475 $X2=0 $Y2=0
cc_2970 N_A_3135_265#_c_3404_n VPWR 0.00593513f $X=18.465 $Y=1.77 $X2=0 $Y2=0
cc_2971 N_A_3135_265#_c_3396_n N_Z_c_9014_n 0.00762343f $X=16.625 $Y=1.4 $X2=0
+ $Y2=0
cc_2972 N_A_3135_265#_c_3400_n N_Z_c_9014_n 0.00704092f $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_2973 N_A_3135_265#_c_3394_n N_Z_c_9057_n 0.00248496f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_2974 N_A_3135_265#_c_3393_n N_Z_c_9060_n 0.00678861f $X=16.155 $Y=1.4 $X2=0
+ $Y2=0
cc_2975 N_A_3135_265#_c_3394_n N_Z_c_9060_n 0.00239476f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_2976 N_A_3135_265#_c_3400_n N_Z_c_9060_n 2.98555e-19 $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_2977 N_A_3135_265#_c_3396_n N_Z_c_9062_n 0.00145542f $X=16.625 $Y=1.4 $X2=0
+ $Y2=0
cc_2978 N_A_3135_265#_c_3398_n N_Z_c_9062_n 0.00597584f $X=17.095 $Y=1.4 $X2=0
+ $Y2=0
cc_2979 N_A_3135_265#_c_3401_n N_Z_c_9062_n 0.00909323f $X=16.715 $Y=1.4 $X2=0
+ $Y2=0
cc_2980 N_A_3135_265#_c_3385_n N_Z_c_9062_n 0.0266078f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_2981 N_A_3135_265#_c_3391_n N_Z_c_9062_n 0.00747617f $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_2982 N_A_3135_265#_c_3392_n N_Z_c_9117_n 0.00834829f $X=15.775 $Y=1.475 $X2=0
+ $Y2=0
cc_2983 N_A_3135_265#_c_3399_n N_Z_c_9119_n 0.00795576f $X=17.185 $Y=1.475 $X2=0
+ $Y2=0
cc_2984 N_A_3135_265#_c_3385_n N_Z_c_9119_n 0.0186685f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_2985 N_A_3135_265#_c_3404_n N_Z_c_9119_n 0.0329704f $X=18.465 $Y=1.77 $X2=0
+ $Y2=0
cc_2986 N_A_3135_265#_c_3391_n N_Z_c_9119_n 2.19754e-19 $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_2987 N_A_3135_265#_c_3395_n Z 0.00372458f $X=16.245 $Y=1.475 $X2=0 $Y2=0
cc_2988 N_A_3135_265#_c_3397_n Z 0.00372248f $X=16.715 $Y=1.475 $X2=0 $Y2=0
cc_2989 N_A_3135_265#_c_3392_n N_Z_c_9135_n 0.0199111f $X=15.775 $Y=1.475 $X2=0
+ $Y2=0
cc_2990 N_A_3135_265#_c_3393_n N_Z_c_9135_n 0.00560592f $X=16.155 $Y=1.4 $X2=0
+ $Y2=0
cc_2991 N_A_3135_265#_c_3394_n N_Z_c_9135_n 0.00474497f $X=15.865 $Y=1.4 $X2=0
+ $Y2=0
cc_2992 N_A_3135_265#_c_3395_n N_Z_c_9135_n 0.0181262f $X=16.245 $Y=1.475 $X2=0
+ $Y2=0
cc_2993 N_A_3135_265#_c_3397_n N_Z_c_9135_n 9.74366e-19 $X=16.715 $Y=1.475 $X2=0
+ $Y2=0
cc_2994 N_A_3135_265#_c_3400_n N_Z_c_9135_n 0.00415268f $X=16.245 $Y=1.4 $X2=0
+ $Y2=0
cc_2995 N_A_3135_265#_c_3395_n N_Z_c_9136_n 9.74366e-19 $X=16.245 $Y=1.475 $X2=0
+ $Y2=0
cc_2996 N_A_3135_265#_c_3397_n N_Z_c_9136_n 0.0181262f $X=16.715 $Y=1.475 $X2=0
+ $Y2=0
cc_2997 N_A_3135_265#_c_3398_n N_Z_c_9136_n 0.00560592f $X=17.095 $Y=1.4 $X2=0
+ $Y2=0
cc_2998 N_A_3135_265#_c_3399_n N_Z_c_9136_n 0.0221748f $X=17.185 $Y=1.475 $X2=0
+ $Y2=0
cc_2999 N_A_3135_265#_c_3401_n N_Z_c_9136_n 0.00181273f $X=16.715 $Y=1.4 $X2=0
+ $Y2=0
cc_3000 N_A_3135_265#_c_3385_n N_Z_c_9136_n 0.00240108f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_3001 N_A_3135_265#_c_3391_n N_Z_c_9136_n 0.00425035f $X=17.505 $Y=1.23 $X2=0
+ $Y2=0
cc_3002 N_A_3135_265#_c_3392_n N_A_2693_297#_c_11159_n 0.00151141f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_3003 N_A_3135_265#_c_3392_n N_A_2693_297#_c_11188_n 0.00307958f $X=15.775
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_3004 N_A_3135_265#_c_3395_n N_A_2693_297#_c_11188_n 0.00307958f $X=16.245
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_3005 N_A_3135_265#_c_3397_n N_A_2693_297#_c_11190_n 0.00307958f $X=16.715
+ $Y=1.475 $X2=0 $Y2=0
cc_3006 N_A_3135_265#_c_3399_n N_A_2693_297#_c_11190_n 0.00307958f $X=17.185
+ $Y=1.475 $X2=0 $Y2=0
cc_3007 N_A_3135_265#_c_3392_n N_A_2693_297#_c_11161_n 0.00554566f $X=15.775
+ $Y=1.475 $X2=0 $Y2=0
cc_3008 N_A_3135_265#_c_3395_n N_A_2693_297#_c_11162_n 0.00210632f $X=16.245
+ $Y=1.475 $X2=0 $Y2=0
cc_3009 N_A_3135_265#_c_3396_n N_A_2693_297#_c_11162_n 0.00251792f $X=16.625
+ $Y=1.4 $X2=0 $Y2=0
cc_3010 N_A_3135_265#_c_3397_n N_A_2693_297#_c_11162_n 0.00210632f $X=16.715
+ $Y=1.475 $X2=0 $Y2=0
cc_3011 N_A_3135_265#_c_3399_n N_A_2693_297#_c_11163_n 0.00499839f $X=17.185
+ $Y=1.475 $X2=0 $Y2=0
cc_3012 N_A_3135_265#_c_3385_n N_A_2693_297#_c_11163_n 0.0218124f $X=18.3
+ $Y=1.23 $X2=0 $Y2=0
cc_3013 N_A_3135_265#_c_3386_n N_A_2693_297#_c_11163_n 5.74251e-19 $X=17.755
+ $Y=1.23 $X2=0 $Y2=0
cc_3014 N_A_3135_265#_c_3391_n N_A_2693_297#_c_11163_n 0.00561627f $X=17.505
+ $Y=1.23 $X2=0 $Y2=0
cc_3015 N_A_3135_265#_c_3385_n N_VGND_c_12723_n 0.0123065f $X=18.3 $Y=1.23 $X2=0
+ $Y2=0
cc_3016 N_A_3135_265#_c_3386_n N_VGND_c_12723_n 2.04129e-19 $X=17.755 $Y=1.23
+ $X2=0 $Y2=0
cc_3017 N_A_3135_265#_c_3387_n N_VGND_c_12811_n 0.0129994f $X=18.465 $Y=0.445
+ $X2=0 $Y2=0
cc_3018 N_A_3135_265#_M1222_s VGND 0.00394793f $X=18.33 $Y=0.235 $X2=0 $Y2=0
cc_3019 N_A_3135_265#_c_3387_n VGND 0.00927134f $X=18.465 $Y=0.445 $X2=0 $Y2=0
cc_3020 N_A_3135_265#_c_3400_n N_A_2695_47#_c_14405_n 7.0477e-19 $X=16.245
+ $Y=1.4 $X2=0 $Y2=0
cc_3021 N_A_3135_265#_c_3385_n N_A_2695_47#_c_14383_n 0.0028695f $X=18.3 $Y=1.23
+ $X2=25.99 $Y2=4.93
cc_3022 N_A_3135_265#_c_3391_n N_A_2695_47#_c_14383_n 0.00589316f $X=17.505
+ $Y=1.23 $X2=25.99 $Y2=4.93
cc_3023 N_A_3135_793#_c_3513_n N_S[10]_c_3746_n 0.00507426f $X=15.865 $Y=4.04
+ $X2=0 $Y2=0
cc_3024 N_A_3135_793#_c_3512_n N_S[10]_c_3749_n 0.00509391f $X=16.155 $Y=4.04
+ $X2=0 $Y2=0
cc_3025 N_A_3135_793#_c_3515_n N_S[10]_c_3751_n 0.00509204f $X=16.625 $Y=4.04
+ $X2=25.905 $Y2=4.845
cc_3026 N_A_3135_793#_c_3517_n N_S[10]_c_3753_n 0.00507688f $X=17.095 $Y=4.04
+ $X2=0 $Y2=0
cc_3027 N_A_3135_793#_c_3506_n N_S[10]_c_3755_n 6.53442e-19 $X=18.425 $Y=4.74
+ $X2=0 $Y2=0
cc_3028 N_A_3135_793#_c_3504_n N_S[10]_c_3757_n 0.0103812f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3029 N_A_3135_793#_c_3505_n N_S[10]_c_3757_n 0.0179529f $X=17.755 $Y=4.21
+ $X2=0 $Y2=0
cc_3030 N_A_3135_793#_c_3524_n N_S[10]_c_3767_n 0.00508008f $X=18.385 $Y=4.045
+ $X2=0 $Y2=0
cc_3031 N_A_3135_793#_c_3510_n N_S[10]_c_3767_n 0.00262132f $X=17.505 $Y=4.21
+ $X2=0 $Y2=0
cc_3032 N_A_3135_793#_c_3504_n N_S[10]_c_3758_n 0.0206368f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3033 N_A_3135_793#_c_3505_n N_S[10]_c_3758_n 0.0175393f $X=17.755 $Y=4.21
+ $X2=0 $Y2=0
cc_3034 N_A_3135_793#_c_3524_n N_S[10]_c_3758_n 0.00255921f $X=18.385 $Y=4.045
+ $X2=0 $Y2=0
cc_3035 N_A_3135_793#_c_3508_n N_S[10]_c_3758_n 0.00322131f $X=18.385 $Y=4.21
+ $X2=0 $Y2=0
cc_3036 N_A_3135_793#_c_3509_n N_S[10]_c_3758_n 0.0085951f $X=18.425 $Y=4.615
+ $X2=0 $Y2=0
cc_3037 N_A_3135_793#_c_3523_n N_S[10]_c_3769_n 0.00970559f $X=18.465 $Y=3.14
+ $X2=0 $Y2=0
cc_3038 N_A_3135_793#_c_3524_n N_S[10]_c_3769_n 0.00254107f $X=18.385 $Y=4.045
+ $X2=0 $Y2=0
cc_3039 N_A_3135_793#_c_3525_n N_S[10]_c_3769_n 0.00216424f $X=18.465 $Y=3.835
+ $X2=0 $Y2=0
cc_3040 N_A_3135_793#_c_3506_n N_S[10]_c_3759_n 9.67113e-19 $X=18.425 $Y=4.74
+ $X2=0 $Y2=0
cc_3041 N_A_3135_793#_c_3507_n N_S[10]_c_3759_n 0.00603996f $X=18.465 $Y=4.995
+ $X2=0 $Y2=0
cc_3042 N_A_3135_793#_c_3506_n N_S[10]_c_3760_n 0.0111895f $X=18.425 $Y=4.74
+ $X2=0 $Y2=0
cc_3043 N_A_3135_793#_c_3509_n N_S[10]_c_3760_n 0.00429801f $X=18.425 $Y=4.615
+ $X2=0 $Y2=0
cc_3044 N_A_3135_793#_c_3524_n N_S[10]_c_3761_n 0.00336772f $X=18.385 $Y=4.045
+ $X2=0 $Y2=0
cc_3045 N_A_3135_793#_c_3506_n N_S[10]_c_3761_n 0.00207203f $X=18.425 $Y=4.74
+ $X2=0 $Y2=0
cc_3046 N_A_3135_793#_c_3525_n N_S[10]_c_3761_n 5.48523e-19 $X=18.465 $Y=3.835
+ $X2=0 $Y2=0
cc_3047 N_A_3135_793#_c_3508_n N_S[10]_c_3761_n 0.00416423f $X=18.385 $Y=4.21
+ $X2=0 $Y2=0
cc_3048 N_A_3135_793#_c_3509_n N_S[10]_c_3761_n 0.00289358f $X=18.425 $Y=4.615
+ $X2=0 $Y2=0
cc_3049 N_A_3135_793#_c_3523_n N_S[10]_c_3771_n 0.00929139f $X=18.465 $Y=3.14
+ $X2=25.99 $Y2=4.8
cc_3050 N_A_3135_793#_c_3524_n N_S[10]_c_3771_n 0.00117303f $X=18.385 $Y=4.045
+ $X2=25.99 $Y2=4.8
cc_3051 N_A_3135_793#_c_3525_n N_S[10]_c_3771_n 0.00304348f $X=18.465 $Y=3.835
+ $X2=25.99 $Y2=4.8
cc_3052 N_A_3135_793#_c_3506_n N_S[10]_c_3765_n 0.00426435f $X=18.425 $Y=4.74
+ $X2=0 $Y2=0
cc_3053 N_A_3135_793#_c_3509_n N_S[10]_c_3765_n 0.00268644f $X=18.425 $Y=4.615
+ $X2=0 $Y2=0
cc_3054 N_A_3135_793#_c_3508_n S[10] 0.0228692f $X=18.385 $Y=4.21 $X2=0 $Y2=0
cc_3055 N_A_3135_793#_c_3509_n S[10] 0.00541767f $X=18.425 $Y=4.615 $X2=0 $Y2=0
cc_3056 N_A_3135_793#_c_3511_n N_VPWR_c_7246_n 0.00324472f $X=15.775 $Y=3.965
+ $X2=0 $Y2=0
cc_3057 N_A_3135_793#_c_3518_n N_VPWR_c_7248_n 0.00367058f $X=17.185 $Y=3.965
+ $X2=0 $Y2=0
cc_3058 N_A_3135_793#_c_3504_n N_VPWR_c_7248_n 0.0193185f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3059 N_A_3135_793#_c_3505_n N_VPWR_c_7248_n 6.4101e-19 $X=17.755 $Y=4.21
+ $X2=0 $Y2=0
cc_3060 N_A_3135_793#_c_3523_n N_VPWR_c_7248_n 0.0316788f $X=18.465 $Y=3.14
+ $X2=0 $Y2=0
cc_3061 N_A_3135_793#_c_3523_n N_VPWR_c_7250_n 0.0356181f $X=18.465 $Y=3.14
+ $X2=0 $Y2=0
cc_3062 N_A_3135_793#_c_3523_n N_VPWR_c_7322_n 0.0233824f $X=18.465 $Y=3.14
+ $X2=0 $Y2=0
cc_3063 N_A_3135_793#_c_3511_n VPWR 0.00473731f $X=15.775 $Y=3.965 $X2=0 $Y2=0
cc_3064 N_A_3135_793#_c_3514_n VPWR 0.00362156f $X=16.245 $Y=3.965 $X2=0 $Y2=0
cc_3065 N_A_3135_793#_c_3516_n VPWR 0.00362156f $X=16.715 $Y=3.965 $X2=0 $Y2=0
cc_3066 N_A_3135_793#_c_3518_n VPWR 0.00473731f $X=17.185 $Y=3.965 $X2=0 $Y2=0
cc_3067 N_A_3135_793#_c_3523_n VPWR 0.00593513f $X=18.465 $Y=3.14 $X2=0 $Y2=0
cc_3068 N_A_3135_793#_c_3515_n N_Z_c_9015_n 0.00762343f $X=16.625 $Y=4.04 $X2=0
+ $Y2=0
cc_3069 N_A_3135_793#_c_3519_n N_Z_c_9015_n 0.00704092f $X=16.245 $Y=4.04 $X2=0
+ $Y2=0
cc_3070 N_A_3135_793#_c_3513_n N_Z_c_9058_n 0.00248496f $X=15.865 $Y=4.04 $X2=0
+ $Y2=0
cc_3071 N_A_3135_793#_c_3512_n N_Z_c_9061_n 0.00678861f $X=16.155 $Y=4.04 $X2=0
+ $Y2=0
cc_3072 N_A_3135_793#_c_3513_n N_Z_c_9061_n 0.00239476f $X=15.865 $Y=4.04 $X2=0
+ $Y2=0
cc_3073 N_A_3135_793#_c_3519_n N_Z_c_9061_n 2.98555e-19 $X=16.245 $Y=4.04 $X2=0
+ $Y2=0
cc_3074 N_A_3135_793#_c_3515_n N_Z_c_9063_n 0.00145542f $X=16.625 $Y=4.04 $X2=0
+ $Y2=0
cc_3075 N_A_3135_793#_c_3517_n N_Z_c_9063_n 0.00597584f $X=17.095 $Y=4.04 $X2=0
+ $Y2=0
cc_3076 N_A_3135_793#_c_3520_n N_Z_c_9063_n 0.00909323f $X=16.715 $Y=4.04 $X2=0
+ $Y2=0
cc_3077 N_A_3135_793#_c_3504_n N_Z_c_9063_n 0.0266078f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3078 N_A_3135_793#_c_3510_n N_Z_c_9063_n 0.00747617f $X=17.505 $Y=4.21 $X2=0
+ $Y2=0
cc_3079 N_A_3135_793#_c_3511_n N_Z_c_9118_n 0.00834829f $X=15.775 $Y=3.965 $X2=0
+ $Y2=0
cc_3080 N_A_3135_793#_c_3518_n N_Z_c_9120_n 0.00795576f $X=17.185 $Y=3.965 $X2=0
+ $Y2=0
cc_3081 N_A_3135_793#_c_3504_n N_Z_c_9120_n 0.0186685f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3082 N_A_3135_793#_c_3523_n N_Z_c_9120_n 0.0329704f $X=18.465 $Y=3.14 $X2=0
+ $Y2=0
cc_3083 N_A_3135_793#_c_3510_n N_Z_c_9120_n 2.19754e-19 $X=17.505 $Y=4.21 $X2=0
+ $Y2=0
cc_3084 N_A_3135_793#_c_3514_n Z 0.00372458f $X=16.245 $Y=3.965 $X2=0 $Y2=0
cc_3085 N_A_3135_793#_c_3516_n Z 0.00372248f $X=16.715 $Y=3.965 $X2=0 $Y2=0
cc_3086 N_A_3135_793#_c_3511_n N_Z_c_9135_n 0.0199111f $X=15.775 $Y=3.965 $X2=0
+ $Y2=0
cc_3087 N_A_3135_793#_c_3512_n N_Z_c_9135_n 0.00560592f $X=16.155 $Y=4.04 $X2=0
+ $Y2=0
cc_3088 N_A_3135_793#_c_3513_n N_Z_c_9135_n 0.00474497f $X=15.865 $Y=4.04 $X2=0
+ $Y2=0
cc_3089 N_A_3135_793#_c_3514_n N_Z_c_9135_n 0.0181262f $X=16.245 $Y=3.965 $X2=0
+ $Y2=0
cc_3090 N_A_3135_793#_c_3516_n N_Z_c_9135_n 9.74366e-19 $X=16.715 $Y=3.965 $X2=0
+ $Y2=0
cc_3091 N_A_3135_793#_c_3519_n N_Z_c_9135_n 0.00415268f $X=16.245 $Y=4.04 $X2=0
+ $Y2=0
cc_3092 N_A_3135_793#_c_3514_n N_Z_c_9136_n 9.74366e-19 $X=16.245 $Y=3.965 $X2=0
+ $Y2=0
cc_3093 N_A_3135_793#_c_3516_n N_Z_c_9136_n 0.0181262f $X=16.715 $Y=3.965 $X2=0
+ $Y2=0
cc_3094 N_A_3135_793#_c_3517_n N_Z_c_9136_n 0.00560592f $X=17.095 $Y=4.04 $X2=0
+ $Y2=0
cc_3095 N_A_3135_793#_c_3518_n N_Z_c_9136_n 0.0221748f $X=17.185 $Y=3.965 $X2=0
+ $Y2=0
cc_3096 N_A_3135_793#_c_3520_n N_Z_c_9136_n 0.00181273f $X=16.715 $Y=4.04 $X2=0
+ $Y2=0
cc_3097 N_A_3135_793#_c_3504_n N_Z_c_9136_n 0.00240108f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3098 N_A_3135_793#_c_3510_n N_Z_c_9136_n 0.00425035f $X=17.505 $Y=4.21 $X2=0
+ $Y2=0
cc_3099 N_A_3135_793#_c_3511_n N_A_2693_591#_c_11287_n 0.00151141f $X=15.775
+ $Y=3.965 $X2=0 $Y2=0
cc_3100 N_A_3135_793#_c_3511_n N_A_2693_591#_c_11316_n 0.00307958f $X=15.775
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_3101 N_A_3135_793#_c_3514_n N_A_2693_591#_c_11316_n 0.00307958f $X=16.245
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_3102 N_A_3135_793#_c_3516_n N_A_2693_591#_c_11318_n 0.00307958f $X=16.715
+ $Y=3.965 $X2=0 $Y2=0
cc_3103 N_A_3135_793#_c_3518_n N_A_2693_591#_c_11318_n 0.00307958f $X=17.185
+ $Y=3.965 $X2=0 $Y2=0
cc_3104 N_A_3135_793#_c_3511_n N_A_2693_591#_c_11289_n 0.00554566f $X=15.775
+ $Y=3.965 $X2=0 $Y2=0
cc_3105 N_A_3135_793#_c_3514_n N_A_2693_591#_c_11290_n 0.00210632f $X=16.245
+ $Y=3.965 $X2=0 $Y2=0
cc_3106 N_A_3135_793#_c_3515_n N_A_2693_591#_c_11290_n 0.00251792f $X=16.625
+ $Y=4.04 $X2=0 $Y2=0
cc_3107 N_A_3135_793#_c_3516_n N_A_2693_591#_c_11290_n 0.00210632f $X=16.715
+ $Y=3.965 $X2=0 $Y2=0
cc_3108 N_A_3135_793#_c_3518_n N_A_2693_591#_c_11291_n 0.00499839f $X=17.185
+ $Y=3.965 $X2=0 $Y2=0
cc_3109 N_A_3135_793#_c_3504_n N_A_2693_591#_c_11291_n 0.0218124f $X=18.3
+ $Y=4.21 $X2=0 $Y2=0
cc_3110 N_A_3135_793#_c_3505_n N_A_2693_591#_c_11291_n 5.74251e-19 $X=17.755
+ $Y=4.21 $X2=0 $Y2=0
cc_3111 N_A_3135_793#_c_3510_n N_A_2693_591#_c_11291_n 0.00561627f $X=17.505
+ $Y=4.21 $X2=0 $Y2=0
cc_3112 N_A_3135_793#_c_3504_n N_VGND_c_12724_n 0.0123065f $X=18.3 $Y=4.21 $X2=0
+ $Y2=0
cc_3113 N_A_3135_793#_c_3505_n N_VGND_c_12724_n 2.04129e-19 $X=17.755 $Y=4.21
+ $X2=0 $Y2=0
cc_3114 N_A_3135_793#_c_3507_n N_VGND_c_12813_n 0.0129994f $X=18.465 $Y=4.995
+ $X2=0 $Y2=0
cc_3115 N_A_3135_793#_M1043_d VGND 0.00394793f $X=18.33 $Y=4.785 $X2=0 $Y2=0
cc_3116 N_A_3135_793#_c_3507_n VGND 0.00927134f $X=18.465 $Y=4.995 $X2=0 $Y2=0
cc_3117 N_A_3135_793#_c_3519_n N_A_2695_911#_c_14484_n 7.0477e-19 $X=16.245
+ $Y=4.04 $X2=0 $Y2=0
cc_3118 N_A_3135_793#_c_3504_n N_A_2695_911#_c_14465_n 0.0028695f $X=18.3
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_3119 N_A_3135_793#_c_3510_n N_A_2695_911#_c_14465_n 0.00589316f $X=17.505
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_3120 N_S[2]_c_3652_n N_S[10]_c_3769_n 0.0130744f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_3121 N_S[2]_c_3645_n N_S[10]_c_3771_n 0.0130744f $X=18.7 $Y=1.55 $X2=25.99
+ $Y2=4.8
cc_3122 N_S[2]_c_3645_n N_S[3]_c_3871_n 0.0215827f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3123 S[2] N_S[3]_c_3871_n 0.00113563f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_3124 N_S[2]_c_3645_n N_S[3]_c_3892_n 0.00113563f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3125 S[2] N_S[3]_c_3892_n 0.0301108f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_3126 N_S[2]_c_3652_n N_VPWR_c_7247_n 0.00950399f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_3127 N_S[2]_c_3645_n N_VPWR_c_7249_n 0.016386f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3128 S[2] N_VPWR_c_7249_n 0.0157609f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_3129 N_S[2]_c_3652_n N_VPWR_c_7322_n 0.0035837f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_3130 N_S[2]_c_3645_n N_VPWR_c_7322_n 0.0035837f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3131 N_S[2]_c_3652_n VPWR 0.00711603f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_3132 N_S[2]_c_3645_n VPWR 0.0070533f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3133 N_S[2]_c_3629_n N_Z_c_9013_n 0.002324f $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_3134 N_S[2]_c_3632_n N_Z_c_9013_n 0.00283489f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_3135 N_S[2]_c_3632_n N_Z_c_9014_n 3.10191e-19 $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_3136 N_S[2]_c_3634_n N_Z_c_9014_n 0.00190704f $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_3137 N_S[2]_c_3632_n N_Z_c_9016_n 6.35774e-19 $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_3138 N_S[2]_c_3634_n N_Z_c_9016_n 0.0077801f $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_3139 N_S[2]_c_3636_n N_Z_c_9016_n 0.0134253f $X=16.96 $Y=0.255 $X2=0 $Y2=0
cc_3140 N_S[2]_c_3629_n N_Z_c_9057_n 0.00443615f $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_3141 N_S[2]_c_3632_n N_Z_c_9057_n 0.00462308f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_3142 N_S[2]_c_3634_n N_Z_c_9057_n 6.35664e-19 $X=16.54 $Y=0.255 $X2=0 $Y2=0
cc_3143 N_S[2]_c_3632_n N_Z_c_9060_n 0.00180363f $X=16.12 $Y=0.255 $X2=0 $Y2=0
cc_3144 N_S[2]_c_3636_n N_Z_c_9062_n 0.00216436f $X=16.96 $Y=0.255 $X2=0 $Y2=0
cc_3145 N_S[2]_c_3652_n N_Z_c_9119_n 0.00478771f $X=18.23 $Y=1.55 $X2=0 $Y2=0
cc_3146 N_S[2]_c_3645_n N_Z_c_9119_n 0.00760321f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3147 S[2] N_Z_c_9119_n 0.010609f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_3148 N_S[2]_c_3629_n N_A_2693_297#_c_11159_n 0.00168571f $X=15.7 $Y=0.255
+ $X2=0 $Y2=0
cc_3149 N_S[2]_c_3652_n N_A_2693_297#_c_11163_n 0.00239129f $X=18.23 $Y=1.55
+ $X2=0 $Y2=0
cc_3150 N_S[2]_c_3629_n N_VGND_c_12721_n 5.5039e-19 $X=15.7 $Y=0.255 $X2=0 $Y2=0
cc_3151 N_S[2]_c_3631_n N_VGND_c_12721_n 0.0028166f $X=15.775 $Y=0.18 $X2=0
+ $Y2=0
cc_3152 N_S[2]_c_3637_n N_VGND_c_12723_n 0.00862298f $X=17.645 $Y=0.18 $X2=0
+ $Y2=0
cc_3153 N_S[2]_c_3639_n N_VGND_c_12723_n 0.00525833f $X=18.13 $Y=0.81 $X2=0
+ $Y2=0
cc_3154 N_S[2]_c_3642_n N_VGND_c_12723_n 0.00173127f $X=18.255 $Y=0.735 $X2=0
+ $Y2=0
cc_3155 N_S[2]_c_3644_n N_VGND_c_12725_n 0.00374526f $X=18.675 $Y=0.735 $X2=0
+ $Y2=0
cc_3156 N_S[2]_c_3645_n N_VGND_c_12725_n 0.00578076f $X=18.7 $Y=1.55 $X2=0 $Y2=0
cc_3157 S[2] N_VGND_c_12725_n 0.0116413f $X=19.005 $Y=1.105 $X2=0 $Y2=0
cc_3158 N_S[2]_c_3631_n N_VGND_c_12807_n 0.0559651f $X=15.775 $Y=0.18 $X2=0
+ $Y2=0
cc_3159 N_S[2]_c_3642_n N_VGND_c_12811_n 0.00542362f $X=18.255 $Y=0.735 $X2=0
+ $Y2=0
cc_3160 N_S[2]_c_3643_n N_VGND_c_12811_n 2.16067e-19 $X=18.6 $Y=0.81 $X2=0 $Y2=0
cc_3161 N_S[2]_c_3644_n N_VGND_c_12811_n 0.00585385f $X=18.675 $Y=0.735 $X2=0
+ $Y2=0
cc_3162 N_S[2]_c_3630_n VGND 0.00642387f $X=16.045 $Y=0.18 $X2=0 $Y2=0
cc_3163 N_S[2]_c_3631_n VGND 0.00591981f $X=15.775 $Y=0.18 $X2=0 $Y2=0
cc_3164 N_S[2]_c_3633_n VGND 0.0064237f $X=16.465 $Y=0.18 $X2=0 $Y2=0
cc_3165 N_S[2]_c_3635_n VGND 0.00642387f $X=16.885 $Y=0.18 $X2=0 $Y2=0
cc_3166 N_S[2]_c_3637_n VGND 0.0345801f $X=17.645 $Y=0.18 $X2=0 $Y2=0
cc_3167 N_S[2]_c_3642_n VGND 0.00990284f $X=18.255 $Y=0.735 $X2=0 $Y2=0
cc_3168 N_S[2]_c_3644_n VGND 0.0119653f $X=18.675 $Y=0.735 $X2=0 $Y2=0
cc_3169 N_S[2]_c_3646_n VGND 0.00366655f $X=16.12 $Y=0.18 $X2=0 $Y2=0
cc_3170 N_S[2]_c_3647_n VGND 0.00366655f $X=16.54 $Y=0.18 $X2=0 $Y2=0
cc_3171 N_S[2]_c_3648_n VGND 0.00366655f $X=16.96 $Y=0.18 $X2=0 $Y2=0
cc_3172 N_S[2]_c_3629_n N_A_2695_47#_c_14378_n 0.00206084f $X=15.7 $Y=0.255
+ $X2=0 $Y2=0
cc_3173 N_S[2]_c_3629_n N_A_2695_47#_c_14380_n 0.0139014f $X=15.7 $Y=0.255 $X2=0
+ $Y2=0
cc_3174 N_S[2]_c_3630_n N_A_2695_47#_c_14380_n 0.00211351f $X=16.045 $Y=0.18
+ $X2=0 $Y2=0
cc_3175 N_S[2]_c_3632_n N_A_2695_47#_c_14380_n 0.0106826f $X=16.12 $Y=0.255
+ $X2=0 $Y2=0
cc_3176 N_S[2]_c_3634_n N_A_2695_47#_c_14382_n 0.0106844f $X=16.54 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_3177 N_S[2]_c_3635_n N_A_2695_47#_c_14382_n 0.00211351f $X=16.885 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_3178 N_S[2]_c_3636_n N_A_2695_47#_c_14382_n 0.0112916f $X=16.96 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_3179 N_S[2]_c_3637_n N_A_2695_47#_c_14382_n 0.00685838f $X=17.645 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_3180 N_S[2]_c_3638_n N_A_2695_47#_c_14382_n 0.00189496f $X=17.72 $Y=0.735
+ $X2=25.99 $Y2=4.8
cc_3181 N_S[2]_c_3638_n N_A_2695_47#_c_14383_n 0.00529837f $X=17.72 $Y=0.735
+ $X2=25.99 $Y2=4.93
cc_3182 N_S[2]_c_3633_n N_A_2695_47#_c_14418_n 0.0034777f $X=16.465 $Y=0.18
+ $X2=0 $Y2=0
cc_3183 N_S[10]_c_3761_n N_S[11]_c_3991_n 0.0215827f $X=18.675 $Y=4.705 $X2=0
+ $Y2=0
cc_3184 S[10] N_S[11]_c_3991_n 0.00113563f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_3185 N_S[10]_c_3761_n N_S[11]_c_4011_n 0.00113563f $X=18.675 $Y=4.705 $X2=0
+ $Y2=0
cc_3186 S[10] N_S[11]_c_4011_n 0.0301108f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_3187 N_S[10]_c_3769_n N_VPWR_c_7248_n 0.00950399f $X=18.23 $Y=3.89 $X2=0
+ $Y2=0
cc_3188 N_S[10]_c_3761_n N_VPWR_c_7250_n 0.00652399f $X=18.675 $Y=4.705 $X2=0
+ $Y2=0
cc_3189 N_S[10]_c_3771_n N_VPWR_c_7250_n 0.00986205f $X=18.7 $Y=3.89 $X2=0 $Y2=0
cc_3190 S[10] N_VPWR_c_7250_n 0.0157609f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_3191 N_S[10]_c_3769_n N_VPWR_c_7322_n 0.0035837f $X=18.23 $Y=3.89 $X2=0 $Y2=0
cc_3192 N_S[10]_c_3771_n N_VPWR_c_7322_n 0.0035837f $X=18.7 $Y=3.89 $X2=0 $Y2=0
cc_3193 N_S[10]_c_3769_n VPWR 0.00711603f $X=18.23 $Y=3.89 $X2=0 $Y2=0
cc_3194 N_S[10]_c_3771_n VPWR 0.0070533f $X=18.7 $Y=3.89 $X2=0 $Y2=0
cc_3195 N_S[10]_c_3749_n N_Z_c_9015_n 3.10191e-19 $X=16.12 $Y=5.185 $X2=0 $Y2=0
cc_3196 N_S[10]_c_3751_n N_Z_c_9015_n 0.00190704f $X=16.54 $Y=5.185 $X2=0 $Y2=0
cc_3197 N_S[10]_c_3749_n N_Z_c_9017_n 6.35774e-19 $X=16.12 $Y=5.185 $X2=0 $Y2=0
cc_3198 N_S[10]_c_3751_n N_Z_c_9017_n 0.0077801f $X=16.54 $Y=5.185 $X2=0 $Y2=0
cc_3199 N_S[10]_c_3753_n N_Z_c_9017_n 0.0134253f $X=16.96 $Y=5.185 $X2=0 $Y2=0
cc_3200 N_S[10]_c_3746_n N_Z_c_9058_n 0.00443615f $X=15.7 $Y=5.185 $X2=0 $Y2=0
cc_3201 N_S[10]_c_3749_n N_Z_c_9058_n 0.00462308f $X=16.12 $Y=5.185 $X2=0 $Y2=0
cc_3202 N_S[10]_c_3746_n N_Z_c_9059_n 0.002324f $X=15.7 $Y=5.185 $X2=0 $Y2=0
cc_3203 N_S[10]_c_3749_n N_Z_c_9059_n 0.00283489f $X=16.12 $Y=5.185 $X2=0 $Y2=0
cc_3204 N_S[10]_c_3751_n N_Z_c_9059_n 6.35664e-19 $X=16.54 $Y=5.185 $X2=0 $Y2=0
cc_3205 N_S[10]_c_3749_n N_Z_c_9061_n 0.00180363f $X=16.12 $Y=5.185 $X2=0 $Y2=0
cc_3206 N_S[10]_c_3753_n N_Z_c_9063_n 0.00216436f $X=16.96 $Y=5.185 $X2=0 $Y2=0
cc_3207 N_S[10]_c_3767_n N_Z_c_9120_n 2.55735e-19 $X=18.23 $Y=3.99 $X2=0 $Y2=0
cc_3208 N_S[10]_c_3769_n N_Z_c_9120_n 0.00453198f $X=18.23 $Y=3.89 $X2=0 $Y2=0
cc_3209 N_S[10]_c_3761_n N_Z_c_9120_n 0.00258545f $X=18.675 $Y=4.705 $X2=0 $Y2=0
cc_3210 N_S[10]_c_3771_n N_Z_c_9120_n 0.00501777f $X=18.7 $Y=3.89 $X2=0 $Y2=0
cc_3211 S[10] N_Z_c_9120_n 0.010609f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_3212 N_S[10]_c_3746_n N_A_2693_591#_c_11287_n 0.00168571f $X=15.7 $Y=5.185
+ $X2=0 $Y2=0
cc_3213 N_S[10]_c_3769_n N_A_2693_591#_c_11291_n 0.00239129f $X=18.23 $Y=3.89
+ $X2=0 $Y2=0
cc_3214 N_S[10]_c_3746_n N_VGND_c_12722_n 5.5039e-19 $X=15.7 $Y=5.185 $X2=0
+ $Y2=0
cc_3215 N_S[10]_c_3748_n N_VGND_c_12722_n 0.0028166f $X=15.775 $Y=5.26 $X2=0
+ $Y2=0
cc_3216 N_S[10]_c_3755_n N_VGND_c_12724_n 0.00862298f $X=17.72 $Y=5.185 $X2=0
+ $Y2=0
cc_3217 N_S[10]_c_3756_n N_VGND_c_12724_n 0.00525833f $X=18.13 $Y=4.63 $X2=0
+ $Y2=0
cc_3218 N_S[10]_c_3759_n N_VGND_c_12724_n 0.00173127f $X=18.255 $Y=4.705 $X2=0
+ $Y2=0
cc_3219 N_S[10]_c_3761_n N_VGND_c_12726_n 0.00952602f $X=18.675 $Y=4.705 $X2=0
+ $Y2=0
cc_3220 S[10] N_VGND_c_12726_n 0.0116413f $X=19.005 $Y=4.165 $X2=0 $Y2=0
cc_3221 N_S[10]_c_3748_n N_VGND_c_12809_n 0.0559651f $X=15.775 $Y=5.26 $X2=0
+ $Y2=0
cc_3222 N_S[10]_c_3759_n N_VGND_c_12813_n 0.00542362f $X=18.255 $Y=4.705 $X2=0
+ $Y2=0
cc_3223 N_S[10]_c_3760_n N_VGND_c_12813_n 2.16067e-19 $X=18.6 $Y=4.63 $X2=0
+ $Y2=0
cc_3224 N_S[10]_c_3761_n N_VGND_c_12813_n 0.00585385f $X=18.675 $Y=4.705 $X2=0
+ $Y2=0
cc_3225 N_S[10]_c_3747_n VGND 0.00642387f $X=16.045 $Y=5.26 $X2=0 $Y2=0
cc_3226 N_S[10]_c_3748_n VGND 0.00591981f $X=15.775 $Y=5.26 $X2=0 $Y2=0
cc_3227 N_S[10]_c_3750_n VGND 0.0064237f $X=16.465 $Y=5.26 $X2=0 $Y2=0
cc_3228 N_S[10]_c_3752_n VGND 0.00642387f $X=16.885 $Y=5.26 $X2=0 $Y2=0
cc_3229 N_S[10]_c_3754_n VGND 0.0345801f $X=17.645 $Y=5.26 $X2=0 $Y2=0
cc_3230 N_S[10]_c_3759_n VGND 0.00990284f $X=18.255 $Y=4.705 $X2=0 $Y2=0
cc_3231 N_S[10]_c_3761_n VGND 0.0119653f $X=18.675 $Y=4.705 $X2=0 $Y2=0
cc_3232 N_S[10]_c_3762_n VGND 0.00366655f $X=16.12 $Y=5.26 $X2=0 $Y2=0
cc_3233 N_S[10]_c_3763_n VGND 0.00366655f $X=16.54 $Y=5.26 $X2=0 $Y2=0
cc_3234 N_S[10]_c_3764_n VGND 0.00366655f $X=16.96 $Y=5.26 $X2=0 $Y2=0
cc_3235 N_S[10]_c_3746_n N_A_2695_911#_c_14460_n 0.00206084f $X=15.7 $Y=5.185
+ $X2=0 $Y2=0
cc_3236 N_S[10]_c_3746_n N_A_2695_911#_c_14462_n 0.0139014f $X=15.7 $Y=5.185
+ $X2=0 $Y2=0
cc_3237 N_S[10]_c_3747_n N_A_2695_911#_c_14462_n 0.00211351f $X=16.045 $Y=5.26
+ $X2=0 $Y2=0
cc_3238 N_S[10]_c_3749_n N_A_2695_911#_c_14462_n 0.0106826f $X=16.12 $Y=5.185
+ $X2=0 $Y2=0
cc_3239 N_S[10]_c_3751_n N_A_2695_911#_c_14464_n 0.0106844f $X=16.54 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_3240 N_S[10]_c_3752_n N_A_2695_911#_c_14464_n 0.00211351f $X=16.885 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_3241 N_S[10]_c_3753_n N_A_2695_911#_c_14464_n 0.0112916f $X=16.96 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_3242 N_S[10]_c_3754_n N_A_2695_911#_c_14464_n 0.00685838f $X=17.645 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_3243 N_S[10]_c_3755_n N_A_2695_911#_c_14464_n 0.00189496f $X=17.72 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_3244 N_S[10]_c_3757_n N_A_2695_911#_c_14465_n 0.00529837f $X=17.795 $Y=4.63
+ $X2=25.99 $Y2=4.8
cc_3245 N_S[10]_c_3750_n N_A_2695_911#_c_14497_n 0.0034777f $X=16.465 $Y=5.26
+ $X2=0 $Y2=0
cc_3246 N_S[3]_c_3872_n N_S[11]_c_4013_n 0.0130744f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_3247 N_S[3]_c_3896_n N_S[11]_c_4017_n 0.0130744f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_3248 N_S[3]_c_3881_n N_A_4006_325#_c_4127_n 0.00507688f $X=21.68 $Y=0.255
+ $X2=25.905 $Y2=0.425
cc_3249 N_S[3]_c_3876_n N_A_4006_325#_c_4119_n 0.00262132f $X=20.41 $Y=1.45
+ $X2=25.905 $Y2=4.845
cc_3250 N_S[3]_c_3883_n N_A_4006_325#_c_4130_n 0.00509204f $X=22.1 $Y=0.255
+ $X2=0 $Y2=0
cc_3251 N_S[3]_c_3887_n N_A_4006_325#_c_4132_n 0.00507426f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_3252 N_S[3]_c_3885_n N_A_4006_325#_c_4135_n 0.00509391f $X=22.52 $Y=0.255
+ $X2=0 $Y2=0
cc_3253 N_S[3]_c_3872_n N_A_4006_325#_c_4136_n 0.0128834f $X=19.94 $Y=1.55 $X2=0
+ $Y2=0
cc_3254 N_S[3]_c_3896_n N_A_4006_325#_c_4136_n 0.0118698f $X=20.41 $Y=1.55 $X2=0
+ $Y2=0
cc_3255 N_S[3]_c_3873_n N_A_4006_325#_c_4120_n 0.00207203f $X=19.965 $Y=0.735
+ $X2=0 $Y2=0
cc_3256 N_S[3]_c_3875_n N_A_4006_325#_c_4120_n 0.00603996f $X=20.385 $Y=0.735
+ $X2=0 $Y2=0
cc_3257 N_S[3]_c_3878_n N_A_4006_325#_c_4120_n 6.53442e-19 $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_3258 N_S[3]_c_3872_n N_A_4006_325#_c_4121_n 0.00289358f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_3259 N_S[3]_c_3874_n N_A_4006_325#_c_4121_n 0.00429801f $X=20.31 $Y=0.81
+ $X2=0 $Y2=0
cc_3260 N_S[3]_c_3876_n N_A_4006_325#_c_4121_n 0.0085951f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_3261 N_S[3]_c_3888_n N_A_4006_325#_c_4121_n 0.00268644f $X=20.41 $Y=0.81
+ $X2=0 $Y2=0
cc_3262 N_S[3]_c_3892_n N_A_4006_325#_c_4121_n 0.00541767f $X=19.9 $Y=1.16 $X2=0
+ $Y2=0
cc_3263 N_S[3]_c_3876_n N_A_4006_325#_c_4122_n 0.0206368f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_3264 N_S[3]_c_3877_n N_A_4006_325#_c_4122_n 0.0103812f $X=20.845 $Y=0.81
+ $X2=0 $Y2=0
cc_3265 N_S[3]_c_3872_n N_A_4006_325#_c_4138_n 0.00454075f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_3266 N_S[3]_c_3876_n N_A_4006_325#_c_4138_n 0.00255921f $X=20.41 $Y=1.45
+ $X2=0 $Y2=0
cc_3267 N_S[3]_c_3896_n N_A_4006_325#_c_4138_n 0.00762115f $X=20.41 $Y=1.55
+ $X2=0 $Y2=0
cc_3268 N_S[3]_c_3874_n N_A_4006_325#_c_4123_n 0.0111895f $X=20.31 $Y=0.81 $X2=0
+ $Y2=0
cc_3269 N_S[3]_c_3875_n N_A_4006_325#_c_4123_n 9.67113e-19 $X=20.385 $Y=0.735
+ $X2=0 $Y2=0
cc_3270 N_S[3]_c_3888_n N_A_4006_325#_c_4123_n 0.00426435f $X=20.41 $Y=0.81
+ $X2=0 $Y2=0
cc_3271 N_S[3]_c_3872_n N_A_4006_325#_c_4124_n 0.00416423f $X=19.94 $Y=1.55
+ $X2=0 $Y2=0
cc_3272 N_S[3]_c_3876_n N_A_4006_325#_c_4124_n 0.00322131f $X=20.41 $Y=1.45
+ $X2=0 $Y2=0
cc_3273 N_S[3]_c_3892_n N_A_4006_325#_c_4124_n 0.0228692f $X=19.9 $Y=1.16 $X2=0
+ $Y2=0
cc_3274 N_S[3]_c_3876_n N_A_4006_325#_c_4125_n 0.0175393f $X=20.41 $Y=1.45 $X2=0
+ $Y2=0
cc_3275 N_S[3]_c_3877_n N_A_4006_325#_c_4125_n 0.0179529f $X=20.845 $Y=0.81
+ $X2=0 $Y2=0
cc_3276 N_S[3]_c_3871_n N_VPWR_c_7252_n 0.00652399f $X=19.84 $Y=1.16 $X2=0 $Y2=0
cc_3277 N_S[3]_c_3872_n N_VPWR_c_7252_n 0.00986205f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_3278 N_S[3]_c_3892_n N_VPWR_c_7252_n 0.0157609f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_3279 N_S[3]_c_3896_n N_VPWR_c_7254_n 0.00950399f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_3280 N_S[3]_c_3872_n N_VPWR_c_7325_n 0.0035837f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_3281 N_S[3]_c_3896_n N_VPWR_c_7325_n 0.0035837f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_3282 N_S[3]_c_3872_n VPWR 0.0070533f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_3283 N_S[3]_c_3896_n VPWR 0.00711603f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_3284 N_S[3]_c_3881_n N_Z_c_9018_n 0.0134253f $X=21.68 $Y=0.255 $X2=0 $Y2=0
cc_3285 N_S[3]_c_3883_n N_Z_c_9018_n 0.0077801f $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_3286 N_S[3]_c_3885_n N_Z_c_9018_n 6.35774e-19 $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_3287 N_S[3]_c_3883_n N_Z_c_9020_n 0.00190704f $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_3288 N_S[3]_c_3885_n N_Z_c_9020_n 3.10191e-19 $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_3289 N_S[3]_c_3885_n N_Z_c_9022_n 0.00283489f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_3290 N_S[3]_c_3887_n N_Z_c_9022_n 0.002324f $X=22.94 $Y=0.255 $X2=0 $Y2=0
cc_3291 N_S[3]_c_3881_n N_Z_c_9064_n 0.00216436f $X=21.68 $Y=0.255 $X2=0 $Y2=0
cc_3292 N_S[3]_c_3885_n N_Z_c_9066_n 0.00180363f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_3293 N_S[3]_c_3883_n N_Z_c_9068_n 6.35664e-19 $X=22.1 $Y=0.255 $X2=0 $Y2=0
cc_3294 N_S[3]_c_3885_n N_Z_c_9068_n 0.00462308f $X=22.52 $Y=0.255 $X2=0 $Y2=0
cc_3295 N_S[3]_c_3887_n N_Z_c_9068_n 0.00443615f $X=22.94 $Y=0.255 $X2=0 $Y2=0
cc_3296 N_S[3]_c_3871_n N_Z_c_9119_n 0.00234109f $X=19.84 $Y=1.16 $X2=0 $Y2=0
cc_3297 N_S[3]_c_3872_n N_Z_c_9119_n 0.0052507f $X=19.94 $Y=1.55 $X2=0 $Y2=0
cc_3298 N_S[3]_c_3896_n N_Z_c_9119_n 0.00478771f $X=20.41 $Y=1.55 $X2=0 $Y2=0
cc_3299 N_S[3]_c_3892_n N_Z_c_9119_n 0.0105931f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_3300 N_S[3]_c_3887_n N_A_4219_311#_c_11416_n 0.00168571f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_3301 N_S[3]_c_3896_n N_A_4219_311#_c_11418_n 0.00239129f $X=20.41 $Y=1.55
+ $X2=0 $Y2=0
cc_3302 N_S[3]_c_3871_n N_VGND_c_12727_n 0.00576464f $X=19.84 $Y=1.16 $X2=0
+ $Y2=0
cc_3303 N_S[3]_c_3873_n N_VGND_c_12727_n 0.00374526f $X=19.965 $Y=0.735 $X2=0
+ $Y2=0
cc_3304 N_S[3]_c_3892_n N_VGND_c_12727_n 0.0116218f $X=19.9 $Y=1.16 $X2=0 $Y2=0
cc_3305 N_S[3]_c_3875_n N_VGND_c_12729_n 0.00173127f $X=20.385 $Y=0.735 $X2=0
+ $Y2=0
cc_3306 N_S[3]_c_3877_n N_VGND_c_12729_n 0.00525833f $X=20.845 $Y=0.81 $X2=0
+ $Y2=0
cc_3307 N_S[3]_c_3880_n N_VGND_c_12729_n 0.00862298f $X=20.995 $Y=0.18 $X2=0
+ $Y2=0
cc_3308 N_S[3]_c_3886_n N_VGND_c_12731_n 0.0028166f $X=22.865 $Y=0.18 $X2=0
+ $Y2=0
cc_3309 N_S[3]_c_3887_n N_VGND_c_12731_n 5.5039e-19 $X=22.94 $Y=0.255 $X2=0
+ $Y2=0
cc_3310 N_S[3]_c_3873_n N_VGND_c_12819_n 0.00585385f $X=19.965 $Y=0.735 $X2=0
+ $Y2=0
cc_3311 N_S[3]_c_3874_n N_VGND_c_12819_n 2.16067e-19 $X=20.31 $Y=0.81 $X2=0
+ $Y2=0
cc_3312 N_S[3]_c_3875_n N_VGND_c_12819_n 0.00542362f $X=20.385 $Y=0.735 $X2=0
+ $Y2=0
cc_3313 N_S[3]_c_3880_n N_VGND_c_12823_n 0.0559651f $X=20.995 $Y=0.18 $X2=0
+ $Y2=0
cc_3314 N_S[3]_c_3873_n VGND 0.0119653f $X=19.965 $Y=0.735 $X2=0 $Y2=0
cc_3315 N_S[3]_c_3875_n VGND 0.00990284f $X=20.385 $Y=0.735 $X2=0 $Y2=0
cc_3316 N_S[3]_c_3879_n VGND 0.0244174f $X=21.605 $Y=0.18 $X2=0 $Y2=0
cc_3317 N_S[3]_c_3880_n VGND 0.0101627f $X=20.995 $Y=0.18 $X2=0 $Y2=0
cc_3318 N_S[3]_c_3882_n VGND 0.00642387f $X=22.025 $Y=0.18 $X2=0 $Y2=0
cc_3319 N_S[3]_c_3884_n VGND 0.0064237f $X=22.445 $Y=0.18 $X2=0 $Y2=0
cc_3320 N_S[3]_c_3886_n VGND 0.0123437f $X=22.865 $Y=0.18 $X2=0 $Y2=0
cc_3321 N_S[3]_c_3889_n VGND 0.00366655f $X=21.68 $Y=0.18 $X2=0 $Y2=0
cc_3322 N_S[3]_c_3890_n VGND 0.00366655f $X=22.1 $Y=0.18 $X2=0 $Y2=0
cc_3323 N_S[3]_c_3891_n VGND 0.00366655f $X=22.52 $Y=0.18 $X2=0 $Y2=0
cc_3324 N_S[3]_c_3878_n N_A_4269_66#_c_14539_n 0.00529837f $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_3325 N_S[3]_c_3881_n N_A_4269_66#_c_14540_n 0.0112916f $X=21.68 $Y=0.255
+ $X2=0 $Y2=0
cc_3326 N_S[3]_c_3882_n N_A_4269_66#_c_14540_n 0.00211351f $X=22.025 $Y=0.18
+ $X2=0 $Y2=0
cc_3327 N_S[3]_c_3883_n N_A_4269_66#_c_14540_n 0.0106844f $X=22.1 $Y=0.255 $X2=0
+ $Y2=0
cc_3328 N_S[3]_c_3878_n N_A_4269_66#_c_14541_n 0.00189496f $X=20.92 $Y=0.735
+ $X2=0 $Y2=0
cc_3329 N_S[3]_c_3879_n N_A_4269_66#_c_14541_n 0.00685838f $X=21.605 $Y=0.18
+ $X2=0 $Y2=0
cc_3330 N_S[3]_c_3885_n N_A_4269_66#_c_14542_n 0.0106826f $X=22.52 $Y=0.255
+ $X2=0 $Y2=0
cc_3331 N_S[3]_c_3886_n N_A_4269_66#_c_14542_n 0.00211351f $X=22.865 $Y=0.18
+ $X2=0 $Y2=0
cc_3332 N_S[3]_c_3887_n N_A_4269_66#_c_14542_n 0.0139014f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_3333 N_S[3]_c_3887_n N_A_4269_66#_c_14545_n 0.00206084f $X=22.94 $Y=0.255
+ $X2=0 $Y2=0
cc_3334 N_S[3]_c_3884_n N_A_4269_66#_c_14558_n 0.0034777f $X=22.445 $Y=0.18
+ $X2=0 $Y2=0
cc_3335 N_S[11]_c_4000_n N_A_4006_599#_c_4243_n 0.00507688f $X=21.68 $Y=5.185
+ $X2=25.905 $Y2=0.425
cc_3336 N_S[11]_c_4015_n N_A_4006_599#_c_4235_n 0.00262132f $X=20.41 $Y=3.99
+ $X2=25.905 $Y2=4.845
cc_3337 N_S[11]_c_4002_n N_A_4006_599#_c_4246_n 0.00509204f $X=22.1 $Y=5.185
+ $X2=0 $Y2=0
cc_3338 N_S[11]_c_4006_n N_A_4006_599#_c_4248_n 0.00507426f $X=22.94 $Y=5.185
+ $X2=0 $Y2=0
cc_3339 N_S[11]_c_4004_n N_A_4006_599#_c_4251_n 0.00509391f $X=22.52 $Y=5.185
+ $X2=0 $Y2=0
cc_3340 N_S[11]_c_4013_n N_A_4006_599#_c_4252_n 0.00929139f $X=19.94 $Y=3.89
+ $X2=0 $Y2=0
cc_3341 N_S[11]_c_4017_n N_A_4006_599#_c_4252_n 0.00970559f $X=20.41 $Y=3.89
+ $X2=0 $Y2=0
cc_3342 N_S[11]_c_3992_n N_A_4006_599#_c_4236_n 0.00207203f $X=19.965 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_3343 N_S[11]_c_3993_n N_A_4006_599#_c_4236_n 0.0111895f $X=20.31 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_3344 N_S[11]_c_3995_n N_A_4006_599#_c_4236_n 9.67113e-19 $X=20.385 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_3345 N_S[11]_c_3997_n N_A_4006_599#_c_4236_n 6.53442e-19 $X=20.92 $Y=5.185
+ $X2=25.99 $Y2=0.51
cc_3346 N_S[11]_c_4007_n N_A_4006_599#_c_4236_n 0.00426435f $X=20.41 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_3347 N_S[11]_c_3995_n N_A_4006_599#_c_4237_n 0.00603996f $X=20.385 $Y=4.705
+ $X2=0 $Y2=0
cc_3348 N_S[11]_c_4013_n N_A_4006_599#_c_4253_n 0.00117303f $X=19.94 $Y=3.89
+ $X2=0 $Y2=0
cc_3349 N_S[11]_c_3992_n N_A_4006_599#_c_4253_n 0.00336772f $X=19.965 $Y=4.705
+ $X2=0 $Y2=0
cc_3350 N_S[11]_c_4015_n N_A_4006_599#_c_4253_n 0.00508008f $X=20.41 $Y=3.99
+ $X2=0 $Y2=0
cc_3351 N_S[11]_c_3994_n N_A_4006_599#_c_4253_n 0.00255921f $X=20.41 $Y=4.555
+ $X2=0 $Y2=0
cc_3352 N_S[11]_c_4017_n N_A_4006_599#_c_4253_n 0.00254107f $X=20.41 $Y=3.89
+ $X2=0 $Y2=0
cc_3353 N_S[11]_c_3994_n N_A_4006_599#_c_4238_n 0.0206368f $X=20.41 $Y=4.555
+ $X2=0 $Y2=0
cc_3354 N_S[11]_c_3996_n N_A_4006_599#_c_4238_n 0.0103812f $X=20.845 $Y=4.63
+ $X2=0 $Y2=0
cc_3355 N_S[11]_c_4013_n N_A_4006_599#_c_4255_n 0.00304348f $X=19.94 $Y=3.89
+ $X2=0 $Y2=0
cc_3356 N_S[11]_c_3992_n N_A_4006_599#_c_4255_n 5.48523e-19 $X=19.965 $Y=4.705
+ $X2=0 $Y2=0
cc_3357 N_S[11]_c_4017_n N_A_4006_599#_c_4255_n 0.00216424f $X=20.41 $Y=3.89
+ $X2=0 $Y2=0
cc_3358 N_S[11]_c_3992_n N_A_4006_599#_c_4239_n 0.00289358f $X=19.965 $Y=4.705
+ $X2=0 $Y2=0
cc_3359 N_S[11]_c_3993_n N_A_4006_599#_c_4239_n 0.00429801f $X=20.31 $Y=4.63
+ $X2=0 $Y2=0
cc_3360 N_S[11]_c_3994_n N_A_4006_599#_c_4239_n 0.0085951f $X=20.41 $Y=4.555
+ $X2=0 $Y2=0
cc_3361 N_S[11]_c_4007_n N_A_4006_599#_c_4239_n 0.00268644f $X=20.41 $Y=4.63
+ $X2=0 $Y2=0
cc_3362 N_S[11]_c_4011_n N_A_4006_599#_c_4239_n 0.00541767f $X=19.9 $Y=4.28
+ $X2=0 $Y2=0
cc_3363 N_S[11]_c_3992_n N_A_4006_599#_c_4240_n 0.00416423f $X=19.965 $Y=4.705
+ $X2=0 $Y2=0
cc_3364 N_S[11]_c_3994_n N_A_4006_599#_c_4240_n 0.00322131f $X=20.41 $Y=4.555
+ $X2=0 $Y2=0
cc_3365 N_S[11]_c_4011_n N_A_4006_599#_c_4240_n 0.0228692f $X=19.9 $Y=4.28 $X2=0
+ $Y2=0
cc_3366 N_S[11]_c_3994_n N_A_4006_599#_c_4241_n 0.0175393f $X=20.41 $Y=4.555
+ $X2=0 $Y2=0
cc_3367 N_S[11]_c_3996_n N_A_4006_599#_c_4241_n 0.0179529f $X=20.845 $Y=4.63
+ $X2=0 $Y2=0
cc_3368 N_S[11]_c_3991_n N_VPWR_c_7253_n 0.00652399f $X=19.84 $Y=4.28 $X2=0
+ $Y2=0
cc_3369 N_S[11]_c_4013_n N_VPWR_c_7253_n 0.00986205f $X=19.94 $Y=3.89 $X2=0
+ $Y2=0
cc_3370 N_S[11]_c_4011_n N_VPWR_c_7253_n 0.0157609f $X=19.9 $Y=4.28 $X2=0 $Y2=0
cc_3371 N_S[11]_c_4017_n N_VPWR_c_7255_n 0.00950399f $X=20.41 $Y=3.89 $X2=0
+ $Y2=0
cc_3372 N_S[11]_c_4013_n N_VPWR_c_7325_n 0.0035837f $X=19.94 $Y=3.89 $X2=0 $Y2=0
cc_3373 N_S[11]_c_4017_n N_VPWR_c_7325_n 0.0035837f $X=20.41 $Y=3.89 $X2=0 $Y2=0
cc_3374 N_S[11]_c_4013_n VPWR 0.0070533f $X=19.94 $Y=3.89 $X2=0 $Y2=0
cc_3375 N_S[11]_c_4017_n VPWR 0.00711603f $X=20.41 $Y=3.89 $X2=0 $Y2=0
cc_3376 N_S[11]_c_4000_n N_Z_c_9019_n 0.0134253f $X=21.68 $Y=5.185 $X2=0 $Y2=0
cc_3377 N_S[11]_c_4002_n N_Z_c_9019_n 0.0077801f $X=22.1 $Y=5.185 $X2=0 $Y2=0
cc_3378 N_S[11]_c_4004_n N_Z_c_9019_n 6.35774e-19 $X=22.52 $Y=5.185 $X2=0 $Y2=0
cc_3379 N_S[11]_c_4002_n N_Z_c_9021_n 0.00190704f $X=22.1 $Y=5.185 $X2=0 $Y2=0
cc_3380 N_S[11]_c_4004_n N_Z_c_9021_n 3.10191e-19 $X=22.52 $Y=5.185 $X2=0 $Y2=0
cc_3381 N_S[11]_c_4000_n N_Z_c_9065_n 0.00216436f $X=21.68 $Y=5.185 $X2=0 $Y2=0
cc_3382 N_S[11]_c_4004_n N_Z_c_9067_n 0.00180363f $X=22.52 $Y=5.185 $X2=0 $Y2=0
cc_3383 N_S[11]_c_4004_n N_Z_c_9069_n 0.00462308f $X=22.52 $Y=5.185 $X2=0 $Y2=0
cc_3384 N_S[11]_c_4006_n N_Z_c_9069_n 0.00443615f $X=22.94 $Y=5.185 $X2=0 $Y2=0
cc_3385 N_S[11]_c_4002_n N_Z_c_9070_n 6.35664e-19 $X=22.1 $Y=5.185 $X2=0 $Y2=0
cc_3386 N_S[11]_c_4004_n N_Z_c_9070_n 0.00283489f $X=22.52 $Y=5.185 $X2=0 $Y2=0
cc_3387 N_S[11]_c_4006_n N_Z_c_9070_n 0.002324f $X=22.94 $Y=5.185 $X2=0 $Y2=0
cc_3388 N_S[11]_c_3991_n N_Z_c_9120_n 0.00234109f $X=19.84 $Y=4.28 $X2=0 $Y2=0
cc_3389 N_S[11]_c_4013_n N_Z_c_9120_n 0.00501777f $X=19.94 $Y=3.89 $X2=0 $Y2=0
cc_3390 N_S[11]_c_3992_n N_Z_c_9120_n 2.32936e-19 $X=19.965 $Y=4.705 $X2=0 $Y2=0
cc_3391 N_S[11]_c_4015_n N_Z_c_9120_n 2.55735e-19 $X=20.41 $Y=3.99 $X2=0 $Y2=0
cc_3392 N_S[11]_c_4017_n N_Z_c_9120_n 0.00453198f $X=20.41 $Y=3.89 $X2=0 $Y2=0
cc_3393 N_S[11]_c_4011_n N_Z_c_9120_n 0.0105931f $X=19.9 $Y=4.28 $X2=0 $Y2=0
cc_3394 N_S[11]_c_4006_n N_A_4219_613#_c_11547_n 0.00168571f $X=22.94 $Y=5.185
+ $X2=0 $Y2=0
cc_3395 N_S[11]_c_4017_n N_A_4219_613#_c_11549_n 0.00239129f $X=20.41 $Y=3.89
+ $X2=0 $Y2=0
cc_3396 N_S[11]_c_3991_n N_VGND_c_12728_n 0.00576464f $X=19.84 $Y=4.28 $X2=0
+ $Y2=0
cc_3397 N_S[11]_c_3992_n N_VGND_c_12728_n 0.00374526f $X=19.965 $Y=4.705 $X2=0
+ $Y2=0
cc_3398 N_S[11]_c_4011_n N_VGND_c_12728_n 0.0116218f $X=19.9 $Y=4.28 $X2=0 $Y2=0
cc_3399 N_S[11]_c_3995_n N_VGND_c_12730_n 0.00173127f $X=20.385 $Y=4.705 $X2=0
+ $Y2=0
cc_3400 N_S[11]_c_3996_n N_VGND_c_12730_n 0.00525833f $X=20.845 $Y=4.63 $X2=0
+ $Y2=0
cc_3401 N_S[11]_c_3997_n N_VGND_c_12730_n 0.00862298f $X=20.92 $Y=5.185 $X2=0
+ $Y2=0
cc_3402 N_S[11]_c_4005_n N_VGND_c_12732_n 0.0028166f $X=22.865 $Y=5.26 $X2=0
+ $Y2=0
cc_3403 N_S[11]_c_4006_n N_VGND_c_12732_n 5.5039e-19 $X=22.94 $Y=5.185 $X2=0
+ $Y2=0
cc_3404 N_S[11]_c_3992_n N_VGND_c_12821_n 0.00585385f $X=19.965 $Y=4.705 $X2=0
+ $Y2=0
cc_3405 N_S[11]_c_3993_n N_VGND_c_12821_n 2.16067e-19 $X=20.31 $Y=4.63 $X2=0
+ $Y2=0
cc_3406 N_S[11]_c_3995_n N_VGND_c_12821_n 0.00542362f $X=20.385 $Y=4.705 $X2=0
+ $Y2=0
cc_3407 N_S[11]_c_3999_n N_VGND_c_12825_n 0.0559651f $X=20.995 $Y=5.26 $X2=0
+ $Y2=0
cc_3408 N_S[11]_c_3992_n VGND 0.0119653f $X=19.965 $Y=4.705 $X2=0 $Y2=0
cc_3409 N_S[11]_c_3995_n VGND 0.00990284f $X=20.385 $Y=4.705 $X2=0 $Y2=0
cc_3410 N_S[11]_c_3998_n VGND 0.0244174f $X=21.605 $Y=5.26 $X2=0 $Y2=0
cc_3411 N_S[11]_c_3999_n VGND 0.0101627f $X=20.995 $Y=5.26 $X2=0 $Y2=0
cc_3412 N_S[11]_c_4001_n VGND 0.00642387f $X=22.025 $Y=5.26 $X2=0 $Y2=0
cc_3413 N_S[11]_c_4003_n VGND 0.0064237f $X=22.445 $Y=5.26 $X2=0 $Y2=0
cc_3414 N_S[11]_c_4005_n VGND 0.0123437f $X=22.865 $Y=5.26 $X2=0 $Y2=0
cc_3415 N_S[11]_c_4008_n VGND 0.00366655f $X=21.68 $Y=5.26 $X2=0 $Y2=0
cc_3416 N_S[11]_c_4009_n VGND 0.00366655f $X=22.1 $Y=5.26 $X2=0 $Y2=0
cc_3417 N_S[11]_c_4010_n VGND 0.00366655f $X=22.52 $Y=5.26 $X2=0 $Y2=0
cc_3418 N_S[11]_c_3996_n N_A_4269_918#_c_14623_n 0.00529837f $X=20.845 $Y=4.63
+ $X2=0 $Y2=0
cc_3419 N_S[11]_c_4000_n N_A_4269_918#_c_14624_n 0.0112916f $X=21.68 $Y=5.185
+ $X2=0 $Y2=0
cc_3420 N_S[11]_c_4001_n N_A_4269_918#_c_14624_n 0.00211351f $X=22.025 $Y=5.26
+ $X2=0 $Y2=0
cc_3421 N_S[11]_c_4002_n N_A_4269_918#_c_14624_n 0.0106844f $X=22.1 $Y=5.185
+ $X2=0 $Y2=0
cc_3422 N_S[11]_c_3997_n N_A_4269_918#_c_14625_n 0.00189496f $X=20.92 $Y=5.185
+ $X2=0 $Y2=0
cc_3423 N_S[11]_c_3998_n N_A_4269_918#_c_14625_n 0.00685838f $X=21.605 $Y=5.26
+ $X2=0 $Y2=0
cc_3424 N_S[11]_c_4004_n N_A_4269_918#_c_14626_n 0.0106826f $X=22.52 $Y=5.185
+ $X2=0 $Y2=0
cc_3425 N_S[11]_c_4005_n N_A_4269_918#_c_14626_n 0.00211351f $X=22.865 $Y=5.26
+ $X2=0 $Y2=0
cc_3426 N_S[11]_c_4006_n N_A_4269_918#_c_14626_n 0.0139014f $X=22.94 $Y=5.185
+ $X2=0 $Y2=0
cc_3427 N_S[11]_c_4006_n N_A_4269_918#_c_14629_n 0.00206084f $X=22.94 $Y=5.185
+ $X2=0 $Y2=0
cc_3428 N_S[11]_c_4003_n N_A_4269_918#_c_14642_n 0.0034777f $X=22.445 $Y=5.26
+ $X2=0 $Y2=0
cc_3429 N_A_4006_325#_c_4126_n N_A_4006_599#_c_4242_n 0.0129371f $X=21.455
+ $Y=1.475 $X2=0 $Y2=0
cc_3430 N_A_4006_325#_c_4129_n N_A_4006_599#_c_4245_n 0.0129371f $X=21.925
+ $Y=1.475 $X2=0 $Y2=0
cc_3431 N_A_4006_325#_c_4131_n N_A_4006_599#_c_4247_n 0.0129371f $X=22.395
+ $Y=1.475 $X2=0 $Y2=0
cc_3432 N_A_4006_325#_c_4133_n N_A_4006_599#_c_4249_n 0.0129371f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_3433 N_A_4006_325#_c_4136_n N_VPWR_c_7252_n 0.0356181f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_3434 N_A_4006_325#_c_4126_n N_VPWR_c_7254_n 0.00367058f $X=21.455 $Y=1.475
+ $X2=0 $Y2=0
cc_3435 N_A_4006_325#_c_4136_n N_VPWR_c_7254_n 0.0316788f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_3436 N_A_4006_325#_c_4122_n N_VPWR_c_7254_n 0.0193185f $X=21.225 $Y=1.23
+ $X2=0 $Y2=0
cc_3437 N_A_4006_325#_c_4125_n N_VPWR_c_7254_n 6.4101e-19 $X=21.135 $Y=1.23
+ $X2=0 $Y2=0
cc_3438 N_A_4006_325#_c_4133_n N_VPWR_c_7256_n 0.00324472f $X=22.865 $Y=1.475
+ $X2=0 $Y2=0
cc_3439 N_A_4006_325#_c_4136_n N_VPWR_c_7325_n 0.0233824f $X=20.175 $Y=1.77
+ $X2=0 $Y2=0
cc_3440 N_A_4006_325#_c_4126_n VPWR 0.00473731f $X=21.455 $Y=1.475 $X2=0 $Y2=0
cc_3441 N_A_4006_325#_c_4129_n VPWR 0.00362156f $X=21.925 $Y=1.475 $X2=0 $Y2=0
cc_3442 N_A_4006_325#_c_4131_n VPWR 0.00362156f $X=22.395 $Y=1.475 $X2=0 $Y2=0
cc_3443 N_A_4006_325#_c_4133_n VPWR 0.00473731f $X=22.865 $Y=1.475 $X2=0 $Y2=0
cc_3444 N_A_4006_325#_c_4136_n VPWR 0.00593513f $X=20.175 $Y=1.77 $X2=0 $Y2=0
cc_3445 N_A_4006_325#_c_4130_n N_Z_c_9020_n 0.00762343f $X=22.305 $Y=1.4 $X2=0
+ $Y2=0
cc_3446 N_A_4006_325#_c_4135_n N_Z_c_9020_n 0.00704092f $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_3447 N_A_4006_325#_c_4127_n N_Z_c_9064_n 0.00597584f $X=21.835 $Y=1.4 $X2=0
+ $Y2=0
cc_3448 N_A_4006_325#_c_4119_n N_Z_c_9064_n 0.00747617f $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_3449 N_A_4006_325#_c_4130_n N_Z_c_9064_n 0.00145542f $X=22.305 $Y=1.4 $X2=0
+ $Y2=0
cc_3450 N_A_4006_325#_c_4134_n N_Z_c_9064_n 0.00909323f $X=21.925 $Y=1.4 $X2=0
+ $Y2=0
cc_3451 N_A_4006_325#_c_4122_n N_Z_c_9064_n 0.0266078f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_3452 N_A_4006_325#_c_4132_n N_Z_c_9066_n 0.00918337f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_3453 N_A_4006_325#_c_4135_n N_Z_c_9066_n 2.98555e-19 $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_3454 N_A_4006_325#_c_4132_n N_Z_c_9068_n 0.00248496f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_3455 N_A_4006_325#_c_4126_n N_Z_c_9119_n 0.00795576f $X=21.455 $Y=1.475 $X2=0
+ $Y2=0
cc_3456 N_A_4006_325#_c_4119_n N_Z_c_9119_n 2.19754e-19 $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_3457 N_A_4006_325#_c_4136_n N_Z_c_9119_n 0.0329704f $X=20.175 $Y=1.77 $X2=0
+ $Y2=0
cc_3458 N_A_4006_325#_c_4122_n N_Z_c_9119_n 0.0186685f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_3459 N_A_4006_325#_c_4133_n N_Z_c_9121_n 0.00834829f $X=22.865 $Y=1.475 $X2=0
+ $Y2=0
cc_3460 N_A_4006_325#_c_4129_n N_Z_c_9494_n 0.00372248f $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_3461 N_A_4006_325#_c_4131_n N_Z_c_9494_n 0.00372458f $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_3462 N_A_4006_325#_c_4126_n N_Z_c_9137_n 0.0221748f $X=21.455 $Y=1.475 $X2=0
+ $Y2=0
cc_3463 N_A_4006_325#_c_4127_n N_Z_c_9137_n 0.00560592f $X=21.835 $Y=1.4 $X2=0
+ $Y2=0
cc_3464 N_A_4006_325#_c_4119_n N_Z_c_9137_n 0.00425035f $X=21.545 $Y=1.4 $X2=0
+ $Y2=0
cc_3465 N_A_4006_325#_c_4129_n N_Z_c_9137_n 0.0181262f $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_3466 N_A_4006_325#_c_4131_n N_Z_c_9137_n 9.74366e-19 $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_3467 N_A_4006_325#_c_4134_n N_Z_c_9137_n 0.00181273f $X=21.925 $Y=1.4 $X2=0
+ $Y2=0
cc_3468 N_A_4006_325#_c_4122_n N_Z_c_9137_n 0.00240108f $X=21.225 $Y=1.23 $X2=0
+ $Y2=0
cc_3469 N_A_4006_325#_c_4129_n N_Z_c_9138_n 9.74366e-19 $X=21.925 $Y=1.475 $X2=0
+ $Y2=0
cc_3470 N_A_4006_325#_c_4131_n N_Z_c_9138_n 0.0181262f $X=22.395 $Y=1.475 $X2=0
+ $Y2=0
cc_3471 N_A_4006_325#_c_4132_n N_Z_c_9138_n 0.0103509f $X=22.775 $Y=1.4 $X2=0
+ $Y2=0
cc_3472 N_A_4006_325#_c_4133_n N_Z_c_9138_n 0.0199111f $X=22.865 $Y=1.475 $X2=0
+ $Y2=0
cc_3473 N_A_4006_325#_c_4135_n N_Z_c_9138_n 0.00415268f $X=22.395 $Y=1.4 $X2=0
+ $Y2=0
cc_3474 N_A_4006_325#_c_4133_n N_A_4219_311#_c_11416_n 0.00151141f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_3475 N_A_4006_325#_c_4126_n N_A_4219_311#_c_11424_n 0.00307958f $X=21.455
+ $Y=1.475 $X2=0 $Y2=0
cc_3476 N_A_4006_325#_c_4129_n N_A_4219_311#_c_11424_n 0.00307958f $X=21.925
+ $Y=1.475 $X2=0 $Y2=0
cc_3477 N_A_4006_325#_c_4131_n N_A_4219_311#_c_11426_n 0.00307958f $X=22.395
+ $Y=1.475 $X2=0 $Y2=0
cc_3478 N_A_4006_325#_c_4133_n N_A_4219_311#_c_11426_n 0.00307958f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_3479 N_A_4006_325#_c_4126_n N_A_4219_311#_c_11418_n 0.00499839f $X=21.455
+ $Y=1.475 $X2=0 $Y2=0
cc_3480 N_A_4006_325#_c_4119_n N_A_4219_311#_c_11418_n 0.00561627f $X=21.545
+ $Y=1.4 $X2=0 $Y2=0
cc_3481 N_A_4006_325#_c_4122_n N_A_4219_311#_c_11418_n 0.0218124f $X=21.225
+ $Y=1.23 $X2=0 $Y2=0
cc_3482 N_A_4006_325#_c_4125_n N_A_4219_311#_c_11418_n 5.74251e-19 $X=21.135
+ $Y=1.23 $X2=0 $Y2=0
cc_3483 N_A_4006_325#_c_4129_n N_A_4219_311#_c_11419_n 0.00210632f $X=21.925
+ $Y=1.475 $X2=0 $Y2=0
cc_3484 N_A_4006_325#_c_4130_n N_A_4219_311#_c_11419_n 0.00251792f $X=22.305
+ $Y=1.4 $X2=0 $Y2=0
cc_3485 N_A_4006_325#_c_4131_n N_A_4219_311#_c_11419_n 0.00210632f $X=22.395
+ $Y=1.475 $X2=0 $Y2=0
cc_3486 N_A_4006_325#_c_4133_n N_A_4219_311#_c_11420_n 0.00554566f $X=22.865
+ $Y=1.475 $X2=0 $Y2=0
cc_3487 N_A_4006_325#_c_4122_n N_VGND_c_12729_n 0.0123065f $X=21.225 $Y=1.23
+ $X2=0 $Y2=0
cc_3488 N_A_4006_325#_c_4125_n N_VGND_c_12729_n 2.04129e-19 $X=21.135 $Y=1.23
+ $X2=0 $Y2=0
cc_3489 N_A_4006_325#_c_4120_n N_VGND_c_12819_n 0.0129994f $X=20.175 $Y=0.445
+ $X2=0 $Y2=0
cc_3490 N_A_4006_325#_M1234_s VGND 0.00394793f $X=20.04 $Y=0.235 $X2=0 $Y2=0
cc_3491 N_A_4006_325#_c_4120_n VGND 0.00927134f $X=20.175 $Y=0.445 $X2=0 $Y2=0
cc_3492 N_A_4006_325#_c_4119_n N_A_4269_66#_c_14539_n 0.00600378f $X=21.545
+ $Y=1.4 $X2=0 $Y2=0
cc_3493 N_A_4006_325#_c_4122_n N_A_4269_66#_c_14539_n 0.0028695f $X=21.225
+ $Y=1.23 $X2=0 $Y2=0
cc_3494 N_A_4006_325#_c_4130_n N_A_4269_66#_c_14561_n 7.0477e-19 $X=22.305
+ $Y=1.4 $X2=0 $Y2=0
cc_3495 N_A_4006_599#_c_4252_n N_VPWR_c_7253_n 0.0356181f $X=20.175 $Y=3.14
+ $X2=0 $Y2=0
cc_3496 N_A_4006_599#_c_4242_n N_VPWR_c_7255_n 0.00367058f $X=21.455 $Y=3.965
+ $X2=0 $Y2=0
cc_3497 N_A_4006_599#_c_4252_n N_VPWR_c_7255_n 0.0316788f $X=20.175 $Y=3.14
+ $X2=0 $Y2=0
cc_3498 N_A_4006_599#_c_4238_n N_VPWR_c_7255_n 0.0193185f $X=21.225 $Y=4.21
+ $X2=0 $Y2=0
cc_3499 N_A_4006_599#_c_4241_n N_VPWR_c_7255_n 6.4101e-19 $X=21.135 $Y=4.21
+ $X2=0 $Y2=0
cc_3500 N_A_4006_599#_c_4249_n N_VPWR_c_7257_n 0.00324472f $X=22.865 $Y=3.965
+ $X2=0 $Y2=0
cc_3501 N_A_4006_599#_c_4252_n N_VPWR_c_7325_n 0.0233824f $X=20.175 $Y=3.14
+ $X2=0 $Y2=0
cc_3502 N_A_4006_599#_c_4242_n VPWR 0.00473731f $X=21.455 $Y=3.965 $X2=0 $Y2=0
cc_3503 N_A_4006_599#_c_4245_n VPWR 0.00362156f $X=21.925 $Y=3.965 $X2=0 $Y2=0
cc_3504 N_A_4006_599#_c_4247_n VPWR 0.00362156f $X=22.395 $Y=3.965 $X2=0 $Y2=0
cc_3505 N_A_4006_599#_c_4249_n VPWR 0.00473731f $X=22.865 $Y=3.965 $X2=0 $Y2=0
cc_3506 N_A_4006_599#_c_4252_n VPWR 0.00593513f $X=20.175 $Y=3.14 $X2=0 $Y2=0
cc_3507 N_A_4006_599#_c_4246_n N_Z_c_9021_n 0.00762343f $X=22.305 $Y=4.04 $X2=0
+ $Y2=0
cc_3508 N_A_4006_599#_c_4251_n N_Z_c_9021_n 0.00704092f $X=22.395 $Y=4.04 $X2=0
+ $Y2=0
cc_3509 N_A_4006_599#_c_4243_n N_Z_c_9065_n 0.00597584f $X=21.835 $Y=4.04 $X2=0
+ $Y2=0
cc_3510 N_A_4006_599#_c_4235_n N_Z_c_9065_n 0.00747617f $X=21.545 $Y=4.04 $X2=0
+ $Y2=0
cc_3511 N_A_4006_599#_c_4246_n N_Z_c_9065_n 0.00145542f $X=22.305 $Y=4.04 $X2=0
+ $Y2=0
cc_3512 N_A_4006_599#_c_4250_n N_Z_c_9065_n 0.00909323f $X=21.925 $Y=4.04 $X2=0
+ $Y2=0
cc_3513 N_A_4006_599#_c_4238_n N_Z_c_9065_n 0.0266078f $X=21.225 $Y=4.21 $X2=0
+ $Y2=0
cc_3514 N_A_4006_599#_c_4248_n N_Z_c_9067_n 0.00918337f $X=22.775 $Y=4.04 $X2=0
+ $Y2=0
cc_3515 N_A_4006_599#_c_4251_n N_Z_c_9067_n 2.98555e-19 $X=22.395 $Y=4.04 $X2=0
+ $Y2=0
cc_3516 N_A_4006_599#_c_4248_n N_Z_c_9069_n 0.00248496f $X=22.775 $Y=4.04 $X2=0
+ $Y2=0
cc_3517 N_A_4006_599#_c_4242_n N_Z_c_9120_n 0.00795576f $X=21.455 $Y=3.965 $X2=0
+ $Y2=0
cc_3518 N_A_4006_599#_c_4235_n N_Z_c_9120_n 2.19754e-19 $X=21.545 $Y=4.04 $X2=0
+ $Y2=0
cc_3519 N_A_4006_599#_c_4252_n N_Z_c_9120_n 0.0329704f $X=20.175 $Y=3.14 $X2=0
+ $Y2=0
cc_3520 N_A_4006_599#_c_4238_n N_Z_c_9120_n 0.0186685f $X=21.225 $Y=4.21 $X2=0
+ $Y2=0
cc_3521 N_A_4006_599#_c_4249_n N_Z_c_9123_n 0.00834829f $X=22.865 $Y=3.965 $X2=0
+ $Y2=0
cc_3522 N_A_4006_599#_c_4245_n N_Z_c_9523_n 0.00372248f $X=21.925 $Y=3.965 $X2=0
+ $Y2=0
cc_3523 N_A_4006_599#_c_4247_n N_Z_c_9523_n 0.00372458f $X=22.395 $Y=3.965 $X2=0
+ $Y2=0
cc_3524 N_A_4006_599#_c_4242_n N_Z_c_9137_n 0.0221748f $X=21.455 $Y=3.965 $X2=0
+ $Y2=0
cc_3525 N_A_4006_599#_c_4243_n N_Z_c_9137_n 0.00560592f $X=21.835 $Y=4.04 $X2=0
+ $Y2=0
cc_3526 N_A_4006_599#_c_4235_n N_Z_c_9137_n 0.00425035f $X=21.545 $Y=4.04 $X2=0
+ $Y2=0
cc_3527 N_A_4006_599#_c_4245_n N_Z_c_9137_n 0.0181262f $X=21.925 $Y=3.965 $X2=0
+ $Y2=0
cc_3528 N_A_4006_599#_c_4247_n N_Z_c_9137_n 9.74366e-19 $X=22.395 $Y=3.965 $X2=0
+ $Y2=0
cc_3529 N_A_4006_599#_c_4250_n N_Z_c_9137_n 0.00181273f $X=21.925 $Y=4.04 $X2=0
+ $Y2=0
cc_3530 N_A_4006_599#_c_4238_n N_Z_c_9137_n 0.00240108f $X=21.225 $Y=4.21 $X2=0
+ $Y2=0
cc_3531 N_A_4006_599#_c_4245_n N_Z_c_9138_n 9.74366e-19 $X=21.925 $Y=3.965 $X2=0
+ $Y2=0
cc_3532 N_A_4006_599#_c_4247_n N_Z_c_9138_n 0.0181262f $X=22.395 $Y=3.965 $X2=0
+ $Y2=0
cc_3533 N_A_4006_599#_c_4248_n N_Z_c_9138_n 0.0103509f $X=22.775 $Y=4.04 $X2=0
+ $Y2=0
cc_3534 N_A_4006_599#_c_4249_n N_Z_c_9138_n 0.0199111f $X=22.865 $Y=3.965 $X2=0
+ $Y2=0
cc_3535 N_A_4006_599#_c_4251_n N_Z_c_9138_n 0.00415268f $X=22.395 $Y=4.04 $X2=0
+ $Y2=0
cc_3536 N_A_4006_599#_c_4249_n N_A_4219_613#_c_11547_n 0.00151141f $X=22.865
+ $Y=3.965 $X2=0 $Y2=0
cc_3537 N_A_4006_599#_c_4242_n N_A_4219_613#_c_11555_n 0.00307958f $X=21.455
+ $Y=3.965 $X2=0 $Y2=0
cc_3538 N_A_4006_599#_c_4245_n N_A_4219_613#_c_11555_n 0.00307958f $X=21.925
+ $Y=3.965 $X2=0 $Y2=0
cc_3539 N_A_4006_599#_c_4247_n N_A_4219_613#_c_11557_n 0.00307958f $X=22.395
+ $Y=3.965 $X2=0 $Y2=0
cc_3540 N_A_4006_599#_c_4249_n N_A_4219_613#_c_11557_n 0.00307958f $X=22.865
+ $Y=3.965 $X2=0 $Y2=0
cc_3541 N_A_4006_599#_c_4242_n N_A_4219_613#_c_11549_n 0.00499839f $X=21.455
+ $Y=3.965 $X2=0 $Y2=0
cc_3542 N_A_4006_599#_c_4235_n N_A_4219_613#_c_11549_n 0.00561627f $X=21.545
+ $Y=4.04 $X2=0 $Y2=0
cc_3543 N_A_4006_599#_c_4238_n N_A_4219_613#_c_11549_n 0.0218124f $X=21.225
+ $Y=4.21 $X2=0 $Y2=0
cc_3544 N_A_4006_599#_c_4241_n N_A_4219_613#_c_11549_n 5.74251e-19 $X=21.135
+ $Y=4.21 $X2=0 $Y2=0
cc_3545 N_A_4006_599#_c_4245_n N_A_4219_613#_c_11550_n 0.00210632f $X=21.925
+ $Y=3.965 $X2=0 $Y2=0
cc_3546 N_A_4006_599#_c_4246_n N_A_4219_613#_c_11550_n 0.00251792f $X=22.305
+ $Y=4.04 $X2=0 $Y2=0
cc_3547 N_A_4006_599#_c_4247_n N_A_4219_613#_c_11550_n 0.00210632f $X=22.395
+ $Y=3.965 $X2=0 $Y2=0
cc_3548 N_A_4006_599#_c_4249_n N_A_4219_613#_c_11551_n 0.00554566f $X=22.865
+ $Y=3.965 $X2=0 $Y2=0
cc_3549 N_A_4006_599#_c_4238_n N_VGND_c_12730_n 0.0123065f $X=21.225 $Y=4.21
+ $X2=0 $Y2=0
cc_3550 N_A_4006_599#_c_4241_n N_VGND_c_12730_n 2.04129e-19 $X=21.135 $Y=4.21
+ $X2=0 $Y2=0
cc_3551 N_A_4006_599#_c_4237_n N_VGND_c_12821_n 0.0129994f $X=20.175 $Y=4.995
+ $X2=0 $Y2=0
cc_3552 N_A_4006_599#_M1054_s VGND 0.00394793f $X=20.04 $Y=4.785 $X2=0 $Y2=0
cc_3553 N_A_4006_599#_c_4237_n VGND 0.00927134f $X=20.175 $Y=4.995 $X2=0 $Y2=0
cc_3554 N_A_4006_599#_c_4235_n N_A_4269_918#_c_14623_n 0.00600378f $X=21.545
+ $Y=4.04 $X2=0 $Y2=0
cc_3555 N_A_4006_599#_c_4238_n N_A_4269_918#_c_14623_n 0.0028695f $X=21.225
+ $Y=4.21 $X2=0 $Y2=0
cc_3556 N_A_4006_599#_c_4246_n N_A_4269_918#_c_14645_n 7.0477e-19 $X=22.305
+ $Y=4.04 $X2=0 $Y2=0
cc_3557 N_D[3]_M1042_g N_D[11]_M1052_g 0.0130744f $X=23.855 $Y=1.985 $X2=0 $Y2=0
cc_3558 N_D[3]_M1089_g N_D[11]_M1101_g 0.0130744f $X=24.325 $Y=1.985 $X2=0 $Y2=0
cc_3559 N_D[3]_M1116_g N_D[11]_M1129_g 0.0130744f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3560 N_D[3]_M1289_g N_D[11]_M1297_g 0.0130744f $X=25.265 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_3561 N_D[3]_M1042_g N_VPWR_c_7256_n 0.00389633f $X=23.855 $Y=1.985 $X2=0
+ $Y2=0
cc_3562 N_D[3]_M1089_g N_VPWR_c_7258_n 0.00208662f $X=24.325 $Y=1.985 $X2=0
+ $Y2=0
cc_3563 N_D[3]_M1116_g N_VPWR_c_7258_n 0.00208662f $X=24.795 $Y=1.985 $X2=0
+ $Y2=0
cc_3564 N_D[3]_M1289_g N_VPWR_c_7260_n 0.00374733f $X=25.265 $Y=1.985 $X2=0
+ $Y2=0
cc_3565 N_D[3]_M1042_g VPWR 0.00573859f $X=23.855 $Y=1.985 $X2=0 $Y2=0
cc_3566 N_D[3]_M1089_g VPWR 0.00445624f $X=24.325 $Y=1.985 $X2=0 $Y2=0
cc_3567 N_D[3]_M1116_g VPWR 0.00445624f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3568 N_D[3]_M1289_g VPWR 0.00691494f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3569 N_D[3]_M1042_g N_VPWR_c_7356_n 0.0035837f $X=23.855 $Y=1.985 $X2=0 $Y2=0
cc_3570 N_D[3]_M1089_g N_VPWR_c_7356_n 0.0035837f $X=24.325 $Y=1.985 $X2=0 $Y2=0
cc_3571 N_D[3]_M1116_g N_VPWR_c_7357_n 0.0035837f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3572 N_D[3]_M1289_g N_VPWR_c_7357_n 0.0035837f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3573 N_D[3]_M1042_g N_Z_c_9121_n 0.00311896f $X=23.855 $Y=1.985 $X2=0 $Y2=0
cc_3574 N_D[3]_M1089_g N_Z_c_9121_n 0.00306964f $X=24.325 $Y=1.985 $X2=0 $Y2=0
cc_3575 N_D[3]_M1116_g N_Z_c_9121_n 0.00306964f $X=24.795 $Y=1.985 $X2=0 $Y2=0
cc_3576 N_D[3]_M1289_g N_Z_c_9121_n 0.00470782f $X=25.265 $Y=1.985 $X2=0 $Y2=0
cc_3577 N_D[3]_c_4367_n N_Z_c_9121_n 0.00846955f $X=25.16 $Y=1.16 $X2=0 $Y2=0
cc_3578 N_D[3]_M1042_g N_A_4219_311#_c_11415_n 0.013247f $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_3579 N_D[3]_M1089_g N_A_4219_311#_c_11437_n 0.00916655f $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_3580 N_D[3]_M1116_g N_A_4219_311#_c_11437_n 0.00916655f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3581 N_D[3]_c_4365_n N_A_4219_311#_c_11437_n 7.15862e-19 $X=24.705 $Y=1.16
+ $X2=0 $Y2=0
cc_3582 N_D[3]_c_4367_n N_A_4219_311#_c_11437_n 0.0387168f $X=25.16 $Y=1.16
+ $X2=0 $Y2=0
cc_3583 N_D[3]_M1042_g N_A_4219_311#_c_11441_n 8.61029e-19 $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_3584 N_D[3]_M1089_g N_A_4219_311#_c_11441_n 5.79575e-19 $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_3585 N_D[3]_c_4366_n N_A_4219_311#_c_11441_n 8.03631e-19 $X=24.415 $Y=1.16
+ $X2=0 $Y2=0
cc_3586 N_D[3]_c_4367_n N_A_4219_311#_c_11441_n 0.0191156f $X=25.16 $Y=1.16
+ $X2=0 $Y2=0
cc_3587 N_D[3]_M1116_g N_A_4219_311#_c_11445_n 5.79575e-19 $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3588 N_D[3]_M1289_g N_A_4219_311#_c_11445_n 0.00215964f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_3589 N_D[3]_c_4367_n N_A_4219_311#_c_11445_n 0.0217153f $X=25.16 $Y=1.16
+ $X2=0 $Y2=0
cc_3590 N_D[3]_c_4368_n N_A_4219_311#_c_11445_n 8.03631e-19 $X=25.265 $Y=1.16
+ $X2=0 $Y2=0
cc_3591 N_D[3]_M1042_g N_A_4219_311#_c_11417_n 0.00232998f $X=23.855 $Y=1.985
+ $X2=25.99 $Y2=0.51
cc_3592 N_D[3]_M1089_g N_A_4219_311#_c_11450_n 0.00232998f $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_3593 N_D[3]_M1116_g N_A_4219_311#_c_11450_n 0.00232998f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3594 N_D[3]_M1042_g N_A_4219_311#_c_11452_n 0.00977623f $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_3595 N_D[3]_M1089_g N_A_4219_311#_c_11452_n 0.00911325f $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_3596 N_D[3]_M1116_g N_A_4219_311#_c_11452_n 7.05028e-19 $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3597 N_D[3]_M1089_g N_A_4219_311#_c_11455_n 7.05028e-19 $X=24.325 $Y=1.985
+ $X2=0 $Y2=0
cc_3598 N_D[3]_M1116_g N_A_4219_311#_c_11455_n 0.00911325f $X=24.795 $Y=1.985
+ $X2=0 $Y2=0
cc_3599 N_D[3]_M1289_g N_A_4219_311#_c_11455_n 0.00847082f $X=25.265 $Y=1.985
+ $X2=0 $Y2=0
cc_3600 N_D[3]_M1042_g N_A_4219_311#_c_11420_n 0.00333758f $X=23.855 $Y=1.985
+ $X2=0 $Y2=0
cc_3601 N_D[3]_M1041_g N_VGND_c_12731_n 0.00321269f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_3602 N_D[3]_M1100_g N_VGND_c_12731_n 2.6376e-19 $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_3603 N_D[3]_M1100_g N_VGND_c_12733_n 0.0019152f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_3604 N_D[3]_M1135_g N_VGND_c_12733_n 0.00166854f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3605 N_D[3]_M1193_g N_VGND_c_12733_n 2.64031e-19 $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3606 N_D[3]_M1193_g N_VGND_c_12735_n 0.00345859f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3607 N_D[3]_M1041_g VGND 0.00702263f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_3608 N_D[3]_M1100_g VGND 0.00624811f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_3609 N_D[3]_M1135_g VGND 0.00593887f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3610 N_D[3]_M1193_g VGND 0.0111368f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3611 N_D[3]_M1041_g N_VGND_c_12878_n 0.00422241f $X=23.88 $Y=0.56 $X2=0 $Y2=0
cc_3612 N_D[3]_M1100_g N_VGND_c_12878_n 0.00430643f $X=24.3 $Y=0.56 $X2=0 $Y2=0
cc_3613 N_D[3]_M1135_g N_VGND_c_12880_n 0.00422241f $X=24.82 $Y=0.56 $X2=0 $Y2=0
cc_3614 N_D[3]_M1193_g N_VGND_c_12880_n 0.00551064f $X=25.24 $Y=0.56 $X2=0 $Y2=0
cc_3615 N_D[3]_M1041_g N_A_4269_66#_c_14543_n 0.00261078f $X=23.88 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_3616 N_D[3]_M1041_g N_A_4269_66#_c_14544_n 0.0121912f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_3617 N_D[3]_M1041_g N_A_4269_66#_c_14564_n 0.00699463f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_3618 N_D[3]_M1100_g N_A_4269_66#_c_14564_n 0.00661764f $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_3619 N_D[3]_M1135_g N_A_4269_66#_c_14564_n 5.22365e-19 $X=24.82 $Y=0.56 $X2=0
+ $Y2=0
cc_3620 N_D[3]_M1100_g N_A_4269_66#_c_14546_n 0.00900364f $X=24.3 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_3621 N_D[3]_M1135_g N_A_4269_66#_c_14546_n 0.00986515f $X=24.82 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_3622 N_D[3]_M1193_g N_A_4269_66#_c_14546_n 0.00228093f $X=25.24 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_3623 N_D[3]_c_4365_n N_A_4269_66#_c_14546_n 0.00463549f $X=24.705 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_3624 N_D[3]_c_4367_n N_A_4269_66#_c_14546_n 0.0608884f $X=25.16 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_3625 N_D[3]_c_4368_n N_A_4269_66#_c_14546_n 0.00208088f $X=25.265 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_3626 N_D[3]_M1100_g N_A_4269_66#_c_14573_n 5.22365e-19 $X=24.3 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_3627 N_D[3]_M1135_g N_A_4269_66#_c_14573_n 0.00661134f $X=24.82 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_3628 N_D[3]_M1193_g N_A_4269_66#_c_14573_n 0.00529286f $X=25.24 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_3629 N_D[3]_M1041_g N_A_4269_66#_c_14547_n 0.00128201f $X=23.88 $Y=0.56 $X2=0
+ $Y2=0
cc_3630 N_D[3]_M1100_g N_A_4269_66#_c_14547_n 8.68782e-19 $X=24.3 $Y=0.56 $X2=0
+ $Y2=0
cc_3631 N_D[3]_c_4366_n N_A_4269_66#_c_14547_n 0.00208088f $X=24.415 $Y=1.16
+ $X2=0 $Y2=0
cc_3632 N_D[3]_c_4367_n N_A_4269_66#_c_14547_n 0.018367f $X=25.16 $Y=1.16 $X2=0
+ $Y2=0
cc_3633 N_D[11]_M1052_g N_VPWR_c_7257_n 0.00389633f $X=23.855 $Y=3.455 $X2=0
+ $Y2=0
cc_3634 N_D[11]_M1101_g N_VPWR_c_7259_n 0.00208662f $X=24.325 $Y=3.455 $X2=0
+ $Y2=0
cc_3635 N_D[11]_M1129_g N_VPWR_c_7259_n 0.00208662f $X=24.795 $Y=3.455 $X2=0
+ $Y2=0
cc_3636 N_D[11]_M1297_g N_VPWR_c_7262_n 0.00374733f $X=25.265 $Y=3.455 $X2=0
+ $Y2=0
cc_3637 N_D[11]_M1052_g VPWR 0.00573859f $X=23.855 $Y=3.455 $X2=0 $Y2=0
cc_3638 N_D[11]_M1101_g VPWR 0.00445624f $X=24.325 $Y=3.455 $X2=0 $Y2=0
cc_3639 N_D[11]_M1129_g VPWR 0.00445624f $X=24.795 $Y=3.455 $X2=0 $Y2=0
cc_3640 N_D[11]_M1297_g VPWR 0.00691494f $X=25.265 $Y=3.455 $X2=0 $Y2=0
cc_3641 N_D[11]_M1052_g N_VPWR_c_7356_n 0.0035837f $X=23.855 $Y=3.455 $X2=0
+ $Y2=0
cc_3642 N_D[11]_M1101_g N_VPWR_c_7356_n 0.0035837f $X=24.325 $Y=3.455 $X2=0
+ $Y2=0
cc_3643 N_D[11]_M1129_g N_VPWR_c_7357_n 0.0035837f $X=24.795 $Y=3.455 $X2=0
+ $Y2=0
cc_3644 N_D[11]_M1297_g N_VPWR_c_7357_n 0.0035837f $X=25.265 $Y=3.455 $X2=0
+ $Y2=0
cc_3645 N_D[11]_M1052_g N_Z_c_9123_n 0.00311896f $X=23.855 $Y=3.455 $X2=0 $Y2=0
cc_3646 N_D[11]_M1101_g N_Z_c_9123_n 0.00306964f $X=24.325 $Y=3.455 $X2=0 $Y2=0
cc_3647 N_D[11]_M1129_g N_Z_c_9123_n 0.00306964f $X=24.795 $Y=3.455 $X2=0 $Y2=0
cc_3648 N_D[11]_M1297_g N_Z_c_9123_n 0.00470782f $X=25.265 $Y=3.455 $X2=0 $Y2=0
cc_3649 N_D[11]_c_4461_n N_Z_c_9123_n 0.00846955f $X=25.16 $Y=4.28 $X2=0 $Y2=0
cc_3650 N_D[11]_M1052_g N_A_4219_613#_c_11546_n 0.013247f $X=23.855 $Y=3.455
+ $X2=0 $Y2=0
cc_3651 N_D[11]_M1101_g N_A_4219_613#_c_11568_n 0.00916655f $X=24.325 $Y=3.455
+ $X2=0 $Y2=0
cc_3652 N_D[11]_M1129_g N_A_4219_613#_c_11568_n 0.00916655f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3653 N_D[11]_c_4459_n N_A_4219_613#_c_11568_n 7.15862e-19 $X=24.705 $Y=4.28
+ $X2=0 $Y2=0
cc_3654 N_D[11]_c_4461_n N_A_4219_613#_c_11568_n 0.0387168f $X=25.16 $Y=4.28
+ $X2=0 $Y2=0
cc_3655 N_D[11]_M1052_g N_A_4219_613#_c_11572_n 8.61029e-19 $X=23.855 $Y=3.455
+ $X2=0 $Y2=0
cc_3656 N_D[11]_M1101_g N_A_4219_613#_c_11572_n 5.79575e-19 $X=24.325 $Y=3.455
+ $X2=0 $Y2=0
cc_3657 N_D[11]_c_4460_n N_A_4219_613#_c_11572_n 8.03631e-19 $X=24.415 $Y=4.28
+ $X2=0 $Y2=0
cc_3658 N_D[11]_c_4461_n N_A_4219_613#_c_11572_n 0.0191156f $X=25.16 $Y=4.28
+ $X2=0 $Y2=0
cc_3659 N_D[11]_M1129_g N_A_4219_613#_c_11576_n 5.79575e-19 $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3660 N_D[11]_M1297_g N_A_4219_613#_c_11576_n 0.00215964f $X=25.265 $Y=3.455
+ $X2=0 $Y2=0
cc_3661 N_D[11]_c_4461_n N_A_4219_613#_c_11576_n 0.0217153f $X=25.16 $Y=4.28
+ $X2=0 $Y2=0
cc_3662 N_D[11]_c_4462_n N_A_4219_613#_c_11576_n 8.03631e-19 $X=25.265 $Y=4.28
+ $X2=0 $Y2=0
cc_3663 N_D[11]_M1052_g N_A_4219_613#_c_11548_n 0.00232998f $X=23.855 $Y=3.455
+ $X2=25.99 $Y2=0.51
cc_3664 N_D[11]_M1101_g N_A_4219_613#_c_11581_n 0.00232998f $X=24.325 $Y=3.455
+ $X2=0 $Y2=0
cc_3665 N_D[11]_M1129_g N_A_4219_613#_c_11581_n 0.00232998f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3666 N_D[11]_M1052_g N_A_4219_613#_c_11551_n 0.00333758f $X=23.855 $Y=3.455
+ $X2=0 $Y2=0
cc_3667 N_D[11]_M1052_g N_A_4219_613#_c_11584_n 0.00977623f $X=23.855 $Y=3.455
+ $X2=0 $Y2=0
cc_3668 N_D[11]_M1101_g N_A_4219_613#_c_11584_n 0.00911325f $X=24.325 $Y=3.455
+ $X2=0 $Y2=0
cc_3669 N_D[11]_M1129_g N_A_4219_613#_c_11584_n 7.05028e-19 $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3670 N_D[11]_M1101_g N_A_4219_613#_c_11587_n 7.05028e-19 $X=24.325 $Y=3.455
+ $X2=0 $Y2=0
cc_3671 N_D[11]_M1129_g N_A_4219_613#_c_11587_n 0.00911325f $X=24.795 $Y=3.455
+ $X2=0 $Y2=0
cc_3672 N_D[11]_M1297_g N_A_4219_613#_c_11587_n 0.00847082f $X=25.265 $Y=3.455
+ $X2=0 $Y2=0
cc_3673 N_D[11]_M1245_g N_VGND_c_12732_n 0.00321269f $X=23.88 $Y=4.88 $X2=0
+ $Y2=0
cc_3674 N_D[11]_M1296_g N_VGND_c_12732_n 2.6376e-19 $X=24.3 $Y=4.88 $X2=0 $Y2=0
cc_3675 N_D[11]_M1296_g N_VGND_c_12734_n 0.0019152f $X=24.3 $Y=4.88 $X2=0 $Y2=0
cc_3676 N_D[11]_M1310_g N_VGND_c_12734_n 0.00166854f $X=24.82 $Y=4.88 $X2=0
+ $Y2=0
cc_3677 N_D[11]_M1311_g N_VGND_c_12734_n 2.64031e-19 $X=25.24 $Y=4.88 $X2=0
+ $Y2=0
cc_3678 N_D[11]_M1311_g N_VGND_c_12737_n 0.00345859f $X=25.24 $Y=4.88 $X2=0
+ $Y2=0
cc_3679 N_D[11]_M1245_g VGND 0.00702263f $X=23.88 $Y=4.88 $X2=0 $Y2=0
cc_3680 N_D[11]_M1296_g VGND 0.00624811f $X=24.3 $Y=4.88 $X2=0 $Y2=0
cc_3681 N_D[11]_M1310_g VGND 0.00593887f $X=24.82 $Y=4.88 $X2=0 $Y2=0
cc_3682 N_D[11]_M1311_g VGND 0.0111368f $X=25.24 $Y=4.88 $X2=0 $Y2=0
cc_3683 N_D[11]_M1245_g N_VGND_c_12879_n 0.00422241f $X=23.88 $Y=4.88 $X2=0
+ $Y2=0
cc_3684 N_D[11]_M1296_g N_VGND_c_12879_n 0.00430643f $X=24.3 $Y=4.88 $X2=0 $Y2=0
cc_3685 N_D[11]_M1310_g N_VGND_c_12881_n 0.00422241f $X=24.82 $Y=4.88 $X2=0
+ $Y2=0
cc_3686 N_D[11]_M1311_g N_VGND_c_12881_n 0.00551064f $X=25.24 $Y=4.88 $X2=0
+ $Y2=0
cc_3687 N_D[11]_M1245_g N_A_4269_918#_c_14627_n 0.00261078f $X=23.88 $Y=4.88
+ $X2=25.99 $Y2=0.51
cc_3688 N_D[11]_M1245_g N_A_4269_918#_c_14628_n 0.0121912f $X=23.88 $Y=4.88
+ $X2=0 $Y2=0
cc_3689 N_D[11]_M1296_g N_A_4269_918#_c_14648_n 0.00900364f $X=24.3 $Y=4.88
+ $X2=0 $Y2=0
cc_3690 N_D[11]_M1310_g N_A_4269_918#_c_14648_n 0.00899636f $X=24.82 $Y=4.88
+ $X2=0 $Y2=0
cc_3691 N_D[11]_c_4459_n N_A_4269_918#_c_14648_n 0.00463549f $X=24.705 $Y=4.28
+ $X2=0 $Y2=0
cc_3692 N_D[11]_c_4461_n N_A_4269_918#_c_14648_n 0.0394855f $X=25.16 $Y=4.28
+ $X2=0 $Y2=0
cc_3693 N_D[11]_M1245_g N_A_4269_918#_c_14630_n 0.00827664f $X=23.88 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_3694 N_D[11]_M1296_g N_A_4269_918#_c_14630_n 0.00748643f $X=24.3 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_3695 N_D[11]_M1310_g N_A_4269_918#_c_14630_n 5.22365e-19 $X=24.82 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_3696 N_D[11]_c_4460_n N_A_4269_918#_c_14630_n 0.00208088f $X=24.415 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_3697 N_D[11]_c_4461_n N_A_4269_918#_c_14630_n 0.018367f $X=25.16 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_3698 N_D[11]_M1296_g N_A_4269_918#_c_14631_n 5.22365e-19 $X=24.3 $Y=4.88
+ $X2=0 $Y2=0
cc_3699 N_D[11]_M1310_g N_A_4269_918#_c_14631_n 0.00748012f $X=24.82 $Y=4.88
+ $X2=0 $Y2=0
cc_3700 N_D[11]_M1311_g N_A_4269_918#_c_14631_n 0.00757379f $X=25.24 $Y=4.88
+ $X2=0 $Y2=0
cc_3701 N_D[11]_c_4461_n N_A_4269_918#_c_14631_n 0.021403f $X=25.16 $Y=4.28
+ $X2=0 $Y2=0
cc_3702 N_D[11]_c_4462_n N_A_4269_918#_c_14631_n 0.00208088f $X=25.265 $Y=4.28
+ $X2=0 $Y2=0
cc_3703 N_D[4]_M1158_g N_D[12]_M1006_g 0.0130744f $X=26.715 $Y=1.985 $X2=0 $Y2=0
cc_3704 N_D[4]_M1194_g N_D[12]_M1165_g 0.0130744f $X=27.185 $Y=1.985 $X2=0 $Y2=0
cc_3705 N_D[4]_M1265_g N_D[12]_M1203_g 0.0130744f $X=27.655 $Y=1.985 $X2=0 $Y2=0
cc_3706 N_D[4]_M1319_g N_D[12]_M1277_g 0.0130744f $X=28.125 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_3707 N_D[4]_M1158_g N_VPWR_c_7264_n 0.00374733f $X=26.715 $Y=1.985 $X2=0
+ $Y2=0
cc_3708 N_D[4]_M1194_g N_VPWR_c_7268_n 0.00208662f $X=27.185 $Y=1.985 $X2=0
+ $Y2=0
cc_3709 N_D[4]_M1265_g N_VPWR_c_7268_n 0.00208662f $X=27.655 $Y=1.985 $X2=0
+ $Y2=0
cc_3710 N_D[4]_M1265_g N_VPWR_c_7270_n 0.0035837f $X=27.655 $Y=1.985 $X2=0 $Y2=0
cc_3711 N_D[4]_M1319_g N_VPWR_c_7270_n 0.0035837f $X=28.125 $Y=1.985 $X2=0 $Y2=0
cc_3712 N_D[4]_M1319_g N_VPWR_c_7271_n 0.00389633f $X=28.125 $Y=1.985 $X2=0
+ $Y2=0
cc_3713 N_D[4]_M1158_g VPWR 0.00691494f $X=26.715 $Y=1.985 $X2=0 $Y2=0
cc_3714 N_D[4]_M1194_g VPWR 0.00445624f $X=27.185 $Y=1.985 $X2=0 $Y2=0
cc_3715 N_D[4]_M1265_g VPWR 0.00445624f $X=27.655 $Y=1.985 $X2=0 $Y2=0
cc_3716 N_D[4]_M1319_g VPWR 0.00573859f $X=28.125 $Y=1.985 $X2=0 $Y2=0
cc_3717 N_D[4]_M1158_g N_VPWR_c_7361_n 0.0035837f $X=26.715 $Y=1.985 $X2=0 $Y2=0
cc_3718 N_D[4]_M1194_g N_VPWR_c_7361_n 0.0035837f $X=27.185 $Y=1.985 $X2=0 $Y2=0
cc_3719 N_D[4]_M1158_g N_Z_c_9121_n 0.00470782f $X=26.715 $Y=1.985 $X2=0 $Y2=0
cc_3720 N_D[4]_M1194_g N_Z_c_9121_n 0.00306964f $X=27.185 $Y=1.985 $X2=0 $Y2=0
cc_3721 N_D[4]_M1265_g N_Z_c_9121_n 0.00306964f $X=27.655 $Y=1.985 $X2=0 $Y2=0
cc_3722 N_D[4]_M1319_g N_Z_c_9121_n 0.00311896f $X=28.125 $Y=1.985 $X2=0 $Y2=0
cc_3723 N_D[4]_c_4553_n N_Z_c_9121_n 0.00846955f $X=27.84 $Y=1.16 $X2=0 $Y2=0
cc_3724 N_D[4]_M1194_g N_A_5361_297#_c_11682_n 0.00916655f $X=27.185 $Y=1.985
+ $X2=0 $Y2=0
cc_3725 N_D[4]_M1265_g N_A_5361_297#_c_11682_n 0.00916655f $X=27.655 $Y=1.985
+ $X2=0 $Y2=0
cc_3726 N_D[4]_c_4551_n N_A_5361_297#_c_11682_n 7.15862e-19 $X=27.565 $Y=1.16
+ $X2=0 $Y2=0
cc_3727 N_D[4]_c_4553_n N_A_5361_297#_c_11682_n 0.0387168f $X=27.84 $Y=1.16
+ $X2=0 $Y2=0
cc_3728 N_D[4]_M1319_g N_A_5361_297#_c_11677_n 0.013247f $X=28.125 $Y=1.985
+ $X2=0 $Y2=0
cc_3729 N_D[4]_M1158_g N_A_5361_297#_c_11687_n 0.00215964f $X=26.715 $Y=1.985
+ $X2=0 $Y2=0
cc_3730 N_D[4]_M1194_g N_A_5361_297#_c_11687_n 5.79575e-19 $X=27.185 $Y=1.985
+ $X2=0 $Y2=0
cc_3731 N_D[4]_c_4552_n N_A_5361_297#_c_11687_n 8.03631e-19 $X=27.275 $Y=1.16
+ $X2=0 $Y2=0
cc_3732 N_D[4]_c_4553_n N_A_5361_297#_c_11687_n 0.0217153f $X=27.84 $Y=1.16
+ $X2=0 $Y2=0
cc_3733 N_D[4]_M1265_g N_A_5361_297#_c_11691_n 5.79575e-19 $X=27.655 $Y=1.985
+ $X2=0 $Y2=0
cc_3734 N_D[4]_M1319_g N_A_5361_297#_c_11691_n 8.61029e-19 $X=28.125 $Y=1.985
+ $X2=0 $Y2=0
cc_3735 N_D[4]_c_4553_n N_A_5361_297#_c_11691_n 0.0191156f $X=27.84 $Y=1.16
+ $X2=0 $Y2=0
cc_3736 N_D[4]_c_4554_n N_A_5361_297#_c_11691_n 8.03631e-19 $X=28.125 $Y=1.16
+ $X2=0 $Y2=0
cc_3737 N_D[4]_M1194_g N_A_5361_297#_c_11695_n 0.00232998f $X=27.185 $Y=1.985
+ $X2=0 $Y2=0
cc_3738 N_D[4]_M1265_g N_A_5361_297#_c_11695_n 0.00232998f $X=27.655 $Y=1.985
+ $X2=0 $Y2=0
cc_3739 N_D[4]_M1319_g N_A_5361_297#_c_11678_n 0.00232998f $X=28.125 $Y=1.985
+ $X2=0 $Y2=0
cc_3740 N_D[4]_M1158_g N_A_5361_297#_c_11698_n 0.00847082f $X=26.715 $Y=1.985
+ $X2=0 $Y2=0
cc_3741 N_D[4]_M1194_g N_A_5361_297#_c_11698_n 0.00911325f $X=27.185 $Y=1.985
+ $X2=0 $Y2=0
cc_3742 N_D[4]_M1265_g N_A_5361_297#_c_11698_n 7.05028e-19 $X=27.655 $Y=1.985
+ $X2=0 $Y2=0
cc_3743 N_D[4]_M1194_g N_A_5361_297#_c_11701_n 7.05028e-19 $X=27.185 $Y=1.985
+ $X2=0 $Y2=0
cc_3744 N_D[4]_M1265_g N_A_5361_297#_c_11701_n 0.00911325f $X=27.655 $Y=1.985
+ $X2=0 $Y2=0
cc_3745 N_D[4]_M1319_g N_A_5361_297#_c_11701_n 0.00977623f $X=28.125 $Y=1.985
+ $X2=0 $Y2=0
cc_3746 N_D[4]_M1319_g N_A_5361_297#_c_11679_n 0.00333758f $X=28.125 $Y=1.985
+ $X2=0 $Y2=0
cc_3747 N_D[4]_M1021_g N_VGND_c_12738_n 0.00345859f $X=26.74 $Y=0.56 $X2=0 $Y2=0
cc_3748 N_D[4]_M1021_g N_VGND_c_12741_n 2.64031e-19 $X=26.74 $Y=0.56 $X2=0 $Y2=0
cc_3749 N_D[4]_M1177_g N_VGND_c_12741_n 0.00166854f $X=27.16 $Y=0.56 $X2=0 $Y2=0
cc_3750 N_D[4]_M1232_g N_VGND_c_12741_n 0.0019152f $X=27.68 $Y=0.56 $X2=0 $Y2=0
cc_3751 N_D[4]_M1232_g N_VGND_c_12743_n 0.00430643f $X=27.68 $Y=0.56 $X2=0 $Y2=0
cc_3752 N_D[4]_M1275_g N_VGND_c_12743_n 0.00422241f $X=28.1 $Y=0.56 $X2=0 $Y2=0
cc_3753 N_D[4]_M1232_g N_VGND_c_12745_n 2.6376e-19 $X=27.68 $Y=0.56 $X2=0 $Y2=0
cc_3754 N_D[4]_M1275_g N_VGND_c_12745_n 0.00321269f $X=28.1 $Y=0.56 $X2=0 $Y2=0
cc_3755 N_D[4]_M1021_g VGND 0.0111368f $X=26.74 $Y=0.56 $X2=0 $Y2=0
cc_3756 N_D[4]_M1177_g VGND 0.00593887f $X=27.16 $Y=0.56 $X2=0 $Y2=0
cc_3757 N_D[4]_M1232_g VGND 0.00624811f $X=27.68 $Y=0.56 $X2=0 $Y2=0
cc_3758 N_D[4]_M1275_g VGND 0.00702263f $X=28.1 $Y=0.56 $X2=0 $Y2=0
cc_3759 N_D[4]_M1021_g N_VGND_c_12885_n 0.00551064f $X=26.74 $Y=0.56 $X2=0 $Y2=0
cc_3760 N_D[4]_M1177_g N_VGND_c_12885_n 0.00422241f $X=27.16 $Y=0.56 $X2=0 $Y2=0
cc_3761 N_D[4]_M1021_g N_A_5363_47#_c_14713_n 0.00529286f $X=26.74 $Y=0.56 $X2=0
+ $Y2=0
cc_3762 N_D[4]_M1177_g N_A_5363_47#_c_14713_n 0.00661134f $X=27.16 $Y=0.56 $X2=0
+ $Y2=0
cc_3763 N_D[4]_M1232_g N_A_5363_47#_c_14713_n 5.22365e-19 $X=27.68 $Y=0.56 $X2=0
+ $Y2=0
cc_3764 N_D[4]_M1177_g N_A_5363_47#_c_14716_n 0.00899636f $X=27.16 $Y=0.56 $X2=0
+ $Y2=0
cc_3765 N_D[4]_M1232_g N_A_5363_47#_c_14716_n 0.00900364f $X=27.68 $Y=0.56 $X2=0
+ $Y2=0
cc_3766 N_D[4]_c_4551_n N_A_5363_47#_c_14716_n 0.00463549f $X=27.565 $Y=1.16
+ $X2=0 $Y2=0
cc_3767 N_D[4]_c_4553_n N_A_5363_47#_c_14716_n 0.0394855f $X=27.84 $Y=1.16 $X2=0
+ $Y2=0
cc_3768 N_D[4]_M1021_g N_A_5363_47#_c_14705_n 0.00228093f $X=26.74 $Y=0.56 $X2=0
+ $Y2=0
cc_3769 N_D[4]_M1177_g N_A_5363_47#_c_14705_n 8.68782e-19 $X=27.16 $Y=0.56 $X2=0
+ $Y2=0
cc_3770 N_D[4]_c_4552_n N_A_5363_47#_c_14705_n 0.00208088f $X=27.275 $Y=1.16
+ $X2=0 $Y2=0
cc_3771 N_D[4]_c_4553_n N_A_5363_47#_c_14705_n 0.021403f $X=27.84 $Y=1.16 $X2=0
+ $Y2=0
cc_3772 N_D[4]_M1177_g N_A_5363_47#_c_14724_n 5.22365e-19 $X=27.16 $Y=0.56 $X2=0
+ $Y2=0
cc_3773 N_D[4]_M1232_g N_A_5363_47#_c_14724_n 0.00661764f $X=27.68 $Y=0.56 $X2=0
+ $Y2=0
cc_3774 N_D[4]_M1275_g N_A_5363_47#_c_14724_n 0.00699463f $X=28.1 $Y=0.56 $X2=0
+ $Y2=0
cc_3775 N_D[4]_M1275_g N_A_5363_47#_c_14706_n 0.0121912f $X=28.1 $Y=0.56 $X2=0
+ $Y2=0
cc_3776 N_D[4]_M1275_g N_A_5363_47#_c_14707_n 0.00261078f $X=28.1 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_3777 N_D[4]_M1232_g N_A_5363_47#_c_14712_n 8.68782e-19 $X=27.68 $Y=0.56 $X2=0
+ $Y2=0
cc_3778 N_D[4]_M1275_g N_A_5363_47#_c_14712_n 0.00128201f $X=28.1 $Y=0.56 $X2=0
+ $Y2=0
cc_3779 N_D[4]_c_4553_n N_A_5363_47#_c_14712_n 0.018367f $X=27.84 $Y=1.16 $X2=0
+ $Y2=0
cc_3780 N_D[4]_c_4554_n N_A_5363_47#_c_14712_n 0.00208088f $X=28.125 $Y=1.16
+ $X2=0 $Y2=0
cc_3781 N_D[12]_M1006_g N_VPWR_c_7266_n 0.00374733f $X=26.715 $Y=3.455 $X2=0
+ $Y2=0
cc_3782 N_D[12]_M1165_g N_VPWR_c_7269_n 0.00208662f $X=27.185 $Y=3.455 $X2=0
+ $Y2=0
cc_3783 N_D[12]_M1203_g N_VPWR_c_7269_n 0.00208662f $X=27.655 $Y=3.455 $X2=0
+ $Y2=0
cc_3784 N_D[12]_M1203_g N_VPWR_c_7270_n 0.0035837f $X=27.655 $Y=3.455 $X2=0
+ $Y2=0
cc_3785 N_D[12]_M1277_g N_VPWR_c_7270_n 0.0035837f $X=28.125 $Y=3.455 $X2=0
+ $Y2=0
cc_3786 N_D[12]_M1277_g N_VPWR_c_7272_n 0.00389633f $X=28.125 $Y=3.455 $X2=0
+ $Y2=0
cc_3787 N_D[12]_M1006_g VPWR 0.00691494f $X=26.715 $Y=3.455 $X2=0 $Y2=0
cc_3788 N_D[12]_M1165_g VPWR 0.00445624f $X=27.185 $Y=3.455 $X2=0 $Y2=0
cc_3789 N_D[12]_M1203_g VPWR 0.00445624f $X=27.655 $Y=3.455 $X2=0 $Y2=0
cc_3790 N_D[12]_M1277_g VPWR 0.00573859f $X=28.125 $Y=3.455 $X2=0 $Y2=0
cc_3791 N_D[12]_M1006_g N_VPWR_c_7361_n 0.0035837f $X=26.715 $Y=3.455 $X2=0
+ $Y2=0
cc_3792 N_D[12]_M1165_g N_VPWR_c_7361_n 0.0035837f $X=27.185 $Y=3.455 $X2=0
+ $Y2=0
cc_3793 N_D[12]_M1006_g N_Z_c_9123_n 0.00470782f $X=26.715 $Y=3.455 $X2=0 $Y2=0
cc_3794 N_D[12]_M1165_g N_Z_c_9123_n 0.00306964f $X=27.185 $Y=3.455 $X2=0 $Y2=0
cc_3795 N_D[12]_M1203_g N_Z_c_9123_n 0.00306964f $X=27.655 $Y=3.455 $X2=0 $Y2=0
cc_3796 N_D[12]_M1277_g N_Z_c_9123_n 0.00311896f $X=28.125 $Y=3.455 $X2=0 $Y2=0
cc_3797 N_D[12]_c_4649_n N_Z_c_9123_n 0.00846955f $X=27.84 $Y=4.28 $X2=0 $Y2=0
cc_3798 N_D[12]_M1165_g N_A_5361_591#_c_11810_n 0.00916655f $X=27.185 $Y=3.455
+ $X2=0 $Y2=0
cc_3799 N_D[12]_M1203_g N_A_5361_591#_c_11810_n 0.00916655f $X=27.655 $Y=3.455
+ $X2=0 $Y2=0
cc_3800 N_D[12]_c_4647_n N_A_5361_591#_c_11810_n 7.15862e-19 $X=27.565 $Y=4.28
+ $X2=0 $Y2=0
cc_3801 N_D[12]_c_4649_n N_A_5361_591#_c_11810_n 0.0387168f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3802 N_D[12]_M1277_g N_A_5361_591#_c_11805_n 0.013247f $X=28.125 $Y=3.455
+ $X2=0 $Y2=0
cc_3803 N_D[12]_M1006_g N_A_5361_591#_c_11815_n 0.00215964f $X=26.715 $Y=3.455
+ $X2=0 $Y2=0
cc_3804 N_D[12]_M1165_g N_A_5361_591#_c_11815_n 5.79575e-19 $X=27.185 $Y=3.455
+ $X2=0 $Y2=0
cc_3805 N_D[12]_c_4648_n N_A_5361_591#_c_11815_n 8.03631e-19 $X=27.275 $Y=4.28
+ $X2=0 $Y2=0
cc_3806 N_D[12]_c_4649_n N_A_5361_591#_c_11815_n 0.0217153f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3807 N_D[12]_M1203_g N_A_5361_591#_c_11819_n 5.79575e-19 $X=27.655 $Y=3.455
+ $X2=0 $Y2=0
cc_3808 N_D[12]_M1277_g N_A_5361_591#_c_11819_n 8.61029e-19 $X=28.125 $Y=3.455
+ $X2=0 $Y2=0
cc_3809 N_D[12]_c_4649_n N_A_5361_591#_c_11819_n 0.0191156f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3810 N_D[12]_c_4650_n N_A_5361_591#_c_11819_n 8.03631e-19 $X=28.125 $Y=4.28
+ $X2=0 $Y2=0
cc_3811 N_D[12]_M1165_g N_A_5361_591#_c_11823_n 0.00232998f $X=27.185 $Y=3.455
+ $X2=0 $Y2=0
cc_3812 N_D[12]_M1203_g N_A_5361_591#_c_11823_n 0.00232998f $X=27.655 $Y=3.455
+ $X2=0 $Y2=0
cc_3813 N_D[12]_M1277_g N_A_5361_591#_c_11806_n 0.00232998f $X=28.125 $Y=3.455
+ $X2=0 $Y2=0
cc_3814 N_D[12]_M1006_g N_A_5361_591#_c_11826_n 0.00847082f $X=26.715 $Y=3.455
+ $X2=0 $Y2=0
cc_3815 N_D[12]_M1165_g N_A_5361_591#_c_11826_n 0.00911325f $X=27.185 $Y=3.455
+ $X2=0 $Y2=0
cc_3816 N_D[12]_M1203_g N_A_5361_591#_c_11826_n 7.05028e-19 $X=27.655 $Y=3.455
+ $X2=0 $Y2=0
cc_3817 N_D[12]_M1165_g N_A_5361_591#_c_11829_n 7.05028e-19 $X=27.185 $Y=3.455
+ $X2=0 $Y2=0
cc_3818 N_D[12]_M1203_g N_A_5361_591#_c_11829_n 0.00911325f $X=27.655 $Y=3.455
+ $X2=0 $Y2=0
cc_3819 N_D[12]_M1277_g N_A_5361_591#_c_11829_n 0.00977623f $X=28.125 $Y=3.455
+ $X2=0 $Y2=0
cc_3820 N_D[12]_M1277_g N_A_5361_591#_c_11807_n 0.00333758f $X=28.125 $Y=3.455
+ $X2=0 $Y2=0
cc_3821 N_D[12]_M1012_g N_VGND_c_12740_n 0.00345859f $X=26.74 $Y=4.88 $X2=0
+ $Y2=0
cc_3822 N_D[12]_M1012_g N_VGND_c_12742_n 2.64031e-19 $X=26.74 $Y=4.88 $X2=0
+ $Y2=0
cc_3823 N_D[12]_M1128_g N_VGND_c_12742_n 0.00166854f $X=27.16 $Y=4.88 $X2=0
+ $Y2=0
cc_3824 N_D[12]_M1187_g N_VGND_c_12742_n 0.0019152f $X=27.68 $Y=4.88 $X2=0 $Y2=0
cc_3825 N_D[12]_M1187_g N_VGND_c_12744_n 0.00430643f $X=27.68 $Y=4.88 $X2=0
+ $Y2=0
cc_3826 N_D[12]_M1267_g N_VGND_c_12744_n 0.00422241f $X=28.1 $Y=4.88 $X2=0 $Y2=0
cc_3827 N_D[12]_M1187_g N_VGND_c_12746_n 2.6376e-19 $X=27.68 $Y=4.88 $X2=0 $Y2=0
cc_3828 N_D[12]_M1267_g N_VGND_c_12746_n 0.00321269f $X=28.1 $Y=4.88 $X2=0 $Y2=0
cc_3829 N_D[12]_M1012_g VGND 0.0111368f $X=26.74 $Y=4.88 $X2=0 $Y2=0
cc_3830 N_D[12]_M1128_g VGND 0.00593887f $X=27.16 $Y=4.88 $X2=0 $Y2=0
cc_3831 N_D[12]_M1187_g VGND 0.00624811f $X=27.68 $Y=4.88 $X2=0 $Y2=0
cc_3832 N_D[12]_M1267_g VGND 0.00702263f $X=28.1 $Y=4.88 $X2=0 $Y2=0
cc_3833 N_D[12]_M1012_g N_VGND_c_12886_n 0.00551064f $X=26.74 $Y=4.88 $X2=0
+ $Y2=0
cc_3834 N_D[12]_M1128_g N_VGND_c_12886_n 0.00422241f $X=27.16 $Y=4.88 $X2=0
+ $Y2=0
cc_3835 N_D[12]_M1128_g N_A_5363_911#_c_14796_n 0.00899636f $X=27.16 $Y=4.88
+ $X2=0 $Y2=0
cc_3836 N_D[12]_M1187_g N_A_5363_911#_c_14796_n 0.00900364f $X=27.68 $Y=4.88
+ $X2=0 $Y2=0
cc_3837 N_D[12]_c_4647_n N_A_5363_911#_c_14796_n 0.00463549f $X=27.565 $Y=4.28
+ $X2=0 $Y2=0
cc_3838 N_D[12]_c_4649_n N_A_5363_911#_c_14796_n 0.0394855f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3839 N_D[12]_M1267_g N_A_5363_911#_c_14788_n 0.0121912f $X=28.1 $Y=4.88 $X2=0
+ $Y2=0
cc_3840 N_D[12]_M1267_g N_A_5363_911#_c_14789_n 0.00261078f $X=28.1 $Y=4.88
+ $X2=0 $Y2=0
cc_3841 N_D[12]_M1012_g N_A_5363_911#_c_14794_n 0.00757379f $X=26.74 $Y=4.88
+ $X2=0 $Y2=0
cc_3842 N_D[12]_M1128_g N_A_5363_911#_c_14794_n 0.00748012f $X=27.16 $Y=4.88
+ $X2=0 $Y2=0
cc_3843 N_D[12]_M1187_g N_A_5363_911#_c_14794_n 5.22365e-19 $X=27.68 $Y=4.88
+ $X2=0 $Y2=0
cc_3844 N_D[12]_c_4648_n N_A_5363_911#_c_14794_n 0.00208088f $X=27.275 $Y=4.28
+ $X2=0 $Y2=0
cc_3845 N_D[12]_c_4649_n N_A_5363_911#_c_14794_n 0.021403f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3846 N_D[12]_M1128_g N_A_5363_911#_c_14795_n 5.22365e-19 $X=27.16 $Y=4.88
+ $X2=0 $Y2=0
cc_3847 N_D[12]_M1187_g N_A_5363_911#_c_14795_n 0.00748643f $X=27.68 $Y=4.88
+ $X2=0 $Y2=0
cc_3848 N_D[12]_M1267_g N_A_5363_911#_c_14795_n 0.00827664f $X=28.1 $Y=4.88
+ $X2=0 $Y2=0
cc_3849 N_D[12]_c_4649_n N_A_5363_911#_c_14795_n 0.018367f $X=27.84 $Y=4.28
+ $X2=0 $Y2=0
cc_3850 N_D[12]_c_4650_n N_A_5363_911#_c_14795_n 0.00208088f $X=28.125 $Y=4.28
+ $X2=0 $Y2=0
cc_3851 N_A_5803_265#_c_4738_n N_A_5803_793#_c_4857_n 0.0129371f $X=29.115
+ $Y=1.475 $X2=0 $Y2=0
cc_3852 N_A_5803_265#_c_4741_n N_A_5803_793#_c_4860_n 0.0129371f $X=29.585
+ $Y=1.475 $X2=0 $Y2=0
cc_3853 N_A_5803_265#_c_4743_n N_A_5803_793#_c_4862_n 0.0129371f $X=30.055
+ $Y=1.475 $X2=0 $Y2=0
cc_3854 N_A_5803_265#_c_4745_n N_A_5803_793#_c_4864_n 0.0129371f $X=30.525
+ $Y=1.475 $X2=0 $Y2=0
cc_3855 N_A_5803_265#_c_4740_n N_S[4]_c_4975_n 0.00507426f $X=29.205 $Y=1.4
+ $X2=0 $Y2=0
cc_3856 N_A_5803_265#_c_4739_n N_S[4]_c_4978_n 0.00509391f $X=29.495 $Y=1.4
+ $X2=0 $Y2=0
cc_3857 N_A_5803_265#_c_4742_n N_S[4]_c_4980_n 0.00509204f $X=29.965 $Y=1.4
+ $X2=25.905 $Y2=4.845
cc_3858 N_A_5803_265#_c_4744_n N_S[4]_c_4982_n 0.00507688f $X=30.435 $Y=1.4
+ $X2=0 $Y2=0
cc_3859 N_A_5803_265#_c_4733_n N_S[4]_c_4984_n 6.53442e-19 $X=31.805 $Y=0.445
+ $X2=0 $Y2=0
cc_3860 N_A_5803_265#_c_4731_n N_S[4]_c_4986_n 0.0103812f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3861 N_A_5803_265#_c_4732_n N_S[4]_c_4986_n 0.0179529f $X=31.095 $Y=1.23
+ $X2=0 $Y2=0
cc_3862 N_A_5803_265#_c_4731_n N_S[4]_c_4987_n 0.0206368f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3863 N_A_5803_265#_c_4732_n N_S[4]_c_4987_n 0.0175393f $X=31.095 $Y=1.23
+ $X2=0 $Y2=0
cc_3864 N_A_5803_265#_c_4734_n N_S[4]_c_4987_n 0.0085951f $X=31.725 $Y=1.065
+ $X2=0 $Y2=0
cc_3865 N_A_5803_265#_c_4736_n N_S[4]_c_4987_n 0.00322131f $X=31.725 $Y=1.23
+ $X2=0 $Y2=0
cc_3866 N_A_5803_265#_c_4752_n N_S[4]_c_4987_n 0.00255921f $X=31.805 $Y=1.605
+ $X2=0 $Y2=0
cc_3867 N_A_5803_265#_c_4737_n N_S[4]_c_4987_n 0.00262132f $X=30.845 $Y=1.23
+ $X2=0 $Y2=0
cc_3868 N_A_5803_265#_c_4750_n N_S[4]_c_4998_n 0.0118698f $X=31.805 $Y=1.77
+ $X2=0 $Y2=0
cc_3869 N_A_5803_265#_c_4752_n N_S[4]_c_4998_n 0.00762115f $X=31.805 $Y=1.605
+ $X2=0 $Y2=0
cc_3870 N_A_5803_265#_c_4733_n N_S[4]_c_4988_n 0.00603996f $X=31.805 $Y=0.445
+ $X2=0 $Y2=0
cc_3871 N_A_5803_265#_c_4735_n N_S[4]_c_4988_n 9.67113e-19 $X=31.765 $Y=0.825
+ $X2=0 $Y2=0
cc_3872 N_A_5803_265#_c_4734_n N_S[4]_c_4989_n 0.00429801f $X=31.725 $Y=1.065
+ $X2=0 $Y2=0
cc_3873 N_A_5803_265#_c_4735_n N_S[4]_c_4989_n 0.0111895f $X=31.765 $Y=0.825
+ $X2=0 $Y2=0
cc_3874 N_A_5803_265#_c_4733_n N_S[4]_c_4990_n 0.00207203f $X=31.805 $Y=0.445
+ $X2=0 $Y2=0
cc_3875 N_A_5803_265#_c_4734_n N_S[4]_c_4991_n 0.00289358f $X=31.725 $Y=1.065
+ $X2=25.99 $Y2=4.8
cc_3876 N_A_5803_265#_c_4750_n N_S[4]_c_4991_n 0.0128834f $X=31.805 $Y=1.77
+ $X2=25.99 $Y2=4.8
cc_3877 N_A_5803_265#_c_4736_n N_S[4]_c_4991_n 0.00416423f $X=31.725 $Y=1.23
+ $X2=25.99 $Y2=4.8
cc_3878 N_A_5803_265#_c_4752_n N_S[4]_c_4991_n 0.00454075f $X=31.805 $Y=1.605
+ $X2=25.99 $Y2=4.8
cc_3879 N_A_5803_265#_c_4734_n N_S[4]_c_4995_n 0.00268644f $X=31.725 $Y=1.065
+ $X2=0 $Y2=0
cc_3880 N_A_5803_265#_c_4735_n N_S[4]_c_4995_n 0.00426435f $X=31.765 $Y=0.825
+ $X2=0 $Y2=0
cc_3881 N_A_5803_265#_c_4734_n S[4] 0.00541767f $X=31.725 $Y=1.065 $X2=0 $Y2=0
cc_3882 N_A_5803_265#_c_4736_n S[4] 0.0228692f $X=31.725 $Y=1.23 $X2=0 $Y2=0
cc_3883 N_A_5803_265#_c_4738_n N_VPWR_c_7271_n 0.00324472f $X=29.115 $Y=1.475
+ $X2=0 $Y2=0
cc_3884 N_A_5803_265#_c_4745_n N_VPWR_c_7273_n 0.00367058f $X=30.525 $Y=1.475
+ $X2=0 $Y2=0
cc_3885 N_A_5803_265#_c_4731_n N_VPWR_c_7273_n 0.0193185f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3886 N_A_5803_265#_c_4732_n N_VPWR_c_7273_n 6.4101e-19 $X=31.095 $Y=1.23
+ $X2=0 $Y2=0
cc_3887 N_A_5803_265#_c_4750_n N_VPWR_c_7273_n 0.0316788f $X=31.805 $Y=1.77
+ $X2=0 $Y2=0
cc_3888 N_A_5803_265#_c_4750_n N_VPWR_c_7275_n 0.0356181f $X=31.805 $Y=1.77
+ $X2=0 $Y2=0
cc_3889 N_A_5803_265#_c_4750_n N_VPWR_c_7331_n 0.0233824f $X=31.805 $Y=1.77
+ $X2=0 $Y2=0
cc_3890 N_A_5803_265#_c_4738_n VPWR 0.00473731f $X=29.115 $Y=1.475 $X2=0 $Y2=0
cc_3891 N_A_5803_265#_c_4741_n VPWR 0.00362156f $X=29.585 $Y=1.475 $X2=0 $Y2=0
cc_3892 N_A_5803_265#_c_4743_n VPWR 0.00362156f $X=30.055 $Y=1.475 $X2=0 $Y2=0
cc_3893 N_A_5803_265#_c_4745_n VPWR 0.00473731f $X=30.525 $Y=1.475 $X2=0 $Y2=0
cc_3894 N_A_5803_265#_c_4750_n VPWR 0.00593513f $X=31.805 $Y=1.77 $X2=0 $Y2=0
cc_3895 N_A_5803_265#_c_4742_n N_Z_c_9024_n 0.00762343f $X=29.965 $Y=1.4 $X2=0
+ $Y2=0
cc_3896 N_A_5803_265#_c_4746_n N_Z_c_9024_n 0.00704092f $X=29.585 $Y=1.4 $X2=0
+ $Y2=0
cc_3897 N_A_5803_265#_c_4740_n N_Z_c_9071_n 0.00248496f $X=29.205 $Y=1.4 $X2=0
+ $Y2=0
cc_3898 N_A_5803_265#_c_4739_n N_Z_c_9074_n 0.00678861f $X=29.495 $Y=1.4 $X2=0
+ $Y2=0
cc_3899 N_A_5803_265#_c_4740_n N_Z_c_9074_n 0.00239476f $X=29.205 $Y=1.4 $X2=0
+ $Y2=0
cc_3900 N_A_5803_265#_c_4746_n N_Z_c_9074_n 2.98555e-19 $X=29.585 $Y=1.4 $X2=0
+ $Y2=0
cc_3901 N_A_5803_265#_c_4742_n N_Z_c_9076_n 0.00145542f $X=29.965 $Y=1.4 $X2=0
+ $Y2=0
cc_3902 N_A_5803_265#_c_4744_n N_Z_c_9076_n 0.00597584f $X=30.435 $Y=1.4 $X2=0
+ $Y2=0
cc_3903 N_A_5803_265#_c_4747_n N_Z_c_9076_n 0.00909323f $X=30.055 $Y=1.4 $X2=0
+ $Y2=0
cc_3904 N_A_5803_265#_c_4731_n N_Z_c_9076_n 0.0266078f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3905 N_A_5803_265#_c_4737_n N_Z_c_9076_n 0.00747617f $X=30.845 $Y=1.23 $X2=0
+ $Y2=0
cc_3906 N_A_5803_265#_c_4738_n N_Z_c_9121_n 0.00834829f $X=29.115 $Y=1.475 $X2=0
+ $Y2=0
cc_3907 N_A_5803_265#_c_4745_n N_Z_c_9125_n 0.00795576f $X=30.525 $Y=1.475 $X2=0
+ $Y2=0
cc_3908 N_A_5803_265#_c_4731_n N_Z_c_9125_n 0.0186685f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3909 N_A_5803_265#_c_4750_n N_Z_c_9125_n 0.0329704f $X=31.805 $Y=1.77 $X2=0
+ $Y2=0
cc_3910 N_A_5803_265#_c_4737_n N_Z_c_9125_n 2.19754e-19 $X=30.845 $Y=1.23 $X2=0
+ $Y2=0
cc_3911 N_A_5803_265#_c_4741_n Z 0.00372458f $X=29.585 $Y=1.475 $X2=0 $Y2=0
cc_3912 N_A_5803_265#_c_4743_n Z 0.00372248f $X=30.055 $Y=1.475 $X2=0 $Y2=0
cc_3913 N_A_5803_265#_c_4738_n N_Z_c_9139_n 0.0199111f $X=29.115 $Y=1.475 $X2=0
+ $Y2=0
cc_3914 N_A_5803_265#_c_4739_n N_Z_c_9139_n 0.00560592f $X=29.495 $Y=1.4 $X2=0
+ $Y2=0
cc_3915 N_A_5803_265#_c_4740_n N_Z_c_9139_n 0.00474497f $X=29.205 $Y=1.4 $X2=0
+ $Y2=0
cc_3916 N_A_5803_265#_c_4741_n N_Z_c_9139_n 0.0181262f $X=29.585 $Y=1.475 $X2=0
+ $Y2=0
cc_3917 N_A_5803_265#_c_4743_n N_Z_c_9139_n 9.74366e-19 $X=30.055 $Y=1.475 $X2=0
+ $Y2=0
cc_3918 N_A_5803_265#_c_4746_n N_Z_c_9139_n 0.00415268f $X=29.585 $Y=1.4 $X2=0
+ $Y2=0
cc_3919 N_A_5803_265#_c_4741_n N_Z_c_9140_n 9.74366e-19 $X=29.585 $Y=1.475 $X2=0
+ $Y2=0
cc_3920 N_A_5803_265#_c_4743_n N_Z_c_9140_n 0.0181262f $X=30.055 $Y=1.475 $X2=0
+ $Y2=0
cc_3921 N_A_5803_265#_c_4744_n N_Z_c_9140_n 0.00560592f $X=30.435 $Y=1.4 $X2=0
+ $Y2=0
cc_3922 N_A_5803_265#_c_4745_n N_Z_c_9140_n 0.0221748f $X=30.525 $Y=1.475 $X2=0
+ $Y2=0
cc_3923 N_A_5803_265#_c_4747_n N_Z_c_9140_n 0.00181273f $X=30.055 $Y=1.4 $X2=0
+ $Y2=0
cc_3924 N_A_5803_265#_c_4731_n N_Z_c_9140_n 0.00240108f $X=31.64 $Y=1.23 $X2=0
+ $Y2=0
cc_3925 N_A_5803_265#_c_4737_n N_Z_c_9140_n 0.00425035f $X=30.845 $Y=1.23 $X2=0
+ $Y2=0
cc_3926 N_A_5803_265#_c_4738_n N_A_5361_297#_c_11677_n 0.00151141f $X=29.115
+ $Y=1.475 $X2=0 $Y2=0
cc_3927 N_A_5803_265#_c_4738_n N_A_5361_297#_c_11706_n 0.00307958f $X=29.115
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_3928 N_A_5803_265#_c_4741_n N_A_5361_297#_c_11706_n 0.00307958f $X=29.585
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_3929 N_A_5803_265#_c_4743_n N_A_5361_297#_c_11708_n 0.00307958f $X=30.055
+ $Y=1.475 $X2=0 $Y2=0
cc_3930 N_A_5803_265#_c_4745_n N_A_5361_297#_c_11708_n 0.00307958f $X=30.525
+ $Y=1.475 $X2=0 $Y2=0
cc_3931 N_A_5803_265#_c_4738_n N_A_5361_297#_c_11679_n 0.00554566f $X=29.115
+ $Y=1.475 $X2=0 $Y2=0
cc_3932 N_A_5803_265#_c_4741_n N_A_5361_297#_c_11680_n 0.00210632f $X=29.585
+ $Y=1.475 $X2=0 $Y2=0
cc_3933 N_A_5803_265#_c_4742_n N_A_5361_297#_c_11680_n 0.00251792f $X=29.965
+ $Y=1.4 $X2=0 $Y2=0
cc_3934 N_A_5803_265#_c_4743_n N_A_5361_297#_c_11680_n 0.00210632f $X=30.055
+ $Y=1.475 $X2=0 $Y2=0
cc_3935 N_A_5803_265#_c_4745_n N_A_5361_297#_c_11681_n 0.00499839f $X=30.525
+ $Y=1.475 $X2=0 $Y2=0
cc_3936 N_A_5803_265#_c_4731_n N_A_5361_297#_c_11681_n 0.0218124f $X=31.64
+ $Y=1.23 $X2=0 $Y2=0
cc_3937 N_A_5803_265#_c_4732_n N_A_5361_297#_c_11681_n 5.74251e-19 $X=31.095
+ $Y=1.23 $X2=0 $Y2=0
cc_3938 N_A_5803_265#_c_4737_n N_A_5361_297#_c_11681_n 0.00561627f $X=30.845
+ $Y=1.23 $X2=0 $Y2=0
cc_3939 N_A_5803_265#_c_4731_n N_VGND_c_12747_n 0.0123065f $X=31.64 $Y=1.23
+ $X2=0 $Y2=0
cc_3940 N_A_5803_265#_c_4732_n N_VGND_c_12747_n 2.04129e-19 $X=31.095 $Y=1.23
+ $X2=0 $Y2=0
cc_3941 N_A_5803_265#_c_4733_n N_VGND_c_12831_n 0.0129994f $X=31.805 $Y=0.445
+ $X2=0 $Y2=0
cc_3942 N_A_5803_265#_M1037_s VGND 0.00394793f $X=31.67 $Y=0.235 $X2=0 $Y2=0
cc_3943 N_A_5803_265#_c_4733_n VGND 0.00927134f $X=31.805 $Y=0.445 $X2=0 $Y2=0
cc_3944 N_A_5803_265#_c_4746_n N_A_5363_47#_c_14733_n 7.0477e-19 $X=29.585
+ $Y=1.4 $X2=0 $Y2=0
cc_3945 N_A_5803_265#_c_4731_n N_A_5363_47#_c_14711_n 0.0028695f $X=31.64
+ $Y=1.23 $X2=25.99 $Y2=4.93
cc_3946 N_A_5803_265#_c_4737_n N_A_5363_47#_c_14711_n 0.00589316f $X=30.845
+ $Y=1.23 $X2=25.99 $Y2=4.93
cc_3947 N_A_5803_793#_c_4859_n N_S[12]_c_5092_n 0.00507426f $X=29.205 $Y=4.04
+ $X2=0 $Y2=0
cc_3948 N_A_5803_793#_c_4858_n N_S[12]_c_5095_n 0.00509391f $X=29.495 $Y=4.04
+ $X2=0 $Y2=0
cc_3949 N_A_5803_793#_c_4861_n N_S[12]_c_5097_n 0.00509204f $X=29.965 $Y=4.04
+ $X2=25.905 $Y2=4.845
cc_3950 N_A_5803_793#_c_4863_n N_S[12]_c_5099_n 0.00507688f $X=30.435 $Y=4.04
+ $X2=0 $Y2=0
cc_3951 N_A_5803_793#_c_4852_n N_S[12]_c_5101_n 6.53442e-19 $X=31.765 $Y=4.74
+ $X2=0 $Y2=0
cc_3952 N_A_5803_793#_c_4850_n N_S[12]_c_5103_n 0.0103812f $X=31.64 $Y=4.21
+ $X2=0 $Y2=0
cc_3953 N_A_5803_793#_c_4851_n N_S[12]_c_5103_n 0.0179529f $X=31.095 $Y=4.21
+ $X2=0 $Y2=0
cc_3954 N_A_5803_793#_c_4870_n N_S[12]_c_5113_n 0.00508008f $X=31.725 $Y=4.045
+ $X2=0 $Y2=0
cc_3955 N_A_5803_793#_c_4856_n N_S[12]_c_5113_n 0.00262132f $X=30.845 $Y=4.21
+ $X2=0 $Y2=0
cc_3956 N_A_5803_793#_c_4850_n N_S[12]_c_5104_n 0.0206368f $X=31.64 $Y=4.21
+ $X2=0 $Y2=0
cc_3957 N_A_5803_793#_c_4851_n N_S[12]_c_5104_n 0.0175393f $X=31.095 $Y=4.21
+ $X2=0 $Y2=0
cc_3958 N_A_5803_793#_c_4870_n N_S[12]_c_5104_n 0.00255921f $X=31.725 $Y=4.045
+ $X2=0 $Y2=0
cc_3959 N_A_5803_793#_c_4854_n N_S[12]_c_5104_n 0.00322131f $X=31.725 $Y=4.21
+ $X2=0 $Y2=0
cc_3960 N_A_5803_793#_c_4855_n N_S[12]_c_5104_n 0.0085951f $X=31.765 $Y=4.615
+ $X2=0 $Y2=0
cc_3961 N_A_5803_793#_c_4869_n N_S[12]_c_5115_n 0.00970559f $X=31.805 $Y=3.14
+ $X2=0 $Y2=0
cc_3962 N_A_5803_793#_c_4870_n N_S[12]_c_5115_n 0.00254107f $X=31.725 $Y=4.045
+ $X2=0 $Y2=0
cc_3963 N_A_5803_793#_c_4871_n N_S[12]_c_5115_n 0.00216424f $X=31.805 $Y=3.835
+ $X2=0 $Y2=0
cc_3964 N_A_5803_793#_c_4852_n N_S[12]_c_5105_n 9.67113e-19 $X=31.765 $Y=4.74
+ $X2=0 $Y2=0
cc_3965 N_A_5803_793#_c_4853_n N_S[12]_c_5105_n 0.00603996f $X=31.805 $Y=4.995
+ $X2=0 $Y2=0
cc_3966 N_A_5803_793#_c_4852_n N_S[12]_c_5106_n 0.0111895f $X=31.765 $Y=4.74
+ $X2=0 $Y2=0
cc_3967 N_A_5803_793#_c_4855_n N_S[12]_c_5106_n 0.00429801f $X=31.765 $Y=4.615
+ $X2=0 $Y2=0
cc_3968 N_A_5803_793#_c_4870_n N_S[12]_c_5107_n 0.00336772f $X=31.725 $Y=4.045
+ $X2=0 $Y2=0
cc_3969 N_A_5803_793#_c_4852_n N_S[12]_c_5107_n 0.00207203f $X=31.765 $Y=4.74
+ $X2=0 $Y2=0
cc_3970 N_A_5803_793#_c_4871_n N_S[12]_c_5107_n 5.48523e-19 $X=31.805 $Y=3.835
+ $X2=0 $Y2=0
cc_3971 N_A_5803_793#_c_4854_n N_S[12]_c_5107_n 0.00416423f $X=31.725 $Y=4.21
+ $X2=0 $Y2=0
cc_3972 N_A_5803_793#_c_4855_n N_S[12]_c_5107_n 0.00289358f $X=31.765 $Y=4.615
+ $X2=0 $Y2=0
cc_3973 N_A_5803_793#_c_4869_n N_S[12]_c_5117_n 0.00929139f $X=31.805 $Y=3.14
+ $X2=25.99 $Y2=4.8
cc_3974 N_A_5803_793#_c_4870_n N_S[12]_c_5117_n 0.00117303f $X=31.725 $Y=4.045
+ $X2=25.99 $Y2=4.8
cc_3975 N_A_5803_793#_c_4871_n N_S[12]_c_5117_n 0.00304348f $X=31.805 $Y=3.835
+ $X2=25.99 $Y2=4.8
cc_3976 N_A_5803_793#_c_4852_n N_S[12]_c_5111_n 0.00426435f $X=31.765 $Y=4.74
+ $X2=0 $Y2=0
cc_3977 N_A_5803_793#_c_4855_n N_S[12]_c_5111_n 0.00268644f $X=31.765 $Y=4.615
+ $X2=0 $Y2=0
cc_3978 N_A_5803_793#_c_4854_n S[12] 0.0228692f $X=31.725 $Y=4.21 $X2=0 $Y2=0
cc_3979 N_A_5803_793#_c_4855_n S[12] 0.00541767f $X=31.765 $Y=4.615 $X2=0 $Y2=0
cc_3980 N_A_5803_793#_c_4857_n N_VPWR_c_7272_n 0.00324472f $X=29.115 $Y=3.965
+ $X2=0 $Y2=0
cc_3981 N_A_5803_793#_c_4864_n N_VPWR_c_7274_n 0.00367058f $X=30.525 $Y=3.965
+ $X2=0 $Y2=0
cc_3982 N_A_5803_793#_c_4850_n N_VPWR_c_7274_n 0.0193185f $X=31.64 $Y=4.21 $X2=0
+ $Y2=0
cc_3983 N_A_5803_793#_c_4851_n N_VPWR_c_7274_n 6.4101e-19 $X=31.095 $Y=4.21
+ $X2=0 $Y2=0
cc_3984 N_A_5803_793#_c_4869_n N_VPWR_c_7274_n 0.0316788f $X=31.805 $Y=3.14
+ $X2=0 $Y2=0
cc_3985 N_A_5803_793#_c_4869_n N_VPWR_c_7276_n 0.0356181f $X=31.805 $Y=3.14
+ $X2=0 $Y2=0
cc_3986 N_A_5803_793#_c_4869_n N_VPWR_c_7331_n 0.0233824f $X=31.805 $Y=3.14
+ $X2=0 $Y2=0
cc_3987 N_A_5803_793#_c_4857_n VPWR 0.00473731f $X=29.115 $Y=3.965 $X2=0 $Y2=0
cc_3988 N_A_5803_793#_c_4860_n VPWR 0.00362156f $X=29.585 $Y=3.965 $X2=0 $Y2=0
cc_3989 N_A_5803_793#_c_4862_n VPWR 0.00362156f $X=30.055 $Y=3.965 $X2=0 $Y2=0
cc_3990 N_A_5803_793#_c_4864_n VPWR 0.00473731f $X=30.525 $Y=3.965 $X2=0 $Y2=0
cc_3991 N_A_5803_793#_c_4869_n VPWR 0.00593513f $X=31.805 $Y=3.14 $X2=0 $Y2=0
cc_3992 N_A_5803_793#_c_4861_n N_Z_c_9025_n 0.00762343f $X=29.965 $Y=4.04 $X2=0
+ $Y2=0
cc_3993 N_A_5803_793#_c_4865_n N_Z_c_9025_n 0.00704092f $X=29.585 $Y=4.04 $X2=0
+ $Y2=0
cc_3994 N_A_5803_793#_c_4859_n N_Z_c_9072_n 0.00248496f $X=29.205 $Y=4.04 $X2=0
+ $Y2=0
cc_3995 N_A_5803_793#_c_4858_n N_Z_c_9075_n 0.00678861f $X=29.495 $Y=4.04 $X2=0
+ $Y2=0
cc_3996 N_A_5803_793#_c_4859_n N_Z_c_9075_n 0.00239476f $X=29.205 $Y=4.04 $X2=0
+ $Y2=0
cc_3997 N_A_5803_793#_c_4865_n N_Z_c_9075_n 2.98555e-19 $X=29.585 $Y=4.04 $X2=0
+ $Y2=0
cc_3998 N_A_5803_793#_c_4861_n N_Z_c_9077_n 0.00145542f $X=29.965 $Y=4.04 $X2=0
+ $Y2=0
cc_3999 N_A_5803_793#_c_4863_n N_Z_c_9077_n 0.00597584f $X=30.435 $Y=4.04 $X2=0
+ $Y2=0
cc_4000 N_A_5803_793#_c_4866_n N_Z_c_9077_n 0.00909323f $X=30.055 $Y=4.04 $X2=0
+ $Y2=0
cc_4001 N_A_5803_793#_c_4850_n N_Z_c_9077_n 0.0266078f $X=31.64 $Y=4.21 $X2=0
+ $Y2=0
cc_4002 N_A_5803_793#_c_4856_n N_Z_c_9077_n 0.00747617f $X=30.845 $Y=4.21 $X2=0
+ $Y2=0
cc_4003 N_A_5803_793#_c_4857_n N_Z_c_9123_n 0.00834829f $X=29.115 $Y=3.965 $X2=0
+ $Y2=0
cc_4004 N_A_5803_793#_c_4864_n N_Z_c_9126_n 0.00795576f $X=30.525 $Y=3.965 $X2=0
+ $Y2=0
cc_4005 N_A_5803_793#_c_4850_n N_Z_c_9126_n 0.0186685f $X=31.64 $Y=4.21 $X2=0
+ $Y2=0
cc_4006 N_A_5803_793#_c_4869_n N_Z_c_9126_n 0.0329704f $X=31.805 $Y=3.14 $X2=0
+ $Y2=0
cc_4007 N_A_5803_793#_c_4856_n N_Z_c_9126_n 2.19754e-19 $X=30.845 $Y=4.21 $X2=0
+ $Y2=0
cc_4008 N_A_5803_793#_c_4860_n Z 0.00372458f $X=29.585 $Y=3.965 $X2=0 $Y2=0
cc_4009 N_A_5803_793#_c_4862_n Z 0.00372248f $X=30.055 $Y=3.965 $X2=0 $Y2=0
cc_4010 N_A_5803_793#_c_4857_n N_Z_c_9139_n 0.0199111f $X=29.115 $Y=3.965 $X2=0
+ $Y2=0
cc_4011 N_A_5803_793#_c_4858_n N_Z_c_9139_n 0.00560592f $X=29.495 $Y=4.04 $X2=0
+ $Y2=0
cc_4012 N_A_5803_793#_c_4859_n N_Z_c_9139_n 0.00474497f $X=29.205 $Y=4.04 $X2=0
+ $Y2=0
cc_4013 N_A_5803_793#_c_4860_n N_Z_c_9139_n 0.0181262f $X=29.585 $Y=3.965 $X2=0
+ $Y2=0
cc_4014 N_A_5803_793#_c_4862_n N_Z_c_9139_n 9.74366e-19 $X=30.055 $Y=3.965 $X2=0
+ $Y2=0
cc_4015 N_A_5803_793#_c_4865_n N_Z_c_9139_n 0.00415268f $X=29.585 $Y=4.04 $X2=0
+ $Y2=0
cc_4016 N_A_5803_793#_c_4860_n N_Z_c_9140_n 9.74366e-19 $X=29.585 $Y=3.965 $X2=0
+ $Y2=0
cc_4017 N_A_5803_793#_c_4862_n N_Z_c_9140_n 0.0181262f $X=30.055 $Y=3.965 $X2=0
+ $Y2=0
cc_4018 N_A_5803_793#_c_4863_n N_Z_c_9140_n 0.00560592f $X=30.435 $Y=4.04 $X2=0
+ $Y2=0
cc_4019 N_A_5803_793#_c_4864_n N_Z_c_9140_n 0.0221748f $X=30.525 $Y=3.965 $X2=0
+ $Y2=0
cc_4020 N_A_5803_793#_c_4866_n N_Z_c_9140_n 0.00181273f $X=30.055 $Y=4.04 $X2=0
+ $Y2=0
cc_4021 N_A_5803_793#_c_4850_n N_Z_c_9140_n 0.00240108f $X=31.64 $Y=4.21 $X2=0
+ $Y2=0
cc_4022 N_A_5803_793#_c_4856_n N_Z_c_9140_n 0.00425035f $X=30.845 $Y=4.21 $X2=0
+ $Y2=0
cc_4023 N_A_5803_793#_c_4857_n N_A_5361_591#_c_11805_n 0.00151141f $X=29.115
+ $Y=3.965 $X2=0 $Y2=0
cc_4024 N_A_5803_793#_c_4857_n N_A_5361_591#_c_11834_n 0.00307958f $X=29.115
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_4025 N_A_5803_793#_c_4860_n N_A_5361_591#_c_11834_n 0.00307958f $X=29.585
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_4026 N_A_5803_793#_c_4862_n N_A_5361_591#_c_11836_n 0.00307958f $X=30.055
+ $Y=3.965 $X2=0 $Y2=0
cc_4027 N_A_5803_793#_c_4864_n N_A_5361_591#_c_11836_n 0.00307958f $X=30.525
+ $Y=3.965 $X2=0 $Y2=0
cc_4028 N_A_5803_793#_c_4857_n N_A_5361_591#_c_11807_n 0.00554566f $X=29.115
+ $Y=3.965 $X2=0 $Y2=0
cc_4029 N_A_5803_793#_c_4860_n N_A_5361_591#_c_11808_n 0.00210632f $X=29.585
+ $Y=3.965 $X2=0 $Y2=0
cc_4030 N_A_5803_793#_c_4861_n N_A_5361_591#_c_11808_n 0.00251792f $X=29.965
+ $Y=4.04 $X2=0 $Y2=0
cc_4031 N_A_5803_793#_c_4862_n N_A_5361_591#_c_11808_n 0.00210632f $X=30.055
+ $Y=3.965 $X2=0 $Y2=0
cc_4032 N_A_5803_793#_c_4864_n N_A_5361_591#_c_11809_n 0.00499839f $X=30.525
+ $Y=3.965 $X2=0 $Y2=0
cc_4033 N_A_5803_793#_c_4850_n N_A_5361_591#_c_11809_n 0.0218124f $X=31.64
+ $Y=4.21 $X2=0 $Y2=0
cc_4034 N_A_5803_793#_c_4851_n N_A_5361_591#_c_11809_n 5.74251e-19 $X=31.095
+ $Y=4.21 $X2=0 $Y2=0
cc_4035 N_A_5803_793#_c_4856_n N_A_5361_591#_c_11809_n 0.00561627f $X=30.845
+ $Y=4.21 $X2=0 $Y2=0
cc_4036 N_A_5803_793#_c_4850_n N_VGND_c_12748_n 0.0123065f $X=31.64 $Y=4.21
+ $X2=0 $Y2=0
cc_4037 N_A_5803_793#_c_4851_n N_VGND_c_12748_n 2.04129e-19 $X=31.095 $Y=4.21
+ $X2=0 $Y2=0
cc_4038 N_A_5803_793#_c_4853_n N_VGND_c_12833_n 0.0129994f $X=31.805 $Y=4.995
+ $X2=0 $Y2=0
cc_4039 N_A_5803_793#_M1188_d VGND 0.00394793f $X=31.67 $Y=4.785 $X2=0 $Y2=0
cc_4040 N_A_5803_793#_c_4853_n VGND 0.00927134f $X=31.805 $Y=4.995 $X2=0 $Y2=0
cc_4041 N_A_5803_793#_c_4865_n N_A_5363_911#_c_14812_n 7.0477e-19 $X=29.585
+ $Y=4.04 $X2=0 $Y2=0
cc_4042 N_A_5803_793#_c_4850_n N_A_5363_911#_c_14793_n 0.0028695f $X=31.64
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_4043 N_A_5803_793#_c_4856_n N_A_5363_911#_c_14793_n 0.00589316f $X=30.845
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_4044 N_S[4]_c_4998_n N_S[12]_c_5115_n 0.0130744f $X=31.57 $Y=1.55 $X2=0 $Y2=0
cc_4045 N_S[4]_c_4991_n N_S[12]_c_5117_n 0.0130744f $X=32.04 $Y=1.55 $X2=25.99
+ $Y2=4.8
cc_4046 N_S[4]_c_4991_n N_S[5]_c_5217_n 0.0215827f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4047 S[4] N_S[5]_c_5217_n 0.00113563f $X=32.345 $Y=1.105 $X2=0 $Y2=0
cc_4048 N_S[4]_c_4991_n N_S[5]_c_5238_n 0.00113563f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4049 S[4] N_S[5]_c_5238_n 0.0301108f $X=32.345 $Y=1.105 $X2=0 $Y2=0
cc_4050 N_S[4]_c_4998_n N_VPWR_c_7273_n 0.00950399f $X=31.57 $Y=1.55 $X2=0 $Y2=0
cc_4051 N_S[4]_c_4991_n N_VPWR_c_7275_n 0.016386f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4052 S[4] N_VPWR_c_7275_n 0.0157609f $X=32.345 $Y=1.105 $X2=0 $Y2=0
cc_4053 N_S[4]_c_4998_n N_VPWR_c_7331_n 0.0035837f $X=31.57 $Y=1.55 $X2=0 $Y2=0
cc_4054 N_S[4]_c_4991_n N_VPWR_c_7331_n 0.0035837f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4055 N_S[4]_c_4998_n VPWR 0.00711603f $X=31.57 $Y=1.55 $X2=0 $Y2=0
cc_4056 N_S[4]_c_4991_n VPWR 0.0070533f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4057 N_S[4]_c_4975_n N_Z_c_9023_n 0.002324f $X=29.04 $Y=0.255 $X2=0 $Y2=0
cc_4058 N_S[4]_c_4978_n N_Z_c_9023_n 0.00283489f $X=29.46 $Y=0.255 $X2=0 $Y2=0
cc_4059 N_S[4]_c_4978_n N_Z_c_9024_n 3.10191e-19 $X=29.46 $Y=0.255 $X2=0 $Y2=0
cc_4060 N_S[4]_c_4980_n N_Z_c_9024_n 0.00190704f $X=29.88 $Y=0.255 $X2=0 $Y2=0
cc_4061 N_S[4]_c_4978_n N_Z_c_9026_n 6.35774e-19 $X=29.46 $Y=0.255 $X2=0 $Y2=0
cc_4062 N_S[4]_c_4980_n N_Z_c_9026_n 0.0077801f $X=29.88 $Y=0.255 $X2=0 $Y2=0
cc_4063 N_S[4]_c_4982_n N_Z_c_9026_n 0.0134253f $X=30.3 $Y=0.255 $X2=0 $Y2=0
cc_4064 N_S[4]_c_4975_n N_Z_c_9071_n 0.00443615f $X=29.04 $Y=0.255 $X2=0 $Y2=0
cc_4065 N_S[4]_c_4978_n N_Z_c_9071_n 0.00462308f $X=29.46 $Y=0.255 $X2=0 $Y2=0
cc_4066 N_S[4]_c_4980_n N_Z_c_9071_n 6.35664e-19 $X=29.88 $Y=0.255 $X2=0 $Y2=0
cc_4067 N_S[4]_c_4978_n N_Z_c_9074_n 0.00180363f $X=29.46 $Y=0.255 $X2=0 $Y2=0
cc_4068 N_S[4]_c_4982_n N_Z_c_9076_n 0.00216436f $X=30.3 $Y=0.255 $X2=0 $Y2=0
cc_4069 N_S[4]_c_4998_n N_Z_c_9125_n 0.00478771f $X=31.57 $Y=1.55 $X2=0 $Y2=0
cc_4070 N_S[4]_c_4991_n N_Z_c_9125_n 0.00760321f $X=32.04 $Y=1.55 $X2=0 $Y2=0
cc_4071 S[4] N_Z_c_9125_n 0.010609f $X=32.345 $Y=1.105 $X2=0 $Y2=0
cc_4072 N_S[4]_c_4975_n N_A_5361_297#_c_11677_n 0.00168571f $X=29.04 $Y=0.255
+ $X2=0 $Y2=0
cc_4073 N_S[4]_c_4998_n N_A_5361_297#_c_11681_n 0.00239129f $X=31.57 $Y=1.55
+ $X2=0 $Y2=0
cc_4074 N_S[4]_c_4975_n N_VGND_c_12745_n 5.5039e-19 $X=29.04 $Y=0.255 $X2=0
+ $Y2=0
cc_4075 N_S[4]_c_4977_n N_VGND_c_12745_n 0.0028166f $X=29.115 $Y=0.18 $X2=0
+ $Y2=0
cc_4076 N_S[4]_c_4983_n N_VGND_c_12747_n 0.00862298f $X=30.985 $Y=0.18 $X2=0
+ $Y2=0
cc_4077 N_S[4]_c_4985_n N_VGND_c_12747_n 0.00525833f $X=31.47 $Y=0.81 $X2=0
+ $Y2=0
cc_4078 N_S[4]_c_4988_n N_VGND_c_12747_n 0.00173127f $X=31.595 $Y=0.735 $X2=0
+ $Y2=0
cc_4079 N_S[4]_c_4990_n N_VGND_c_12749_n 0.00374526f $X=32.015 $Y=0.735 $X2=0
+ $Y2=0
cc_4080 N_S[4]_c_4991_n N_VGND_c_12749_n 0.00578076f $X=32.04 $Y=1.55 $X2=0
+ $Y2=0
cc_4081 S[4] N_VGND_c_12749_n 0.0116413f $X=32.345 $Y=1.105 $X2=0 $Y2=0
cc_4082 N_S[4]_c_4977_n N_VGND_c_12827_n 0.0559651f $X=29.115 $Y=0.18 $X2=0
+ $Y2=0
cc_4083 N_S[4]_c_4988_n N_VGND_c_12831_n 0.00542362f $X=31.595 $Y=0.735 $X2=0
+ $Y2=0
cc_4084 N_S[4]_c_4989_n N_VGND_c_12831_n 2.16067e-19 $X=31.94 $Y=0.81 $X2=0
+ $Y2=0
cc_4085 N_S[4]_c_4990_n N_VGND_c_12831_n 0.00585385f $X=32.015 $Y=0.735 $X2=0
+ $Y2=0
cc_4086 N_S[4]_c_4976_n VGND 0.00642387f $X=29.385 $Y=0.18 $X2=0 $Y2=0
cc_4087 N_S[4]_c_4977_n VGND 0.00591981f $X=29.115 $Y=0.18 $X2=0 $Y2=0
cc_4088 N_S[4]_c_4979_n VGND 0.0064237f $X=29.805 $Y=0.18 $X2=0 $Y2=0
cc_4089 N_S[4]_c_4981_n VGND 0.00642387f $X=30.225 $Y=0.18 $X2=0 $Y2=0
cc_4090 N_S[4]_c_4983_n VGND 0.0345801f $X=30.985 $Y=0.18 $X2=0 $Y2=0
cc_4091 N_S[4]_c_4988_n VGND 0.00990284f $X=31.595 $Y=0.735 $X2=0 $Y2=0
cc_4092 N_S[4]_c_4990_n VGND 0.0119653f $X=32.015 $Y=0.735 $X2=0 $Y2=0
cc_4093 N_S[4]_c_4992_n VGND 0.00366655f $X=29.46 $Y=0.18 $X2=0 $Y2=0
cc_4094 N_S[4]_c_4993_n VGND 0.00366655f $X=29.88 $Y=0.18 $X2=0 $Y2=0
cc_4095 N_S[4]_c_4994_n VGND 0.00366655f $X=30.3 $Y=0.18 $X2=0 $Y2=0
cc_4096 N_S[4]_c_4975_n N_A_5363_47#_c_14706_n 0.00206084f $X=29.04 $Y=0.255
+ $X2=0 $Y2=0
cc_4097 N_S[4]_c_4975_n N_A_5363_47#_c_14708_n 0.0139014f $X=29.04 $Y=0.255
+ $X2=0 $Y2=0
cc_4098 N_S[4]_c_4976_n N_A_5363_47#_c_14708_n 0.00211351f $X=29.385 $Y=0.18
+ $X2=0 $Y2=0
cc_4099 N_S[4]_c_4978_n N_A_5363_47#_c_14708_n 0.0106826f $X=29.46 $Y=0.255
+ $X2=0 $Y2=0
cc_4100 N_S[4]_c_4980_n N_A_5363_47#_c_14710_n 0.0106844f $X=29.88 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_4101 N_S[4]_c_4981_n N_A_5363_47#_c_14710_n 0.00211351f $X=30.225 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_4102 N_S[4]_c_4982_n N_A_5363_47#_c_14710_n 0.0112916f $X=30.3 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_4103 N_S[4]_c_4983_n N_A_5363_47#_c_14710_n 0.00685838f $X=30.985 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_4104 N_S[4]_c_4984_n N_A_5363_47#_c_14710_n 0.00189496f $X=31.06 $Y=0.735
+ $X2=25.99 $Y2=4.8
cc_4105 N_S[4]_c_4984_n N_A_5363_47#_c_14711_n 0.00529837f $X=31.06 $Y=0.735
+ $X2=25.99 $Y2=4.93
cc_4106 N_S[4]_c_4979_n N_A_5363_47#_c_14746_n 0.0034777f $X=29.805 $Y=0.18
+ $X2=0 $Y2=0
cc_4107 N_S[12]_c_5107_n N_S[13]_c_5337_n 0.0215827f $X=32.015 $Y=4.705 $X2=0
+ $Y2=0
cc_4108 S[12] N_S[13]_c_5337_n 0.00113563f $X=32.345 $Y=4.165 $X2=0 $Y2=0
cc_4109 N_S[12]_c_5107_n N_S[13]_c_5357_n 0.00113563f $X=32.015 $Y=4.705 $X2=0
+ $Y2=0
cc_4110 S[12] N_S[13]_c_5357_n 0.0301108f $X=32.345 $Y=4.165 $X2=0 $Y2=0
cc_4111 N_S[12]_c_5115_n N_VPWR_c_7274_n 0.00950399f $X=31.57 $Y=3.89 $X2=0
+ $Y2=0
cc_4112 N_S[12]_c_5107_n N_VPWR_c_7276_n 0.00652399f $X=32.015 $Y=4.705 $X2=0
+ $Y2=0
cc_4113 N_S[12]_c_5117_n N_VPWR_c_7276_n 0.00986205f $X=32.04 $Y=3.89 $X2=0
+ $Y2=0
cc_4114 S[12] N_VPWR_c_7276_n 0.0157609f $X=32.345 $Y=4.165 $X2=0 $Y2=0
cc_4115 N_S[12]_c_5115_n N_VPWR_c_7331_n 0.0035837f $X=31.57 $Y=3.89 $X2=0 $Y2=0
cc_4116 N_S[12]_c_5117_n N_VPWR_c_7331_n 0.0035837f $X=32.04 $Y=3.89 $X2=0 $Y2=0
cc_4117 N_S[12]_c_5115_n VPWR 0.00711603f $X=31.57 $Y=3.89 $X2=0 $Y2=0
cc_4118 N_S[12]_c_5117_n VPWR 0.0070533f $X=32.04 $Y=3.89 $X2=0 $Y2=0
cc_4119 N_S[12]_c_5095_n N_Z_c_9025_n 3.10191e-19 $X=29.46 $Y=5.185 $X2=0 $Y2=0
cc_4120 N_S[12]_c_5097_n N_Z_c_9025_n 0.00190704f $X=29.88 $Y=5.185 $X2=0 $Y2=0
cc_4121 N_S[12]_c_5095_n N_Z_c_9027_n 6.35774e-19 $X=29.46 $Y=5.185 $X2=0 $Y2=0
cc_4122 N_S[12]_c_5097_n N_Z_c_9027_n 0.0077801f $X=29.88 $Y=5.185 $X2=0 $Y2=0
cc_4123 N_S[12]_c_5099_n N_Z_c_9027_n 0.0134253f $X=30.3 $Y=5.185 $X2=0 $Y2=0
cc_4124 N_S[12]_c_5092_n N_Z_c_9072_n 0.00443615f $X=29.04 $Y=5.185 $X2=0 $Y2=0
cc_4125 N_S[12]_c_5095_n N_Z_c_9072_n 0.00462308f $X=29.46 $Y=5.185 $X2=0 $Y2=0
cc_4126 N_S[12]_c_5092_n N_Z_c_9073_n 0.002324f $X=29.04 $Y=5.185 $X2=0 $Y2=0
cc_4127 N_S[12]_c_5095_n N_Z_c_9073_n 0.00283489f $X=29.46 $Y=5.185 $X2=0 $Y2=0
cc_4128 N_S[12]_c_5097_n N_Z_c_9073_n 6.35664e-19 $X=29.88 $Y=5.185 $X2=0 $Y2=0
cc_4129 N_S[12]_c_5095_n N_Z_c_9075_n 0.00180363f $X=29.46 $Y=5.185 $X2=0 $Y2=0
cc_4130 N_S[12]_c_5099_n N_Z_c_9077_n 0.00216436f $X=30.3 $Y=5.185 $X2=0 $Y2=0
cc_4131 N_S[12]_c_5113_n N_Z_c_9126_n 2.55735e-19 $X=31.57 $Y=3.99 $X2=0 $Y2=0
cc_4132 N_S[12]_c_5115_n N_Z_c_9126_n 0.00453198f $X=31.57 $Y=3.89 $X2=0 $Y2=0
cc_4133 N_S[12]_c_5107_n N_Z_c_9126_n 0.00258545f $X=32.015 $Y=4.705 $X2=0 $Y2=0
cc_4134 N_S[12]_c_5117_n N_Z_c_9126_n 0.00501777f $X=32.04 $Y=3.89 $X2=0 $Y2=0
cc_4135 S[12] N_Z_c_9126_n 0.010609f $X=32.345 $Y=4.165 $X2=0 $Y2=0
cc_4136 N_S[12]_c_5092_n N_A_5361_591#_c_11805_n 0.00168571f $X=29.04 $Y=5.185
+ $X2=0 $Y2=0
cc_4137 N_S[12]_c_5115_n N_A_5361_591#_c_11809_n 0.00239129f $X=31.57 $Y=3.89
+ $X2=0 $Y2=0
cc_4138 N_S[12]_c_5092_n N_VGND_c_12746_n 5.5039e-19 $X=29.04 $Y=5.185 $X2=0
+ $Y2=0
cc_4139 N_S[12]_c_5094_n N_VGND_c_12746_n 0.0028166f $X=29.115 $Y=5.26 $X2=0
+ $Y2=0
cc_4140 N_S[12]_c_5101_n N_VGND_c_12748_n 0.00862298f $X=31.06 $Y=5.185 $X2=0
+ $Y2=0
cc_4141 N_S[12]_c_5102_n N_VGND_c_12748_n 0.00525833f $X=31.47 $Y=4.63 $X2=0
+ $Y2=0
cc_4142 N_S[12]_c_5105_n N_VGND_c_12748_n 0.00173127f $X=31.595 $Y=4.705 $X2=0
+ $Y2=0
cc_4143 N_S[12]_c_5107_n N_VGND_c_12750_n 0.00952602f $X=32.015 $Y=4.705 $X2=0
+ $Y2=0
cc_4144 S[12] N_VGND_c_12750_n 0.0116413f $X=32.345 $Y=4.165 $X2=0 $Y2=0
cc_4145 N_S[12]_c_5094_n N_VGND_c_12829_n 0.0559651f $X=29.115 $Y=5.26 $X2=0
+ $Y2=0
cc_4146 N_S[12]_c_5105_n N_VGND_c_12833_n 0.00542362f $X=31.595 $Y=4.705 $X2=0
+ $Y2=0
cc_4147 N_S[12]_c_5106_n N_VGND_c_12833_n 2.16067e-19 $X=31.94 $Y=4.63 $X2=0
+ $Y2=0
cc_4148 N_S[12]_c_5107_n N_VGND_c_12833_n 0.00585385f $X=32.015 $Y=4.705 $X2=0
+ $Y2=0
cc_4149 N_S[12]_c_5093_n VGND 0.00642387f $X=29.385 $Y=5.26 $X2=0 $Y2=0
cc_4150 N_S[12]_c_5094_n VGND 0.00591981f $X=29.115 $Y=5.26 $X2=0 $Y2=0
cc_4151 N_S[12]_c_5096_n VGND 0.0064237f $X=29.805 $Y=5.26 $X2=0 $Y2=0
cc_4152 N_S[12]_c_5098_n VGND 0.00642387f $X=30.225 $Y=5.26 $X2=0 $Y2=0
cc_4153 N_S[12]_c_5100_n VGND 0.0345801f $X=30.985 $Y=5.26 $X2=0 $Y2=0
cc_4154 N_S[12]_c_5105_n VGND 0.00990284f $X=31.595 $Y=4.705 $X2=0 $Y2=0
cc_4155 N_S[12]_c_5107_n VGND 0.0119653f $X=32.015 $Y=4.705 $X2=0 $Y2=0
cc_4156 N_S[12]_c_5108_n VGND 0.00366655f $X=29.46 $Y=5.26 $X2=0 $Y2=0
cc_4157 N_S[12]_c_5109_n VGND 0.00366655f $X=29.88 $Y=5.26 $X2=0 $Y2=0
cc_4158 N_S[12]_c_5110_n VGND 0.00366655f $X=30.3 $Y=5.26 $X2=0 $Y2=0
cc_4159 N_S[12]_c_5092_n N_A_5363_911#_c_14788_n 0.00206084f $X=29.04 $Y=5.185
+ $X2=0 $Y2=0
cc_4160 N_S[12]_c_5092_n N_A_5363_911#_c_14790_n 0.0139014f $X=29.04 $Y=5.185
+ $X2=0 $Y2=0
cc_4161 N_S[12]_c_5093_n N_A_5363_911#_c_14790_n 0.00211351f $X=29.385 $Y=5.26
+ $X2=0 $Y2=0
cc_4162 N_S[12]_c_5095_n N_A_5363_911#_c_14790_n 0.0106826f $X=29.46 $Y=5.185
+ $X2=0 $Y2=0
cc_4163 N_S[12]_c_5097_n N_A_5363_911#_c_14792_n 0.0106844f $X=29.88 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_4164 N_S[12]_c_5098_n N_A_5363_911#_c_14792_n 0.00211351f $X=30.225 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_4165 N_S[12]_c_5099_n N_A_5363_911#_c_14792_n 0.0112916f $X=30.3 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_4166 N_S[12]_c_5100_n N_A_5363_911#_c_14792_n 0.00685838f $X=30.985 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_4167 N_S[12]_c_5101_n N_A_5363_911#_c_14792_n 0.00189496f $X=31.06 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_4168 N_S[12]_c_5103_n N_A_5363_911#_c_14793_n 0.00529837f $X=31.135 $Y=4.63
+ $X2=25.99 $Y2=4.8
cc_4169 N_S[12]_c_5096_n N_A_5363_911#_c_14825_n 0.0034777f $X=29.805 $Y=5.26
+ $X2=0 $Y2=0
cc_4170 N_S[5]_c_5218_n N_S[13]_c_5359_n 0.0130744f $X=33.28 $Y=1.55 $X2=0 $Y2=0
cc_4171 N_S[5]_c_5242_n N_S[13]_c_5363_n 0.0130744f $X=33.75 $Y=1.55 $X2=0 $Y2=0
cc_4172 N_S[5]_c_5227_n N_A_6674_325#_c_5473_n 0.00507688f $X=35.02 $Y=0.255
+ $X2=25.905 $Y2=0.425
cc_4173 N_S[5]_c_5222_n N_A_6674_325#_c_5465_n 0.00262132f $X=33.75 $Y=1.45
+ $X2=25.905 $Y2=4.845
cc_4174 N_S[5]_c_5229_n N_A_6674_325#_c_5476_n 0.00509204f $X=35.44 $Y=0.255
+ $X2=0 $Y2=0
cc_4175 N_S[5]_c_5233_n N_A_6674_325#_c_5478_n 0.00507426f $X=36.28 $Y=0.255
+ $X2=0 $Y2=0
cc_4176 N_S[5]_c_5231_n N_A_6674_325#_c_5481_n 0.00509391f $X=35.86 $Y=0.255
+ $X2=0 $Y2=0
cc_4177 N_S[5]_c_5218_n N_A_6674_325#_c_5482_n 0.0128834f $X=33.28 $Y=1.55 $X2=0
+ $Y2=0
cc_4178 N_S[5]_c_5242_n N_A_6674_325#_c_5482_n 0.0118698f $X=33.75 $Y=1.55 $X2=0
+ $Y2=0
cc_4179 N_S[5]_c_5219_n N_A_6674_325#_c_5466_n 0.00207203f $X=33.305 $Y=0.735
+ $X2=0 $Y2=0
cc_4180 N_S[5]_c_5221_n N_A_6674_325#_c_5466_n 0.00603996f $X=33.725 $Y=0.735
+ $X2=0 $Y2=0
cc_4181 N_S[5]_c_5224_n N_A_6674_325#_c_5466_n 6.53442e-19 $X=34.26 $Y=0.735
+ $X2=0 $Y2=0
cc_4182 N_S[5]_c_5218_n N_A_6674_325#_c_5467_n 0.00289358f $X=33.28 $Y=1.55
+ $X2=0 $Y2=0
cc_4183 N_S[5]_c_5220_n N_A_6674_325#_c_5467_n 0.00429801f $X=33.65 $Y=0.81
+ $X2=0 $Y2=0
cc_4184 N_S[5]_c_5222_n N_A_6674_325#_c_5467_n 0.0085951f $X=33.75 $Y=1.45 $X2=0
+ $Y2=0
cc_4185 N_S[5]_c_5234_n N_A_6674_325#_c_5467_n 0.00268644f $X=33.75 $Y=0.81
+ $X2=0 $Y2=0
cc_4186 N_S[5]_c_5238_n N_A_6674_325#_c_5467_n 0.00541767f $X=33.24 $Y=1.16
+ $X2=0 $Y2=0
cc_4187 N_S[5]_c_5222_n N_A_6674_325#_c_5468_n 0.0206368f $X=33.75 $Y=1.45 $X2=0
+ $Y2=0
cc_4188 N_S[5]_c_5223_n N_A_6674_325#_c_5468_n 0.0103812f $X=34.185 $Y=0.81
+ $X2=0 $Y2=0
cc_4189 N_S[5]_c_5218_n N_A_6674_325#_c_5484_n 0.00454075f $X=33.28 $Y=1.55
+ $X2=0 $Y2=0
cc_4190 N_S[5]_c_5222_n N_A_6674_325#_c_5484_n 0.00255921f $X=33.75 $Y=1.45
+ $X2=0 $Y2=0
cc_4191 N_S[5]_c_5242_n N_A_6674_325#_c_5484_n 0.00762115f $X=33.75 $Y=1.55
+ $X2=0 $Y2=0
cc_4192 N_S[5]_c_5220_n N_A_6674_325#_c_5469_n 0.0111895f $X=33.65 $Y=0.81 $X2=0
+ $Y2=0
cc_4193 N_S[5]_c_5221_n N_A_6674_325#_c_5469_n 9.67113e-19 $X=33.725 $Y=0.735
+ $X2=0 $Y2=0
cc_4194 N_S[5]_c_5234_n N_A_6674_325#_c_5469_n 0.00426435f $X=33.75 $Y=0.81
+ $X2=0 $Y2=0
cc_4195 N_S[5]_c_5218_n N_A_6674_325#_c_5470_n 0.00416423f $X=33.28 $Y=1.55
+ $X2=0 $Y2=0
cc_4196 N_S[5]_c_5222_n N_A_6674_325#_c_5470_n 0.00322131f $X=33.75 $Y=1.45
+ $X2=0 $Y2=0
cc_4197 N_S[5]_c_5238_n N_A_6674_325#_c_5470_n 0.0228692f $X=33.24 $Y=1.16 $X2=0
+ $Y2=0
cc_4198 N_S[5]_c_5222_n N_A_6674_325#_c_5471_n 0.0175393f $X=33.75 $Y=1.45 $X2=0
+ $Y2=0
cc_4199 N_S[5]_c_5223_n N_A_6674_325#_c_5471_n 0.0179529f $X=34.185 $Y=0.81
+ $X2=0 $Y2=0
cc_4200 N_S[5]_c_5217_n N_VPWR_c_7278_n 0.00652399f $X=33.18 $Y=1.16 $X2=0 $Y2=0
cc_4201 N_S[5]_c_5218_n N_VPWR_c_7278_n 0.00986205f $X=33.28 $Y=1.55 $X2=0 $Y2=0
cc_4202 N_S[5]_c_5238_n N_VPWR_c_7278_n 0.0157609f $X=33.24 $Y=1.16 $X2=0 $Y2=0
cc_4203 N_S[5]_c_5242_n N_VPWR_c_7280_n 0.00950399f $X=33.75 $Y=1.55 $X2=0 $Y2=0
cc_4204 N_S[5]_c_5218_n N_VPWR_c_7334_n 0.0035837f $X=33.28 $Y=1.55 $X2=0 $Y2=0
cc_4205 N_S[5]_c_5242_n N_VPWR_c_7334_n 0.0035837f $X=33.75 $Y=1.55 $X2=0 $Y2=0
cc_4206 N_S[5]_c_5218_n VPWR 0.0070533f $X=33.28 $Y=1.55 $X2=0 $Y2=0
cc_4207 N_S[5]_c_5242_n VPWR 0.00711603f $X=33.75 $Y=1.55 $X2=0 $Y2=0
cc_4208 N_S[5]_c_5227_n N_Z_c_9028_n 0.0134253f $X=35.02 $Y=0.255 $X2=0 $Y2=0
cc_4209 N_S[5]_c_5229_n N_Z_c_9028_n 0.0077801f $X=35.44 $Y=0.255 $X2=0 $Y2=0
cc_4210 N_S[5]_c_5231_n N_Z_c_9028_n 6.35774e-19 $X=35.86 $Y=0.255 $X2=0 $Y2=0
cc_4211 N_S[5]_c_5229_n N_Z_c_9030_n 0.00190704f $X=35.44 $Y=0.255 $X2=0 $Y2=0
cc_4212 N_S[5]_c_5231_n N_Z_c_9030_n 3.10191e-19 $X=35.86 $Y=0.255 $X2=0 $Y2=0
cc_4213 N_S[5]_c_5231_n N_Z_c_9032_n 0.00283489f $X=35.86 $Y=0.255 $X2=0 $Y2=0
cc_4214 N_S[5]_c_5233_n N_Z_c_9032_n 0.002324f $X=36.28 $Y=0.255 $X2=0 $Y2=0
cc_4215 N_S[5]_c_5227_n N_Z_c_9078_n 0.00216436f $X=35.02 $Y=0.255 $X2=0 $Y2=0
cc_4216 N_S[5]_c_5231_n N_Z_c_9080_n 0.00180363f $X=35.86 $Y=0.255 $X2=0 $Y2=0
cc_4217 N_S[5]_c_5229_n N_Z_c_9082_n 6.35664e-19 $X=35.44 $Y=0.255 $X2=0 $Y2=0
cc_4218 N_S[5]_c_5231_n N_Z_c_9082_n 0.00462308f $X=35.86 $Y=0.255 $X2=0 $Y2=0
cc_4219 N_S[5]_c_5233_n N_Z_c_9082_n 0.00443615f $X=36.28 $Y=0.255 $X2=0 $Y2=0
cc_4220 N_S[5]_c_5217_n N_Z_c_9125_n 0.00234109f $X=33.18 $Y=1.16 $X2=0 $Y2=0
cc_4221 N_S[5]_c_5218_n N_Z_c_9125_n 0.0052507f $X=33.28 $Y=1.55 $X2=0 $Y2=0
cc_4222 N_S[5]_c_5242_n N_Z_c_9125_n 0.00478771f $X=33.75 $Y=1.55 $X2=0 $Y2=0
cc_4223 N_S[5]_c_5238_n N_Z_c_9125_n 0.0105931f $X=33.24 $Y=1.16 $X2=0 $Y2=0
cc_4224 N_S[5]_c_5233_n N_A_6887_311#_c_11934_n 0.00168571f $X=36.28 $Y=0.255
+ $X2=0 $Y2=0
cc_4225 N_S[5]_c_5242_n N_A_6887_311#_c_11936_n 0.00239129f $X=33.75 $Y=1.55
+ $X2=0 $Y2=0
cc_4226 N_S[5]_c_5217_n N_VGND_c_12751_n 0.00576464f $X=33.18 $Y=1.16 $X2=0
+ $Y2=0
cc_4227 N_S[5]_c_5219_n N_VGND_c_12751_n 0.00374526f $X=33.305 $Y=0.735 $X2=0
+ $Y2=0
cc_4228 N_S[5]_c_5238_n N_VGND_c_12751_n 0.0116218f $X=33.24 $Y=1.16 $X2=0 $Y2=0
cc_4229 N_S[5]_c_5221_n N_VGND_c_12753_n 0.00173127f $X=33.725 $Y=0.735 $X2=0
+ $Y2=0
cc_4230 N_S[5]_c_5223_n N_VGND_c_12753_n 0.00525833f $X=34.185 $Y=0.81 $X2=0
+ $Y2=0
cc_4231 N_S[5]_c_5226_n N_VGND_c_12753_n 0.00862298f $X=34.335 $Y=0.18 $X2=0
+ $Y2=0
cc_4232 N_S[5]_c_5232_n N_VGND_c_12755_n 0.0028166f $X=36.205 $Y=0.18 $X2=0
+ $Y2=0
cc_4233 N_S[5]_c_5233_n N_VGND_c_12755_n 5.5039e-19 $X=36.28 $Y=0.255 $X2=0
+ $Y2=0
cc_4234 N_S[5]_c_5219_n N_VGND_c_12839_n 0.00585385f $X=33.305 $Y=0.735 $X2=0
+ $Y2=0
cc_4235 N_S[5]_c_5220_n N_VGND_c_12839_n 2.16067e-19 $X=33.65 $Y=0.81 $X2=0
+ $Y2=0
cc_4236 N_S[5]_c_5221_n N_VGND_c_12839_n 0.00542362f $X=33.725 $Y=0.735 $X2=0
+ $Y2=0
cc_4237 N_S[5]_c_5226_n N_VGND_c_12843_n 0.0559651f $X=34.335 $Y=0.18 $X2=0
+ $Y2=0
cc_4238 N_S[5]_c_5219_n VGND 0.0119653f $X=33.305 $Y=0.735 $X2=0 $Y2=0
cc_4239 N_S[5]_c_5221_n VGND 0.00990284f $X=33.725 $Y=0.735 $X2=0 $Y2=0
cc_4240 N_S[5]_c_5225_n VGND 0.0244174f $X=34.945 $Y=0.18 $X2=0 $Y2=0
cc_4241 N_S[5]_c_5226_n VGND 0.0101627f $X=34.335 $Y=0.18 $X2=0 $Y2=0
cc_4242 N_S[5]_c_5228_n VGND 0.00642387f $X=35.365 $Y=0.18 $X2=0 $Y2=0
cc_4243 N_S[5]_c_5230_n VGND 0.0064237f $X=35.785 $Y=0.18 $X2=0 $Y2=0
cc_4244 N_S[5]_c_5232_n VGND 0.0123437f $X=36.205 $Y=0.18 $X2=0 $Y2=0
cc_4245 N_S[5]_c_5235_n VGND 0.00366655f $X=35.02 $Y=0.18 $X2=0 $Y2=0
cc_4246 N_S[5]_c_5236_n VGND 0.00366655f $X=35.44 $Y=0.18 $X2=0 $Y2=0
cc_4247 N_S[5]_c_5237_n VGND 0.00366655f $X=35.86 $Y=0.18 $X2=0 $Y2=0
cc_4248 N_S[5]_c_5224_n N_A_6937_66#_c_14867_n 0.00529837f $X=34.26 $Y=0.735
+ $X2=0 $Y2=0
cc_4249 N_S[5]_c_5227_n N_A_6937_66#_c_14868_n 0.0112916f $X=35.02 $Y=0.255
+ $X2=0 $Y2=0
cc_4250 N_S[5]_c_5228_n N_A_6937_66#_c_14868_n 0.00211351f $X=35.365 $Y=0.18
+ $X2=0 $Y2=0
cc_4251 N_S[5]_c_5229_n N_A_6937_66#_c_14868_n 0.0106844f $X=35.44 $Y=0.255
+ $X2=0 $Y2=0
cc_4252 N_S[5]_c_5224_n N_A_6937_66#_c_14869_n 0.00189496f $X=34.26 $Y=0.735
+ $X2=0 $Y2=0
cc_4253 N_S[5]_c_5225_n N_A_6937_66#_c_14869_n 0.00685838f $X=34.945 $Y=0.18
+ $X2=0 $Y2=0
cc_4254 N_S[5]_c_5231_n N_A_6937_66#_c_14870_n 0.0106826f $X=35.86 $Y=0.255
+ $X2=0 $Y2=0
cc_4255 N_S[5]_c_5232_n N_A_6937_66#_c_14870_n 0.00211351f $X=36.205 $Y=0.18
+ $X2=0 $Y2=0
cc_4256 N_S[5]_c_5233_n N_A_6937_66#_c_14870_n 0.0139014f $X=36.28 $Y=0.255
+ $X2=0 $Y2=0
cc_4257 N_S[5]_c_5233_n N_A_6937_66#_c_14873_n 0.00206084f $X=36.28 $Y=0.255
+ $X2=0 $Y2=0
cc_4258 N_S[5]_c_5230_n N_A_6937_66#_c_14886_n 0.0034777f $X=35.785 $Y=0.18
+ $X2=0 $Y2=0
cc_4259 N_S[13]_c_5346_n N_A_6674_599#_c_5589_n 0.00507688f $X=35.02 $Y=5.185
+ $X2=25.905 $Y2=0.425
cc_4260 N_S[13]_c_5361_n N_A_6674_599#_c_5581_n 0.00262132f $X=33.75 $Y=3.99
+ $X2=25.905 $Y2=4.845
cc_4261 N_S[13]_c_5348_n N_A_6674_599#_c_5592_n 0.00509204f $X=35.44 $Y=5.185
+ $X2=0 $Y2=0
cc_4262 N_S[13]_c_5352_n N_A_6674_599#_c_5594_n 0.00507426f $X=36.28 $Y=5.185
+ $X2=0 $Y2=0
cc_4263 N_S[13]_c_5350_n N_A_6674_599#_c_5597_n 0.00509391f $X=35.86 $Y=5.185
+ $X2=0 $Y2=0
cc_4264 N_S[13]_c_5359_n N_A_6674_599#_c_5598_n 0.00929139f $X=33.28 $Y=3.89
+ $X2=0 $Y2=0
cc_4265 N_S[13]_c_5363_n N_A_6674_599#_c_5598_n 0.00970559f $X=33.75 $Y=3.89
+ $X2=0 $Y2=0
cc_4266 N_S[13]_c_5338_n N_A_6674_599#_c_5582_n 0.00207203f $X=33.305 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_4267 N_S[13]_c_5339_n N_A_6674_599#_c_5582_n 0.0111895f $X=33.65 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_4268 N_S[13]_c_5341_n N_A_6674_599#_c_5582_n 9.67113e-19 $X=33.725 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_4269 N_S[13]_c_5343_n N_A_6674_599#_c_5582_n 6.53442e-19 $X=34.26 $Y=5.185
+ $X2=25.99 $Y2=0.51
cc_4270 N_S[13]_c_5353_n N_A_6674_599#_c_5582_n 0.00426435f $X=33.75 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_4271 N_S[13]_c_5341_n N_A_6674_599#_c_5583_n 0.00603996f $X=33.725 $Y=4.705
+ $X2=0 $Y2=0
cc_4272 N_S[13]_c_5359_n N_A_6674_599#_c_5599_n 0.00117303f $X=33.28 $Y=3.89
+ $X2=0 $Y2=0
cc_4273 N_S[13]_c_5338_n N_A_6674_599#_c_5599_n 0.00336772f $X=33.305 $Y=4.705
+ $X2=0 $Y2=0
cc_4274 N_S[13]_c_5361_n N_A_6674_599#_c_5599_n 0.00508008f $X=33.75 $Y=3.99
+ $X2=0 $Y2=0
cc_4275 N_S[13]_c_5340_n N_A_6674_599#_c_5599_n 0.00255921f $X=33.75 $Y=4.555
+ $X2=0 $Y2=0
cc_4276 N_S[13]_c_5363_n N_A_6674_599#_c_5599_n 0.00254107f $X=33.75 $Y=3.89
+ $X2=0 $Y2=0
cc_4277 N_S[13]_c_5340_n N_A_6674_599#_c_5584_n 0.0206368f $X=33.75 $Y=4.555
+ $X2=0 $Y2=0
cc_4278 N_S[13]_c_5342_n N_A_6674_599#_c_5584_n 0.0103812f $X=34.185 $Y=4.63
+ $X2=0 $Y2=0
cc_4279 N_S[13]_c_5359_n N_A_6674_599#_c_5601_n 0.00304348f $X=33.28 $Y=3.89
+ $X2=0 $Y2=0
cc_4280 N_S[13]_c_5338_n N_A_6674_599#_c_5601_n 5.48523e-19 $X=33.305 $Y=4.705
+ $X2=0 $Y2=0
cc_4281 N_S[13]_c_5363_n N_A_6674_599#_c_5601_n 0.00216424f $X=33.75 $Y=3.89
+ $X2=0 $Y2=0
cc_4282 N_S[13]_c_5338_n N_A_6674_599#_c_5585_n 0.00289358f $X=33.305 $Y=4.705
+ $X2=0 $Y2=0
cc_4283 N_S[13]_c_5339_n N_A_6674_599#_c_5585_n 0.00429801f $X=33.65 $Y=4.63
+ $X2=0 $Y2=0
cc_4284 N_S[13]_c_5340_n N_A_6674_599#_c_5585_n 0.0085951f $X=33.75 $Y=4.555
+ $X2=0 $Y2=0
cc_4285 N_S[13]_c_5353_n N_A_6674_599#_c_5585_n 0.00268644f $X=33.75 $Y=4.63
+ $X2=0 $Y2=0
cc_4286 N_S[13]_c_5357_n N_A_6674_599#_c_5585_n 0.00541767f $X=33.24 $Y=4.28
+ $X2=0 $Y2=0
cc_4287 N_S[13]_c_5338_n N_A_6674_599#_c_5586_n 0.00416423f $X=33.305 $Y=4.705
+ $X2=0 $Y2=0
cc_4288 N_S[13]_c_5340_n N_A_6674_599#_c_5586_n 0.00322131f $X=33.75 $Y=4.555
+ $X2=0 $Y2=0
cc_4289 N_S[13]_c_5357_n N_A_6674_599#_c_5586_n 0.0228692f $X=33.24 $Y=4.28
+ $X2=0 $Y2=0
cc_4290 N_S[13]_c_5340_n N_A_6674_599#_c_5587_n 0.0175393f $X=33.75 $Y=4.555
+ $X2=0 $Y2=0
cc_4291 N_S[13]_c_5342_n N_A_6674_599#_c_5587_n 0.0179529f $X=34.185 $Y=4.63
+ $X2=0 $Y2=0
cc_4292 N_S[13]_c_5337_n N_VPWR_c_7279_n 0.00652399f $X=33.18 $Y=4.28 $X2=0
+ $Y2=0
cc_4293 N_S[13]_c_5359_n N_VPWR_c_7279_n 0.00986205f $X=33.28 $Y=3.89 $X2=0
+ $Y2=0
cc_4294 N_S[13]_c_5357_n N_VPWR_c_7279_n 0.0157609f $X=33.24 $Y=4.28 $X2=0 $Y2=0
cc_4295 N_S[13]_c_5363_n N_VPWR_c_7281_n 0.00950399f $X=33.75 $Y=3.89 $X2=0
+ $Y2=0
cc_4296 N_S[13]_c_5359_n N_VPWR_c_7334_n 0.0035837f $X=33.28 $Y=3.89 $X2=0 $Y2=0
cc_4297 N_S[13]_c_5363_n N_VPWR_c_7334_n 0.0035837f $X=33.75 $Y=3.89 $X2=0 $Y2=0
cc_4298 N_S[13]_c_5359_n VPWR 0.0070533f $X=33.28 $Y=3.89 $X2=0 $Y2=0
cc_4299 N_S[13]_c_5363_n VPWR 0.00711603f $X=33.75 $Y=3.89 $X2=0 $Y2=0
cc_4300 N_S[13]_c_5346_n N_Z_c_9029_n 0.0134253f $X=35.02 $Y=5.185 $X2=0 $Y2=0
cc_4301 N_S[13]_c_5348_n N_Z_c_9029_n 0.0077801f $X=35.44 $Y=5.185 $X2=0 $Y2=0
cc_4302 N_S[13]_c_5350_n N_Z_c_9029_n 6.35774e-19 $X=35.86 $Y=5.185 $X2=0 $Y2=0
cc_4303 N_S[13]_c_5348_n N_Z_c_9031_n 0.00190704f $X=35.44 $Y=5.185 $X2=0 $Y2=0
cc_4304 N_S[13]_c_5350_n N_Z_c_9031_n 3.10191e-19 $X=35.86 $Y=5.185 $X2=0 $Y2=0
cc_4305 N_S[13]_c_5346_n N_Z_c_9079_n 0.00216436f $X=35.02 $Y=5.185 $X2=0 $Y2=0
cc_4306 N_S[13]_c_5350_n N_Z_c_9081_n 0.00180363f $X=35.86 $Y=5.185 $X2=0 $Y2=0
cc_4307 N_S[13]_c_5350_n N_Z_c_9083_n 0.00462308f $X=35.86 $Y=5.185 $X2=0 $Y2=0
cc_4308 N_S[13]_c_5352_n N_Z_c_9083_n 0.00443615f $X=36.28 $Y=5.185 $X2=0 $Y2=0
cc_4309 N_S[13]_c_5348_n N_Z_c_9084_n 6.35664e-19 $X=35.44 $Y=5.185 $X2=0 $Y2=0
cc_4310 N_S[13]_c_5350_n N_Z_c_9084_n 0.00283489f $X=35.86 $Y=5.185 $X2=0 $Y2=0
cc_4311 N_S[13]_c_5352_n N_Z_c_9084_n 0.002324f $X=36.28 $Y=5.185 $X2=0 $Y2=0
cc_4312 N_S[13]_c_5337_n N_Z_c_9126_n 0.00234109f $X=33.18 $Y=4.28 $X2=0 $Y2=0
cc_4313 N_S[13]_c_5359_n N_Z_c_9126_n 0.00501777f $X=33.28 $Y=3.89 $X2=0 $Y2=0
cc_4314 N_S[13]_c_5338_n N_Z_c_9126_n 2.32936e-19 $X=33.305 $Y=4.705 $X2=0 $Y2=0
cc_4315 N_S[13]_c_5361_n N_Z_c_9126_n 2.55735e-19 $X=33.75 $Y=3.99 $X2=0 $Y2=0
cc_4316 N_S[13]_c_5363_n N_Z_c_9126_n 0.00453198f $X=33.75 $Y=3.89 $X2=0 $Y2=0
cc_4317 N_S[13]_c_5357_n N_Z_c_9126_n 0.0105931f $X=33.24 $Y=4.28 $X2=0 $Y2=0
cc_4318 N_S[13]_c_5352_n N_A_6887_613#_c_12065_n 0.00168571f $X=36.28 $Y=5.185
+ $X2=0 $Y2=0
cc_4319 N_S[13]_c_5363_n N_A_6887_613#_c_12067_n 0.00239129f $X=33.75 $Y=3.89
+ $X2=0 $Y2=0
cc_4320 N_S[13]_c_5337_n N_VGND_c_12752_n 0.00576464f $X=33.18 $Y=4.28 $X2=0
+ $Y2=0
cc_4321 N_S[13]_c_5338_n N_VGND_c_12752_n 0.00374526f $X=33.305 $Y=4.705 $X2=0
+ $Y2=0
cc_4322 N_S[13]_c_5357_n N_VGND_c_12752_n 0.0116218f $X=33.24 $Y=4.28 $X2=0
+ $Y2=0
cc_4323 N_S[13]_c_5341_n N_VGND_c_12754_n 0.00173127f $X=33.725 $Y=4.705 $X2=0
+ $Y2=0
cc_4324 N_S[13]_c_5342_n N_VGND_c_12754_n 0.00525833f $X=34.185 $Y=4.63 $X2=0
+ $Y2=0
cc_4325 N_S[13]_c_5343_n N_VGND_c_12754_n 0.00862298f $X=34.26 $Y=5.185 $X2=0
+ $Y2=0
cc_4326 N_S[13]_c_5351_n N_VGND_c_12756_n 0.0028166f $X=36.205 $Y=5.26 $X2=0
+ $Y2=0
cc_4327 N_S[13]_c_5352_n N_VGND_c_12756_n 5.5039e-19 $X=36.28 $Y=5.185 $X2=0
+ $Y2=0
cc_4328 N_S[13]_c_5338_n N_VGND_c_12841_n 0.00585385f $X=33.305 $Y=4.705 $X2=0
+ $Y2=0
cc_4329 N_S[13]_c_5339_n N_VGND_c_12841_n 2.16067e-19 $X=33.65 $Y=4.63 $X2=0
+ $Y2=0
cc_4330 N_S[13]_c_5341_n N_VGND_c_12841_n 0.00542362f $X=33.725 $Y=4.705 $X2=0
+ $Y2=0
cc_4331 N_S[13]_c_5345_n N_VGND_c_12845_n 0.0559651f $X=34.335 $Y=5.26 $X2=0
+ $Y2=0
cc_4332 N_S[13]_c_5338_n VGND 0.0119653f $X=33.305 $Y=4.705 $X2=0 $Y2=0
cc_4333 N_S[13]_c_5341_n VGND 0.00990284f $X=33.725 $Y=4.705 $X2=0 $Y2=0
cc_4334 N_S[13]_c_5344_n VGND 0.0244174f $X=34.945 $Y=5.26 $X2=0 $Y2=0
cc_4335 N_S[13]_c_5345_n VGND 0.0101627f $X=34.335 $Y=5.26 $X2=0 $Y2=0
cc_4336 N_S[13]_c_5347_n VGND 0.00642387f $X=35.365 $Y=5.26 $X2=0 $Y2=0
cc_4337 N_S[13]_c_5349_n VGND 0.0064237f $X=35.785 $Y=5.26 $X2=0 $Y2=0
cc_4338 N_S[13]_c_5351_n VGND 0.0123437f $X=36.205 $Y=5.26 $X2=0 $Y2=0
cc_4339 N_S[13]_c_5354_n VGND 0.00366655f $X=35.02 $Y=5.26 $X2=0 $Y2=0
cc_4340 N_S[13]_c_5355_n VGND 0.00366655f $X=35.44 $Y=5.26 $X2=0 $Y2=0
cc_4341 N_S[13]_c_5356_n VGND 0.00366655f $X=35.86 $Y=5.26 $X2=0 $Y2=0
cc_4342 N_S[13]_c_5342_n N_A_6937_918#_c_14951_n 0.00529837f $X=34.185 $Y=4.63
+ $X2=0 $Y2=0
cc_4343 N_S[13]_c_5346_n N_A_6937_918#_c_14952_n 0.0112916f $X=35.02 $Y=5.185
+ $X2=0 $Y2=0
cc_4344 N_S[13]_c_5347_n N_A_6937_918#_c_14952_n 0.00211351f $X=35.365 $Y=5.26
+ $X2=0 $Y2=0
cc_4345 N_S[13]_c_5348_n N_A_6937_918#_c_14952_n 0.0106844f $X=35.44 $Y=5.185
+ $X2=0 $Y2=0
cc_4346 N_S[13]_c_5343_n N_A_6937_918#_c_14953_n 0.00189496f $X=34.26 $Y=5.185
+ $X2=0 $Y2=0
cc_4347 N_S[13]_c_5344_n N_A_6937_918#_c_14953_n 0.00685838f $X=34.945 $Y=5.26
+ $X2=0 $Y2=0
cc_4348 N_S[13]_c_5350_n N_A_6937_918#_c_14954_n 0.0106826f $X=35.86 $Y=5.185
+ $X2=0 $Y2=0
cc_4349 N_S[13]_c_5351_n N_A_6937_918#_c_14954_n 0.00211351f $X=36.205 $Y=5.26
+ $X2=0 $Y2=0
cc_4350 N_S[13]_c_5352_n N_A_6937_918#_c_14954_n 0.0139014f $X=36.28 $Y=5.185
+ $X2=0 $Y2=0
cc_4351 N_S[13]_c_5352_n N_A_6937_918#_c_14957_n 0.00206084f $X=36.28 $Y=5.185
+ $X2=0 $Y2=0
cc_4352 N_S[13]_c_5349_n N_A_6937_918#_c_14970_n 0.0034777f $X=35.785 $Y=5.26
+ $X2=0 $Y2=0
cc_4353 N_A_6674_325#_c_5472_n N_A_6674_599#_c_5588_n 0.0129371f $X=34.795
+ $Y=1.475 $X2=0 $Y2=0
cc_4354 N_A_6674_325#_c_5475_n N_A_6674_599#_c_5591_n 0.0129371f $X=35.265
+ $Y=1.475 $X2=0 $Y2=0
cc_4355 N_A_6674_325#_c_5477_n N_A_6674_599#_c_5593_n 0.0129371f $X=35.735
+ $Y=1.475 $X2=0 $Y2=0
cc_4356 N_A_6674_325#_c_5479_n N_A_6674_599#_c_5595_n 0.0129371f $X=36.205
+ $Y=1.475 $X2=0 $Y2=0
cc_4357 N_A_6674_325#_c_5482_n N_VPWR_c_7278_n 0.0356181f $X=33.515 $Y=1.77
+ $X2=0 $Y2=0
cc_4358 N_A_6674_325#_c_5472_n N_VPWR_c_7280_n 0.00367058f $X=34.795 $Y=1.475
+ $X2=0 $Y2=0
cc_4359 N_A_6674_325#_c_5482_n N_VPWR_c_7280_n 0.0316788f $X=33.515 $Y=1.77
+ $X2=0 $Y2=0
cc_4360 N_A_6674_325#_c_5468_n N_VPWR_c_7280_n 0.0193185f $X=34.565 $Y=1.23
+ $X2=0 $Y2=0
cc_4361 N_A_6674_325#_c_5471_n N_VPWR_c_7280_n 6.4101e-19 $X=34.475 $Y=1.23
+ $X2=0 $Y2=0
cc_4362 N_A_6674_325#_c_5479_n N_VPWR_c_7282_n 0.00324472f $X=36.205 $Y=1.475
+ $X2=0 $Y2=0
cc_4363 N_A_6674_325#_c_5482_n N_VPWR_c_7334_n 0.0233824f $X=33.515 $Y=1.77
+ $X2=0 $Y2=0
cc_4364 N_A_6674_325#_c_5472_n VPWR 0.00473731f $X=34.795 $Y=1.475 $X2=0 $Y2=0
cc_4365 N_A_6674_325#_c_5475_n VPWR 0.00362156f $X=35.265 $Y=1.475 $X2=0 $Y2=0
cc_4366 N_A_6674_325#_c_5477_n VPWR 0.00362156f $X=35.735 $Y=1.475 $X2=0 $Y2=0
cc_4367 N_A_6674_325#_c_5479_n VPWR 0.00473731f $X=36.205 $Y=1.475 $X2=0 $Y2=0
cc_4368 N_A_6674_325#_c_5482_n VPWR 0.00593513f $X=33.515 $Y=1.77 $X2=0 $Y2=0
cc_4369 N_A_6674_325#_c_5476_n N_Z_c_9030_n 0.00762343f $X=35.645 $Y=1.4 $X2=0
+ $Y2=0
cc_4370 N_A_6674_325#_c_5481_n N_Z_c_9030_n 0.00704092f $X=35.735 $Y=1.4 $X2=0
+ $Y2=0
cc_4371 N_A_6674_325#_c_5473_n N_Z_c_9078_n 0.00597584f $X=35.175 $Y=1.4 $X2=0
+ $Y2=0
cc_4372 N_A_6674_325#_c_5465_n N_Z_c_9078_n 0.00747617f $X=34.885 $Y=1.4 $X2=0
+ $Y2=0
cc_4373 N_A_6674_325#_c_5476_n N_Z_c_9078_n 0.00145542f $X=35.645 $Y=1.4 $X2=0
+ $Y2=0
cc_4374 N_A_6674_325#_c_5480_n N_Z_c_9078_n 0.00909323f $X=35.265 $Y=1.4 $X2=0
+ $Y2=0
cc_4375 N_A_6674_325#_c_5468_n N_Z_c_9078_n 0.0266078f $X=34.565 $Y=1.23 $X2=0
+ $Y2=0
cc_4376 N_A_6674_325#_c_5478_n N_Z_c_9080_n 0.00918337f $X=36.115 $Y=1.4 $X2=0
+ $Y2=0
cc_4377 N_A_6674_325#_c_5481_n N_Z_c_9080_n 2.98555e-19 $X=35.735 $Y=1.4 $X2=0
+ $Y2=0
cc_4378 N_A_6674_325#_c_5478_n N_Z_c_9082_n 0.00248496f $X=36.115 $Y=1.4 $X2=0
+ $Y2=0
cc_4379 N_A_6674_325#_c_5472_n N_Z_c_9125_n 0.00795576f $X=34.795 $Y=1.475 $X2=0
+ $Y2=0
cc_4380 N_A_6674_325#_c_5465_n N_Z_c_9125_n 2.19754e-19 $X=34.885 $Y=1.4 $X2=0
+ $Y2=0
cc_4381 N_A_6674_325#_c_5482_n N_Z_c_9125_n 0.0329704f $X=33.515 $Y=1.77 $X2=0
+ $Y2=0
cc_4382 N_A_6674_325#_c_5468_n N_Z_c_9125_n 0.0186685f $X=34.565 $Y=1.23 $X2=0
+ $Y2=0
cc_4383 N_A_6674_325#_c_5479_n N_Z_c_9127_n 0.00834829f $X=36.205 $Y=1.475 $X2=0
+ $Y2=0
cc_4384 N_A_6674_325#_c_5475_n N_Z_c_9700_n 0.00372248f $X=35.265 $Y=1.475 $X2=0
+ $Y2=0
cc_4385 N_A_6674_325#_c_5477_n N_Z_c_9700_n 0.00372458f $X=35.735 $Y=1.475 $X2=0
+ $Y2=0
cc_4386 N_A_6674_325#_c_5472_n N_Z_c_9141_n 0.0221748f $X=34.795 $Y=1.475 $X2=0
+ $Y2=0
cc_4387 N_A_6674_325#_c_5473_n N_Z_c_9141_n 0.00560592f $X=35.175 $Y=1.4 $X2=0
+ $Y2=0
cc_4388 N_A_6674_325#_c_5465_n N_Z_c_9141_n 0.00425035f $X=34.885 $Y=1.4 $X2=0
+ $Y2=0
cc_4389 N_A_6674_325#_c_5475_n N_Z_c_9141_n 0.0181262f $X=35.265 $Y=1.475 $X2=0
+ $Y2=0
cc_4390 N_A_6674_325#_c_5477_n N_Z_c_9141_n 9.74366e-19 $X=35.735 $Y=1.475 $X2=0
+ $Y2=0
cc_4391 N_A_6674_325#_c_5480_n N_Z_c_9141_n 0.00181273f $X=35.265 $Y=1.4 $X2=0
+ $Y2=0
cc_4392 N_A_6674_325#_c_5468_n N_Z_c_9141_n 0.00240108f $X=34.565 $Y=1.23 $X2=0
+ $Y2=0
cc_4393 N_A_6674_325#_c_5475_n N_Z_c_9142_n 9.74366e-19 $X=35.265 $Y=1.475 $X2=0
+ $Y2=0
cc_4394 N_A_6674_325#_c_5477_n N_Z_c_9142_n 0.0181262f $X=35.735 $Y=1.475 $X2=0
+ $Y2=0
cc_4395 N_A_6674_325#_c_5478_n N_Z_c_9142_n 0.0103509f $X=36.115 $Y=1.4 $X2=0
+ $Y2=0
cc_4396 N_A_6674_325#_c_5479_n N_Z_c_9142_n 0.0199111f $X=36.205 $Y=1.475 $X2=0
+ $Y2=0
cc_4397 N_A_6674_325#_c_5481_n N_Z_c_9142_n 0.00415268f $X=35.735 $Y=1.4 $X2=0
+ $Y2=0
cc_4398 N_A_6674_325#_c_5479_n N_A_6887_311#_c_11934_n 0.00151141f $X=36.205
+ $Y=1.475 $X2=0 $Y2=0
cc_4399 N_A_6674_325#_c_5472_n N_A_6887_311#_c_11942_n 0.00307958f $X=34.795
+ $Y=1.475 $X2=0 $Y2=0
cc_4400 N_A_6674_325#_c_5475_n N_A_6887_311#_c_11942_n 0.00307958f $X=35.265
+ $Y=1.475 $X2=0 $Y2=0
cc_4401 N_A_6674_325#_c_5477_n N_A_6887_311#_c_11944_n 0.00307958f $X=35.735
+ $Y=1.475 $X2=0 $Y2=0
cc_4402 N_A_6674_325#_c_5479_n N_A_6887_311#_c_11944_n 0.00307958f $X=36.205
+ $Y=1.475 $X2=0 $Y2=0
cc_4403 N_A_6674_325#_c_5472_n N_A_6887_311#_c_11936_n 0.00499839f $X=34.795
+ $Y=1.475 $X2=0 $Y2=0
cc_4404 N_A_6674_325#_c_5465_n N_A_6887_311#_c_11936_n 0.00561627f $X=34.885
+ $Y=1.4 $X2=0 $Y2=0
cc_4405 N_A_6674_325#_c_5468_n N_A_6887_311#_c_11936_n 0.0218124f $X=34.565
+ $Y=1.23 $X2=0 $Y2=0
cc_4406 N_A_6674_325#_c_5471_n N_A_6887_311#_c_11936_n 5.74251e-19 $X=34.475
+ $Y=1.23 $X2=0 $Y2=0
cc_4407 N_A_6674_325#_c_5475_n N_A_6887_311#_c_11937_n 0.00210632f $X=35.265
+ $Y=1.475 $X2=0 $Y2=0
cc_4408 N_A_6674_325#_c_5476_n N_A_6887_311#_c_11937_n 0.00251792f $X=35.645
+ $Y=1.4 $X2=0 $Y2=0
cc_4409 N_A_6674_325#_c_5477_n N_A_6887_311#_c_11937_n 0.00210632f $X=35.735
+ $Y=1.475 $X2=0 $Y2=0
cc_4410 N_A_6674_325#_c_5479_n N_A_6887_311#_c_11938_n 0.00554566f $X=36.205
+ $Y=1.475 $X2=0 $Y2=0
cc_4411 N_A_6674_325#_c_5468_n N_VGND_c_12753_n 0.0123065f $X=34.565 $Y=1.23
+ $X2=0 $Y2=0
cc_4412 N_A_6674_325#_c_5471_n N_VGND_c_12753_n 2.04129e-19 $X=34.475 $Y=1.23
+ $X2=0 $Y2=0
cc_4413 N_A_6674_325#_c_5466_n N_VGND_c_12839_n 0.0129994f $X=33.515 $Y=0.445
+ $X2=0 $Y2=0
cc_4414 N_A_6674_325#_M1126_s VGND 0.00394793f $X=33.38 $Y=0.235 $X2=0 $Y2=0
cc_4415 N_A_6674_325#_c_5466_n VGND 0.00927134f $X=33.515 $Y=0.445 $X2=0 $Y2=0
cc_4416 N_A_6674_325#_c_5465_n N_A_6937_66#_c_14867_n 0.00600378f $X=34.885
+ $Y=1.4 $X2=0 $Y2=0
cc_4417 N_A_6674_325#_c_5468_n N_A_6937_66#_c_14867_n 0.0028695f $X=34.565
+ $Y=1.23 $X2=0 $Y2=0
cc_4418 N_A_6674_325#_c_5476_n N_A_6937_66#_c_14889_n 7.0477e-19 $X=35.645
+ $Y=1.4 $X2=0 $Y2=0
cc_4419 N_A_6674_599#_c_5598_n N_VPWR_c_7279_n 0.0356181f $X=33.515 $Y=3.14
+ $X2=0 $Y2=0
cc_4420 N_A_6674_599#_c_5588_n N_VPWR_c_7281_n 0.00367058f $X=34.795 $Y=3.965
+ $X2=0 $Y2=0
cc_4421 N_A_6674_599#_c_5598_n N_VPWR_c_7281_n 0.0316788f $X=33.515 $Y=3.14
+ $X2=0 $Y2=0
cc_4422 N_A_6674_599#_c_5584_n N_VPWR_c_7281_n 0.0193185f $X=34.565 $Y=4.21
+ $X2=0 $Y2=0
cc_4423 N_A_6674_599#_c_5587_n N_VPWR_c_7281_n 6.4101e-19 $X=34.475 $Y=4.21
+ $X2=0 $Y2=0
cc_4424 N_A_6674_599#_c_5595_n N_VPWR_c_7283_n 0.00324472f $X=36.205 $Y=3.965
+ $X2=0 $Y2=0
cc_4425 N_A_6674_599#_c_5598_n N_VPWR_c_7334_n 0.0233824f $X=33.515 $Y=3.14
+ $X2=0 $Y2=0
cc_4426 N_A_6674_599#_c_5588_n VPWR 0.00473731f $X=34.795 $Y=3.965 $X2=0 $Y2=0
cc_4427 N_A_6674_599#_c_5591_n VPWR 0.00362156f $X=35.265 $Y=3.965 $X2=0 $Y2=0
cc_4428 N_A_6674_599#_c_5593_n VPWR 0.00362156f $X=35.735 $Y=3.965 $X2=0 $Y2=0
cc_4429 N_A_6674_599#_c_5595_n VPWR 0.00473731f $X=36.205 $Y=3.965 $X2=0 $Y2=0
cc_4430 N_A_6674_599#_c_5598_n VPWR 0.00593513f $X=33.515 $Y=3.14 $X2=0 $Y2=0
cc_4431 N_A_6674_599#_c_5592_n N_Z_c_9031_n 0.00762343f $X=35.645 $Y=4.04 $X2=0
+ $Y2=0
cc_4432 N_A_6674_599#_c_5597_n N_Z_c_9031_n 0.00704092f $X=35.735 $Y=4.04 $X2=0
+ $Y2=0
cc_4433 N_A_6674_599#_c_5589_n N_Z_c_9079_n 0.00597584f $X=35.175 $Y=4.04 $X2=0
+ $Y2=0
cc_4434 N_A_6674_599#_c_5581_n N_Z_c_9079_n 0.00747617f $X=34.885 $Y=4.04 $X2=0
+ $Y2=0
cc_4435 N_A_6674_599#_c_5592_n N_Z_c_9079_n 0.00145542f $X=35.645 $Y=4.04 $X2=0
+ $Y2=0
cc_4436 N_A_6674_599#_c_5596_n N_Z_c_9079_n 0.00909323f $X=35.265 $Y=4.04 $X2=0
+ $Y2=0
cc_4437 N_A_6674_599#_c_5584_n N_Z_c_9079_n 0.0266078f $X=34.565 $Y=4.21 $X2=0
+ $Y2=0
cc_4438 N_A_6674_599#_c_5594_n N_Z_c_9081_n 0.00918337f $X=36.115 $Y=4.04 $X2=0
+ $Y2=0
cc_4439 N_A_6674_599#_c_5597_n N_Z_c_9081_n 2.98555e-19 $X=35.735 $Y=4.04 $X2=0
+ $Y2=0
cc_4440 N_A_6674_599#_c_5594_n N_Z_c_9083_n 0.00248496f $X=36.115 $Y=4.04 $X2=0
+ $Y2=0
cc_4441 N_A_6674_599#_c_5588_n N_Z_c_9126_n 0.00795576f $X=34.795 $Y=3.965 $X2=0
+ $Y2=0
cc_4442 N_A_6674_599#_c_5581_n N_Z_c_9126_n 2.19754e-19 $X=34.885 $Y=4.04 $X2=0
+ $Y2=0
cc_4443 N_A_6674_599#_c_5598_n N_Z_c_9126_n 0.0329704f $X=33.515 $Y=3.14 $X2=0
+ $Y2=0
cc_4444 N_A_6674_599#_c_5584_n N_Z_c_9126_n 0.0186685f $X=34.565 $Y=4.21 $X2=0
+ $Y2=0
cc_4445 N_A_6674_599#_c_5595_n N_Z_c_9128_n 0.00834829f $X=36.205 $Y=3.965 $X2=0
+ $Y2=0
cc_4446 N_A_6674_599#_c_5591_n N_Z_c_9729_n 0.00372248f $X=35.265 $Y=3.965 $X2=0
+ $Y2=0
cc_4447 N_A_6674_599#_c_5593_n N_Z_c_9729_n 0.00372458f $X=35.735 $Y=3.965 $X2=0
+ $Y2=0
cc_4448 N_A_6674_599#_c_5588_n N_Z_c_9141_n 0.0221748f $X=34.795 $Y=3.965 $X2=0
+ $Y2=0
cc_4449 N_A_6674_599#_c_5589_n N_Z_c_9141_n 0.00560592f $X=35.175 $Y=4.04 $X2=0
+ $Y2=0
cc_4450 N_A_6674_599#_c_5581_n N_Z_c_9141_n 0.00425035f $X=34.885 $Y=4.04 $X2=0
+ $Y2=0
cc_4451 N_A_6674_599#_c_5591_n N_Z_c_9141_n 0.0181262f $X=35.265 $Y=3.965 $X2=0
+ $Y2=0
cc_4452 N_A_6674_599#_c_5593_n N_Z_c_9141_n 9.74366e-19 $X=35.735 $Y=3.965 $X2=0
+ $Y2=0
cc_4453 N_A_6674_599#_c_5596_n N_Z_c_9141_n 0.00181273f $X=35.265 $Y=4.04 $X2=0
+ $Y2=0
cc_4454 N_A_6674_599#_c_5584_n N_Z_c_9141_n 0.00240108f $X=34.565 $Y=4.21 $X2=0
+ $Y2=0
cc_4455 N_A_6674_599#_c_5591_n N_Z_c_9142_n 9.74366e-19 $X=35.265 $Y=3.965 $X2=0
+ $Y2=0
cc_4456 N_A_6674_599#_c_5593_n N_Z_c_9142_n 0.0181262f $X=35.735 $Y=3.965 $X2=0
+ $Y2=0
cc_4457 N_A_6674_599#_c_5594_n N_Z_c_9142_n 0.0103509f $X=36.115 $Y=4.04 $X2=0
+ $Y2=0
cc_4458 N_A_6674_599#_c_5595_n N_Z_c_9142_n 0.0199111f $X=36.205 $Y=3.965 $X2=0
+ $Y2=0
cc_4459 N_A_6674_599#_c_5597_n N_Z_c_9142_n 0.00415268f $X=35.735 $Y=4.04 $X2=0
+ $Y2=0
cc_4460 N_A_6674_599#_c_5595_n N_A_6887_613#_c_12065_n 0.00151141f $X=36.205
+ $Y=3.965 $X2=0 $Y2=0
cc_4461 N_A_6674_599#_c_5588_n N_A_6887_613#_c_12073_n 0.00307958f $X=34.795
+ $Y=3.965 $X2=0 $Y2=0
cc_4462 N_A_6674_599#_c_5591_n N_A_6887_613#_c_12073_n 0.00307958f $X=35.265
+ $Y=3.965 $X2=0 $Y2=0
cc_4463 N_A_6674_599#_c_5593_n N_A_6887_613#_c_12075_n 0.00307958f $X=35.735
+ $Y=3.965 $X2=0 $Y2=0
cc_4464 N_A_6674_599#_c_5595_n N_A_6887_613#_c_12075_n 0.00307958f $X=36.205
+ $Y=3.965 $X2=0 $Y2=0
cc_4465 N_A_6674_599#_c_5588_n N_A_6887_613#_c_12067_n 0.00499839f $X=34.795
+ $Y=3.965 $X2=0 $Y2=0
cc_4466 N_A_6674_599#_c_5581_n N_A_6887_613#_c_12067_n 0.00561627f $X=34.885
+ $Y=4.04 $X2=0 $Y2=0
cc_4467 N_A_6674_599#_c_5584_n N_A_6887_613#_c_12067_n 0.0218124f $X=34.565
+ $Y=4.21 $X2=0 $Y2=0
cc_4468 N_A_6674_599#_c_5587_n N_A_6887_613#_c_12067_n 5.74251e-19 $X=34.475
+ $Y=4.21 $X2=0 $Y2=0
cc_4469 N_A_6674_599#_c_5591_n N_A_6887_613#_c_12068_n 0.00210632f $X=35.265
+ $Y=3.965 $X2=0 $Y2=0
cc_4470 N_A_6674_599#_c_5592_n N_A_6887_613#_c_12068_n 0.00251792f $X=35.645
+ $Y=4.04 $X2=0 $Y2=0
cc_4471 N_A_6674_599#_c_5593_n N_A_6887_613#_c_12068_n 0.00210632f $X=35.735
+ $Y=3.965 $X2=0 $Y2=0
cc_4472 N_A_6674_599#_c_5595_n N_A_6887_613#_c_12069_n 0.00554566f $X=36.205
+ $Y=3.965 $X2=0 $Y2=0
cc_4473 N_A_6674_599#_c_5584_n N_VGND_c_12754_n 0.0123065f $X=34.565 $Y=4.21
+ $X2=0 $Y2=0
cc_4474 N_A_6674_599#_c_5587_n N_VGND_c_12754_n 2.04129e-19 $X=34.475 $Y=4.21
+ $X2=0 $Y2=0
cc_4475 N_A_6674_599#_c_5583_n N_VGND_c_12841_n 0.0129994f $X=33.515 $Y=4.995
+ $X2=0 $Y2=0
cc_4476 N_A_6674_599#_M1060_s VGND 0.00394793f $X=33.38 $Y=4.785 $X2=0 $Y2=0
cc_4477 N_A_6674_599#_c_5583_n VGND 0.00927134f $X=33.515 $Y=4.995 $X2=0 $Y2=0
cc_4478 N_A_6674_599#_c_5581_n N_A_6937_918#_c_14951_n 0.00600378f $X=34.885
+ $Y=4.04 $X2=0 $Y2=0
cc_4479 N_A_6674_599#_c_5584_n N_A_6937_918#_c_14951_n 0.0028695f $X=34.565
+ $Y=4.21 $X2=0 $Y2=0
cc_4480 N_A_6674_599#_c_5592_n N_A_6937_918#_c_14973_n 7.0477e-19 $X=35.645
+ $Y=4.04 $X2=0 $Y2=0
cc_4481 N_D[5]_M1088_g N_D[13]_M1102_g 0.0130744f $X=37.195 $Y=1.985 $X2=0 $Y2=0
cc_4482 N_D[5]_M1183_g N_D[13]_M1186_g 0.0130744f $X=37.665 $Y=1.985 $X2=0 $Y2=0
cc_4483 N_D[5]_M1217_g N_D[13]_M1224_g 0.0130744f $X=38.135 $Y=1.985 $X2=0 $Y2=0
cc_4484 N_D[5]_M1255_g N_D[13]_M1264_g 0.0130744f $X=38.605 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_4485 N_D[5]_M1088_g N_VPWR_c_7282_n 0.00389633f $X=37.195 $Y=1.985 $X2=0
+ $Y2=0
cc_4486 N_D[5]_M1183_g N_VPWR_c_7284_n 0.00208662f $X=37.665 $Y=1.985 $X2=0
+ $Y2=0
cc_4487 N_D[5]_M1217_g N_VPWR_c_7284_n 0.00208662f $X=38.135 $Y=1.985 $X2=0
+ $Y2=0
cc_4488 N_D[5]_M1255_g N_VPWR_c_7286_n 0.00374733f $X=38.605 $Y=1.985 $X2=0
+ $Y2=0
cc_4489 N_D[5]_M1088_g VPWR 0.00573859f $X=37.195 $Y=1.985 $X2=0 $Y2=0
cc_4490 N_D[5]_M1183_g VPWR 0.00445624f $X=37.665 $Y=1.985 $X2=0 $Y2=0
cc_4491 N_D[5]_M1217_g VPWR 0.00445624f $X=38.135 $Y=1.985 $X2=0 $Y2=0
cc_4492 N_D[5]_M1255_g VPWR 0.00691494f $X=38.605 $Y=1.985 $X2=0 $Y2=0
cc_4493 N_D[5]_M1088_g N_VPWR_c_7363_n 0.0035837f $X=37.195 $Y=1.985 $X2=0 $Y2=0
cc_4494 N_D[5]_M1183_g N_VPWR_c_7363_n 0.0035837f $X=37.665 $Y=1.985 $X2=0 $Y2=0
cc_4495 N_D[5]_M1217_g N_VPWR_c_7364_n 0.0035837f $X=38.135 $Y=1.985 $X2=0 $Y2=0
cc_4496 N_D[5]_M1255_g N_VPWR_c_7364_n 0.0035837f $X=38.605 $Y=1.985 $X2=0 $Y2=0
cc_4497 N_D[5]_M1088_g N_Z_c_9127_n 0.00311896f $X=37.195 $Y=1.985 $X2=0 $Y2=0
cc_4498 N_D[5]_M1183_g N_Z_c_9127_n 0.00306964f $X=37.665 $Y=1.985 $X2=0 $Y2=0
cc_4499 N_D[5]_M1217_g N_Z_c_9127_n 0.00306964f $X=38.135 $Y=1.985 $X2=0 $Y2=0
cc_4500 N_D[5]_M1255_g N_Z_c_9127_n 0.00470782f $X=38.605 $Y=1.985 $X2=0 $Y2=0
cc_4501 N_D[5]_c_5713_n N_Z_c_9127_n 0.00846955f $X=38.5 $Y=1.16 $X2=0 $Y2=0
cc_4502 N_D[5]_M1088_g N_A_6887_311#_c_11933_n 0.013247f $X=37.195 $Y=1.985
+ $X2=0 $Y2=0
cc_4503 N_D[5]_M1183_g N_A_6887_311#_c_11955_n 0.00916655f $X=37.665 $Y=1.985
+ $X2=0 $Y2=0
cc_4504 N_D[5]_M1217_g N_A_6887_311#_c_11955_n 0.00916655f $X=38.135 $Y=1.985
+ $X2=0 $Y2=0
cc_4505 N_D[5]_c_5711_n N_A_6887_311#_c_11955_n 7.15862e-19 $X=38.045 $Y=1.16
+ $X2=0 $Y2=0
cc_4506 N_D[5]_c_5713_n N_A_6887_311#_c_11955_n 0.0387168f $X=38.5 $Y=1.16 $X2=0
+ $Y2=0
cc_4507 N_D[5]_M1088_g N_A_6887_311#_c_11959_n 8.61029e-19 $X=37.195 $Y=1.985
+ $X2=0 $Y2=0
cc_4508 N_D[5]_M1183_g N_A_6887_311#_c_11959_n 5.79575e-19 $X=37.665 $Y=1.985
+ $X2=0 $Y2=0
cc_4509 N_D[5]_c_5712_n N_A_6887_311#_c_11959_n 8.03631e-19 $X=37.755 $Y=1.16
+ $X2=0 $Y2=0
cc_4510 N_D[5]_c_5713_n N_A_6887_311#_c_11959_n 0.0191156f $X=38.5 $Y=1.16 $X2=0
+ $Y2=0
cc_4511 N_D[5]_M1217_g N_A_6887_311#_c_11963_n 5.79575e-19 $X=38.135 $Y=1.985
+ $X2=0 $Y2=0
cc_4512 N_D[5]_M1255_g N_A_6887_311#_c_11963_n 0.00215964f $X=38.605 $Y=1.985
+ $X2=0 $Y2=0
cc_4513 N_D[5]_c_5713_n N_A_6887_311#_c_11963_n 0.0217153f $X=38.5 $Y=1.16 $X2=0
+ $Y2=0
cc_4514 N_D[5]_c_5714_n N_A_6887_311#_c_11963_n 8.03631e-19 $X=38.605 $Y=1.16
+ $X2=0 $Y2=0
cc_4515 N_D[5]_M1088_g N_A_6887_311#_c_11935_n 0.00232998f $X=37.195 $Y=1.985
+ $X2=25.99 $Y2=0.51
cc_4516 N_D[5]_M1183_g N_A_6887_311#_c_11968_n 0.00232998f $X=37.665 $Y=1.985
+ $X2=0 $Y2=0
cc_4517 N_D[5]_M1217_g N_A_6887_311#_c_11968_n 0.00232998f $X=38.135 $Y=1.985
+ $X2=0 $Y2=0
cc_4518 N_D[5]_M1088_g N_A_6887_311#_c_11970_n 0.00977623f $X=37.195 $Y=1.985
+ $X2=0 $Y2=0
cc_4519 N_D[5]_M1183_g N_A_6887_311#_c_11970_n 0.00911325f $X=37.665 $Y=1.985
+ $X2=0 $Y2=0
cc_4520 N_D[5]_M1217_g N_A_6887_311#_c_11970_n 7.05028e-19 $X=38.135 $Y=1.985
+ $X2=0 $Y2=0
cc_4521 N_D[5]_M1183_g N_A_6887_311#_c_11973_n 7.05028e-19 $X=37.665 $Y=1.985
+ $X2=0 $Y2=0
cc_4522 N_D[5]_M1217_g N_A_6887_311#_c_11973_n 0.00911325f $X=38.135 $Y=1.985
+ $X2=0 $Y2=0
cc_4523 N_D[5]_M1255_g N_A_6887_311#_c_11973_n 0.00847082f $X=38.605 $Y=1.985
+ $X2=0 $Y2=0
cc_4524 N_D[5]_M1088_g N_A_6887_311#_c_11938_n 0.00333758f $X=37.195 $Y=1.985
+ $X2=0 $Y2=0
cc_4525 N_D[5]_M1029_g N_VGND_c_12755_n 0.00321269f $X=37.22 $Y=0.56 $X2=0 $Y2=0
cc_4526 N_D[5]_M1057_g N_VGND_c_12755_n 2.6376e-19 $X=37.64 $Y=0.56 $X2=0 $Y2=0
cc_4527 N_D[5]_M1057_g N_VGND_c_12757_n 0.0019152f $X=37.64 $Y=0.56 $X2=0 $Y2=0
cc_4528 N_D[5]_M1247_g N_VGND_c_12757_n 0.00166854f $X=38.16 $Y=0.56 $X2=0 $Y2=0
cc_4529 N_D[5]_M1262_g N_VGND_c_12757_n 2.64031e-19 $X=38.58 $Y=0.56 $X2=0 $Y2=0
cc_4530 N_D[5]_M1262_g N_VGND_c_12759_n 0.00345859f $X=38.58 $Y=0.56 $X2=0 $Y2=0
cc_4531 N_D[5]_M1029_g VGND 0.00702263f $X=37.22 $Y=0.56 $X2=0 $Y2=0
cc_4532 N_D[5]_M1057_g VGND 0.00624811f $X=37.64 $Y=0.56 $X2=0 $Y2=0
cc_4533 N_D[5]_M1247_g VGND 0.00593887f $X=38.16 $Y=0.56 $X2=0 $Y2=0
cc_4534 N_D[5]_M1262_g VGND 0.0111368f $X=38.58 $Y=0.56 $X2=0 $Y2=0
cc_4535 N_D[5]_M1029_g N_VGND_c_12887_n 0.00422241f $X=37.22 $Y=0.56 $X2=0 $Y2=0
cc_4536 N_D[5]_M1057_g N_VGND_c_12887_n 0.00430643f $X=37.64 $Y=0.56 $X2=0 $Y2=0
cc_4537 N_D[5]_M1247_g N_VGND_c_12889_n 0.00422241f $X=38.16 $Y=0.56 $X2=0 $Y2=0
cc_4538 N_D[5]_M1262_g N_VGND_c_12889_n 0.00551064f $X=38.58 $Y=0.56 $X2=0 $Y2=0
cc_4539 N_D[5]_M1029_g N_A_6937_66#_c_14871_n 0.00261078f $X=37.22 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_4540 N_D[5]_M1029_g N_A_6937_66#_c_14872_n 0.0121912f $X=37.22 $Y=0.56 $X2=0
+ $Y2=0
cc_4541 N_D[5]_M1029_g N_A_6937_66#_c_14892_n 0.00699463f $X=37.22 $Y=0.56 $X2=0
+ $Y2=0
cc_4542 N_D[5]_M1057_g N_A_6937_66#_c_14892_n 0.00661764f $X=37.64 $Y=0.56 $X2=0
+ $Y2=0
cc_4543 N_D[5]_M1247_g N_A_6937_66#_c_14892_n 5.22365e-19 $X=38.16 $Y=0.56 $X2=0
+ $Y2=0
cc_4544 N_D[5]_M1057_g N_A_6937_66#_c_14874_n 0.00900364f $X=37.64 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_4545 N_D[5]_M1247_g N_A_6937_66#_c_14874_n 0.00986515f $X=38.16 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_4546 N_D[5]_M1262_g N_A_6937_66#_c_14874_n 0.00228093f $X=38.58 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_4547 N_D[5]_c_5711_n N_A_6937_66#_c_14874_n 0.00463549f $X=38.045 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_4548 N_D[5]_c_5713_n N_A_6937_66#_c_14874_n 0.0608884f $X=38.5 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_4549 N_D[5]_c_5714_n N_A_6937_66#_c_14874_n 0.00208088f $X=38.605 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_4550 N_D[5]_M1057_g N_A_6937_66#_c_14901_n 5.22365e-19 $X=37.64 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_4551 N_D[5]_M1247_g N_A_6937_66#_c_14901_n 0.00661134f $X=38.16 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_4552 N_D[5]_M1262_g N_A_6937_66#_c_14901_n 0.00529286f $X=38.58 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_4553 N_D[5]_M1029_g N_A_6937_66#_c_14875_n 0.00128201f $X=37.22 $Y=0.56 $X2=0
+ $Y2=0
cc_4554 N_D[5]_M1057_g N_A_6937_66#_c_14875_n 8.68782e-19 $X=37.64 $Y=0.56 $X2=0
+ $Y2=0
cc_4555 N_D[5]_c_5712_n N_A_6937_66#_c_14875_n 0.00208088f $X=37.755 $Y=1.16
+ $X2=0 $Y2=0
cc_4556 N_D[5]_c_5713_n N_A_6937_66#_c_14875_n 0.018367f $X=38.5 $Y=1.16 $X2=0
+ $Y2=0
cc_4557 N_D[13]_M1102_g N_VPWR_c_7283_n 0.00389633f $X=37.195 $Y=3.455 $X2=0
+ $Y2=0
cc_4558 N_D[13]_M1186_g N_VPWR_c_7285_n 0.00208662f $X=37.665 $Y=3.455 $X2=0
+ $Y2=0
cc_4559 N_D[13]_M1224_g N_VPWR_c_7285_n 0.00208662f $X=38.135 $Y=3.455 $X2=0
+ $Y2=0
cc_4560 N_D[13]_M1264_g N_VPWR_c_7287_n 0.00374733f $X=38.605 $Y=3.455 $X2=0
+ $Y2=0
cc_4561 N_D[13]_M1102_g VPWR 0.00573859f $X=37.195 $Y=3.455 $X2=0 $Y2=0
cc_4562 N_D[13]_M1186_g VPWR 0.00445624f $X=37.665 $Y=3.455 $X2=0 $Y2=0
cc_4563 N_D[13]_M1224_g VPWR 0.00445624f $X=38.135 $Y=3.455 $X2=0 $Y2=0
cc_4564 N_D[13]_M1264_g VPWR 0.00691494f $X=38.605 $Y=3.455 $X2=0 $Y2=0
cc_4565 N_D[13]_M1102_g N_VPWR_c_7363_n 0.0035837f $X=37.195 $Y=3.455 $X2=0
+ $Y2=0
cc_4566 N_D[13]_M1186_g N_VPWR_c_7363_n 0.0035837f $X=37.665 $Y=3.455 $X2=0
+ $Y2=0
cc_4567 N_D[13]_M1224_g N_VPWR_c_7364_n 0.0035837f $X=38.135 $Y=3.455 $X2=0
+ $Y2=0
cc_4568 N_D[13]_M1264_g N_VPWR_c_7364_n 0.0035837f $X=38.605 $Y=3.455 $X2=0
+ $Y2=0
cc_4569 N_D[13]_M1102_g N_Z_c_9128_n 0.00311896f $X=37.195 $Y=3.455 $X2=0 $Y2=0
cc_4570 N_D[13]_M1186_g N_Z_c_9128_n 0.00306964f $X=37.665 $Y=3.455 $X2=0 $Y2=0
cc_4571 N_D[13]_M1224_g N_Z_c_9128_n 0.00306964f $X=38.135 $Y=3.455 $X2=0 $Y2=0
cc_4572 N_D[13]_M1264_g N_Z_c_9128_n 0.00470782f $X=38.605 $Y=3.455 $X2=0 $Y2=0
cc_4573 N_D[13]_c_5806_n N_Z_c_9128_n 0.00846955f $X=38.5 $Y=4.28 $X2=0 $Y2=0
cc_4574 N_D[13]_M1102_g N_A_6887_613#_c_12064_n 0.013247f $X=37.195 $Y=3.455
+ $X2=0 $Y2=0
cc_4575 N_D[13]_M1186_g N_A_6887_613#_c_12086_n 0.00916655f $X=37.665 $Y=3.455
+ $X2=0 $Y2=0
cc_4576 N_D[13]_M1224_g N_A_6887_613#_c_12086_n 0.00916655f $X=38.135 $Y=3.455
+ $X2=0 $Y2=0
cc_4577 N_D[13]_c_5804_n N_A_6887_613#_c_12086_n 7.15862e-19 $X=38.045 $Y=4.28
+ $X2=0 $Y2=0
cc_4578 N_D[13]_c_5806_n N_A_6887_613#_c_12086_n 0.0387168f $X=38.5 $Y=4.28
+ $X2=0 $Y2=0
cc_4579 N_D[13]_M1102_g N_A_6887_613#_c_12090_n 8.61029e-19 $X=37.195 $Y=3.455
+ $X2=0 $Y2=0
cc_4580 N_D[13]_M1186_g N_A_6887_613#_c_12090_n 5.79575e-19 $X=37.665 $Y=3.455
+ $X2=0 $Y2=0
cc_4581 N_D[13]_c_5805_n N_A_6887_613#_c_12090_n 8.03631e-19 $X=37.755 $Y=4.28
+ $X2=0 $Y2=0
cc_4582 N_D[13]_c_5806_n N_A_6887_613#_c_12090_n 0.0191156f $X=38.5 $Y=4.28
+ $X2=0 $Y2=0
cc_4583 N_D[13]_M1224_g N_A_6887_613#_c_12094_n 5.79575e-19 $X=38.135 $Y=3.455
+ $X2=0 $Y2=0
cc_4584 N_D[13]_M1264_g N_A_6887_613#_c_12094_n 0.00215964f $X=38.605 $Y=3.455
+ $X2=0 $Y2=0
cc_4585 N_D[13]_c_5806_n N_A_6887_613#_c_12094_n 0.0217153f $X=38.5 $Y=4.28
+ $X2=0 $Y2=0
cc_4586 N_D[13]_c_5807_n N_A_6887_613#_c_12094_n 8.03631e-19 $X=38.605 $Y=4.28
+ $X2=0 $Y2=0
cc_4587 N_D[13]_M1102_g N_A_6887_613#_c_12066_n 0.00232998f $X=37.195 $Y=3.455
+ $X2=25.99 $Y2=0.51
cc_4588 N_D[13]_M1186_g N_A_6887_613#_c_12099_n 0.00232998f $X=37.665 $Y=3.455
+ $X2=0 $Y2=0
cc_4589 N_D[13]_M1224_g N_A_6887_613#_c_12099_n 0.00232998f $X=38.135 $Y=3.455
+ $X2=0 $Y2=0
cc_4590 N_D[13]_M1102_g N_A_6887_613#_c_12069_n 0.00333758f $X=37.195 $Y=3.455
+ $X2=0 $Y2=0
cc_4591 N_D[13]_M1102_g N_A_6887_613#_c_12102_n 0.00977623f $X=37.195 $Y=3.455
+ $X2=0 $Y2=0
cc_4592 N_D[13]_M1186_g N_A_6887_613#_c_12102_n 0.00911325f $X=37.665 $Y=3.455
+ $X2=0 $Y2=0
cc_4593 N_D[13]_M1224_g N_A_6887_613#_c_12102_n 7.05028e-19 $X=38.135 $Y=3.455
+ $X2=0 $Y2=0
cc_4594 N_D[13]_M1186_g N_A_6887_613#_c_12105_n 7.05028e-19 $X=37.665 $Y=3.455
+ $X2=0 $Y2=0
cc_4595 N_D[13]_M1224_g N_A_6887_613#_c_12105_n 0.00911325f $X=38.135 $Y=3.455
+ $X2=0 $Y2=0
cc_4596 N_D[13]_M1264_g N_A_6887_613#_c_12105_n 0.00847082f $X=38.605 $Y=3.455
+ $X2=0 $Y2=0
cc_4597 N_D[13]_M1132_g N_VGND_c_12756_n 0.00321269f $X=37.22 $Y=4.88 $X2=0
+ $Y2=0
cc_4598 N_D[13]_M1136_g N_VGND_c_12756_n 2.6376e-19 $X=37.64 $Y=4.88 $X2=0 $Y2=0
cc_4599 N_D[13]_M1136_g N_VGND_c_12758_n 0.0019152f $X=37.64 $Y=4.88 $X2=0 $Y2=0
cc_4600 N_D[13]_M1274_g N_VGND_c_12758_n 0.00166854f $X=38.16 $Y=4.88 $X2=0
+ $Y2=0
cc_4601 N_D[13]_M1298_g N_VGND_c_12758_n 2.64031e-19 $X=38.58 $Y=4.88 $X2=0
+ $Y2=0
cc_4602 N_D[13]_M1298_g N_VGND_c_12760_n 0.00345859f $X=38.58 $Y=4.88 $X2=0
+ $Y2=0
cc_4603 N_D[13]_M1132_g VGND 0.00702263f $X=37.22 $Y=4.88 $X2=0 $Y2=0
cc_4604 N_D[13]_M1136_g VGND 0.00624811f $X=37.64 $Y=4.88 $X2=0 $Y2=0
cc_4605 N_D[13]_M1274_g VGND 0.00593887f $X=38.16 $Y=4.88 $X2=0 $Y2=0
cc_4606 N_D[13]_M1298_g VGND 0.0111368f $X=38.58 $Y=4.88 $X2=0 $Y2=0
cc_4607 N_D[13]_M1132_g N_VGND_c_12888_n 0.00422241f $X=37.22 $Y=4.88 $X2=0
+ $Y2=0
cc_4608 N_D[13]_M1136_g N_VGND_c_12888_n 0.00430643f $X=37.64 $Y=4.88 $X2=0
+ $Y2=0
cc_4609 N_D[13]_M1274_g N_VGND_c_12890_n 0.00422241f $X=38.16 $Y=4.88 $X2=0
+ $Y2=0
cc_4610 N_D[13]_M1298_g N_VGND_c_12890_n 0.00551064f $X=38.58 $Y=4.88 $X2=0
+ $Y2=0
cc_4611 N_D[13]_M1132_g N_A_6937_918#_c_14955_n 0.00261078f $X=37.22 $Y=4.88
+ $X2=25.99 $Y2=0.51
cc_4612 N_D[13]_M1132_g N_A_6937_918#_c_14956_n 0.0121912f $X=37.22 $Y=4.88
+ $X2=0 $Y2=0
cc_4613 N_D[13]_M1136_g N_A_6937_918#_c_14976_n 0.00900364f $X=37.64 $Y=4.88
+ $X2=0 $Y2=0
cc_4614 N_D[13]_M1274_g N_A_6937_918#_c_14976_n 0.00899636f $X=38.16 $Y=4.88
+ $X2=0 $Y2=0
cc_4615 N_D[13]_c_5804_n N_A_6937_918#_c_14976_n 0.00463549f $X=38.045 $Y=4.28
+ $X2=0 $Y2=0
cc_4616 N_D[13]_c_5806_n N_A_6937_918#_c_14976_n 0.0394855f $X=38.5 $Y=4.28
+ $X2=0 $Y2=0
cc_4617 N_D[13]_M1132_g N_A_6937_918#_c_14958_n 0.00827664f $X=37.22 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_4618 N_D[13]_M1136_g N_A_6937_918#_c_14958_n 0.00748643f $X=37.64 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_4619 N_D[13]_M1274_g N_A_6937_918#_c_14958_n 5.22365e-19 $X=38.16 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_4620 N_D[13]_c_5805_n N_A_6937_918#_c_14958_n 0.00208088f $X=37.755 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_4621 N_D[13]_c_5806_n N_A_6937_918#_c_14958_n 0.018367f $X=38.5 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_4622 N_D[13]_M1136_g N_A_6937_918#_c_14959_n 5.22365e-19 $X=37.64 $Y=4.88
+ $X2=0 $Y2=0
cc_4623 N_D[13]_M1274_g N_A_6937_918#_c_14959_n 0.00748012f $X=38.16 $Y=4.88
+ $X2=0 $Y2=0
cc_4624 N_D[13]_M1298_g N_A_6937_918#_c_14959_n 0.00757379f $X=38.58 $Y=4.88
+ $X2=0 $Y2=0
cc_4625 N_D[13]_c_5806_n N_A_6937_918#_c_14959_n 0.021403f $X=38.5 $Y=4.28 $X2=0
+ $Y2=0
cc_4626 N_D[13]_c_5807_n N_A_6937_918#_c_14959_n 0.00208088f $X=38.605 $Y=4.28
+ $X2=0 $Y2=0
cc_4627 N_D[6]_M1099_g N_D[14]_M1109_g 0.0130744f $X=39.595 $Y=1.985 $X2=0 $Y2=0
cc_4628 N_D[6]_M1176_g N_D[14]_M1184_g 0.0130744f $X=40.065 $Y=1.985 $X2=0 $Y2=0
cc_4629 N_D[6]_M1246_g N_D[14]_M1251_g 0.0130744f $X=40.535 $Y=1.985 $X2=0 $Y2=0
cc_4630 N_D[6]_M1282_g N_D[14]_M1293_g 0.0130744f $X=41.005 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_4631 N_D[6]_M1099_g N_VPWR_c_7289_n 0.00374733f $X=39.595 $Y=1.985 $X2=0
+ $Y2=0
cc_4632 N_D[6]_M1176_g N_VPWR_c_7291_n 0.00208662f $X=40.065 $Y=1.985 $X2=0
+ $Y2=0
cc_4633 N_D[6]_M1246_g N_VPWR_c_7291_n 0.00208662f $X=40.535 $Y=1.985 $X2=0
+ $Y2=0
cc_4634 N_D[6]_M1246_g N_VPWR_c_7293_n 0.0035837f $X=40.535 $Y=1.985 $X2=0 $Y2=0
cc_4635 N_D[6]_M1282_g N_VPWR_c_7293_n 0.0035837f $X=41.005 $Y=1.985 $X2=0 $Y2=0
cc_4636 N_D[6]_M1282_g N_VPWR_c_7294_n 0.00389633f $X=41.005 $Y=1.985 $X2=0
+ $Y2=0
cc_4637 N_D[6]_M1099_g VPWR 0.00691494f $X=39.595 $Y=1.985 $X2=0 $Y2=0
cc_4638 N_D[6]_M1176_g VPWR 0.00445624f $X=40.065 $Y=1.985 $X2=0 $Y2=0
cc_4639 N_D[6]_M1246_g VPWR 0.00445624f $X=40.535 $Y=1.985 $X2=0 $Y2=0
cc_4640 N_D[6]_M1282_g VPWR 0.00573859f $X=41.005 $Y=1.985 $X2=0 $Y2=0
cc_4641 N_D[6]_M1099_g N_VPWR_c_7365_n 0.0035837f $X=39.595 $Y=1.985 $X2=0 $Y2=0
cc_4642 N_D[6]_M1176_g N_VPWR_c_7365_n 0.0035837f $X=40.065 $Y=1.985 $X2=0 $Y2=0
cc_4643 N_D[6]_M1099_g N_Z_c_9127_n 0.00470782f $X=39.595 $Y=1.985 $X2=0 $Y2=0
cc_4644 N_D[6]_M1176_g N_Z_c_9127_n 0.00306964f $X=40.065 $Y=1.985 $X2=0 $Y2=0
cc_4645 N_D[6]_M1246_g N_Z_c_9127_n 0.00306964f $X=40.535 $Y=1.985 $X2=0 $Y2=0
cc_4646 N_D[6]_M1282_g N_Z_c_9127_n 0.00311896f $X=41.005 $Y=1.985 $X2=0 $Y2=0
cc_4647 N_D[6]_c_5897_n N_Z_c_9127_n 0.00846955f $X=40.72 $Y=1.16 $X2=0 $Y2=0
cc_4648 N_D[6]_M1176_g N_A_7937_297#_c_12200_n 0.00916655f $X=40.065 $Y=1.985
+ $X2=0 $Y2=0
cc_4649 N_D[6]_M1246_g N_A_7937_297#_c_12200_n 0.00916655f $X=40.535 $Y=1.985
+ $X2=0 $Y2=0
cc_4650 N_D[6]_c_5895_n N_A_7937_297#_c_12200_n 7.15862e-19 $X=40.445 $Y=1.16
+ $X2=0 $Y2=0
cc_4651 N_D[6]_c_5897_n N_A_7937_297#_c_12200_n 0.0387168f $X=40.72 $Y=1.16
+ $X2=0 $Y2=0
cc_4652 N_D[6]_M1282_g N_A_7937_297#_c_12195_n 0.013247f $X=41.005 $Y=1.985
+ $X2=0 $Y2=0
cc_4653 N_D[6]_M1099_g N_A_7937_297#_c_12205_n 0.00215964f $X=39.595 $Y=1.985
+ $X2=0 $Y2=0
cc_4654 N_D[6]_M1176_g N_A_7937_297#_c_12205_n 5.79575e-19 $X=40.065 $Y=1.985
+ $X2=0 $Y2=0
cc_4655 N_D[6]_c_5896_n N_A_7937_297#_c_12205_n 8.03631e-19 $X=40.155 $Y=1.16
+ $X2=0 $Y2=0
cc_4656 N_D[6]_c_5897_n N_A_7937_297#_c_12205_n 0.0217153f $X=40.72 $Y=1.16
+ $X2=0 $Y2=0
cc_4657 N_D[6]_M1246_g N_A_7937_297#_c_12209_n 5.79575e-19 $X=40.535 $Y=1.985
+ $X2=0 $Y2=0
cc_4658 N_D[6]_M1282_g N_A_7937_297#_c_12209_n 8.61029e-19 $X=41.005 $Y=1.985
+ $X2=0 $Y2=0
cc_4659 N_D[6]_c_5897_n N_A_7937_297#_c_12209_n 0.0191156f $X=40.72 $Y=1.16
+ $X2=0 $Y2=0
cc_4660 N_D[6]_c_5898_n N_A_7937_297#_c_12209_n 8.03631e-19 $X=41.005 $Y=1.16
+ $X2=0 $Y2=0
cc_4661 N_D[6]_M1176_g N_A_7937_297#_c_12213_n 0.00232998f $X=40.065 $Y=1.985
+ $X2=0 $Y2=0
cc_4662 N_D[6]_M1246_g N_A_7937_297#_c_12213_n 0.00232998f $X=40.535 $Y=1.985
+ $X2=0 $Y2=0
cc_4663 N_D[6]_M1282_g N_A_7937_297#_c_12196_n 0.00232998f $X=41.005 $Y=1.985
+ $X2=0 $Y2=0
cc_4664 N_D[6]_M1099_g N_A_7937_297#_c_12216_n 0.00847082f $X=39.595 $Y=1.985
+ $X2=0 $Y2=0
cc_4665 N_D[6]_M1176_g N_A_7937_297#_c_12216_n 0.00911325f $X=40.065 $Y=1.985
+ $X2=0 $Y2=0
cc_4666 N_D[6]_M1246_g N_A_7937_297#_c_12216_n 7.05028e-19 $X=40.535 $Y=1.985
+ $X2=0 $Y2=0
cc_4667 N_D[6]_M1176_g N_A_7937_297#_c_12219_n 7.05028e-19 $X=40.065 $Y=1.985
+ $X2=0 $Y2=0
cc_4668 N_D[6]_M1246_g N_A_7937_297#_c_12219_n 0.00911325f $X=40.535 $Y=1.985
+ $X2=0 $Y2=0
cc_4669 N_D[6]_M1282_g N_A_7937_297#_c_12219_n 0.00977623f $X=41.005 $Y=1.985
+ $X2=0 $Y2=0
cc_4670 N_D[6]_M1282_g N_A_7937_297#_c_12197_n 0.00333758f $X=41.005 $Y=1.985
+ $X2=0 $Y2=0
cc_4671 N_D[6]_M1069_g N_VGND_c_12763_n 0.00345859f $X=39.62 $Y=0.56 $X2=0 $Y2=0
cc_4672 N_D[6]_M1069_g N_VGND_c_12765_n 2.64031e-19 $X=39.62 $Y=0.56 $X2=0 $Y2=0
cc_4673 N_D[6]_M1122_g N_VGND_c_12765_n 0.00166854f $X=40.04 $Y=0.56 $X2=0 $Y2=0
cc_4674 N_D[6]_M1147_g N_VGND_c_12765_n 0.0019152f $X=40.56 $Y=0.56 $X2=0 $Y2=0
cc_4675 N_D[6]_M1147_g N_VGND_c_12767_n 0.00430643f $X=40.56 $Y=0.56 $X2=0 $Y2=0
cc_4676 N_D[6]_M1258_g N_VGND_c_12767_n 0.00422241f $X=40.98 $Y=0.56 $X2=0 $Y2=0
cc_4677 N_D[6]_M1147_g N_VGND_c_12769_n 2.6376e-19 $X=40.56 $Y=0.56 $X2=0 $Y2=0
cc_4678 N_D[6]_M1258_g N_VGND_c_12769_n 0.00321269f $X=40.98 $Y=0.56 $X2=0 $Y2=0
cc_4679 N_D[6]_M1069_g VGND 0.0111368f $X=39.62 $Y=0.56 $X2=0 $Y2=0
cc_4680 N_D[6]_M1122_g VGND 0.00593887f $X=40.04 $Y=0.56 $X2=0 $Y2=0
cc_4681 N_D[6]_M1147_g VGND 0.00624811f $X=40.56 $Y=0.56 $X2=0 $Y2=0
cc_4682 N_D[6]_M1258_g VGND 0.00702263f $X=40.98 $Y=0.56 $X2=0 $Y2=0
cc_4683 N_D[6]_M1069_g N_VGND_c_12891_n 0.00551064f $X=39.62 $Y=0.56 $X2=0 $Y2=0
cc_4684 N_D[6]_M1122_g N_VGND_c_12891_n 0.00422241f $X=40.04 $Y=0.56 $X2=0 $Y2=0
cc_4685 N_D[6]_M1069_g N_A_7939_47#_c_15041_n 0.00529286f $X=39.62 $Y=0.56 $X2=0
+ $Y2=0
cc_4686 N_D[6]_M1122_g N_A_7939_47#_c_15041_n 0.00661134f $X=40.04 $Y=0.56 $X2=0
+ $Y2=0
cc_4687 N_D[6]_M1147_g N_A_7939_47#_c_15041_n 5.22365e-19 $X=40.56 $Y=0.56 $X2=0
+ $Y2=0
cc_4688 N_D[6]_M1122_g N_A_7939_47#_c_15044_n 0.00899636f $X=40.04 $Y=0.56 $X2=0
+ $Y2=0
cc_4689 N_D[6]_M1147_g N_A_7939_47#_c_15044_n 0.00900364f $X=40.56 $Y=0.56 $X2=0
+ $Y2=0
cc_4690 N_D[6]_c_5895_n N_A_7939_47#_c_15044_n 0.00463549f $X=40.445 $Y=1.16
+ $X2=0 $Y2=0
cc_4691 N_D[6]_c_5897_n N_A_7939_47#_c_15044_n 0.0394855f $X=40.72 $Y=1.16 $X2=0
+ $Y2=0
cc_4692 N_D[6]_M1069_g N_A_7939_47#_c_15033_n 0.00228093f $X=39.62 $Y=0.56 $X2=0
+ $Y2=0
cc_4693 N_D[6]_M1122_g N_A_7939_47#_c_15033_n 8.68782e-19 $X=40.04 $Y=0.56 $X2=0
+ $Y2=0
cc_4694 N_D[6]_c_5896_n N_A_7939_47#_c_15033_n 0.00208088f $X=40.155 $Y=1.16
+ $X2=0 $Y2=0
cc_4695 N_D[6]_c_5897_n N_A_7939_47#_c_15033_n 0.021403f $X=40.72 $Y=1.16 $X2=0
+ $Y2=0
cc_4696 N_D[6]_M1122_g N_A_7939_47#_c_15052_n 5.22365e-19 $X=40.04 $Y=0.56 $X2=0
+ $Y2=0
cc_4697 N_D[6]_M1147_g N_A_7939_47#_c_15052_n 0.00661764f $X=40.56 $Y=0.56 $X2=0
+ $Y2=0
cc_4698 N_D[6]_M1258_g N_A_7939_47#_c_15052_n 0.00699463f $X=40.98 $Y=0.56 $X2=0
+ $Y2=0
cc_4699 N_D[6]_M1258_g N_A_7939_47#_c_15034_n 0.0121912f $X=40.98 $Y=0.56 $X2=0
+ $Y2=0
cc_4700 N_D[6]_M1258_g N_A_7939_47#_c_15035_n 0.00261078f $X=40.98 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_4701 N_D[6]_M1147_g N_A_7939_47#_c_15040_n 8.68782e-19 $X=40.56 $Y=0.56 $X2=0
+ $Y2=0
cc_4702 N_D[6]_M1258_g N_A_7939_47#_c_15040_n 0.00128201f $X=40.98 $Y=0.56 $X2=0
+ $Y2=0
cc_4703 N_D[6]_c_5897_n N_A_7939_47#_c_15040_n 0.018367f $X=40.72 $Y=1.16 $X2=0
+ $Y2=0
cc_4704 N_D[6]_c_5898_n N_A_7939_47#_c_15040_n 0.00208088f $X=41.005 $Y=1.16
+ $X2=0 $Y2=0
cc_4705 N_D[14]_M1109_g N_VPWR_c_7290_n 0.00374733f $X=39.595 $Y=3.455 $X2=0
+ $Y2=0
cc_4706 N_D[14]_M1184_g N_VPWR_c_7292_n 0.00208662f $X=40.065 $Y=3.455 $X2=0
+ $Y2=0
cc_4707 N_D[14]_M1251_g N_VPWR_c_7292_n 0.00208662f $X=40.535 $Y=3.455 $X2=0
+ $Y2=0
cc_4708 N_D[14]_M1251_g N_VPWR_c_7293_n 0.0035837f $X=40.535 $Y=3.455 $X2=0
+ $Y2=0
cc_4709 N_D[14]_M1293_g N_VPWR_c_7293_n 0.0035837f $X=41.005 $Y=3.455 $X2=0
+ $Y2=0
cc_4710 N_D[14]_M1293_g N_VPWR_c_7295_n 0.00389633f $X=41.005 $Y=3.455 $X2=0
+ $Y2=0
cc_4711 N_D[14]_M1109_g VPWR 0.00691494f $X=39.595 $Y=3.455 $X2=0 $Y2=0
cc_4712 N_D[14]_M1184_g VPWR 0.00445624f $X=40.065 $Y=3.455 $X2=0 $Y2=0
cc_4713 N_D[14]_M1251_g VPWR 0.00445624f $X=40.535 $Y=3.455 $X2=0 $Y2=0
cc_4714 N_D[14]_M1293_g VPWR 0.00573859f $X=41.005 $Y=3.455 $X2=0 $Y2=0
cc_4715 N_D[14]_M1109_g N_VPWR_c_7365_n 0.0035837f $X=39.595 $Y=3.455 $X2=0
+ $Y2=0
cc_4716 N_D[14]_M1184_g N_VPWR_c_7365_n 0.0035837f $X=40.065 $Y=3.455 $X2=0
+ $Y2=0
cc_4717 N_D[14]_M1109_g N_Z_c_9128_n 0.00470782f $X=39.595 $Y=3.455 $X2=0 $Y2=0
cc_4718 N_D[14]_M1184_g N_Z_c_9128_n 0.00306964f $X=40.065 $Y=3.455 $X2=0 $Y2=0
cc_4719 N_D[14]_M1251_g N_Z_c_9128_n 0.00306964f $X=40.535 $Y=3.455 $X2=0 $Y2=0
cc_4720 N_D[14]_M1293_g N_Z_c_9128_n 0.00311896f $X=41.005 $Y=3.455 $X2=0 $Y2=0
cc_4721 N_D[14]_c_5992_n N_Z_c_9128_n 0.00846955f $X=40.72 $Y=4.28 $X2=0 $Y2=0
cc_4722 N_D[14]_M1184_g N_A_7937_591#_c_12328_n 0.00916655f $X=40.065 $Y=3.455
+ $X2=0 $Y2=0
cc_4723 N_D[14]_M1251_g N_A_7937_591#_c_12328_n 0.00916655f $X=40.535 $Y=3.455
+ $X2=0 $Y2=0
cc_4724 N_D[14]_c_5990_n N_A_7937_591#_c_12328_n 7.15862e-19 $X=40.445 $Y=4.28
+ $X2=0 $Y2=0
cc_4725 N_D[14]_c_5992_n N_A_7937_591#_c_12328_n 0.0387168f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4726 N_D[14]_M1293_g N_A_7937_591#_c_12323_n 0.013247f $X=41.005 $Y=3.455
+ $X2=0 $Y2=0
cc_4727 N_D[14]_M1109_g N_A_7937_591#_c_12333_n 0.00215964f $X=39.595 $Y=3.455
+ $X2=0 $Y2=0
cc_4728 N_D[14]_M1184_g N_A_7937_591#_c_12333_n 5.79575e-19 $X=40.065 $Y=3.455
+ $X2=0 $Y2=0
cc_4729 N_D[14]_c_5991_n N_A_7937_591#_c_12333_n 8.03631e-19 $X=40.155 $Y=4.28
+ $X2=0 $Y2=0
cc_4730 N_D[14]_c_5992_n N_A_7937_591#_c_12333_n 0.0217153f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4731 N_D[14]_M1251_g N_A_7937_591#_c_12337_n 5.79575e-19 $X=40.535 $Y=3.455
+ $X2=0 $Y2=0
cc_4732 N_D[14]_M1293_g N_A_7937_591#_c_12337_n 8.61029e-19 $X=41.005 $Y=3.455
+ $X2=0 $Y2=0
cc_4733 N_D[14]_c_5992_n N_A_7937_591#_c_12337_n 0.0191156f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4734 N_D[14]_c_5993_n N_A_7937_591#_c_12337_n 8.03631e-19 $X=41.005 $Y=4.28
+ $X2=0 $Y2=0
cc_4735 N_D[14]_M1184_g N_A_7937_591#_c_12341_n 0.00232998f $X=40.065 $Y=3.455
+ $X2=0 $Y2=0
cc_4736 N_D[14]_M1251_g N_A_7937_591#_c_12341_n 0.00232998f $X=40.535 $Y=3.455
+ $X2=0 $Y2=0
cc_4737 N_D[14]_M1293_g N_A_7937_591#_c_12324_n 0.00232998f $X=41.005 $Y=3.455
+ $X2=0 $Y2=0
cc_4738 N_D[14]_M1109_g N_A_7937_591#_c_12344_n 0.00847082f $X=39.595 $Y=3.455
+ $X2=0 $Y2=0
cc_4739 N_D[14]_M1184_g N_A_7937_591#_c_12344_n 0.00911325f $X=40.065 $Y=3.455
+ $X2=0 $Y2=0
cc_4740 N_D[14]_M1251_g N_A_7937_591#_c_12344_n 7.05028e-19 $X=40.535 $Y=3.455
+ $X2=0 $Y2=0
cc_4741 N_D[14]_M1184_g N_A_7937_591#_c_12347_n 7.05028e-19 $X=40.065 $Y=3.455
+ $X2=0 $Y2=0
cc_4742 N_D[14]_M1251_g N_A_7937_591#_c_12347_n 0.00911325f $X=40.535 $Y=3.455
+ $X2=0 $Y2=0
cc_4743 N_D[14]_M1293_g N_A_7937_591#_c_12347_n 0.00977623f $X=41.005 $Y=3.455
+ $X2=0 $Y2=0
cc_4744 N_D[14]_M1293_g N_A_7937_591#_c_12325_n 0.00333758f $X=41.005 $Y=3.455
+ $X2=0 $Y2=0
cc_4745 N_D[14]_M1004_g N_VGND_c_12764_n 0.00345859f $X=39.62 $Y=4.88 $X2=0
+ $Y2=0
cc_4746 N_D[14]_M1004_g N_VGND_c_12766_n 2.64031e-19 $X=39.62 $Y=4.88 $X2=0
+ $Y2=0
cc_4747 N_D[14]_M1179_g N_VGND_c_12766_n 0.00166854f $X=40.04 $Y=4.88 $X2=0
+ $Y2=0
cc_4748 N_D[14]_M1189_g N_VGND_c_12766_n 0.0019152f $X=40.56 $Y=4.88 $X2=0 $Y2=0
cc_4749 N_D[14]_M1189_g N_VGND_c_12768_n 0.00430643f $X=40.56 $Y=4.88 $X2=0
+ $Y2=0
cc_4750 N_D[14]_M1305_g N_VGND_c_12768_n 0.00422241f $X=40.98 $Y=4.88 $X2=0
+ $Y2=0
cc_4751 N_D[14]_M1189_g N_VGND_c_12770_n 2.6376e-19 $X=40.56 $Y=4.88 $X2=0 $Y2=0
cc_4752 N_D[14]_M1305_g N_VGND_c_12770_n 0.00321269f $X=40.98 $Y=4.88 $X2=0
+ $Y2=0
cc_4753 N_D[14]_M1004_g VGND 0.0111368f $X=39.62 $Y=4.88 $X2=0 $Y2=0
cc_4754 N_D[14]_M1179_g VGND 0.00593887f $X=40.04 $Y=4.88 $X2=0 $Y2=0
cc_4755 N_D[14]_M1189_g VGND 0.00624811f $X=40.56 $Y=4.88 $X2=0 $Y2=0
cc_4756 N_D[14]_M1305_g VGND 0.00702263f $X=40.98 $Y=4.88 $X2=0 $Y2=0
cc_4757 N_D[14]_M1004_g N_VGND_c_12892_n 0.00551064f $X=39.62 $Y=4.88 $X2=0
+ $Y2=0
cc_4758 N_D[14]_M1179_g N_VGND_c_12892_n 0.00422241f $X=40.04 $Y=4.88 $X2=0
+ $Y2=0
cc_4759 N_D[14]_M1179_g N_A_7939_911#_c_15124_n 0.00899636f $X=40.04 $Y=4.88
+ $X2=0 $Y2=0
cc_4760 N_D[14]_M1189_g N_A_7939_911#_c_15124_n 0.00900364f $X=40.56 $Y=4.88
+ $X2=0 $Y2=0
cc_4761 N_D[14]_c_5990_n N_A_7939_911#_c_15124_n 0.00463549f $X=40.445 $Y=4.28
+ $X2=0 $Y2=0
cc_4762 N_D[14]_c_5992_n N_A_7939_911#_c_15124_n 0.0394855f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4763 N_D[14]_M1305_g N_A_7939_911#_c_15116_n 0.0121912f $X=40.98 $Y=4.88
+ $X2=0 $Y2=0
cc_4764 N_D[14]_M1305_g N_A_7939_911#_c_15117_n 0.00261078f $X=40.98 $Y=4.88
+ $X2=0 $Y2=0
cc_4765 N_D[14]_M1004_g N_A_7939_911#_c_15122_n 0.00757379f $X=39.62 $Y=4.88
+ $X2=0 $Y2=0
cc_4766 N_D[14]_M1179_g N_A_7939_911#_c_15122_n 0.00748012f $X=40.04 $Y=4.88
+ $X2=0 $Y2=0
cc_4767 N_D[14]_M1189_g N_A_7939_911#_c_15122_n 5.22365e-19 $X=40.56 $Y=4.88
+ $X2=0 $Y2=0
cc_4768 N_D[14]_c_5991_n N_A_7939_911#_c_15122_n 0.00208088f $X=40.155 $Y=4.28
+ $X2=0 $Y2=0
cc_4769 N_D[14]_c_5992_n N_A_7939_911#_c_15122_n 0.021403f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4770 N_D[14]_M1179_g N_A_7939_911#_c_15123_n 5.22365e-19 $X=40.04 $Y=4.88
+ $X2=0 $Y2=0
cc_4771 N_D[14]_M1189_g N_A_7939_911#_c_15123_n 0.00748643f $X=40.56 $Y=4.88
+ $X2=0 $Y2=0
cc_4772 N_D[14]_M1305_g N_A_7939_911#_c_15123_n 0.00827664f $X=40.98 $Y=4.88
+ $X2=0 $Y2=0
cc_4773 N_D[14]_c_5992_n N_A_7939_911#_c_15123_n 0.018367f $X=40.72 $Y=4.28
+ $X2=0 $Y2=0
cc_4774 N_D[14]_c_5993_n N_A_7939_911#_c_15123_n 0.00208088f $X=41.005 $Y=4.28
+ $X2=0 $Y2=0
cc_4775 N_A_8379_265#_c_6080_n N_A_8379_793#_c_6199_n 0.0129371f $X=41.995
+ $Y=1.475 $X2=0 $Y2=0
cc_4776 N_A_8379_265#_c_6083_n N_A_8379_793#_c_6202_n 0.0129371f $X=42.465
+ $Y=1.475 $X2=0 $Y2=0
cc_4777 N_A_8379_265#_c_6085_n N_A_8379_793#_c_6204_n 0.0129371f $X=42.935
+ $Y=1.475 $X2=0 $Y2=0
cc_4778 N_A_8379_265#_c_6087_n N_A_8379_793#_c_6206_n 0.0129371f $X=43.405
+ $Y=1.475 $X2=0 $Y2=0
cc_4779 N_A_8379_265#_c_6082_n N_S[6]_c_6317_n 0.00507426f $X=42.085 $Y=1.4
+ $X2=0 $Y2=0
cc_4780 N_A_8379_265#_c_6081_n N_S[6]_c_6320_n 0.00509391f $X=42.375 $Y=1.4
+ $X2=0 $Y2=0
cc_4781 N_A_8379_265#_c_6084_n N_S[6]_c_6322_n 0.00509204f $X=42.845 $Y=1.4
+ $X2=25.905 $Y2=4.845
cc_4782 N_A_8379_265#_c_6086_n N_S[6]_c_6324_n 0.00507688f $X=43.315 $Y=1.4
+ $X2=0 $Y2=0
cc_4783 N_A_8379_265#_c_6075_n N_S[6]_c_6326_n 6.53442e-19 $X=44.685 $Y=0.445
+ $X2=0 $Y2=0
cc_4784 N_A_8379_265#_c_6073_n N_S[6]_c_6328_n 0.0103812f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4785 N_A_8379_265#_c_6074_n N_S[6]_c_6328_n 0.0179529f $X=43.975 $Y=1.23
+ $X2=0 $Y2=0
cc_4786 N_A_8379_265#_c_6073_n N_S[6]_c_6329_n 0.0206368f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4787 N_A_8379_265#_c_6074_n N_S[6]_c_6329_n 0.0175393f $X=43.975 $Y=1.23
+ $X2=0 $Y2=0
cc_4788 N_A_8379_265#_c_6076_n N_S[6]_c_6329_n 0.0085951f $X=44.605 $Y=1.065
+ $X2=0 $Y2=0
cc_4789 N_A_8379_265#_c_6078_n N_S[6]_c_6329_n 0.00322131f $X=44.605 $Y=1.23
+ $X2=0 $Y2=0
cc_4790 N_A_8379_265#_c_6094_n N_S[6]_c_6329_n 0.00255921f $X=44.685 $Y=1.605
+ $X2=0 $Y2=0
cc_4791 N_A_8379_265#_c_6079_n N_S[6]_c_6329_n 0.00262132f $X=43.725 $Y=1.23
+ $X2=0 $Y2=0
cc_4792 N_A_8379_265#_c_6092_n N_S[6]_c_6340_n 0.0118698f $X=44.685 $Y=1.77
+ $X2=0 $Y2=0
cc_4793 N_A_8379_265#_c_6094_n N_S[6]_c_6340_n 0.00762115f $X=44.685 $Y=1.605
+ $X2=0 $Y2=0
cc_4794 N_A_8379_265#_c_6075_n N_S[6]_c_6330_n 0.00603996f $X=44.685 $Y=0.445
+ $X2=0 $Y2=0
cc_4795 N_A_8379_265#_c_6077_n N_S[6]_c_6330_n 9.67113e-19 $X=44.645 $Y=0.825
+ $X2=0 $Y2=0
cc_4796 N_A_8379_265#_c_6076_n N_S[6]_c_6331_n 0.00429801f $X=44.605 $Y=1.065
+ $X2=0 $Y2=0
cc_4797 N_A_8379_265#_c_6077_n N_S[6]_c_6331_n 0.0111895f $X=44.645 $Y=0.825
+ $X2=0 $Y2=0
cc_4798 N_A_8379_265#_c_6075_n N_S[6]_c_6332_n 0.00207203f $X=44.685 $Y=0.445
+ $X2=0 $Y2=0
cc_4799 N_A_8379_265#_c_6076_n N_S[6]_c_6333_n 0.00289358f $X=44.605 $Y=1.065
+ $X2=25.99 $Y2=4.8
cc_4800 N_A_8379_265#_c_6092_n N_S[6]_c_6333_n 0.0128834f $X=44.685 $Y=1.77
+ $X2=25.99 $Y2=4.8
cc_4801 N_A_8379_265#_c_6078_n N_S[6]_c_6333_n 0.00416423f $X=44.605 $Y=1.23
+ $X2=25.99 $Y2=4.8
cc_4802 N_A_8379_265#_c_6094_n N_S[6]_c_6333_n 0.00454075f $X=44.685 $Y=1.605
+ $X2=25.99 $Y2=4.8
cc_4803 N_A_8379_265#_c_6076_n N_S[6]_c_6337_n 0.00268644f $X=44.605 $Y=1.065
+ $X2=0 $Y2=0
cc_4804 N_A_8379_265#_c_6077_n N_S[6]_c_6337_n 0.00426435f $X=44.645 $Y=0.825
+ $X2=0 $Y2=0
cc_4805 N_A_8379_265#_c_6076_n S[6] 0.00541767f $X=44.605 $Y=1.065 $X2=0 $Y2=0
cc_4806 N_A_8379_265#_c_6078_n S[6] 0.0228692f $X=44.605 $Y=1.23 $X2=0 $Y2=0
cc_4807 N_A_8379_265#_c_6080_n N_VPWR_c_7294_n 0.00324472f $X=41.995 $Y=1.475
+ $X2=0 $Y2=0
cc_4808 N_A_8379_265#_c_6087_n N_VPWR_c_7296_n 0.00367058f $X=43.405 $Y=1.475
+ $X2=0 $Y2=0
cc_4809 N_A_8379_265#_c_6073_n N_VPWR_c_7296_n 0.0193185f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4810 N_A_8379_265#_c_6074_n N_VPWR_c_7296_n 6.4101e-19 $X=43.975 $Y=1.23
+ $X2=0 $Y2=0
cc_4811 N_A_8379_265#_c_6092_n N_VPWR_c_7296_n 0.0316788f $X=44.685 $Y=1.77
+ $X2=0 $Y2=0
cc_4812 N_A_8379_265#_c_6092_n N_VPWR_c_7298_n 0.0356181f $X=44.685 $Y=1.77
+ $X2=0 $Y2=0
cc_4813 N_A_8379_265#_c_6092_n N_VPWR_c_7340_n 0.0233824f $X=44.685 $Y=1.77
+ $X2=0 $Y2=0
cc_4814 N_A_8379_265#_c_6080_n VPWR 0.00473731f $X=41.995 $Y=1.475 $X2=0 $Y2=0
cc_4815 N_A_8379_265#_c_6083_n VPWR 0.00362156f $X=42.465 $Y=1.475 $X2=0 $Y2=0
cc_4816 N_A_8379_265#_c_6085_n VPWR 0.00362156f $X=42.935 $Y=1.475 $X2=0 $Y2=0
cc_4817 N_A_8379_265#_c_6087_n VPWR 0.00473731f $X=43.405 $Y=1.475 $X2=0 $Y2=0
cc_4818 N_A_8379_265#_c_6092_n VPWR 0.00593513f $X=44.685 $Y=1.77 $X2=0 $Y2=0
cc_4819 N_A_8379_265#_c_6084_n N_Z_c_9034_n 0.00762343f $X=42.845 $Y=1.4 $X2=0
+ $Y2=0
cc_4820 N_A_8379_265#_c_6088_n N_Z_c_9034_n 0.00704092f $X=42.465 $Y=1.4 $X2=0
+ $Y2=0
cc_4821 N_A_8379_265#_c_6082_n N_Z_c_9085_n 0.00248496f $X=42.085 $Y=1.4 $X2=0
+ $Y2=0
cc_4822 N_A_8379_265#_c_6081_n N_Z_c_9088_n 0.00678861f $X=42.375 $Y=1.4 $X2=0
+ $Y2=0
cc_4823 N_A_8379_265#_c_6082_n N_Z_c_9088_n 0.00239476f $X=42.085 $Y=1.4 $X2=0
+ $Y2=0
cc_4824 N_A_8379_265#_c_6088_n N_Z_c_9088_n 2.98555e-19 $X=42.465 $Y=1.4 $X2=0
+ $Y2=0
cc_4825 N_A_8379_265#_c_6084_n N_Z_c_9090_n 0.00145542f $X=42.845 $Y=1.4 $X2=0
+ $Y2=0
cc_4826 N_A_8379_265#_c_6086_n N_Z_c_9090_n 0.00597584f $X=43.315 $Y=1.4 $X2=0
+ $Y2=0
cc_4827 N_A_8379_265#_c_6089_n N_Z_c_9090_n 0.00909323f $X=42.935 $Y=1.4 $X2=0
+ $Y2=0
cc_4828 N_A_8379_265#_c_6073_n N_Z_c_9090_n 0.0266078f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4829 N_A_8379_265#_c_6079_n N_Z_c_9090_n 0.00747617f $X=43.725 $Y=1.23 $X2=0
+ $Y2=0
cc_4830 N_A_8379_265#_c_6080_n N_Z_c_9127_n 0.00834829f $X=41.995 $Y=1.475 $X2=0
+ $Y2=0
cc_4831 N_A_8379_265#_c_6087_n N_Z_c_9129_n 0.00795576f $X=43.405 $Y=1.475 $X2=0
+ $Y2=0
cc_4832 N_A_8379_265#_c_6073_n N_Z_c_9129_n 0.0186685f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4833 N_A_8379_265#_c_6092_n N_Z_c_9129_n 0.0329704f $X=44.685 $Y=1.77 $X2=0
+ $Y2=0
cc_4834 N_A_8379_265#_c_6079_n N_Z_c_9129_n 2.19754e-19 $X=43.725 $Y=1.23 $X2=0
+ $Y2=0
cc_4835 N_A_8379_265#_c_6083_n Z 0.00372458f $X=42.465 $Y=1.475 $X2=0 $Y2=0
cc_4836 N_A_8379_265#_c_6085_n Z 0.00372248f $X=42.935 $Y=1.475 $X2=0 $Y2=0
cc_4837 N_A_8379_265#_c_6080_n N_Z_c_9143_n 0.0199111f $X=41.995 $Y=1.475 $X2=0
+ $Y2=0
cc_4838 N_A_8379_265#_c_6081_n N_Z_c_9143_n 0.00560592f $X=42.375 $Y=1.4 $X2=0
+ $Y2=0
cc_4839 N_A_8379_265#_c_6082_n N_Z_c_9143_n 0.00474497f $X=42.085 $Y=1.4 $X2=0
+ $Y2=0
cc_4840 N_A_8379_265#_c_6083_n N_Z_c_9143_n 0.0181262f $X=42.465 $Y=1.475 $X2=0
+ $Y2=0
cc_4841 N_A_8379_265#_c_6085_n N_Z_c_9143_n 9.74366e-19 $X=42.935 $Y=1.475 $X2=0
+ $Y2=0
cc_4842 N_A_8379_265#_c_6088_n N_Z_c_9143_n 0.00415268f $X=42.465 $Y=1.4 $X2=0
+ $Y2=0
cc_4843 N_A_8379_265#_c_6083_n N_Z_c_9144_n 9.74366e-19 $X=42.465 $Y=1.475 $X2=0
+ $Y2=0
cc_4844 N_A_8379_265#_c_6085_n N_Z_c_9144_n 0.0181262f $X=42.935 $Y=1.475 $X2=0
+ $Y2=0
cc_4845 N_A_8379_265#_c_6086_n N_Z_c_9144_n 0.00560592f $X=43.315 $Y=1.4 $X2=0
+ $Y2=0
cc_4846 N_A_8379_265#_c_6087_n N_Z_c_9144_n 0.0221748f $X=43.405 $Y=1.475 $X2=0
+ $Y2=0
cc_4847 N_A_8379_265#_c_6089_n N_Z_c_9144_n 0.00181273f $X=42.935 $Y=1.4 $X2=0
+ $Y2=0
cc_4848 N_A_8379_265#_c_6073_n N_Z_c_9144_n 0.00240108f $X=44.52 $Y=1.23 $X2=0
+ $Y2=0
cc_4849 N_A_8379_265#_c_6079_n N_Z_c_9144_n 0.00425035f $X=43.725 $Y=1.23 $X2=0
+ $Y2=0
cc_4850 N_A_8379_265#_c_6080_n N_A_7937_297#_c_12195_n 0.00151141f $X=41.995
+ $Y=1.475 $X2=0 $Y2=0
cc_4851 N_A_8379_265#_c_6080_n N_A_7937_297#_c_12224_n 0.00307958f $X=41.995
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_4852 N_A_8379_265#_c_6083_n N_A_7937_297#_c_12224_n 0.00307958f $X=42.465
+ $Y=1.475 $X2=25.99 $Y2=0.51
cc_4853 N_A_8379_265#_c_6085_n N_A_7937_297#_c_12226_n 0.00307958f $X=42.935
+ $Y=1.475 $X2=0 $Y2=0
cc_4854 N_A_8379_265#_c_6087_n N_A_7937_297#_c_12226_n 0.00307958f $X=43.405
+ $Y=1.475 $X2=0 $Y2=0
cc_4855 N_A_8379_265#_c_6080_n N_A_7937_297#_c_12197_n 0.00554566f $X=41.995
+ $Y=1.475 $X2=0 $Y2=0
cc_4856 N_A_8379_265#_c_6083_n N_A_7937_297#_c_12198_n 0.00210632f $X=42.465
+ $Y=1.475 $X2=0 $Y2=0
cc_4857 N_A_8379_265#_c_6084_n N_A_7937_297#_c_12198_n 0.00251792f $X=42.845
+ $Y=1.4 $X2=0 $Y2=0
cc_4858 N_A_8379_265#_c_6085_n N_A_7937_297#_c_12198_n 0.00210632f $X=42.935
+ $Y=1.475 $X2=0 $Y2=0
cc_4859 N_A_8379_265#_c_6087_n N_A_7937_297#_c_12199_n 0.00499839f $X=43.405
+ $Y=1.475 $X2=0 $Y2=0
cc_4860 N_A_8379_265#_c_6073_n N_A_7937_297#_c_12199_n 0.0218124f $X=44.52
+ $Y=1.23 $X2=0 $Y2=0
cc_4861 N_A_8379_265#_c_6074_n N_A_7937_297#_c_12199_n 5.74251e-19 $X=43.975
+ $Y=1.23 $X2=0 $Y2=0
cc_4862 N_A_8379_265#_c_6079_n N_A_7937_297#_c_12199_n 0.00561627f $X=43.725
+ $Y=1.23 $X2=0 $Y2=0
cc_4863 N_A_8379_265#_c_6073_n N_VGND_c_12771_n 0.0123065f $X=44.52 $Y=1.23
+ $X2=0 $Y2=0
cc_4864 N_A_8379_265#_c_6074_n N_VGND_c_12771_n 2.04129e-19 $X=43.975 $Y=1.23
+ $X2=0 $Y2=0
cc_4865 N_A_8379_265#_c_6075_n N_VGND_c_12851_n 0.0129994f $X=44.685 $Y=0.445
+ $X2=0 $Y2=0
cc_4866 N_A_8379_265#_M1009_d VGND 0.00394793f $X=44.55 $Y=0.235 $X2=0 $Y2=0
cc_4867 N_A_8379_265#_c_6075_n VGND 0.00927134f $X=44.685 $Y=0.445 $X2=0 $Y2=0
cc_4868 N_A_8379_265#_c_6088_n N_A_7939_47#_c_15061_n 7.0477e-19 $X=42.465
+ $Y=1.4 $X2=0 $Y2=0
cc_4869 N_A_8379_265#_c_6073_n N_A_7939_47#_c_15039_n 0.0028695f $X=44.52
+ $Y=1.23 $X2=25.99 $Y2=4.93
cc_4870 N_A_8379_265#_c_6079_n N_A_7939_47#_c_15039_n 0.00589316f $X=43.725
+ $Y=1.23 $X2=25.99 $Y2=4.93
cc_4871 N_A_8379_793#_c_6201_n N_S[14]_c_6434_n 0.00507426f $X=42.085 $Y=4.04
+ $X2=0 $Y2=0
cc_4872 N_A_8379_793#_c_6200_n N_S[14]_c_6437_n 0.00509391f $X=42.375 $Y=4.04
+ $X2=0 $Y2=0
cc_4873 N_A_8379_793#_c_6203_n N_S[14]_c_6439_n 0.00509204f $X=42.845 $Y=4.04
+ $X2=25.905 $Y2=4.845
cc_4874 N_A_8379_793#_c_6205_n N_S[14]_c_6441_n 0.00507688f $X=43.315 $Y=4.04
+ $X2=0 $Y2=0
cc_4875 N_A_8379_793#_c_6194_n N_S[14]_c_6443_n 6.53442e-19 $X=44.645 $Y=4.74
+ $X2=0 $Y2=0
cc_4876 N_A_8379_793#_c_6192_n N_S[14]_c_6445_n 0.0103812f $X=44.52 $Y=4.21
+ $X2=0 $Y2=0
cc_4877 N_A_8379_793#_c_6193_n N_S[14]_c_6445_n 0.0179529f $X=43.975 $Y=4.21
+ $X2=0 $Y2=0
cc_4878 N_A_8379_793#_c_6212_n N_S[14]_c_6455_n 0.00508008f $X=44.605 $Y=4.045
+ $X2=0 $Y2=0
cc_4879 N_A_8379_793#_c_6198_n N_S[14]_c_6455_n 0.00262132f $X=43.725 $Y=4.21
+ $X2=0 $Y2=0
cc_4880 N_A_8379_793#_c_6192_n N_S[14]_c_6446_n 0.0206368f $X=44.52 $Y=4.21
+ $X2=0 $Y2=0
cc_4881 N_A_8379_793#_c_6193_n N_S[14]_c_6446_n 0.0175393f $X=43.975 $Y=4.21
+ $X2=0 $Y2=0
cc_4882 N_A_8379_793#_c_6212_n N_S[14]_c_6446_n 0.00255921f $X=44.605 $Y=4.045
+ $X2=0 $Y2=0
cc_4883 N_A_8379_793#_c_6196_n N_S[14]_c_6446_n 0.00322131f $X=44.605 $Y=4.21
+ $X2=0 $Y2=0
cc_4884 N_A_8379_793#_c_6197_n N_S[14]_c_6446_n 0.0085951f $X=44.645 $Y=4.615
+ $X2=0 $Y2=0
cc_4885 N_A_8379_793#_c_6211_n N_S[14]_c_6457_n 0.00970559f $X=44.685 $Y=3.14
+ $X2=0 $Y2=0
cc_4886 N_A_8379_793#_c_6212_n N_S[14]_c_6457_n 0.00254107f $X=44.605 $Y=4.045
+ $X2=0 $Y2=0
cc_4887 N_A_8379_793#_c_6213_n N_S[14]_c_6457_n 0.00216424f $X=44.685 $Y=3.835
+ $X2=0 $Y2=0
cc_4888 N_A_8379_793#_c_6194_n N_S[14]_c_6447_n 9.67113e-19 $X=44.645 $Y=4.74
+ $X2=0 $Y2=0
cc_4889 N_A_8379_793#_c_6195_n N_S[14]_c_6447_n 0.00603996f $X=44.685 $Y=4.995
+ $X2=0 $Y2=0
cc_4890 N_A_8379_793#_c_6194_n N_S[14]_c_6448_n 0.0111895f $X=44.645 $Y=4.74
+ $X2=0 $Y2=0
cc_4891 N_A_8379_793#_c_6197_n N_S[14]_c_6448_n 0.00429801f $X=44.645 $Y=4.615
+ $X2=0 $Y2=0
cc_4892 N_A_8379_793#_c_6212_n N_S[14]_c_6449_n 0.00336772f $X=44.605 $Y=4.045
+ $X2=0 $Y2=0
cc_4893 N_A_8379_793#_c_6194_n N_S[14]_c_6449_n 0.00207203f $X=44.645 $Y=4.74
+ $X2=0 $Y2=0
cc_4894 N_A_8379_793#_c_6213_n N_S[14]_c_6449_n 5.48523e-19 $X=44.685 $Y=3.835
+ $X2=0 $Y2=0
cc_4895 N_A_8379_793#_c_6196_n N_S[14]_c_6449_n 0.00416423f $X=44.605 $Y=4.21
+ $X2=0 $Y2=0
cc_4896 N_A_8379_793#_c_6197_n N_S[14]_c_6449_n 0.00289358f $X=44.645 $Y=4.615
+ $X2=0 $Y2=0
cc_4897 N_A_8379_793#_c_6211_n N_S[14]_c_6459_n 0.00929139f $X=44.685 $Y=3.14
+ $X2=25.99 $Y2=4.8
cc_4898 N_A_8379_793#_c_6212_n N_S[14]_c_6459_n 0.00117303f $X=44.605 $Y=4.045
+ $X2=25.99 $Y2=4.8
cc_4899 N_A_8379_793#_c_6213_n N_S[14]_c_6459_n 0.00304348f $X=44.685 $Y=3.835
+ $X2=25.99 $Y2=4.8
cc_4900 N_A_8379_793#_c_6194_n N_S[14]_c_6453_n 0.00426435f $X=44.645 $Y=4.74
+ $X2=0 $Y2=0
cc_4901 N_A_8379_793#_c_6197_n N_S[14]_c_6453_n 0.00268644f $X=44.645 $Y=4.615
+ $X2=0 $Y2=0
cc_4902 N_A_8379_793#_c_6196_n S[14] 0.0228692f $X=44.605 $Y=4.21 $X2=0 $Y2=0
cc_4903 N_A_8379_793#_c_6197_n S[14] 0.00541767f $X=44.645 $Y=4.615 $X2=0 $Y2=0
cc_4904 N_A_8379_793#_c_6199_n N_VPWR_c_7295_n 0.00324472f $X=41.995 $Y=3.965
+ $X2=0 $Y2=0
cc_4905 N_A_8379_793#_c_6206_n N_VPWR_c_7297_n 0.00367058f $X=43.405 $Y=3.965
+ $X2=0 $Y2=0
cc_4906 N_A_8379_793#_c_6192_n N_VPWR_c_7297_n 0.0193185f $X=44.52 $Y=4.21 $X2=0
+ $Y2=0
cc_4907 N_A_8379_793#_c_6193_n N_VPWR_c_7297_n 6.4101e-19 $X=43.975 $Y=4.21
+ $X2=0 $Y2=0
cc_4908 N_A_8379_793#_c_6211_n N_VPWR_c_7297_n 0.0316788f $X=44.685 $Y=3.14
+ $X2=0 $Y2=0
cc_4909 N_A_8379_793#_c_6211_n N_VPWR_c_7299_n 0.0356181f $X=44.685 $Y=3.14
+ $X2=0 $Y2=0
cc_4910 N_A_8379_793#_c_6211_n N_VPWR_c_7340_n 0.0233824f $X=44.685 $Y=3.14
+ $X2=0 $Y2=0
cc_4911 N_A_8379_793#_c_6199_n VPWR 0.00473731f $X=41.995 $Y=3.965 $X2=0 $Y2=0
cc_4912 N_A_8379_793#_c_6202_n VPWR 0.00362156f $X=42.465 $Y=3.965 $X2=0 $Y2=0
cc_4913 N_A_8379_793#_c_6204_n VPWR 0.00362156f $X=42.935 $Y=3.965 $X2=0 $Y2=0
cc_4914 N_A_8379_793#_c_6206_n VPWR 0.00473731f $X=43.405 $Y=3.965 $X2=0 $Y2=0
cc_4915 N_A_8379_793#_c_6211_n VPWR 0.00593513f $X=44.685 $Y=3.14 $X2=0 $Y2=0
cc_4916 N_A_8379_793#_c_6203_n N_Z_c_9035_n 0.00762343f $X=42.845 $Y=4.04 $X2=0
+ $Y2=0
cc_4917 N_A_8379_793#_c_6207_n N_Z_c_9035_n 0.00704092f $X=42.465 $Y=4.04 $X2=0
+ $Y2=0
cc_4918 N_A_8379_793#_c_6201_n N_Z_c_9086_n 0.00248496f $X=42.085 $Y=4.04 $X2=0
+ $Y2=0
cc_4919 N_A_8379_793#_c_6200_n N_Z_c_9089_n 0.00678861f $X=42.375 $Y=4.04 $X2=0
+ $Y2=0
cc_4920 N_A_8379_793#_c_6201_n N_Z_c_9089_n 0.00239476f $X=42.085 $Y=4.04 $X2=0
+ $Y2=0
cc_4921 N_A_8379_793#_c_6207_n N_Z_c_9089_n 2.98555e-19 $X=42.465 $Y=4.04 $X2=0
+ $Y2=0
cc_4922 N_A_8379_793#_c_6203_n N_Z_c_9091_n 0.00145542f $X=42.845 $Y=4.04 $X2=0
+ $Y2=0
cc_4923 N_A_8379_793#_c_6205_n N_Z_c_9091_n 0.00597584f $X=43.315 $Y=4.04 $X2=0
+ $Y2=0
cc_4924 N_A_8379_793#_c_6208_n N_Z_c_9091_n 0.00909323f $X=42.935 $Y=4.04 $X2=0
+ $Y2=0
cc_4925 N_A_8379_793#_c_6192_n N_Z_c_9091_n 0.0266078f $X=44.52 $Y=4.21 $X2=0
+ $Y2=0
cc_4926 N_A_8379_793#_c_6198_n N_Z_c_9091_n 0.00747617f $X=43.725 $Y=4.21 $X2=0
+ $Y2=0
cc_4927 N_A_8379_793#_c_6199_n N_Z_c_9128_n 0.00834829f $X=41.995 $Y=3.965 $X2=0
+ $Y2=0
cc_4928 N_A_8379_793#_c_6206_n N_Z_c_9130_n 0.00795576f $X=43.405 $Y=3.965 $X2=0
+ $Y2=0
cc_4929 N_A_8379_793#_c_6192_n N_Z_c_9130_n 0.0186685f $X=44.52 $Y=4.21 $X2=0
+ $Y2=0
cc_4930 N_A_8379_793#_c_6211_n N_Z_c_9130_n 0.0329704f $X=44.685 $Y=3.14 $X2=0
+ $Y2=0
cc_4931 N_A_8379_793#_c_6198_n N_Z_c_9130_n 2.19754e-19 $X=43.725 $Y=4.21 $X2=0
+ $Y2=0
cc_4932 N_A_8379_793#_c_6202_n Z 0.00372458f $X=42.465 $Y=3.965 $X2=0 $Y2=0
cc_4933 N_A_8379_793#_c_6204_n Z 0.00372248f $X=42.935 $Y=3.965 $X2=0 $Y2=0
cc_4934 N_A_8379_793#_c_6199_n N_Z_c_9143_n 0.0199111f $X=41.995 $Y=3.965 $X2=0
+ $Y2=0
cc_4935 N_A_8379_793#_c_6200_n N_Z_c_9143_n 0.00560592f $X=42.375 $Y=4.04 $X2=0
+ $Y2=0
cc_4936 N_A_8379_793#_c_6201_n N_Z_c_9143_n 0.00474497f $X=42.085 $Y=4.04 $X2=0
+ $Y2=0
cc_4937 N_A_8379_793#_c_6202_n N_Z_c_9143_n 0.0181262f $X=42.465 $Y=3.965 $X2=0
+ $Y2=0
cc_4938 N_A_8379_793#_c_6204_n N_Z_c_9143_n 9.74366e-19 $X=42.935 $Y=3.965 $X2=0
+ $Y2=0
cc_4939 N_A_8379_793#_c_6207_n N_Z_c_9143_n 0.00415268f $X=42.465 $Y=4.04 $X2=0
+ $Y2=0
cc_4940 N_A_8379_793#_c_6202_n N_Z_c_9144_n 9.74366e-19 $X=42.465 $Y=3.965 $X2=0
+ $Y2=0
cc_4941 N_A_8379_793#_c_6204_n N_Z_c_9144_n 0.0181262f $X=42.935 $Y=3.965 $X2=0
+ $Y2=0
cc_4942 N_A_8379_793#_c_6205_n N_Z_c_9144_n 0.00560592f $X=43.315 $Y=4.04 $X2=0
+ $Y2=0
cc_4943 N_A_8379_793#_c_6206_n N_Z_c_9144_n 0.0221748f $X=43.405 $Y=3.965 $X2=0
+ $Y2=0
cc_4944 N_A_8379_793#_c_6208_n N_Z_c_9144_n 0.00181273f $X=42.935 $Y=4.04 $X2=0
+ $Y2=0
cc_4945 N_A_8379_793#_c_6192_n N_Z_c_9144_n 0.00240108f $X=44.52 $Y=4.21 $X2=0
+ $Y2=0
cc_4946 N_A_8379_793#_c_6198_n N_Z_c_9144_n 0.00425035f $X=43.725 $Y=4.21 $X2=0
+ $Y2=0
cc_4947 N_A_8379_793#_c_6199_n N_A_7937_591#_c_12323_n 0.00151141f $X=41.995
+ $Y=3.965 $X2=0 $Y2=0
cc_4948 N_A_8379_793#_c_6199_n N_A_7937_591#_c_12352_n 0.00307958f $X=41.995
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_4949 N_A_8379_793#_c_6202_n N_A_7937_591#_c_12352_n 0.00307958f $X=42.465
+ $Y=3.965 $X2=25.99 $Y2=0.51
cc_4950 N_A_8379_793#_c_6204_n N_A_7937_591#_c_12354_n 0.00307958f $X=42.935
+ $Y=3.965 $X2=0 $Y2=0
cc_4951 N_A_8379_793#_c_6206_n N_A_7937_591#_c_12354_n 0.00307958f $X=43.405
+ $Y=3.965 $X2=0 $Y2=0
cc_4952 N_A_8379_793#_c_6199_n N_A_7937_591#_c_12325_n 0.00554566f $X=41.995
+ $Y=3.965 $X2=0 $Y2=0
cc_4953 N_A_8379_793#_c_6202_n N_A_7937_591#_c_12326_n 0.00210632f $X=42.465
+ $Y=3.965 $X2=0 $Y2=0
cc_4954 N_A_8379_793#_c_6203_n N_A_7937_591#_c_12326_n 0.00251792f $X=42.845
+ $Y=4.04 $X2=0 $Y2=0
cc_4955 N_A_8379_793#_c_6204_n N_A_7937_591#_c_12326_n 0.00210632f $X=42.935
+ $Y=3.965 $X2=0 $Y2=0
cc_4956 N_A_8379_793#_c_6206_n N_A_7937_591#_c_12327_n 0.00499839f $X=43.405
+ $Y=3.965 $X2=0 $Y2=0
cc_4957 N_A_8379_793#_c_6192_n N_A_7937_591#_c_12327_n 0.0218124f $X=44.52
+ $Y=4.21 $X2=0 $Y2=0
cc_4958 N_A_8379_793#_c_6193_n N_A_7937_591#_c_12327_n 5.74251e-19 $X=43.975
+ $Y=4.21 $X2=0 $Y2=0
cc_4959 N_A_8379_793#_c_6198_n N_A_7937_591#_c_12327_n 0.00561627f $X=43.725
+ $Y=4.21 $X2=0 $Y2=0
cc_4960 N_A_8379_793#_c_6192_n N_VGND_c_12772_n 0.0123065f $X=44.52 $Y=4.21
+ $X2=0 $Y2=0
cc_4961 N_A_8379_793#_c_6193_n N_VGND_c_12772_n 2.04129e-19 $X=43.975 $Y=4.21
+ $X2=0 $Y2=0
cc_4962 N_A_8379_793#_c_6195_n N_VGND_c_12853_n 0.0129994f $X=44.685 $Y=4.995
+ $X2=0 $Y2=0
cc_4963 N_A_8379_793#_M1028_d VGND 0.00394793f $X=44.55 $Y=4.785 $X2=0 $Y2=0
cc_4964 N_A_8379_793#_c_6195_n VGND 0.00927134f $X=44.685 $Y=4.995 $X2=0 $Y2=0
cc_4965 N_A_8379_793#_c_6207_n N_A_7939_911#_c_15140_n 7.0477e-19 $X=42.465
+ $Y=4.04 $X2=0 $Y2=0
cc_4966 N_A_8379_793#_c_6192_n N_A_7939_911#_c_15121_n 0.0028695f $X=44.52
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_4967 N_A_8379_793#_c_6198_n N_A_7939_911#_c_15121_n 0.00589316f $X=43.725
+ $Y=4.21 $X2=25.99 $Y2=4.8
cc_4968 N_S[6]_c_6340_n N_S[14]_c_6457_n 0.0130744f $X=44.45 $Y=1.55 $X2=0 $Y2=0
cc_4969 N_S[6]_c_6333_n N_S[14]_c_6459_n 0.0130744f $X=44.92 $Y=1.55 $X2=25.99
+ $Y2=4.8
cc_4970 N_S[6]_c_6333_n N_S[7]_c_6559_n 0.0215827f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4971 S[6] N_S[7]_c_6559_n 0.00113563f $X=45.225 $Y=1.105 $X2=0 $Y2=0
cc_4972 N_S[6]_c_6333_n N_S[7]_c_6580_n 0.00113563f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4973 S[6] N_S[7]_c_6580_n 0.0301108f $X=45.225 $Y=1.105 $X2=0 $Y2=0
cc_4974 N_S[6]_c_6340_n N_VPWR_c_7296_n 0.00950399f $X=44.45 $Y=1.55 $X2=0 $Y2=0
cc_4975 N_S[6]_c_6333_n N_VPWR_c_7298_n 0.016386f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4976 S[6] N_VPWR_c_7298_n 0.0157609f $X=45.225 $Y=1.105 $X2=0 $Y2=0
cc_4977 N_S[6]_c_6340_n N_VPWR_c_7340_n 0.0035837f $X=44.45 $Y=1.55 $X2=0 $Y2=0
cc_4978 N_S[6]_c_6333_n N_VPWR_c_7340_n 0.0035837f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4979 N_S[6]_c_6340_n VPWR 0.00711603f $X=44.45 $Y=1.55 $X2=0 $Y2=0
cc_4980 N_S[6]_c_6333_n VPWR 0.0070533f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4981 N_S[6]_c_6317_n N_Z_c_9033_n 0.002324f $X=41.92 $Y=0.255 $X2=0 $Y2=0
cc_4982 N_S[6]_c_6320_n N_Z_c_9033_n 0.00283489f $X=42.34 $Y=0.255 $X2=0 $Y2=0
cc_4983 N_S[6]_c_6320_n N_Z_c_9034_n 3.10191e-19 $X=42.34 $Y=0.255 $X2=0 $Y2=0
cc_4984 N_S[6]_c_6322_n N_Z_c_9034_n 0.00190704f $X=42.76 $Y=0.255 $X2=0 $Y2=0
cc_4985 N_S[6]_c_6320_n N_Z_c_9036_n 6.35774e-19 $X=42.34 $Y=0.255 $X2=0 $Y2=0
cc_4986 N_S[6]_c_6322_n N_Z_c_9036_n 0.0077801f $X=42.76 $Y=0.255 $X2=0 $Y2=0
cc_4987 N_S[6]_c_6324_n N_Z_c_9036_n 0.0134253f $X=43.18 $Y=0.255 $X2=0 $Y2=0
cc_4988 N_S[6]_c_6317_n N_Z_c_9085_n 0.00443615f $X=41.92 $Y=0.255 $X2=0 $Y2=0
cc_4989 N_S[6]_c_6320_n N_Z_c_9085_n 0.00462308f $X=42.34 $Y=0.255 $X2=0 $Y2=0
cc_4990 N_S[6]_c_6322_n N_Z_c_9085_n 6.35664e-19 $X=42.76 $Y=0.255 $X2=0 $Y2=0
cc_4991 N_S[6]_c_6320_n N_Z_c_9088_n 0.00180363f $X=42.34 $Y=0.255 $X2=0 $Y2=0
cc_4992 N_S[6]_c_6324_n N_Z_c_9090_n 0.00216436f $X=43.18 $Y=0.255 $X2=0 $Y2=0
cc_4993 N_S[6]_c_6340_n N_Z_c_9129_n 0.00478771f $X=44.45 $Y=1.55 $X2=0 $Y2=0
cc_4994 N_S[6]_c_6333_n N_Z_c_9129_n 0.00760321f $X=44.92 $Y=1.55 $X2=0 $Y2=0
cc_4995 S[6] N_Z_c_9129_n 0.010609f $X=45.225 $Y=1.105 $X2=0 $Y2=0
cc_4996 N_S[6]_c_6317_n N_A_7937_297#_c_12195_n 0.00168571f $X=41.92 $Y=0.255
+ $X2=0 $Y2=0
cc_4997 N_S[6]_c_6340_n N_A_7937_297#_c_12199_n 0.00239129f $X=44.45 $Y=1.55
+ $X2=0 $Y2=0
cc_4998 N_S[6]_c_6317_n N_VGND_c_12769_n 5.5039e-19 $X=41.92 $Y=0.255 $X2=0
+ $Y2=0
cc_4999 N_S[6]_c_6319_n N_VGND_c_12769_n 0.0028166f $X=41.995 $Y=0.18 $X2=0
+ $Y2=0
cc_5000 N_S[6]_c_6325_n N_VGND_c_12771_n 0.00862298f $X=43.865 $Y=0.18 $X2=0
+ $Y2=0
cc_5001 N_S[6]_c_6327_n N_VGND_c_12771_n 0.00525833f $X=44.35 $Y=0.81 $X2=0
+ $Y2=0
cc_5002 N_S[6]_c_6330_n N_VGND_c_12771_n 0.00173127f $X=44.475 $Y=0.735 $X2=0
+ $Y2=0
cc_5003 N_S[6]_c_6332_n N_VGND_c_12773_n 0.00374526f $X=44.895 $Y=0.735 $X2=0
+ $Y2=0
cc_5004 N_S[6]_c_6333_n N_VGND_c_12773_n 0.00578076f $X=44.92 $Y=1.55 $X2=0
+ $Y2=0
cc_5005 S[6] N_VGND_c_12773_n 0.0116413f $X=45.225 $Y=1.105 $X2=0 $Y2=0
cc_5006 N_S[6]_c_6319_n N_VGND_c_12847_n 0.0559651f $X=41.995 $Y=0.18 $X2=0
+ $Y2=0
cc_5007 N_S[6]_c_6330_n N_VGND_c_12851_n 0.00542362f $X=44.475 $Y=0.735 $X2=0
+ $Y2=0
cc_5008 N_S[6]_c_6331_n N_VGND_c_12851_n 2.16067e-19 $X=44.82 $Y=0.81 $X2=0
+ $Y2=0
cc_5009 N_S[6]_c_6332_n N_VGND_c_12851_n 0.00585385f $X=44.895 $Y=0.735 $X2=0
+ $Y2=0
cc_5010 N_S[6]_c_6318_n VGND 0.00642387f $X=42.265 $Y=0.18 $X2=0 $Y2=0
cc_5011 N_S[6]_c_6319_n VGND 0.00591981f $X=41.995 $Y=0.18 $X2=0 $Y2=0
cc_5012 N_S[6]_c_6321_n VGND 0.0064237f $X=42.685 $Y=0.18 $X2=0 $Y2=0
cc_5013 N_S[6]_c_6323_n VGND 0.00642387f $X=43.105 $Y=0.18 $X2=0 $Y2=0
cc_5014 N_S[6]_c_6325_n VGND 0.0345801f $X=43.865 $Y=0.18 $X2=0 $Y2=0
cc_5015 N_S[6]_c_6330_n VGND 0.00990284f $X=44.475 $Y=0.735 $X2=0 $Y2=0
cc_5016 N_S[6]_c_6332_n VGND 0.0119653f $X=44.895 $Y=0.735 $X2=0 $Y2=0
cc_5017 N_S[6]_c_6334_n VGND 0.00366655f $X=42.34 $Y=0.18 $X2=0 $Y2=0
cc_5018 N_S[6]_c_6335_n VGND 0.00366655f $X=42.76 $Y=0.18 $X2=0 $Y2=0
cc_5019 N_S[6]_c_6336_n VGND 0.00366655f $X=43.18 $Y=0.18 $X2=0 $Y2=0
cc_5020 N_S[6]_c_6317_n N_A_7939_47#_c_15034_n 0.00206084f $X=41.92 $Y=0.255
+ $X2=0 $Y2=0
cc_5021 N_S[6]_c_6317_n N_A_7939_47#_c_15036_n 0.0139014f $X=41.92 $Y=0.255
+ $X2=0 $Y2=0
cc_5022 N_S[6]_c_6318_n N_A_7939_47#_c_15036_n 0.00211351f $X=42.265 $Y=0.18
+ $X2=0 $Y2=0
cc_5023 N_S[6]_c_6320_n N_A_7939_47#_c_15036_n 0.0106826f $X=42.34 $Y=0.255
+ $X2=0 $Y2=0
cc_5024 N_S[6]_c_6322_n N_A_7939_47#_c_15038_n 0.0106844f $X=42.76 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_5025 N_S[6]_c_6323_n N_A_7939_47#_c_15038_n 0.00211351f $X=43.105 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_5026 N_S[6]_c_6324_n N_A_7939_47#_c_15038_n 0.0112916f $X=43.18 $Y=0.255
+ $X2=25.99 $Y2=4.8
cc_5027 N_S[6]_c_6325_n N_A_7939_47#_c_15038_n 0.00685838f $X=43.865 $Y=0.18
+ $X2=25.99 $Y2=4.8
cc_5028 N_S[6]_c_6326_n N_A_7939_47#_c_15038_n 0.00189496f $X=43.94 $Y=0.735
+ $X2=25.99 $Y2=4.8
cc_5029 N_S[6]_c_6326_n N_A_7939_47#_c_15039_n 0.00529837f $X=43.94 $Y=0.735
+ $X2=25.99 $Y2=4.93
cc_5030 N_S[6]_c_6321_n N_A_7939_47#_c_15074_n 0.0034777f $X=42.685 $Y=0.18
+ $X2=0 $Y2=0
cc_5031 N_S[14]_c_6449_n N_S[15]_c_6679_n 0.0215827f $X=44.895 $Y=4.705 $X2=0
+ $Y2=0
cc_5032 S[14] N_S[15]_c_6679_n 0.00113563f $X=45.225 $Y=4.165 $X2=0 $Y2=0
cc_5033 N_S[14]_c_6449_n N_S[15]_c_6699_n 0.00113563f $X=44.895 $Y=4.705 $X2=0
+ $Y2=0
cc_5034 S[14] N_S[15]_c_6699_n 0.0301108f $X=45.225 $Y=4.165 $X2=0 $Y2=0
cc_5035 N_S[14]_c_6457_n N_VPWR_c_7297_n 0.00950399f $X=44.45 $Y=3.89 $X2=0
+ $Y2=0
cc_5036 N_S[14]_c_6449_n N_VPWR_c_7299_n 0.00652399f $X=44.895 $Y=4.705 $X2=0
+ $Y2=0
cc_5037 N_S[14]_c_6459_n N_VPWR_c_7299_n 0.00986205f $X=44.92 $Y=3.89 $X2=0
+ $Y2=0
cc_5038 S[14] N_VPWR_c_7299_n 0.0157609f $X=45.225 $Y=4.165 $X2=0 $Y2=0
cc_5039 N_S[14]_c_6457_n N_VPWR_c_7340_n 0.0035837f $X=44.45 $Y=3.89 $X2=0 $Y2=0
cc_5040 N_S[14]_c_6459_n N_VPWR_c_7340_n 0.0035837f $X=44.92 $Y=3.89 $X2=0 $Y2=0
cc_5041 N_S[14]_c_6457_n VPWR 0.00711603f $X=44.45 $Y=3.89 $X2=0 $Y2=0
cc_5042 N_S[14]_c_6459_n VPWR 0.0070533f $X=44.92 $Y=3.89 $X2=0 $Y2=0
cc_5043 N_S[14]_c_6437_n N_Z_c_9035_n 3.10191e-19 $X=42.34 $Y=5.185 $X2=0 $Y2=0
cc_5044 N_S[14]_c_6439_n N_Z_c_9035_n 0.00190704f $X=42.76 $Y=5.185 $X2=0 $Y2=0
cc_5045 N_S[14]_c_6437_n N_Z_c_9037_n 6.35774e-19 $X=42.34 $Y=5.185 $X2=0 $Y2=0
cc_5046 N_S[14]_c_6439_n N_Z_c_9037_n 0.0077801f $X=42.76 $Y=5.185 $X2=0 $Y2=0
cc_5047 N_S[14]_c_6441_n N_Z_c_9037_n 0.0134253f $X=43.18 $Y=5.185 $X2=0 $Y2=0
cc_5048 N_S[14]_c_6434_n N_Z_c_9086_n 0.00443615f $X=41.92 $Y=5.185 $X2=0 $Y2=0
cc_5049 N_S[14]_c_6437_n N_Z_c_9086_n 0.00462308f $X=42.34 $Y=5.185 $X2=0 $Y2=0
cc_5050 N_S[14]_c_6434_n N_Z_c_9087_n 0.002324f $X=41.92 $Y=5.185 $X2=0 $Y2=0
cc_5051 N_S[14]_c_6437_n N_Z_c_9087_n 0.00283489f $X=42.34 $Y=5.185 $X2=0 $Y2=0
cc_5052 N_S[14]_c_6439_n N_Z_c_9087_n 6.35664e-19 $X=42.76 $Y=5.185 $X2=0 $Y2=0
cc_5053 N_S[14]_c_6437_n N_Z_c_9089_n 0.00180363f $X=42.34 $Y=5.185 $X2=0 $Y2=0
cc_5054 N_S[14]_c_6441_n N_Z_c_9091_n 0.00216436f $X=43.18 $Y=5.185 $X2=0 $Y2=0
cc_5055 N_S[14]_c_6455_n N_Z_c_9130_n 2.55735e-19 $X=44.45 $Y=3.99 $X2=0 $Y2=0
cc_5056 N_S[14]_c_6457_n N_Z_c_9130_n 0.00453198f $X=44.45 $Y=3.89 $X2=0 $Y2=0
cc_5057 N_S[14]_c_6449_n N_Z_c_9130_n 0.00258545f $X=44.895 $Y=4.705 $X2=0 $Y2=0
cc_5058 N_S[14]_c_6459_n N_Z_c_9130_n 0.00501777f $X=44.92 $Y=3.89 $X2=0 $Y2=0
cc_5059 S[14] N_Z_c_9130_n 0.010609f $X=45.225 $Y=4.165 $X2=0 $Y2=0
cc_5060 N_S[14]_c_6434_n N_A_7937_591#_c_12323_n 0.00168571f $X=41.92 $Y=5.185
+ $X2=0 $Y2=0
cc_5061 N_S[14]_c_6457_n N_A_7937_591#_c_12327_n 0.00239129f $X=44.45 $Y=3.89
+ $X2=0 $Y2=0
cc_5062 N_S[14]_c_6434_n N_VGND_c_12770_n 5.5039e-19 $X=41.92 $Y=5.185 $X2=0
+ $Y2=0
cc_5063 N_S[14]_c_6436_n N_VGND_c_12770_n 0.0028166f $X=41.995 $Y=5.26 $X2=0
+ $Y2=0
cc_5064 N_S[14]_c_6443_n N_VGND_c_12772_n 0.00862298f $X=43.94 $Y=5.185 $X2=0
+ $Y2=0
cc_5065 N_S[14]_c_6444_n N_VGND_c_12772_n 0.00525833f $X=44.35 $Y=4.63 $X2=0
+ $Y2=0
cc_5066 N_S[14]_c_6447_n N_VGND_c_12772_n 0.00173127f $X=44.475 $Y=4.705 $X2=0
+ $Y2=0
cc_5067 N_S[14]_c_6449_n N_VGND_c_12774_n 0.00952602f $X=44.895 $Y=4.705 $X2=0
+ $Y2=0
cc_5068 S[14] N_VGND_c_12774_n 0.0116413f $X=45.225 $Y=4.165 $X2=0 $Y2=0
cc_5069 N_S[14]_c_6436_n N_VGND_c_12849_n 0.0559651f $X=41.995 $Y=5.26 $X2=0
+ $Y2=0
cc_5070 N_S[14]_c_6447_n N_VGND_c_12853_n 0.00542362f $X=44.475 $Y=4.705 $X2=0
+ $Y2=0
cc_5071 N_S[14]_c_6448_n N_VGND_c_12853_n 2.16067e-19 $X=44.82 $Y=4.63 $X2=0
+ $Y2=0
cc_5072 N_S[14]_c_6449_n N_VGND_c_12853_n 0.00585385f $X=44.895 $Y=4.705 $X2=0
+ $Y2=0
cc_5073 N_S[14]_c_6435_n VGND 0.00642387f $X=42.265 $Y=5.26 $X2=0 $Y2=0
cc_5074 N_S[14]_c_6436_n VGND 0.00591981f $X=41.995 $Y=5.26 $X2=0 $Y2=0
cc_5075 N_S[14]_c_6438_n VGND 0.0064237f $X=42.685 $Y=5.26 $X2=0 $Y2=0
cc_5076 N_S[14]_c_6440_n VGND 0.00642387f $X=43.105 $Y=5.26 $X2=0 $Y2=0
cc_5077 N_S[14]_c_6442_n VGND 0.0345801f $X=43.865 $Y=5.26 $X2=0 $Y2=0
cc_5078 N_S[14]_c_6447_n VGND 0.00990284f $X=44.475 $Y=4.705 $X2=0 $Y2=0
cc_5079 N_S[14]_c_6449_n VGND 0.0119653f $X=44.895 $Y=4.705 $X2=0 $Y2=0
cc_5080 N_S[14]_c_6450_n VGND 0.00366655f $X=42.34 $Y=5.26 $X2=0 $Y2=0
cc_5081 N_S[14]_c_6451_n VGND 0.00366655f $X=42.76 $Y=5.26 $X2=0 $Y2=0
cc_5082 N_S[14]_c_6452_n VGND 0.00366655f $X=43.18 $Y=5.26 $X2=0 $Y2=0
cc_5083 N_S[14]_c_6434_n N_A_7939_911#_c_15116_n 0.00206084f $X=41.92 $Y=5.185
+ $X2=0 $Y2=0
cc_5084 N_S[14]_c_6434_n N_A_7939_911#_c_15118_n 0.0139014f $X=41.92 $Y=5.185
+ $X2=0 $Y2=0
cc_5085 N_S[14]_c_6435_n N_A_7939_911#_c_15118_n 0.00211351f $X=42.265 $Y=5.26
+ $X2=0 $Y2=0
cc_5086 N_S[14]_c_6437_n N_A_7939_911#_c_15118_n 0.0106826f $X=42.34 $Y=5.185
+ $X2=0 $Y2=0
cc_5087 N_S[14]_c_6439_n N_A_7939_911#_c_15120_n 0.0106844f $X=42.76 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_5088 N_S[14]_c_6440_n N_A_7939_911#_c_15120_n 0.00211351f $X=43.105 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_5089 N_S[14]_c_6441_n N_A_7939_911#_c_15120_n 0.0112916f $X=43.18 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_5090 N_S[14]_c_6442_n N_A_7939_911#_c_15120_n 0.00685838f $X=43.865 $Y=5.26
+ $X2=25.99 $Y2=0.64
cc_5091 N_S[14]_c_6443_n N_A_7939_911#_c_15120_n 0.00189496f $X=43.94 $Y=5.185
+ $X2=25.99 $Y2=0.64
cc_5092 N_S[14]_c_6445_n N_A_7939_911#_c_15121_n 0.00529837f $X=44.015 $Y=4.63
+ $X2=25.99 $Y2=4.8
cc_5093 N_S[14]_c_6438_n N_A_7939_911#_c_15153_n 0.0034777f $X=42.685 $Y=5.26
+ $X2=0 $Y2=0
cc_5094 N_S[7]_c_6560_n N_S[15]_c_6701_n 0.0130744f $X=46.16 $Y=1.55 $X2=0 $Y2=0
cc_5095 N_S[7]_c_6584_n N_S[15]_c_6705_n 0.0130744f $X=46.63 $Y=1.55 $X2=0 $Y2=0
cc_5096 N_S[7]_c_6569_n N_A_9250_325#_c_6815_n 0.00507688f $X=47.9 $Y=0.255
+ $X2=25.905 $Y2=0.425
cc_5097 N_S[7]_c_6564_n N_A_9250_325#_c_6807_n 0.00262132f $X=46.63 $Y=1.45
+ $X2=25.905 $Y2=4.845
cc_5098 N_S[7]_c_6571_n N_A_9250_325#_c_6818_n 0.00509204f $X=48.32 $Y=0.255
+ $X2=0 $Y2=0
cc_5099 N_S[7]_c_6575_n N_A_9250_325#_c_6820_n 0.00507426f $X=49.16 $Y=0.255
+ $X2=0 $Y2=0
cc_5100 N_S[7]_c_6573_n N_A_9250_325#_c_6823_n 0.00509391f $X=48.74 $Y=0.255
+ $X2=0 $Y2=0
cc_5101 N_S[7]_c_6560_n N_A_9250_325#_c_6824_n 0.0128834f $X=46.16 $Y=1.55 $X2=0
+ $Y2=0
cc_5102 N_S[7]_c_6584_n N_A_9250_325#_c_6824_n 0.0118698f $X=46.63 $Y=1.55 $X2=0
+ $Y2=0
cc_5103 N_S[7]_c_6561_n N_A_9250_325#_c_6808_n 0.00207203f $X=46.185 $Y=0.735
+ $X2=0 $Y2=0
cc_5104 N_S[7]_c_6563_n N_A_9250_325#_c_6808_n 0.00603996f $X=46.605 $Y=0.735
+ $X2=0 $Y2=0
cc_5105 N_S[7]_c_6566_n N_A_9250_325#_c_6808_n 6.53442e-19 $X=47.14 $Y=0.735
+ $X2=0 $Y2=0
cc_5106 N_S[7]_c_6560_n N_A_9250_325#_c_6809_n 0.00289358f $X=46.16 $Y=1.55
+ $X2=0 $Y2=0
cc_5107 N_S[7]_c_6562_n N_A_9250_325#_c_6809_n 0.00429801f $X=46.53 $Y=0.81
+ $X2=0 $Y2=0
cc_5108 N_S[7]_c_6564_n N_A_9250_325#_c_6809_n 0.0085951f $X=46.63 $Y=1.45 $X2=0
+ $Y2=0
cc_5109 N_S[7]_c_6576_n N_A_9250_325#_c_6809_n 0.00268644f $X=46.63 $Y=0.81
+ $X2=0 $Y2=0
cc_5110 N_S[7]_c_6580_n N_A_9250_325#_c_6809_n 0.00541767f $X=46.12 $Y=1.16
+ $X2=0 $Y2=0
cc_5111 N_S[7]_c_6564_n N_A_9250_325#_c_6810_n 0.0206368f $X=46.63 $Y=1.45 $X2=0
+ $Y2=0
cc_5112 N_S[7]_c_6565_n N_A_9250_325#_c_6810_n 0.0103812f $X=47.065 $Y=0.81
+ $X2=0 $Y2=0
cc_5113 N_S[7]_c_6560_n N_A_9250_325#_c_6826_n 0.00454075f $X=46.16 $Y=1.55
+ $X2=0 $Y2=0
cc_5114 N_S[7]_c_6564_n N_A_9250_325#_c_6826_n 0.00255921f $X=46.63 $Y=1.45
+ $X2=0 $Y2=0
cc_5115 N_S[7]_c_6584_n N_A_9250_325#_c_6826_n 0.00762115f $X=46.63 $Y=1.55
+ $X2=0 $Y2=0
cc_5116 N_S[7]_c_6562_n N_A_9250_325#_c_6811_n 0.0111895f $X=46.53 $Y=0.81 $X2=0
+ $Y2=0
cc_5117 N_S[7]_c_6563_n N_A_9250_325#_c_6811_n 9.67113e-19 $X=46.605 $Y=0.735
+ $X2=0 $Y2=0
cc_5118 N_S[7]_c_6576_n N_A_9250_325#_c_6811_n 0.00426435f $X=46.63 $Y=0.81
+ $X2=0 $Y2=0
cc_5119 N_S[7]_c_6560_n N_A_9250_325#_c_6812_n 0.00416423f $X=46.16 $Y=1.55
+ $X2=0 $Y2=0
cc_5120 N_S[7]_c_6564_n N_A_9250_325#_c_6812_n 0.00322131f $X=46.63 $Y=1.45
+ $X2=0 $Y2=0
cc_5121 N_S[7]_c_6580_n N_A_9250_325#_c_6812_n 0.0228692f $X=46.12 $Y=1.16 $X2=0
+ $Y2=0
cc_5122 N_S[7]_c_6564_n N_A_9250_325#_c_6813_n 0.0175393f $X=46.63 $Y=1.45 $X2=0
+ $Y2=0
cc_5123 N_S[7]_c_6565_n N_A_9250_325#_c_6813_n 0.0179529f $X=47.065 $Y=0.81
+ $X2=0 $Y2=0
cc_5124 N_S[7]_c_6559_n N_VPWR_c_7301_n 0.00652399f $X=46.06 $Y=1.16 $X2=0 $Y2=0
cc_5125 N_S[7]_c_6560_n N_VPWR_c_7301_n 0.00986205f $X=46.16 $Y=1.55 $X2=0 $Y2=0
cc_5126 N_S[7]_c_6580_n N_VPWR_c_7301_n 0.0157609f $X=46.12 $Y=1.16 $X2=0 $Y2=0
cc_5127 N_S[7]_c_6584_n N_VPWR_c_7303_n 0.00950399f $X=46.63 $Y=1.55 $X2=0 $Y2=0
cc_5128 N_S[7]_c_6560_n N_VPWR_c_7343_n 0.0035837f $X=46.16 $Y=1.55 $X2=0 $Y2=0
cc_5129 N_S[7]_c_6584_n N_VPWR_c_7343_n 0.0035837f $X=46.63 $Y=1.55 $X2=0 $Y2=0
cc_5130 N_S[7]_c_6560_n VPWR 0.0070533f $X=46.16 $Y=1.55 $X2=0 $Y2=0
cc_5131 N_S[7]_c_6584_n VPWR 0.00711603f $X=46.63 $Y=1.55 $X2=0 $Y2=0
cc_5132 N_S[7]_c_6569_n N_Z_c_9038_n 0.0134253f $X=47.9 $Y=0.255 $X2=0 $Y2=0
cc_5133 N_S[7]_c_6571_n N_Z_c_9038_n 0.0077801f $X=48.32 $Y=0.255 $X2=0 $Y2=0
cc_5134 N_S[7]_c_6573_n N_Z_c_9038_n 6.35774e-19 $X=48.74 $Y=0.255 $X2=0 $Y2=0
cc_5135 N_S[7]_c_6571_n N_Z_c_9040_n 0.00190704f $X=48.32 $Y=0.255 $X2=0 $Y2=0
cc_5136 N_S[7]_c_6573_n N_Z_c_9040_n 3.10191e-19 $X=48.74 $Y=0.255 $X2=0 $Y2=0
cc_5137 N_S[7]_c_6573_n N_Z_c_9042_n 0.00283489f $X=48.74 $Y=0.255 $X2=0 $Y2=0
cc_5138 N_S[7]_c_6575_n N_Z_c_9042_n 0.002324f $X=49.16 $Y=0.255 $X2=0 $Y2=0
cc_5139 N_S[7]_c_6569_n N_Z_c_9092_n 0.00216436f $X=47.9 $Y=0.255 $X2=0 $Y2=0
cc_5140 N_S[7]_c_6573_n N_Z_c_9094_n 0.00180363f $X=48.74 $Y=0.255 $X2=0 $Y2=0
cc_5141 N_S[7]_c_6571_n N_Z_c_9096_n 6.35664e-19 $X=48.32 $Y=0.255 $X2=0 $Y2=0
cc_5142 N_S[7]_c_6573_n N_Z_c_9096_n 0.00462308f $X=48.74 $Y=0.255 $X2=0 $Y2=0
cc_5143 N_S[7]_c_6575_n N_Z_c_9096_n 0.00443615f $X=49.16 $Y=0.255 $X2=0 $Y2=0
cc_5144 N_S[7]_c_6559_n N_Z_c_9129_n 0.00234109f $X=46.06 $Y=1.16 $X2=0 $Y2=0
cc_5145 N_S[7]_c_6560_n N_Z_c_9129_n 0.0052507f $X=46.16 $Y=1.55 $X2=0 $Y2=0
cc_5146 N_S[7]_c_6584_n N_Z_c_9129_n 0.00478771f $X=46.63 $Y=1.55 $X2=0 $Y2=0
cc_5147 N_S[7]_c_6580_n N_Z_c_9129_n 0.0105931f $X=46.12 $Y=1.16 $X2=0 $Y2=0
cc_5148 N_S[7]_c_6575_n N_A_9463_311#_c_12452_n 0.00168571f $X=49.16 $Y=0.255
+ $X2=0 $Y2=0
cc_5149 N_S[7]_c_6584_n N_A_9463_311#_c_12454_n 0.00239129f $X=46.63 $Y=1.55
+ $X2=0 $Y2=0
cc_5150 N_S[7]_c_6559_n N_VGND_c_12775_n 0.00576464f $X=46.06 $Y=1.16 $X2=0
+ $Y2=0
cc_5151 N_S[7]_c_6561_n N_VGND_c_12775_n 0.00374526f $X=46.185 $Y=0.735 $X2=0
+ $Y2=0
cc_5152 N_S[7]_c_6580_n N_VGND_c_12775_n 0.0116218f $X=46.12 $Y=1.16 $X2=0 $Y2=0
cc_5153 N_S[7]_c_6563_n N_VGND_c_12777_n 0.00173127f $X=46.605 $Y=0.735 $X2=0
+ $Y2=0
cc_5154 N_S[7]_c_6565_n N_VGND_c_12777_n 0.00525833f $X=47.065 $Y=0.81 $X2=0
+ $Y2=0
cc_5155 N_S[7]_c_6568_n N_VGND_c_12777_n 0.00862298f $X=47.215 $Y=0.18 $X2=0
+ $Y2=0
cc_5156 N_S[7]_c_6574_n N_VGND_c_12779_n 0.0028166f $X=49.085 $Y=0.18 $X2=0
+ $Y2=0
cc_5157 N_S[7]_c_6575_n N_VGND_c_12779_n 5.5039e-19 $X=49.16 $Y=0.255 $X2=0
+ $Y2=0
cc_5158 N_S[7]_c_6561_n N_VGND_c_12859_n 0.00585385f $X=46.185 $Y=0.735 $X2=0
+ $Y2=0
cc_5159 N_S[7]_c_6562_n N_VGND_c_12859_n 2.16067e-19 $X=46.53 $Y=0.81 $X2=0
+ $Y2=0
cc_5160 N_S[7]_c_6563_n N_VGND_c_12859_n 0.00542362f $X=46.605 $Y=0.735 $X2=0
+ $Y2=0
cc_5161 N_S[7]_c_6568_n N_VGND_c_12863_n 0.0559651f $X=47.215 $Y=0.18 $X2=0
+ $Y2=0
cc_5162 N_S[7]_c_6561_n VGND 0.0119653f $X=46.185 $Y=0.735 $X2=0 $Y2=0
cc_5163 N_S[7]_c_6563_n VGND 0.00990284f $X=46.605 $Y=0.735 $X2=0 $Y2=0
cc_5164 N_S[7]_c_6567_n VGND 0.0244174f $X=47.825 $Y=0.18 $X2=0 $Y2=0
cc_5165 N_S[7]_c_6568_n VGND 0.0101627f $X=47.215 $Y=0.18 $X2=0 $Y2=0
cc_5166 N_S[7]_c_6570_n VGND 0.00642387f $X=48.245 $Y=0.18 $X2=0 $Y2=0
cc_5167 N_S[7]_c_6572_n VGND 0.0064237f $X=48.665 $Y=0.18 $X2=0 $Y2=0
cc_5168 N_S[7]_c_6574_n VGND 0.0123437f $X=49.085 $Y=0.18 $X2=0 $Y2=0
cc_5169 N_S[7]_c_6577_n VGND 0.00366655f $X=47.9 $Y=0.18 $X2=0 $Y2=0
cc_5170 N_S[7]_c_6578_n VGND 0.00366655f $X=48.32 $Y=0.18 $X2=0 $Y2=0
cc_5171 N_S[7]_c_6579_n VGND 0.00366655f $X=48.74 $Y=0.18 $X2=0 $Y2=0
cc_5172 N_S[7]_c_6566_n N_A_9513_66#_c_15195_n 0.00529837f $X=47.14 $Y=0.735
+ $X2=0 $Y2=0
cc_5173 N_S[7]_c_6569_n N_A_9513_66#_c_15196_n 0.0112916f $X=47.9 $Y=0.255 $X2=0
+ $Y2=0
cc_5174 N_S[7]_c_6570_n N_A_9513_66#_c_15196_n 0.00211351f $X=48.245 $Y=0.18
+ $X2=0 $Y2=0
cc_5175 N_S[7]_c_6571_n N_A_9513_66#_c_15196_n 0.0106844f $X=48.32 $Y=0.255
+ $X2=0 $Y2=0
cc_5176 N_S[7]_c_6566_n N_A_9513_66#_c_15197_n 0.00189496f $X=47.14 $Y=0.735
+ $X2=0 $Y2=0
cc_5177 N_S[7]_c_6567_n N_A_9513_66#_c_15197_n 0.00685838f $X=47.825 $Y=0.18
+ $X2=0 $Y2=0
cc_5178 N_S[7]_c_6573_n N_A_9513_66#_c_15198_n 0.0106826f $X=48.74 $Y=0.255
+ $X2=0 $Y2=0
cc_5179 N_S[7]_c_6574_n N_A_9513_66#_c_15198_n 0.00211351f $X=49.085 $Y=0.18
+ $X2=0 $Y2=0
cc_5180 N_S[7]_c_6575_n N_A_9513_66#_c_15198_n 0.0139014f $X=49.16 $Y=0.255
+ $X2=0 $Y2=0
cc_5181 N_S[7]_c_6575_n N_A_9513_66#_c_15201_n 0.00206084f $X=49.16 $Y=0.255
+ $X2=0 $Y2=0
cc_5182 N_S[7]_c_6572_n N_A_9513_66#_c_15214_n 0.0034777f $X=48.665 $Y=0.18
+ $X2=0 $Y2=0
cc_5183 N_S[15]_c_6688_n N_A_9250_599#_c_6930_n 0.00507688f $X=47.9 $Y=5.185
+ $X2=25.905 $Y2=0.425
cc_5184 N_S[15]_c_6703_n N_A_9250_599#_c_6922_n 0.00262132f $X=46.63 $Y=3.99
+ $X2=25.905 $Y2=4.845
cc_5185 N_S[15]_c_6690_n N_A_9250_599#_c_6933_n 0.00509204f $X=48.32 $Y=5.185
+ $X2=0 $Y2=0
cc_5186 N_S[15]_c_6694_n N_A_9250_599#_c_6935_n 0.00507426f $X=49.16 $Y=5.185
+ $X2=0 $Y2=0
cc_5187 N_S[15]_c_6692_n N_A_9250_599#_c_6938_n 0.00509391f $X=48.74 $Y=5.185
+ $X2=0 $Y2=0
cc_5188 N_S[15]_c_6701_n N_A_9250_599#_c_6939_n 0.00929139f $X=46.16 $Y=3.89
+ $X2=0 $Y2=0
cc_5189 N_S[15]_c_6705_n N_A_9250_599#_c_6939_n 0.00970559f $X=46.63 $Y=3.89
+ $X2=0 $Y2=0
cc_5190 N_S[15]_c_6680_n N_A_9250_599#_c_6923_n 0.00207203f $X=46.185 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_5191 N_S[15]_c_6681_n N_A_9250_599#_c_6923_n 0.0111895f $X=46.53 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_5192 N_S[15]_c_6683_n N_A_9250_599#_c_6923_n 9.67113e-19 $X=46.605 $Y=4.705
+ $X2=25.99 $Y2=0.51
cc_5193 N_S[15]_c_6685_n N_A_9250_599#_c_6923_n 6.53442e-19 $X=47.14 $Y=5.185
+ $X2=25.99 $Y2=0.51
cc_5194 N_S[15]_c_6695_n N_A_9250_599#_c_6923_n 0.00426435f $X=46.63 $Y=4.63
+ $X2=25.99 $Y2=0.51
cc_5195 N_S[15]_c_6683_n N_A_9250_599#_c_6924_n 0.00603996f $X=46.605 $Y=4.705
+ $X2=0 $Y2=0
cc_5196 N_S[15]_c_6701_n N_A_9250_599#_c_6940_n 0.00117303f $X=46.16 $Y=3.89
+ $X2=0 $Y2=0
cc_5197 N_S[15]_c_6680_n N_A_9250_599#_c_6940_n 0.00336772f $X=46.185 $Y=4.705
+ $X2=0 $Y2=0
cc_5198 N_S[15]_c_6703_n N_A_9250_599#_c_6940_n 0.00508008f $X=46.63 $Y=3.99
+ $X2=0 $Y2=0
cc_5199 N_S[15]_c_6682_n N_A_9250_599#_c_6940_n 0.00255921f $X=46.63 $Y=4.555
+ $X2=0 $Y2=0
cc_5200 N_S[15]_c_6705_n N_A_9250_599#_c_6940_n 0.00254107f $X=46.63 $Y=3.89
+ $X2=0 $Y2=0
cc_5201 N_S[15]_c_6682_n N_A_9250_599#_c_6925_n 0.0206368f $X=46.63 $Y=4.555
+ $X2=0 $Y2=0
cc_5202 N_S[15]_c_6684_n N_A_9250_599#_c_6925_n 0.0103812f $X=47.065 $Y=4.63
+ $X2=0 $Y2=0
cc_5203 N_S[15]_c_6701_n N_A_9250_599#_c_6942_n 0.00304348f $X=46.16 $Y=3.89
+ $X2=0 $Y2=0
cc_5204 N_S[15]_c_6680_n N_A_9250_599#_c_6942_n 5.48523e-19 $X=46.185 $Y=4.705
+ $X2=0 $Y2=0
cc_5205 N_S[15]_c_6705_n N_A_9250_599#_c_6942_n 0.00216424f $X=46.63 $Y=3.89
+ $X2=0 $Y2=0
cc_5206 N_S[15]_c_6680_n N_A_9250_599#_c_6926_n 0.00289358f $X=46.185 $Y=4.705
+ $X2=0 $Y2=0
cc_5207 N_S[15]_c_6681_n N_A_9250_599#_c_6926_n 0.00429801f $X=46.53 $Y=4.63
+ $X2=0 $Y2=0
cc_5208 N_S[15]_c_6682_n N_A_9250_599#_c_6926_n 0.0085951f $X=46.63 $Y=4.555
+ $X2=0 $Y2=0
cc_5209 N_S[15]_c_6695_n N_A_9250_599#_c_6926_n 0.00268644f $X=46.63 $Y=4.63
+ $X2=0 $Y2=0
cc_5210 N_S[15]_c_6699_n N_A_9250_599#_c_6926_n 0.00541767f $X=46.12 $Y=4.28
+ $X2=0 $Y2=0
cc_5211 N_S[15]_c_6680_n N_A_9250_599#_c_6927_n 0.00416423f $X=46.185 $Y=4.705
+ $X2=0 $Y2=0
cc_5212 N_S[15]_c_6682_n N_A_9250_599#_c_6927_n 0.00322131f $X=46.63 $Y=4.555
+ $X2=0 $Y2=0
cc_5213 N_S[15]_c_6699_n N_A_9250_599#_c_6927_n 0.0228692f $X=46.12 $Y=4.28
+ $X2=0 $Y2=0
cc_5214 N_S[15]_c_6682_n N_A_9250_599#_c_6928_n 0.0175393f $X=46.63 $Y=4.555
+ $X2=0 $Y2=0
cc_5215 N_S[15]_c_6684_n N_A_9250_599#_c_6928_n 0.0179529f $X=47.065 $Y=4.63
+ $X2=0 $Y2=0
cc_5216 N_S[15]_c_6679_n N_VPWR_c_7302_n 0.00652399f $X=46.06 $Y=4.28 $X2=0
+ $Y2=0
cc_5217 N_S[15]_c_6701_n N_VPWR_c_7302_n 0.00986205f $X=46.16 $Y=3.89 $X2=0
+ $Y2=0
cc_5218 N_S[15]_c_6699_n N_VPWR_c_7302_n 0.0157609f $X=46.12 $Y=4.28 $X2=0 $Y2=0
cc_5219 N_S[15]_c_6705_n N_VPWR_c_7304_n 0.00950399f $X=46.63 $Y=3.89 $X2=0
+ $Y2=0
cc_5220 N_S[15]_c_6701_n N_VPWR_c_7343_n 0.0035837f $X=46.16 $Y=3.89 $X2=0 $Y2=0
cc_5221 N_S[15]_c_6705_n N_VPWR_c_7343_n 0.0035837f $X=46.63 $Y=3.89 $X2=0 $Y2=0
cc_5222 N_S[15]_c_6701_n VPWR 0.0070533f $X=46.16 $Y=3.89 $X2=0 $Y2=0
cc_5223 N_S[15]_c_6705_n VPWR 0.00711603f $X=46.63 $Y=3.89 $X2=0 $Y2=0
cc_5224 N_S[15]_c_6688_n N_Z_c_9039_n 0.0134253f $X=47.9 $Y=5.185 $X2=0 $Y2=0
cc_5225 N_S[15]_c_6690_n N_Z_c_9039_n 0.0077801f $X=48.32 $Y=5.185 $X2=0 $Y2=0
cc_5226 N_S[15]_c_6692_n N_Z_c_9039_n 6.35774e-19 $X=48.74 $Y=5.185 $X2=0 $Y2=0
cc_5227 N_S[15]_c_6690_n N_Z_c_9041_n 0.00190704f $X=48.32 $Y=5.185 $X2=0 $Y2=0
cc_5228 N_S[15]_c_6692_n N_Z_c_9041_n 3.10191e-19 $X=48.74 $Y=5.185 $X2=0 $Y2=0
cc_5229 N_S[15]_c_6688_n N_Z_c_9093_n 0.00216436f $X=47.9 $Y=5.185 $X2=0 $Y2=0
cc_5230 N_S[15]_c_6692_n N_Z_c_9095_n 0.00180363f $X=48.74 $Y=5.185 $X2=0 $Y2=0
cc_5231 N_S[15]_c_6692_n N_Z_c_9097_n 0.00462308f $X=48.74 $Y=5.185 $X2=0 $Y2=0
cc_5232 N_S[15]_c_6694_n N_Z_c_9097_n 0.00443615f $X=49.16 $Y=5.185 $X2=0 $Y2=0
cc_5233 N_S[15]_c_6690_n N_Z_c_9098_n 6.35664e-19 $X=48.32 $Y=5.185 $X2=0 $Y2=0
cc_5234 N_S[15]_c_6692_n N_Z_c_9098_n 0.00283489f $X=48.74 $Y=5.185 $X2=0 $Y2=0
cc_5235 N_S[15]_c_6694_n N_Z_c_9098_n 0.002324f $X=49.16 $Y=5.185 $X2=0 $Y2=0
cc_5236 N_S[15]_c_6679_n N_Z_c_9130_n 0.00234109f $X=46.06 $Y=4.28 $X2=0 $Y2=0
cc_5237 N_S[15]_c_6701_n N_Z_c_9130_n 0.00501777f $X=46.16 $Y=3.89 $X2=0 $Y2=0
cc_5238 N_S[15]_c_6680_n N_Z_c_9130_n 2.32936e-19 $X=46.185 $Y=4.705 $X2=0 $Y2=0
cc_5239 N_S[15]_c_6703_n N_Z_c_9130_n 2.55735e-19 $X=46.63 $Y=3.99 $X2=0 $Y2=0
cc_5240 N_S[15]_c_6705_n N_Z_c_9130_n 0.00453198f $X=46.63 $Y=3.89 $X2=0 $Y2=0
cc_5241 N_S[15]_c_6699_n N_Z_c_9130_n 0.0105931f $X=46.12 $Y=4.28 $X2=0 $Y2=0
cc_5242 N_S[15]_c_6694_n N_A_9463_613#_c_12571_n 0.00168571f $X=49.16 $Y=5.185
+ $X2=0 $Y2=0
cc_5243 N_S[15]_c_6705_n N_A_9463_613#_c_12573_n 0.00239129f $X=46.63 $Y=3.89
+ $X2=0 $Y2=0
cc_5244 N_S[15]_c_6679_n N_VGND_c_12776_n 0.00576464f $X=46.06 $Y=4.28 $X2=0
+ $Y2=0
cc_5245 N_S[15]_c_6680_n N_VGND_c_12776_n 0.00374526f $X=46.185 $Y=4.705 $X2=0
+ $Y2=0
cc_5246 N_S[15]_c_6699_n N_VGND_c_12776_n 0.0116218f $X=46.12 $Y=4.28 $X2=0
+ $Y2=0
cc_5247 N_S[15]_c_6683_n N_VGND_c_12778_n 0.00173127f $X=46.605 $Y=4.705 $X2=0
+ $Y2=0
cc_5248 N_S[15]_c_6684_n N_VGND_c_12778_n 0.00525833f $X=47.065 $Y=4.63 $X2=0
+ $Y2=0
cc_5249 N_S[15]_c_6685_n N_VGND_c_12778_n 0.00862298f $X=47.14 $Y=5.185 $X2=0
+ $Y2=0
cc_5250 N_S[15]_c_6693_n N_VGND_c_12780_n 0.0028166f $X=49.085 $Y=5.26 $X2=0
+ $Y2=0
cc_5251 N_S[15]_c_6694_n N_VGND_c_12780_n 5.5039e-19 $X=49.16 $Y=5.185 $X2=0
+ $Y2=0
cc_5252 N_S[15]_c_6680_n N_VGND_c_12861_n 0.00585385f $X=46.185 $Y=4.705 $X2=0
+ $Y2=0
cc_5253 N_S[15]_c_6681_n N_VGND_c_12861_n 2.16067e-19 $X=46.53 $Y=4.63 $X2=0
+ $Y2=0
cc_5254 N_S[15]_c_6683_n N_VGND_c_12861_n 0.00542362f $X=46.605 $Y=4.705 $X2=0
+ $Y2=0
cc_5255 N_S[15]_c_6687_n N_VGND_c_12865_n 0.0559651f $X=47.215 $Y=5.26 $X2=0
+ $Y2=0
cc_5256 N_S[15]_c_6680_n VGND 0.0119653f $X=46.185 $Y=4.705 $X2=0 $Y2=0
cc_5257 N_S[15]_c_6683_n VGND 0.00990284f $X=46.605 $Y=4.705 $X2=0 $Y2=0
cc_5258 N_S[15]_c_6686_n VGND 0.0244174f $X=47.825 $Y=5.26 $X2=0 $Y2=0
cc_5259 N_S[15]_c_6687_n VGND 0.0101627f $X=47.215 $Y=5.26 $X2=0 $Y2=0
cc_5260 N_S[15]_c_6689_n VGND 0.00642387f $X=48.245 $Y=5.26 $X2=0 $Y2=0
cc_5261 N_S[15]_c_6691_n VGND 0.0064237f $X=48.665 $Y=5.26 $X2=0 $Y2=0
cc_5262 N_S[15]_c_6693_n VGND 0.0123437f $X=49.085 $Y=5.26 $X2=0 $Y2=0
cc_5263 N_S[15]_c_6696_n VGND 0.00366655f $X=47.9 $Y=5.26 $X2=0 $Y2=0
cc_5264 N_S[15]_c_6697_n VGND 0.00366655f $X=48.32 $Y=5.26 $X2=0 $Y2=0
cc_5265 N_S[15]_c_6698_n VGND 0.00366655f $X=48.74 $Y=5.26 $X2=0 $Y2=0
cc_5266 N_S[15]_c_6684_n N_A_9513_918#_c_15279_n 0.00529837f $X=47.065 $Y=4.63
+ $X2=0 $Y2=0
cc_5267 N_S[15]_c_6688_n N_A_9513_918#_c_15280_n 0.0112916f $X=47.9 $Y=5.185
+ $X2=0 $Y2=0
cc_5268 N_S[15]_c_6689_n N_A_9513_918#_c_15280_n 0.00211351f $X=48.245 $Y=5.26
+ $X2=0 $Y2=0
cc_5269 N_S[15]_c_6690_n N_A_9513_918#_c_15280_n 0.0106844f $X=48.32 $Y=5.185
+ $X2=0 $Y2=0
cc_5270 N_S[15]_c_6685_n N_A_9513_918#_c_15281_n 0.00189496f $X=47.14 $Y=5.185
+ $X2=0 $Y2=0
cc_5271 N_S[15]_c_6686_n N_A_9513_918#_c_15281_n 0.00685838f $X=47.825 $Y=5.26
+ $X2=0 $Y2=0
cc_5272 N_S[15]_c_6692_n N_A_9513_918#_c_15282_n 0.0106826f $X=48.74 $Y=5.185
+ $X2=0 $Y2=0
cc_5273 N_S[15]_c_6693_n N_A_9513_918#_c_15282_n 0.00211351f $X=49.085 $Y=5.26
+ $X2=0 $Y2=0
cc_5274 N_S[15]_c_6694_n N_A_9513_918#_c_15282_n 0.0139014f $X=49.16 $Y=5.185
+ $X2=0 $Y2=0
cc_5275 N_S[15]_c_6694_n N_A_9513_918#_c_15285_n 0.00206084f $X=49.16 $Y=5.185
+ $X2=0 $Y2=0
cc_5276 N_S[15]_c_6691_n N_A_9513_918#_c_15298_n 0.0034777f $X=48.665 $Y=5.26
+ $X2=0 $Y2=0
cc_5277 N_A_9250_325#_c_6814_n N_A_9250_599#_c_6929_n 0.0129371f $X=47.675
+ $Y=1.475 $X2=0 $Y2=0
cc_5278 N_A_9250_325#_c_6817_n N_A_9250_599#_c_6932_n 0.0129371f $X=48.145
+ $Y=1.475 $X2=0 $Y2=0
cc_5279 N_A_9250_325#_c_6819_n N_A_9250_599#_c_6934_n 0.0129371f $X=48.615
+ $Y=1.475 $X2=0 $Y2=0
cc_5280 N_A_9250_325#_c_6821_n N_A_9250_599#_c_6936_n 0.0129371f $X=49.085
+ $Y=1.475 $X2=0 $Y2=0
cc_5281 N_A_9250_325#_c_6824_n N_VPWR_c_7301_n 0.0356181f $X=46.395 $Y=1.77
+ $X2=0 $Y2=0
cc_5282 N_A_9250_325#_c_6814_n N_VPWR_c_7303_n 0.00367058f $X=47.675 $Y=1.475
+ $X2=0 $Y2=0
cc_5283 N_A_9250_325#_c_6824_n N_VPWR_c_7303_n 0.0316788f $X=46.395 $Y=1.77
+ $X2=0 $Y2=0
cc_5284 N_A_9250_325#_c_6810_n N_VPWR_c_7303_n 0.0193185f $X=47.445 $Y=1.23
+ $X2=0 $Y2=0
cc_5285 N_A_9250_325#_c_6813_n N_VPWR_c_7303_n 6.4101e-19 $X=47.355 $Y=1.23
+ $X2=0 $Y2=0
cc_5286 N_A_9250_325#_c_6821_n N_VPWR_c_7305_n 0.00331565f $X=49.085 $Y=1.475
+ $X2=0 $Y2=0
cc_5287 N_A_9250_325#_c_6824_n N_VPWR_c_7343_n 0.0233824f $X=46.395 $Y=1.77
+ $X2=0 $Y2=0
cc_5288 N_A_9250_325#_c_6814_n VPWR 0.00473731f $X=47.675 $Y=1.475 $X2=0 $Y2=0
cc_5289 N_A_9250_325#_c_6817_n VPWR 0.00362156f $X=48.145 $Y=1.475 $X2=0 $Y2=0
cc_5290 N_A_9250_325#_c_6819_n VPWR 0.00362156f $X=48.615 $Y=1.475 $X2=0 $Y2=0
cc_5291 N_A_9250_325#_c_6821_n VPWR 0.00473731f $X=49.085 $Y=1.475 $X2=0 $Y2=0
cc_5292 N_A_9250_325#_c_6824_n VPWR 0.00593513f $X=46.395 $Y=1.77 $X2=0 $Y2=0
cc_5293 N_A_9250_325#_c_6818_n N_Z_c_9040_n 0.00762343f $X=48.525 $Y=1.4 $X2=0
+ $Y2=0
cc_5294 N_A_9250_325#_c_6823_n N_Z_c_9040_n 0.00704092f $X=48.615 $Y=1.4 $X2=0
+ $Y2=0
cc_5295 N_A_9250_325#_c_6815_n N_Z_c_9092_n 0.00597584f $X=48.055 $Y=1.4 $X2=0
+ $Y2=0
cc_5296 N_A_9250_325#_c_6807_n N_Z_c_9092_n 0.00747617f $X=47.765 $Y=1.4 $X2=0
+ $Y2=0
cc_5297 N_A_9250_325#_c_6818_n N_Z_c_9092_n 0.00145542f $X=48.525 $Y=1.4 $X2=0
+ $Y2=0
cc_5298 N_A_9250_325#_c_6822_n N_Z_c_9092_n 0.00909323f $X=48.145 $Y=1.4 $X2=0
+ $Y2=0
cc_5299 N_A_9250_325#_c_6810_n N_Z_c_9092_n 0.0266078f $X=47.445 $Y=1.23 $X2=0
+ $Y2=0
cc_5300 N_A_9250_325#_c_6820_n N_Z_c_9094_n 0.00918337f $X=48.995 $Y=1.4 $X2=0
+ $Y2=0
cc_5301 N_A_9250_325#_c_6823_n N_Z_c_9094_n 2.98555e-19 $X=48.615 $Y=1.4 $X2=0
+ $Y2=0
cc_5302 N_A_9250_325#_c_6820_n N_Z_c_9096_n 0.00248496f $X=48.995 $Y=1.4 $X2=0
+ $Y2=0
cc_5303 N_A_9250_325#_c_6814_n N_Z_c_9129_n 0.00795576f $X=47.675 $Y=1.475 $X2=0
+ $Y2=0
cc_5304 N_A_9250_325#_c_6807_n N_Z_c_9129_n 2.19754e-19 $X=47.765 $Y=1.4 $X2=0
+ $Y2=0
cc_5305 N_A_9250_325#_c_6824_n N_Z_c_9129_n 0.0329704f $X=46.395 $Y=1.77 $X2=0
+ $Y2=0
cc_5306 N_A_9250_325#_c_6810_n N_Z_c_9129_n 0.0186685f $X=47.445 $Y=1.23 $X2=0
+ $Y2=0
cc_5307 N_A_9250_325#_c_6817_n N_Z_c_9905_n 0.00372248f $X=48.145 $Y=1.475 $X2=0
+ $Y2=0
cc_5308 N_A_9250_325#_c_6819_n N_Z_c_9905_n 0.00372458f $X=48.615 $Y=1.475 $X2=0
+ $Y2=0
cc_5309 N_A_9250_325#_c_6814_n N_Z_c_9145_n 0.0221748f $X=47.675 $Y=1.475 $X2=0
+ $Y2=0
cc_5310 N_A_9250_325#_c_6815_n N_Z_c_9145_n 0.00560592f $X=48.055 $Y=1.4 $X2=0
+ $Y2=0
cc_5311 N_A_9250_325#_c_6807_n N_Z_c_9145_n 0.00425035f $X=47.765 $Y=1.4 $X2=0
+ $Y2=0
cc_5312 N_A_9250_325#_c_6817_n N_Z_c_9145_n 0.0181262f $X=48.145 $Y=1.475 $X2=0
+ $Y2=0
cc_5313 N_A_9250_325#_c_6819_n N_Z_c_9145_n 9.74366e-19 $X=48.615 $Y=1.475 $X2=0
+ $Y2=0
cc_5314 N_A_9250_325#_c_6822_n N_Z_c_9145_n 0.00181273f $X=48.145 $Y=1.4 $X2=0
+ $Y2=0
cc_5315 N_A_9250_325#_c_6810_n N_Z_c_9145_n 0.00240108f $X=47.445 $Y=1.23 $X2=0
+ $Y2=0
cc_5316 N_A_9250_325#_c_6817_n N_Z_c_9146_n 9.74366e-19 $X=48.145 $Y=1.475 $X2=0
+ $Y2=0
cc_5317 N_A_9250_325#_c_6819_n N_Z_c_9146_n 0.0181262f $X=48.615 $Y=1.475 $X2=0
+ $Y2=0
cc_5318 N_A_9250_325#_c_6820_n N_Z_c_9146_n 0.0103509f $X=48.995 $Y=1.4 $X2=0
+ $Y2=0
cc_5319 N_A_9250_325#_c_6821_n N_Z_c_9146_n 0.020403f $X=49.085 $Y=1.475 $X2=0
+ $Y2=0
cc_5320 N_A_9250_325#_c_6823_n N_Z_c_9146_n 0.00415268f $X=48.615 $Y=1.4 $X2=0
+ $Y2=0
cc_5321 N_A_9250_325#_c_6821_n N_A_9463_311#_c_12452_n 0.00151141f $X=49.085
+ $Y=1.475 $X2=0 $Y2=0
cc_5322 N_A_9250_325#_c_6814_n N_A_9463_311#_c_12460_n 0.00307958f $X=47.675
+ $Y=1.475 $X2=0 $Y2=0
cc_5323 N_A_9250_325#_c_6817_n N_A_9463_311#_c_12460_n 0.00307958f $X=48.145
+ $Y=1.475 $X2=0 $Y2=0
cc_5324 N_A_9250_325#_c_6819_n N_A_9463_311#_c_12462_n 0.00307958f $X=48.615
+ $Y=1.475 $X2=0 $Y2=0
cc_5325 N_A_9250_325#_c_6821_n N_A_9463_311#_c_12462_n 0.00799829f $X=49.085
+ $Y=1.475 $X2=0 $Y2=0
cc_5326 N_A_9250_325#_c_6814_n N_A_9463_311#_c_12454_n 0.00499839f $X=47.675
+ $Y=1.475 $X2=0 $Y2=0
cc_5327 N_A_9250_325#_c_6807_n N_A_9463_311#_c_12454_n 0.00561627f $X=47.765
+ $Y=1.4 $X2=0 $Y2=0
cc_5328 N_A_9250_325#_c_6810_n N_A_9463_311#_c_12454_n 0.0218124f $X=47.445
+ $Y=1.23 $X2=0 $Y2=0
cc_5329 N_A_9250_325#_c_6813_n N_A_9463_311#_c_12454_n 5.74251e-19 $X=47.355
+ $Y=1.23 $X2=0 $Y2=0
cc_5330 N_A_9250_325#_c_6817_n N_A_9463_311#_c_12455_n 0.00210632f $X=48.145
+ $Y=1.475 $X2=0 $Y2=0
cc_5331 N_A_9250_325#_c_6818_n N_A_9463_311#_c_12455_n 0.00251792f $X=48.525
+ $Y=1.4 $X2=0 $Y2=0
cc_5332 N_A_9250_325#_c_6819_n N_A_9463_311#_c_12455_n 0.00210632f $X=48.615
+ $Y=1.475 $X2=0 $Y2=0
cc_5333 N_A_9250_325#_c_6821_n N_A_9463_311#_c_12456_n 0.00546785f $X=49.085
+ $Y=1.475 $X2=0 $Y2=0
cc_5334 N_A_9250_325#_c_6810_n N_VGND_c_12777_n 0.0123065f $X=47.445 $Y=1.23
+ $X2=0 $Y2=0
cc_5335 N_A_9250_325#_c_6813_n N_VGND_c_12777_n 2.04129e-19 $X=47.355 $Y=1.23
+ $X2=0 $Y2=0
cc_5336 N_A_9250_325#_c_6808_n N_VGND_c_12859_n 0.0129994f $X=46.395 $Y=0.445
+ $X2=0 $Y2=0
cc_5337 N_A_9250_325#_M1141_d VGND 0.00394793f $X=46.26 $Y=0.235 $X2=0 $Y2=0
cc_5338 N_A_9250_325#_c_6808_n VGND 0.00927134f $X=46.395 $Y=0.445 $X2=0 $Y2=0
cc_5339 N_A_9250_325#_c_6807_n N_A_9513_66#_c_15195_n 0.00600378f $X=47.765
+ $Y=1.4 $X2=0 $Y2=0
cc_5340 N_A_9250_325#_c_6810_n N_A_9513_66#_c_15195_n 0.0028695f $X=47.445
+ $Y=1.23 $X2=0 $Y2=0
cc_5341 N_A_9250_325#_c_6818_n N_A_9513_66#_c_15217_n 7.0477e-19 $X=48.525
+ $Y=1.4 $X2=0 $Y2=0
cc_5342 N_A_9250_599#_c_6939_n N_VPWR_c_7302_n 0.0356181f $X=46.395 $Y=3.14
+ $X2=0 $Y2=0
cc_5343 N_A_9250_599#_c_6929_n N_VPWR_c_7304_n 0.00367058f $X=47.675 $Y=3.965
+ $X2=0 $Y2=0
cc_5344 N_A_9250_599#_c_6939_n N_VPWR_c_7304_n 0.0316788f $X=46.395 $Y=3.14
+ $X2=0 $Y2=0
cc_5345 N_A_9250_599#_c_6925_n N_VPWR_c_7304_n 0.0193185f $X=47.445 $Y=4.21
+ $X2=0 $Y2=0
cc_5346 N_A_9250_599#_c_6928_n N_VPWR_c_7304_n 6.4101e-19 $X=47.355 $Y=4.21
+ $X2=0 $Y2=0
cc_5347 N_A_9250_599#_c_6936_n N_VPWR_c_7306_n 0.00331565f $X=49.085 $Y=3.965
+ $X2=0 $Y2=0
cc_5348 N_A_9250_599#_c_6939_n N_VPWR_c_7343_n 0.0233824f $X=46.395 $Y=3.14
+ $X2=0 $Y2=0
cc_5349 N_A_9250_599#_c_6929_n VPWR 0.00473731f $X=47.675 $Y=3.965 $X2=0 $Y2=0
cc_5350 N_A_9250_599#_c_6932_n VPWR 0.00362156f $X=48.145 $Y=3.965 $X2=0 $Y2=0
cc_5351 N_A_9250_599#_c_6934_n VPWR 0.00362156f $X=48.615 $Y=3.965 $X2=0 $Y2=0
cc_5352 N_A_9250_599#_c_6936_n VPWR 0.00473731f $X=49.085 $Y=3.965 $X2=0 $Y2=0
cc_5353 N_A_9250_599#_c_6939_n VPWR 0.00593513f $X=46.395 $Y=3.14 $X2=0 $Y2=0
cc_5354 N_A_9250_599#_c_6933_n N_Z_c_9041_n 0.00762343f $X=48.525 $Y=4.04 $X2=0
+ $Y2=0
cc_5355 N_A_9250_599#_c_6938_n N_Z_c_9041_n 0.00704092f $X=48.615 $Y=4.04 $X2=0
+ $Y2=0
cc_5356 N_A_9250_599#_c_6930_n N_Z_c_9093_n 0.00597584f $X=48.055 $Y=4.04 $X2=0
+ $Y2=0
cc_5357 N_A_9250_599#_c_6922_n N_Z_c_9093_n 0.00747617f $X=47.765 $Y=4.04 $X2=0
+ $Y2=0
cc_5358 N_A_9250_599#_c_6933_n N_Z_c_9093_n 0.00145542f $X=48.525 $Y=4.04 $X2=0
+ $Y2=0
cc_5359 N_A_9250_599#_c_6937_n N_Z_c_9093_n 0.00909323f $X=48.145 $Y=4.04 $X2=0
+ $Y2=0
cc_5360 N_A_9250_599#_c_6925_n N_Z_c_9093_n 0.0266078f $X=47.445 $Y=4.21 $X2=0
+ $Y2=0
cc_5361 N_A_9250_599#_c_6935_n N_Z_c_9095_n 0.00918337f $X=48.995 $Y=4.04 $X2=0
+ $Y2=0
cc_5362 N_A_9250_599#_c_6938_n N_Z_c_9095_n 2.98555e-19 $X=48.615 $Y=4.04 $X2=0
+ $Y2=0
cc_5363 N_A_9250_599#_c_6935_n N_Z_c_9097_n 0.00248496f $X=48.995 $Y=4.04 $X2=0
+ $Y2=0
cc_5364 N_A_9250_599#_c_6929_n N_Z_c_9130_n 0.00795576f $X=47.675 $Y=3.965 $X2=0
+ $Y2=0
cc_5365 N_A_9250_599#_c_6922_n N_Z_c_9130_n 2.19754e-19 $X=47.765 $Y=4.04 $X2=0
+ $Y2=0
cc_5366 N_A_9250_599#_c_6939_n N_Z_c_9130_n 0.0329704f $X=46.395 $Y=3.14 $X2=0
+ $Y2=0
cc_5367 N_A_9250_599#_c_6925_n N_Z_c_9130_n 0.0186685f $X=47.445 $Y=4.21 $X2=0
+ $Y2=0
cc_5368 N_A_9250_599#_c_6932_n N_Z_c_9933_n 0.00372248f $X=48.145 $Y=3.965 $X2=0
+ $Y2=0
cc_5369 N_A_9250_599#_c_6934_n N_Z_c_9933_n 0.00372458f $X=48.615 $Y=3.965 $X2=0
+ $Y2=0
cc_5370 N_A_9250_599#_c_6929_n N_Z_c_9145_n 0.0221748f $X=47.675 $Y=3.965 $X2=0
+ $Y2=0
cc_5371 N_A_9250_599#_c_6930_n N_Z_c_9145_n 0.00560592f $X=48.055 $Y=4.04 $X2=0
+ $Y2=0
cc_5372 N_A_9250_599#_c_6922_n N_Z_c_9145_n 0.00425035f $X=47.765 $Y=4.04 $X2=0
+ $Y2=0
cc_5373 N_A_9250_599#_c_6932_n N_Z_c_9145_n 0.0181262f $X=48.145 $Y=3.965 $X2=0
+ $Y2=0
cc_5374 N_A_9250_599#_c_6934_n N_Z_c_9145_n 9.74366e-19 $X=48.615 $Y=3.965 $X2=0
+ $Y2=0
cc_5375 N_A_9250_599#_c_6937_n N_Z_c_9145_n 0.00181273f $X=48.145 $Y=4.04 $X2=0
+ $Y2=0
cc_5376 N_A_9250_599#_c_6925_n N_Z_c_9145_n 0.00240108f $X=47.445 $Y=4.21 $X2=0
+ $Y2=0
cc_5377 N_A_9250_599#_c_6932_n N_Z_c_9146_n 9.74366e-19 $X=48.145 $Y=3.965 $X2=0
+ $Y2=0
cc_5378 N_A_9250_599#_c_6934_n N_Z_c_9146_n 0.0181262f $X=48.615 $Y=3.965 $X2=0
+ $Y2=0
cc_5379 N_A_9250_599#_c_6935_n N_Z_c_9146_n 0.0103509f $X=48.995 $Y=4.04 $X2=0
+ $Y2=0
cc_5380 N_A_9250_599#_c_6936_n N_Z_c_9146_n 0.020403f $X=49.085 $Y=3.965 $X2=0
+ $Y2=0
cc_5381 N_A_9250_599#_c_6938_n N_Z_c_9146_n 0.00415268f $X=48.615 $Y=4.04 $X2=0
+ $Y2=0
cc_5382 N_A_9250_599#_c_6936_n N_A_9463_613#_c_12571_n 0.00151141f $X=49.085
+ $Y=3.965 $X2=0 $Y2=0
cc_5383 N_A_9250_599#_c_6929_n N_A_9463_613#_c_12579_n 0.00307958f $X=47.675
+ $Y=3.965 $X2=0 $Y2=0
cc_5384 N_A_9250_599#_c_6932_n N_A_9463_613#_c_12579_n 0.00307958f $X=48.145
+ $Y=3.965 $X2=0 $Y2=0
cc_5385 N_A_9250_599#_c_6934_n N_A_9463_613#_c_12581_n 0.00307958f $X=48.615
+ $Y=3.965 $X2=0 $Y2=0
cc_5386 N_A_9250_599#_c_6936_n N_A_9463_613#_c_12581_n 0.00799829f $X=49.085
+ $Y=3.965 $X2=0 $Y2=0
cc_5387 N_A_9250_599#_c_6929_n N_A_9463_613#_c_12573_n 0.00499839f $X=47.675
+ $Y=3.965 $X2=0 $Y2=0
cc_5388 N_A_9250_599#_c_6922_n N_A_9463_613#_c_12573_n 0.00561627f $X=47.765
+ $Y=4.04 $X2=0 $Y2=0
cc_5389 N_A_9250_599#_c_6925_n N_A_9463_613#_c_12573_n 0.0218124f $X=47.445
+ $Y=4.21 $X2=0 $Y2=0
cc_5390 N_A_9250_599#_c_6928_n N_A_9463_613#_c_12573_n 5.74251e-19 $X=47.355
+ $Y=4.21 $X2=0 $Y2=0
cc_5391 N_A_9250_599#_c_6932_n N_A_9463_613#_c_12574_n 0.00210632f $X=48.145
+ $Y=3.965 $X2=0 $Y2=0
cc_5392 N_A_9250_599#_c_6933_n N_A_9463_613#_c_12574_n 0.00251792f $X=48.525
+ $Y=4.04 $X2=0 $Y2=0
cc_5393 N_A_9250_599#_c_6934_n N_A_9463_613#_c_12574_n 0.00210632f $X=48.615
+ $Y=3.965 $X2=0 $Y2=0
cc_5394 N_A_9250_599#_c_6936_n N_A_9463_613#_c_12575_n 0.00546785f $X=49.085
+ $Y=3.965 $X2=0 $Y2=0
cc_5395 N_A_9250_599#_c_6925_n N_VGND_c_12778_n 0.0123065f $X=47.445 $Y=4.21
+ $X2=0 $Y2=0
cc_5396 N_A_9250_599#_c_6928_n N_VGND_c_12778_n 2.04129e-19 $X=47.355 $Y=4.21
+ $X2=0 $Y2=0
cc_5397 N_A_9250_599#_c_6924_n N_VGND_c_12861_n 0.0129994f $X=46.395 $Y=4.995
+ $X2=0 $Y2=0
cc_5398 N_A_9250_599#_M1174_d VGND 0.00394793f $X=46.26 $Y=4.785 $X2=0 $Y2=0
cc_5399 N_A_9250_599#_c_6924_n VGND 0.00927134f $X=46.395 $Y=4.995 $X2=0 $Y2=0
cc_5400 N_A_9250_599#_c_6922_n N_A_9513_918#_c_15279_n 0.00600378f $X=47.765
+ $Y=4.04 $X2=0 $Y2=0
cc_5401 N_A_9250_599#_c_6925_n N_A_9513_918#_c_15279_n 0.0028695f $X=47.445
+ $Y=4.21 $X2=0 $Y2=0
cc_5402 N_A_9250_599#_c_6933_n N_A_9513_918#_c_15301_n 7.0477e-19 $X=48.525
+ $Y=4.04 $X2=0 $Y2=0
cc_5403 N_D[7]_M1040_g N_D[15]_M1056_g 0.0130744f $X=50.075 $Y=1.985 $X2=0 $Y2=0
cc_5404 N_D[7]_M1087_g N_D[15]_M1103_g 0.0130744f $X=50.545 $Y=1.985 $X2=0 $Y2=0
cc_5405 N_D[7]_M1131_g N_D[15]_M1145_g 0.0130744f $X=51.015 $Y=1.985 $X2=0 $Y2=0
cc_5406 N_D[7]_M1151_g N_D[15]_M1156_g 0.0130744f $X=51.485 $Y=1.985 $X2=25.99
+ $Y2=0.51
cc_5407 N_D[7]_M1040_g N_VPWR_c_7305_n 0.00374733f $X=50.075 $Y=1.985 $X2=0
+ $Y2=0
cc_5408 N_D[7]_M1087_g N_VPWR_c_7307_n 0.00193762f $X=50.545 $Y=1.985 $X2=0
+ $Y2=0
cc_5409 N_D[7]_M1131_g N_VPWR_c_7307_n 0.00193762f $X=51.015 $Y=1.985 $X2=0
+ $Y2=0
cc_5410 N_D[7]_M1151_g N_VPWR_c_7309_n 0.00354866f $X=51.485 $Y=1.985 $X2=0
+ $Y2=0
cc_5411 N_D[7]_M1040_g VPWR 0.00573859f $X=50.075 $Y=1.985 $X2=0 $Y2=0
cc_5412 N_D[7]_M1087_g VPWR 0.00445624f $X=50.545 $Y=1.985 $X2=0 $Y2=0
cc_5413 N_D[7]_M1131_g VPWR 0.00445624f $X=51.015 $Y=1.985 $X2=0 $Y2=0
cc_5414 N_D[7]_M1151_g VPWR 0.0112159f $X=51.485 $Y=1.985 $X2=0 $Y2=0
cc_5415 N_D[7]_M1040_g N_VPWR_c_7367_n 0.0035837f $X=50.075 $Y=1.985 $X2=0 $Y2=0
cc_5416 N_D[7]_M1087_g N_VPWR_c_7367_n 0.0035837f $X=50.545 $Y=1.985 $X2=0 $Y2=0
cc_5417 N_D[7]_M1131_g N_VPWR_c_7368_n 0.0035837f $X=51.015 $Y=1.985 $X2=0 $Y2=0
cc_5418 N_D[7]_M1151_g N_VPWR_c_7368_n 0.0035837f $X=51.485 $Y=1.985 $X2=0 $Y2=0
cc_5419 N_D[7]_M1040_g N_A_9463_311#_c_12451_n 0.0143215f $X=50.075 $Y=1.985
+ $X2=0 $Y2=0
cc_5420 N_D[7]_M1087_g N_A_9463_311#_c_12473_n 0.0102411f $X=50.545 $Y=1.985
+ $X2=0 $Y2=0
cc_5421 N_D[7]_M1131_g N_A_9463_311#_c_12473_n 0.0102411f $X=51.015 $Y=1.985
+ $X2=0 $Y2=0
cc_5422 N_D[7]_c_7051_n N_A_9463_311#_c_12473_n 7.15862e-19 $X=50.925 $Y=1.16
+ $X2=0 $Y2=0
cc_5423 N_D[7]_c_7053_n N_A_9463_311#_c_12473_n 0.0405252f $X=51.38 $Y=1.16
+ $X2=0 $Y2=0
cc_5424 N_D[7]_M1040_g N_A_9463_311#_c_12477_n 8.61029e-19 $X=50.075 $Y=1.985
+ $X2=0 $Y2=0
cc_5425 N_D[7]_M1087_g N_A_9463_311#_c_12477_n 5.79575e-19 $X=50.545 $Y=1.985
+ $X2=0 $Y2=0
cc_5426 N_D[7]_c_7052_n N_A_9463_311#_c_12477_n 8.03631e-19 $X=50.635 $Y=1.16
+ $X2=0 $Y2=0
cc_5427 N_D[7]_c_7053_n N_A_9463_311#_c_12477_n 0.0199757f $X=51.38 $Y=1.16
+ $X2=0 $Y2=0
cc_5428 N_D[7]_M1131_g N_A_9463_311#_c_12481_n 5.79575e-19 $X=51.015 $Y=1.985
+ $X2=0 $Y2=0
cc_5429 N_D[7]_M1151_g N_A_9463_311#_c_12481_n 0.00215964f $X=51.485 $Y=1.985
+ $X2=0 $Y2=0
cc_5430 N_D[7]_c_7053_n N_A_9463_311#_c_12481_n 0.022724f $X=51.38 $Y=1.16 $X2=0
+ $Y2=0
cc_5431 N_D[7]_c_7054_n N_A_9463_311#_c_12481_n 8.03631e-19 $X=51.485 $Y=1.16
+ $X2=0 $Y2=0
cc_5432 N_D[7]_M1040_g N_A_9463_311#_c_12453_n 0.00316234f $X=50.075 $Y=1.985
+ $X2=25.99 $Y2=0.51
cc_5433 N_D[7]_M1087_g N_A_9463_311#_c_12486_n 0.00316234f $X=50.545 $Y=1.985
+ $X2=0 $Y2=0
cc_5434 N_D[7]_M1131_g N_A_9463_311#_c_12486_n 0.00316234f $X=51.015 $Y=1.985
+ $X2=0 $Y2=0
cc_5435 N_D[7]_M1040_g N_A_9463_311#_c_12488_n 0.0104026f $X=50.075 $Y=1.985
+ $X2=0 $Y2=0
cc_5436 N_D[7]_M1087_g N_A_9463_311#_c_12488_n 0.0095928f $X=50.545 $Y=1.985
+ $X2=0 $Y2=0
cc_5437 N_D[7]_M1131_g N_A_9463_311#_c_12488_n 6.38147e-19 $X=51.015 $Y=1.985
+ $X2=0 $Y2=0
cc_5438 N_D[7]_M1087_g N_A_9463_311#_c_12491_n 6.38147e-19 $X=50.545 $Y=1.985
+ $X2=0 $Y2=0
cc_5439 N_D[7]_M1131_g N_A_9463_311#_c_12491_n 0.0095928f $X=51.015 $Y=1.985
+ $X2=0 $Y2=0
cc_5440 N_D[7]_M1151_g N_A_9463_311#_c_12491_n 0.00896273f $X=51.485 $Y=1.985
+ $X2=0 $Y2=0
cc_5441 N_D[7]_M1040_g N_A_9463_311#_c_12456_n 0.0035027f $X=50.075 $Y=1.985
+ $X2=0 $Y2=0
cc_5442 N_D[7]_M1068_g N_VGND_c_12779_n 0.00321269f $X=50.1 $Y=0.56 $X2=0 $Y2=0
cc_5443 N_D[7]_M1115_g N_VGND_c_12779_n 2.6376e-19 $X=50.52 $Y=0.56 $X2=0 $Y2=0
cc_5444 N_D[7]_M1115_g N_VGND_c_12781_n 0.0019152f $X=50.52 $Y=0.56 $X2=0 $Y2=0
cc_5445 N_D[7]_M1216_g N_VGND_c_12781_n 0.00166854f $X=51.04 $Y=0.56 $X2=0 $Y2=0
cc_5446 N_D[7]_M1281_g N_VGND_c_12781_n 2.64031e-19 $X=51.46 $Y=0.56 $X2=0 $Y2=0
cc_5447 N_D[7]_M1281_g N_VGND_c_12784_n 0.00345859f $X=51.46 $Y=0.56 $X2=0 $Y2=0
cc_5448 N_D[7]_M1068_g VGND 0.00702263f $X=50.1 $Y=0.56 $X2=0 $Y2=0
cc_5449 N_D[7]_M1115_g VGND 0.00624811f $X=50.52 $Y=0.56 $X2=0 $Y2=0
cc_5450 N_D[7]_M1216_g VGND 0.00593887f $X=51.04 $Y=0.56 $X2=0 $Y2=0
cc_5451 N_D[7]_M1281_g VGND 0.0107845f $X=51.46 $Y=0.56 $X2=0 $Y2=0
cc_5452 N_D[7]_M1068_g N_VGND_c_12893_n 0.00422241f $X=50.1 $Y=0.56 $X2=0 $Y2=0
cc_5453 N_D[7]_M1115_g N_VGND_c_12893_n 0.00430643f $X=50.52 $Y=0.56 $X2=0 $Y2=0
cc_5454 N_D[7]_M1216_g N_VGND_c_12895_n 0.00422241f $X=51.04 $Y=0.56 $X2=0 $Y2=0
cc_5455 N_D[7]_M1281_g N_VGND_c_12895_n 0.00551064f $X=51.46 $Y=0.56 $X2=0 $Y2=0
cc_5456 N_D[7]_M1068_g N_A_9513_66#_c_15199_n 0.00261078f $X=50.1 $Y=0.56
+ $X2=25.99 $Y2=0.51
cc_5457 N_D[7]_M1068_g N_A_9513_66#_c_15200_n 0.0121912f $X=50.1 $Y=0.56 $X2=0
+ $Y2=0
cc_5458 N_D[7]_M1068_g N_A_9513_66#_c_15220_n 0.00699463f $X=50.1 $Y=0.56 $X2=0
+ $Y2=0
cc_5459 N_D[7]_M1115_g N_A_9513_66#_c_15220_n 0.00661764f $X=50.52 $Y=0.56 $X2=0
+ $Y2=0
cc_5460 N_D[7]_M1216_g N_A_9513_66#_c_15220_n 5.22365e-19 $X=51.04 $Y=0.56 $X2=0
+ $Y2=0
cc_5461 N_D[7]_M1115_g N_A_9513_66#_c_15202_n 0.00900364f $X=50.52 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_5462 N_D[7]_M1216_g N_A_9513_66#_c_15202_n 0.00986515f $X=51.04 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_5463 N_D[7]_M1281_g N_A_9513_66#_c_15202_n 0.00228093f $X=51.46 $Y=0.56
+ $X2=25.99 $Y2=4.8
cc_5464 N_D[7]_c_7051_n N_A_9513_66#_c_15202_n 0.00463549f $X=50.925 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_5465 N_D[7]_c_7053_n N_A_9513_66#_c_15202_n 0.0608884f $X=51.38 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_5466 N_D[7]_c_7054_n N_A_9513_66#_c_15202_n 0.00208088f $X=51.485 $Y=1.16
+ $X2=25.99 $Y2=4.8
cc_5467 N_D[7]_M1115_g N_A_9513_66#_c_15229_n 5.22365e-19 $X=50.52 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_5468 N_D[7]_M1216_g N_A_9513_66#_c_15229_n 0.00661134f $X=51.04 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_5469 N_D[7]_M1281_g N_A_9513_66#_c_15229_n 0.00529286f $X=51.46 $Y=0.56
+ $X2=25.99 $Y2=4.93
cc_5470 N_D[7]_M1068_g N_A_9513_66#_c_15203_n 0.00128201f $X=50.1 $Y=0.56 $X2=0
+ $Y2=0
cc_5471 N_D[7]_M1115_g N_A_9513_66#_c_15203_n 8.68782e-19 $X=50.52 $Y=0.56 $X2=0
+ $Y2=0
cc_5472 N_D[7]_c_7052_n N_A_9513_66#_c_15203_n 0.00208088f $X=50.635 $Y=1.16
+ $X2=0 $Y2=0
cc_5473 N_D[7]_c_7053_n N_A_9513_66#_c_15203_n 0.018367f $X=51.38 $Y=1.16 $X2=0
+ $Y2=0
cc_5474 N_D[15]_M1056_g N_VPWR_c_7306_n 0.00374733f $X=50.075 $Y=3.455 $X2=0
+ $Y2=0
cc_5475 N_D[15]_M1103_g N_VPWR_c_7308_n 0.00193762f $X=50.545 $Y=3.455 $X2=0
+ $Y2=0
cc_5476 N_D[15]_M1145_g N_VPWR_c_7308_n 0.00193762f $X=51.015 $Y=3.455 $X2=0
+ $Y2=0
cc_5477 N_D[15]_M1156_g N_VPWR_c_7310_n 0.00354866f $X=51.485 $Y=3.455 $X2=0
+ $Y2=0
cc_5478 N_D[15]_M1056_g VPWR 0.00573859f $X=50.075 $Y=3.455 $X2=0 $Y2=0
cc_5479 N_D[15]_M1103_g VPWR 0.00445624f $X=50.545 $Y=3.455 $X2=0 $Y2=0
cc_5480 N_D[15]_M1145_g VPWR 0.00445624f $X=51.015 $Y=3.455 $X2=0 $Y2=0
cc_5481 N_D[15]_M1156_g VPWR 0.0112159f $X=51.485 $Y=3.455 $X2=0 $Y2=0
cc_5482 N_D[15]_M1056_g N_VPWR_c_7367_n 0.0035837f $X=50.075 $Y=3.455 $X2=0
+ $Y2=0
cc_5483 N_D[15]_M1103_g N_VPWR_c_7367_n 0.0035837f $X=50.545 $Y=3.455 $X2=0
+ $Y2=0
cc_5484 N_D[15]_M1145_g N_VPWR_c_7368_n 0.0035837f $X=51.015 $Y=3.455 $X2=0
+ $Y2=0
cc_5485 N_D[15]_M1156_g N_VPWR_c_7368_n 0.0035837f $X=51.485 $Y=3.455 $X2=0
+ $Y2=0
cc_5486 N_D[15]_M1056_g N_A_9463_613#_c_12570_n 0.0143215f $X=50.075 $Y=3.455
+ $X2=0 $Y2=0
cc_5487 N_D[15]_M1103_g N_A_9463_613#_c_12592_n 0.0102411f $X=50.545 $Y=3.455
+ $X2=0 $Y2=0
cc_5488 N_D[15]_M1145_g N_A_9463_613#_c_12592_n 0.0102411f $X=51.015 $Y=3.455
+ $X2=0 $Y2=0
cc_5489 N_D[15]_c_7139_n N_A_9463_613#_c_12592_n 7.15862e-19 $X=50.925 $Y=4.28
+ $X2=0 $Y2=0
cc_5490 N_D[15]_c_7141_n N_A_9463_613#_c_12592_n 0.0405252f $X=51.38 $Y=4.28
+ $X2=0 $Y2=0
cc_5491 N_D[15]_M1056_g N_A_9463_613#_c_12596_n 8.61029e-19 $X=50.075 $Y=3.455
+ $X2=0 $Y2=0
cc_5492 N_D[15]_M1103_g N_A_9463_613#_c_12596_n 5.79575e-19 $X=50.545 $Y=3.455
+ $X2=0 $Y2=0
cc_5493 N_D[15]_c_7140_n N_A_9463_613#_c_12596_n 8.03631e-19 $X=50.635 $Y=4.28
+ $X2=0 $Y2=0
cc_5494 N_D[15]_c_7141_n N_A_9463_613#_c_12596_n 0.0199757f $X=51.38 $Y=4.28
+ $X2=0 $Y2=0
cc_5495 N_D[15]_M1145_g N_A_9463_613#_c_12600_n 5.79575e-19 $X=51.015 $Y=3.455
+ $X2=0 $Y2=0
cc_5496 N_D[15]_M1156_g N_A_9463_613#_c_12600_n 0.00215964f $X=51.485 $Y=3.455
+ $X2=0 $Y2=0
cc_5497 N_D[15]_c_7141_n N_A_9463_613#_c_12600_n 0.022724f $X=51.38 $Y=4.28
+ $X2=0 $Y2=0
cc_5498 N_D[15]_c_7142_n N_A_9463_613#_c_12600_n 8.03631e-19 $X=51.485 $Y=4.28
+ $X2=0 $Y2=0
cc_5499 N_D[15]_M1056_g N_A_9463_613#_c_12572_n 0.00316234f $X=50.075 $Y=3.455
+ $X2=25.99 $Y2=0.51
cc_5500 N_D[15]_M1103_g N_A_9463_613#_c_12605_n 0.00316234f $X=50.545 $Y=3.455
+ $X2=0 $Y2=0
cc_5501 N_D[15]_M1145_g N_A_9463_613#_c_12605_n 0.00316234f $X=51.015 $Y=3.455
+ $X2=0 $Y2=0
cc_5502 N_D[15]_M1056_g N_A_9463_613#_c_12575_n 0.0035027f $X=50.075 $Y=3.455
+ $X2=0 $Y2=0
cc_5503 N_D[15]_M1056_g N_A_9463_613#_c_12608_n 0.0104026f $X=50.075 $Y=3.455
+ $X2=0 $Y2=0
cc_5504 N_D[15]_M1103_g N_A_9463_613#_c_12608_n 0.0095928f $X=50.545 $Y=3.455
+ $X2=0 $Y2=0
cc_5505 N_D[15]_M1145_g N_A_9463_613#_c_12608_n 6.38147e-19 $X=51.015 $Y=3.455
+ $X2=0 $Y2=0
cc_5506 N_D[15]_M1103_g N_A_9463_613#_c_12611_n 6.38147e-19 $X=50.545 $Y=3.455
+ $X2=0 $Y2=0
cc_5507 N_D[15]_M1145_g N_A_9463_613#_c_12611_n 0.0095928f $X=51.015 $Y=3.455
+ $X2=0 $Y2=0
cc_5508 N_D[15]_M1156_g N_A_9463_613#_c_12611_n 0.00896273f $X=51.485 $Y=3.455
+ $X2=0 $Y2=0
cc_5509 N_D[15]_M1073_g N_VGND_c_12780_n 0.00321269f $X=50.1 $Y=4.88 $X2=0 $Y2=0
cc_5510 N_D[15]_M1144_g N_VGND_c_12780_n 2.6376e-19 $X=50.52 $Y=4.88 $X2=0 $Y2=0
cc_5511 N_D[15]_M1144_g N_VGND_c_12782_n 0.0019152f $X=50.52 $Y=4.88 $X2=0 $Y2=0
cc_5512 N_D[15]_M1190_g N_VGND_c_12782_n 0.00166854f $X=51.04 $Y=4.88 $X2=0
+ $Y2=0
cc_5513 N_D[15]_M1278_g N_VGND_c_12782_n 2.64031e-19 $X=51.46 $Y=4.88 $X2=0
+ $Y2=0
cc_5514 N_D[15]_M1278_g N_VGND_c_12786_n 0.00345859f $X=51.46 $Y=4.88 $X2=0
+ $Y2=0
cc_5515 N_D[15]_M1073_g VGND 0.00702263f $X=50.1 $Y=4.88 $X2=0 $Y2=0
cc_5516 N_D[15]_M1144_g VGND 0.00624811f $X=50.52 $Y=4.88 $X2=0 $Y2=0
cc_5517 N_D[15]_M1190_g VGND 0.00593887f $X=51.04 $Y=4.88 $X2=0 $Y2=0
cc_5518 N_D[15]_M1278_g VGND 0.0107845f $X=51.46 $Y=4.88 $X2=0 $Y2=0
cc_5519 N_D[15]_M1073_g N_VGND_c_12894_n 0.00422241f $X=50.1 $Y=4.88 $X2=0 $Y2=0
cc_5520 N_D[15]_M1144_g N_VGND_c_12894_n 0.00430643f $X=50.52 $Y=4.88 $X2=0
+ $Y2=0
cc_5521 N_D[15]_M1190_g N_VGND_c_12896_n 0.00422241f $X=51.04 $Y=4.88 $X2=0
+ $Y2=0
cc_5522 N_D[15]_M1278_g N_VGND_c_12896_n 0.00551064f $X=51.46 $Y=4.88 $X2=0
+ $Y2=0
cc_5523 N_D[15]_M1073_g N_A_9513_918#_c_15283_n 0.00261078f $X=50.1 $Y=4.88
+ $X2=25.99 $Y2=0.51
cc_5524 N_D[15]_M1073_g N_A_9513_918#_c_15284_n 0.0121912f $X=50.1 $Y=4.88 $X2=0
+ $Y2=0
cc_5525 N_D[15]_M1144_g N_A_9513_918#_c_15304_n 0.00900364f $X=50.52 $Y=4.88
+ $X2=0 $Y2=0
cc_5526 N_D[15]_M1190_g N_A_9513_918#_c_15304_n 0.00899636f $X=51.04 $Y=4.88
+ $X2=0 $Y2=0
cc_5527 N_D[15]_c_7139_n N_A_9513_918#_c_15304_n 0.00463549f $X=50.925 $Y=4.28
+ $X2=0 $Y2=0
cc_5528 N_D[15]_c_7141_n N_A_9513_918#_c_15304_n 0.0394855f $X=51.38 $Y=4.28
+ $X2=0 $Y2=0
cc_5529 N_D[15]_M1073_g N_A_9513_918#_c_15286_n 0.00827664f $X=50.1 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_5530 N_D[15]_M1144_g N_A_9513_918#_c_15286_n 0.00748643f $X=50.52 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_5531 N_D[15]_M1190_g N_A_9513_918#_c_15286_n 5.22365e-19 $X=51.04 $Y=4.88
+ $X2=25.99 $Y2=4.93
cc_5532 N_D[15]_c_7140_n N_A_9513_918#_c_15286_n 0.00208088f $X=50.635 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_5533 N_D[15]_c_7141_n N_A_9513_918#_c_15286_n 0.018367f $X=51.38 $Y=4.28
+ $X2=25.99 $Y2=4.93
cc_5534 N_D[15]_M1144_g N_A_9513_918#_c_15287_n 5.22365e-19 $X=50.52 $Y=4.88
+ $X2=0 $Y2=0
cc_5535 N_D[15]_M1190_g N_A_9513_918#_c_15287_n 0.00748012f $X=51.04 $Y=4.88
+ $X2=0 $Y2=0
cc_5536 N_D[15]_M1278_g N_A_9513_918#_c_15287_n 0.00757379f $X=51.46 $Y=4.88
+ $X2=0 $Y2=0
cc_5537 N_D[15]_c_7141_n N_A_9513_918#_c_15287_n 0.021403f $X=51.38 $Y=4.28
+ $X2=0 $Y2=0
cc_5538 N_D[15]_c_7142_n N_A_9513_918#_c_15287_n 0.00208088f $X=51.485 $Y=4.28
+ $X2=0 $Y2=0
cc_5539 VPWR N_A_117_297#_M1014_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_5540 VPWR N_A_117_297#_M1208_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_5541 N_VPWR_M1146_d N_A_117_297#_c_8776_n 0.00346031f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_5542 N_VPWR_c_7219_n N_A_117_297#_c_8776_n 0.0138552f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_5543 N_VPWR_M1294_d N_A_117_297#_c_8771_n 0.00732532f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_5544 N_VPWR_c_7222_n N_A_117_297#_c_8771_n 0.0175034f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_5545 N_VPWR_M1146_d N_A_117_297#_c_8789_n 2.7385e-19 $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_5546 N_VPWR_c_7219_n N_A_117_297#_c_8789_n 0.0156895f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_5547 N_VPWR_c_7221_n N_A_117_297#_c_8789_n 8.30334e-19 $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5548 VPWR N_A_117_297#_c_8789_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5549 N_VPWR_c_7350_n N_A_117_297#_c_8789_n 8.30334e-19 $X=1.065 $Y=2.72 $X2=0
+ $Y2=0
cc_5550 N_VPWR_c_7217_n N_A_117_297#_c_8825_n 0.00167228f $X=0.26 $Y=1.66
+ $X2=25.99 $Y2=1.87
cc_5551 N_VPWR_c_7219_n N_A_117_297#_c_8825_n 6.68271e-19 $X=1.2 $Y=2 $X2=25.99
+ $Y2=1.87
cc_5552 VPWR N_A_117_297#_c_8825_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5553 N_VPWR_c_7221_n N_A_117_297#_c_8772_n 8.30334e-19 $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5554 N_VPWR_c_7222_n N_A_117_297#_c_8772_n 0.0160196f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_5555 VPWR N_A_117_297#_c_8772_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5556 N_VPWR_c_7351_n N_A_117_297#_c_8772_n 0.00115812f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_5557 N_VPWR_c_7219_n N_A_117_297#_c_8832_n 6.68271e-19 $X=1.2 $Y=2 $X2=25.99
+ $Y2=2.21
cc_5558 N_VPWR_c_7222_n N_A_117_297#_c_8832_n 6.68271e-19 $X=2.14 $Y=2 $X2=25.99
+ $Y2=2.21
cc_5559 VPWR N_A_117_297#_c_8832_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5560 VPWR N_A_117_297#_c_8800_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5561 N_VPWR_c_7222_n N_A_117_297#_c_8836_n 6.69936e-19 $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_5562 VPWR N_A_117_297#_c_8836_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5563 VPWR N_A_117_297#_c_8802_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5564 VPWR N_A_117_297#_c_8839_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5565 N_VPWR_c_7219_n N_A_117_297#_c_8792_n 0.0254588f $X=1.2 $Y=2 $X2=25.99
+ $Y2=3.57
cc_5566 VPWR N_A_117_297#_c_8792_n 0.00345059f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.57
cc_5567 N_VPWR_c_7350_n N_A_117_297#_c_8792_n 0.0189467f $X=1.065 $Y=2.72
+ $X2=25.99 $Y2=3.57
cc_5568 N_VPWR_c_7219_n N_A_117_297#_c_8795_n 0.0254588f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_5569 N_VPWR_c_7221_n N_A_117_297#_c_8795_n 0.0189467f $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5570 N_VPWR_c_7222_n N_A_117_297#_c_8795_n 0.0254588f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_5571 VPWR N_A_117_297#_c_8795_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5572 N_VPWR_c_7224_n N_A_117_297#_c_8847_n 0.00167067f $X=5.115 $Y=1.77 $X2=0
+ $Y2=0
cc_5573 VPWR N_A_117_297#_c_8847_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5574 N_VPWR_c_7222_n N_A_117_297#_c_8773_n 0.0403522f $X=2.14 $Y=2 $X2=0
+ $Y2=0
cc_5575 VPWR N_A_117_297#_c_8773_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5576 N_VPWR_c_7351_n N_A_117_297#_c_8773_n 0.0213652f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_5577 VPWR N_A_117_297#_c_8774_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5578 N_VPWR_c_7224_n N_A_117_297#_c_8775_n 0.0505494f $X=5.115 $Y=1.77 $X2=0
+ $Y2=0
cc_5579 N_VPWR_c_7311_n N_A_117_297#_c_8775_n 0.0213652f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_5580 VPWR N_A_117_297#_c_8775_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5581 VPWR N_A_117_591#_M1023_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_5582 VPWR N_A_117_591#_M1221_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_5583 N_VPWR_M1155_d N_A_117_591#_c_8892_n 0.00346031f $X=1.055 $Y=2.955 $X2=0
+ $Y2=0
cc_5584 N_VPWR_c_7220_n N_A_117_591#_c_8892_n 0.0138552f $X=1.2 $Y=3.1 $X2=0
+ $Y2=0
cc_5585 N_VPWR_M1304_d N_A_117_591#_c_8887_n 0.00732532f $X=1.995 $Y=2.955 $X2=0
+ $Y2=0
cc_5586 N_VPWR_c_7223_n N_A_117_591#_c_8887_n 0.0175034f $X=2.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5587 N_VPWR_M1155_d N_A_117_591#_c_8905_n 2.7385e-19 $X=1.055 $Y=2.955 $X2=0
+ $Y2=0
cc_5588 N_VPWR_c_7220_n N_A_117_591#_c_8905_n 0.0156895f $X=1.2 $Y=3.1 $X2=0
+ $Y2=0
cc_5589 N_VPWR_c_7221_n N_A_117_591#_c_8905_n 8.30334e-19 $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5590 VPWR N_A_117_591#_c_8905_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5591 N_VPWR_c_7350_n N_A_117_591#_c_8905_n 8.30334e-19 $X=1.065 $Y=2.72 $X2=0
+ $Y2=0
cc_5592 N_VPWR_c_7218_n N_A_117_591#_c_8941_n 0.00167228f $X=0.26 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_5593 N_VPWR_c_7220_n N_A_117_591#_c_8941_n 6.68271e-19 $X=1.2 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_5594 VPWR N_A_117_591#_c_8941_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5595 N_VPWR_c_7221_n N_A_117_591#_c_8888_n 8.30334e-19 $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5596 N_VPWR_c_7223_n N_A_117_591#_c_8888_n 0.0160196f $X=2.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5597 VPWR N_A_117_591#_c_8888_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5598 N_VPWR_c_7351_n N_A_117_591#_c_8888_n 0.00115812f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_5599 N_VPWR_c_7220_n N_A_117_591#_c_8948_n 6.68271e-19 $X=1.2 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_5600 N_VPWR_c_7223_n N_A_117_591#_c_8948_n 6.68271e-19 $X=2.14 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_5601 VPWR N_A_117_591#_c_8948_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5602 VPWR N_A_117_591#_c_8916_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5603 N_VPWR_c_7223_n N_A_117_591#_c_8952_n 6.69936e-19 $X=2.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5604 VPWR N_A_117_591#_c_8952_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5605 VPWR N_A_117_591#_c_8918_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5606 VPWR N_A_117_591#_c_8955_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5607 N_VPWR_c_7225_n N_A_117_591#_c_8956_n 0.00167067f $X=5.115 $Y=3.14 $X2=0
+ $Y2=0
cc_5608 VPWR N_A_117_591#_c_8956_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5609 N_VPWR_c_7220_n N_A_117_591#_c_8908_n 0.0254588f $X=1.2 $Y=3.1 $X2=0
+ $Y2=0
cc_5610 VPWR N_A_117_591#_c_8908_n 0.00345059f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5611 N_VPWR_c_7350_n N_A_117_591#_c_8908_n 0.0189467f $X=1.065 $Y=2.72 $X2=0
+ $Y2=0
cc_5612 N_VPWR_c_7220_n N_A_117_591#_c_8911_n 0.0254588f $X=1.2 $Y=3.1 $X2=0
+ $Y2=0
cc_5613 N_VPWR_c_7221_n N_A_117_591#_c_8911_n 0.0189467f $X=2.005 $Y=2.72 $X2=0
+ $Y2=0
cc_5614 N_VPWR_c_7223_n N_A_117_591#_c_8911_n 0.0254588f $X=2.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5615 VPWR N_A_117_591#_c_8911_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5616 N_VPWR_c_7223_n N_A_117_591#_c_8889_n 0.0403522f $X=2.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5617 VPWR N_A_117_591#_c_8889_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5618 N_VPWR_c_7351_n N_A_117_591#_c_8889_n 0.0213652f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_5619 VPWR N_A_117_591#_c_8890_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5620 N_VPWR_c_7225_n N_A_117_591#_c_8891_n 0.0505494f $X=5.115 $Y=3.14 $X2=0
+ $Y2=0
cc_5621 N_VPWR_c_7311_n N_A_117_591#_c_8891_n 0.0213652f $X=4.95 $Y=2.72 $X2=0
+ $Y2=0
cc_5622 VPWR N_A_117_591#_c_8891_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5623 N_VPWR_M1018_d N_Z_c_9115_n 8.15553e-19 $X=4.99 $Y=1.625 $X2=0 $Y2=0
cc_5624 N_VPWR_M1061_d N_Z_c_9115_n 2.0504e-19 $X=5.91 $Y=1.625 $X2=0 $Y2=0
cc_5625 N_VPWR_M1133_d N_Z_c_9115_n 2.0504e-19 $X=6.7 $Y=1.625 $X2=0 $Y2=0
cc_5626 N_VPWR_M1180_d N_Z_c_9115_n 8.15553e-19 $X=7.62 $Y=1.625 $X2=0 $Y2=0
cc_5627 N_VPWR_c_7224_n N_Z_c_9115_n 0.0196216f $X=5.115 $Y=1.77 $X2=0 $Y2=0
cc_5628 N_VPWR_c_7226_n N_Z_c_9115_n 0.0222682f $X=6.055 $Y=1.77 $X2=0 $Y2=0
cc_5629 N_VPWR_c_7229_n N_Z_c_9115_n 0.0222682f $X=6.825 $Y=1.77 $X2=0 $Y2=0
cc_5630 N_VPWR_c_7231_n N_Z_c_9115_n 0.0196216f $X=7.765 $Y=1.77 $X2=0 $Y2=0
cc_5631 VPWR N_Z_c_9115_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5632 N_VPWR_M1123_d N_Z_c_9116_n 8.15553e-19 $X=4.99 $Y=2.995 $X2=0 $Y2=0
cc_5633 N_VPWR_M1172_d N_Z_c_9116_n 2.0504e-19 $X=5.91 $Y=2.995 $X2=0 $Y2=0
cc_5634 N_VPWR_M1225_d N_Z_c_9116_n 2.0504e-19 $X=6.7 $Y=2.995 $X2=0 $Y2=0
cc_5635 N_VPWR_M1266_d N_Z_c_9116_n 8.15553e-19 $X=7.62 $Y=2.995 $X2=0 $Y2=0
cc_5636 N_VPWR_c_7225_n N_Z_c_9116_n 0.0196216f $X=5.115 $Y=3.14 $X2=0 $Y2=0
cc_5637 N_VPWR_c_7227_n N_Z_c_9116_n 0.0222682f $X=6.055 $Y=3.14 $X2=0 $Y2=0
cc_5638 N_VPWR_c_7230_n N_Z_c_9116_n 0.0222682f $X=6.825 $Y=3.14 $X2=0 $Y2=0
cc_5639 N_VPWR_c_7232_n N_Z_c_9116_n 0.0196216f $X=7.765 $Y=3.14 $X2=0 $Y2=0
cc_5640 VPWR N_Z_c_9116_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5641 N_VPWR_M1002_s N_Z_c_9117_n 0.00213438f $X=10.615 $Y=1.485 $X2=0 $Y2=0
cc_5642 N_VPWR_M1038_s N_Z_c_9117_n 0.00236137f $X=11.535 $Y=1.485 $X2=0 $Y2=0
cc_5643 N_VPWR_M1271_s N_Z_c_9117_n 2.0504e-19 $X=12.475 $Y=1.485 $X2=0 $Y2=0
cc_5644 N_VPWR_M1020_s N_Z_c_9117_n 2.0504e-19 $X=13.015 $Y=1.485 $X2=0 $Y2=0
cc_5645 N_VPWR_M1067_s N_Z_c_9117_n 0.00236137f $X=13.935 $Y=1.485 $X2=0 $Y2=0
cc_5646 N_VPWR_M1301_s N_Z_c_9117_n 0.00213438f $X=14.875 $Y=1.485 $X2=0 $Y2=0
cc_5647 N_VPWR_c_7233_n N_Z_c_9117_n 0.0106064f $X=10.74 $Y=2 $X2=0 $Y2=0
cc_5648 N_VPWR_c_7235_n N_Z_c_9117_n 0.010348f $X=11.68 $Y=2 $X2=0 $Y2=0
cc_5649 N_VPWR_c_7237_n N_Z_c_9117_n 0.0276847f $X=12.62 $Y=1.66 $X2=0 $Y2=0
cc_5650 N_VPWR_c_7240_n N_Z_c_9117_n 0.0276847f $X=13.14 $Y=1.66 $X2=0 $Y2=0
cc_5651 N_VPWR_c_7242_n N_Z_c_9117_n 0.010348f $X=14.08 $Y=2 $X2=0 $Y2=0
cc_5652 N_VPWR_c_7245_n N_Z_c_9117_n 0.0106064f $X=15.02 $Y=2 $X2=0 $Y2=0
cc_5653 VPWR N_Z_c_9117_n 0.0537526f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5654 N_VPWR_M1011_s N_Z_c_9118_n 0.00213438f $X=10.615 $Y=2.955 $X2=0 $Y2=0
cc_5655 N_VPWR_M1051_s N_Z_c_9118_n 0.00236137f $X=11.535 $Y=2.955 $X2=0 $Y2=0
cc_5656 N_VPWR_M1285_s N_Z_c_9118_n 2.0504e-19 $X=12.475 $Y=2.955 $X2=0 $Y2=0
cc_5657 N_VPWR_M1024_s N_Z_c_9118_n 2.0504e-19 $X=13.015 $Y=2.955 $X2=0 $Y2=0
cc_5658 N_VPWR_M1076_s N_Z_c_9118_n 0.00236137f $X=13.935 $Y=2.955 $X2=0 $Y2=0
cc_5659 N_VPWR_M1309_s N_Z_c_9118_n 0.00213438f $X=14.875 $Y=2.955 $X2=0 $Y2=0
cc_5660 N_VPWR_c_7234_n N_Z_c_9118_n 0.0106064f $X=10.74 $Y=3.1 $X2=0 $Y2=0
cc_5661 N_VPWR_c_7236_n N_Z_c_9118_n 0.010348f $X=11.68 $Y=3.1 $X2=0 $Y2=0
cc_5662 N_VPWR_c_7238_n N_Z_c_9118_n 0.0276847f $X=12.62 $Y=3.1 $X2=0 $Y2=0
cc_5663 N_VPWR_c_7241_n N_Z_c_9118_n 0.0276847f $X=13.14 $Y=3.1 $X2=0 $Y2=0
cc_5664 N_VPWR_c_7243_n N_Z_c_9118_n 0.010348f $X=14.08 $Y=3.1 $X2=0 $Y2=0
cc_5665 N_VPWR_c_7246_n N_Z_c_9118_n 0.0106064f $X=15.02 $Y=3.1 $X2=0 $Y2=0
cc_5666 VPWR N_Z_c_9118_n 0.0537526f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5667 N_VPWR_M1065_s N_Z_c_9119_n 8.15553e-19 $X=17.87 $Y=1.625 $X2=0 $Y2=0
cc_5668 N_VPWR_M1308_s N_Z_c_9119_n 2.0504e-19 $X=18.79 $Y=1.625 $X2=0 $Y2=0
cc_5669 N_VPWR_M1150_s N_Z_c_9119_n 2.0504e-19 $X=19.58 $Y=1.625 $X2=0 $Y2=0
cc_5670 N_VPWR_M1280_s N_Z_c_9119_n 8.15553e-19 $X=20.5 $Y=1.625 $X2=0 $Y2=0
cc_5671 N_VPWR_c_7247_n N_Z_c_9119_n 0.0196216f $X=17.995 $Y=1.77 $X2=0 $Y2=0
cc_5672 N_VPWR_c_7249_n N_Z_c_9119_n 0.0222682f $X=18.935 $Y=1.77 $X2=0 $Y2=0
cc_5673 N_VPWR_c_7252_n N_Z_c_9119_n 0.0222682f $X=19.705 $Y=1.77 $X2=0 $Y2=0
cc_5674 N_VPWR_c_7254_n N_Z_c_9119_n 0.0196216f $X=20.645 $Y=1.77 $X2=0 $Y2=0
cc_5675 VPWR N_Z_c_9119_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5676 N_VPWR_M1083_d N_Z_c_9120_n 8.15553e-19 $X=17.87 $Y=2.995 $X2=0 $Y2=0
cc_5677 N_VPWR_M1173_d N_Z_c_9120_n 2.0504e-19 $X=18.79 $Y=2.995 $X2=0 $Y2=0
cc_5678 N_VPWR_M1066_d N_Z_c_9120_n 2.0504e-19 $X=19.58 $Y=2.995 $X2=0 $Y2=0
cc_5679 N_VPWR_M1237_d N_Z_c_9120_n 8.15553e-19 $X=20.5 $Y=2.995 $X2=0 $Y2=0
cc_5680 N_VPWR_c_7248_n N_Z_c_9120_n 0.0196216f $X=17.995 $Y=3.14 $X2=0 $Y2=0
cc_5681 N_VPWR_c_7250_n N_Z_c_9120_n 0.0222682f $X=18.935 $Y=3.14 $X2=0 $Y2=0
cc_5682 N_VPWR_c_7253_n N_Z_c_9120_n 0.0222682f $X=19.705 $Y=3.14 $X2=0 $Y2=0
cc_5683 N_VPWR_c_7255_n N_Z_c_9120_n 0.0196216f $X=20.645 $Y=3.14 $X2=0 $Y2=0
cc_5684 VPWR N_Z_c_9120_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5685 N_VPWR_M1042_d N_Z_c_9121_n 0.00213438f $X=23.495 $Y=1.485 $X2=0 $Y2=0
cc_5686 N_VPWR_M1089_d N_Z_c_9121_n 0.00236137f $X=24.415 $Y=1.485 $X2=0 $Y2=0
cc_5687 N_VPWR_M1289_d N_Z_c_9121_n 2.0504e-19 $X=25.355 $Y=1.485 $X2=0 $Y2=0
cc_5688 N_VPWR_M1158_d N_Z_c_9121_n 2.0504e-19 $X=26.355 $Y=1.485 $X2=0 $Y2=0
cc_5689 N_VPWR_M1194_d N_Z_c_9121_n 0.00236137f $X=27.275 $Y=1.485 $X2=0 $Y2=0
cc_5690 N_VPWR_M1319_d N_Z_c_9121_n 0.00213438f $X=28.215 $Y=1.485 $X2=0 $Y2=0
cc_5691 N_VPWR_c_7256_n N_Z_c_9121_n 0.0106064f $X=23.62 $Y=2 $X2=0 $Y2=0
cc_5692 N_VPWR_c_7258_n N_Z_c_9121_n 0.010348f $X=24.56 $Y=2 $X2=0 $Y2=0
cc_5693 N_VPWR_c_7260_n N_Z_c_9121_n 0.0274858f $X=25.5 $Y=1.66 $X2=0 $Y2=0
cc_5694 N_VPWR_c_7264_n N_Z_c_9121_n 0.0274858f $X=26.48 $Y=1.66 $X2=0 $Y2=0
cc_5695 N_VPWR_c_7268_n N_Z_c_9121_n 0.010348f $X=27.42 $Y=2 $X2=0 $Y2=0
cc_5696 N_VPWR_c_7271_n N_Z_c_9121_n 0.0106064f $X=28.36 $Y=2 $X2=0 $Y2=0
cc_5697 VPWR N_Z_c_9121_n 0.0762799f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5698 N_VPWR_M1052_d N_Z_c_9123_n 0.00213438f $X=23.495 $Y=2.955 $X2=0 $Y2=0
cc_5699 N_VPWR_M1101_d N_Z_c_9123_n 0.00236137f $X=24.415 $Y=2.955 $X2=0 $Y2=0
cc_5700 N_VPWR_M1297_d N_Z_c_9123_n 2.0504e-19 $X=25.355 $Y=2.955 $X2=0 $Y2=0
cc_5701 N_VPWR_M1006_s N_Z_c_9123_n 2.0504e-19 $X=26.355 $Y=2.955 $X2=0 $Y2=0
cc_5702 N_VPWR_M1165_s N_Z_c_9123_n 0.00236137f $X=27.275 $Y=2.955 $X2=0 $Y2=0
cc_5703 N_VPWR_M1277_s N_Z_c_9123_n 0.00213438f $X=28.215 $Y=2.955 $X2=0 $Y2=0
cc_5704 N_VPWR_c_7257_n N_Z_c_9123_n 0.0106064f $X=23.62 $Y=3.1 $X2=0 $Y2=0
cc_5705 N_VPWR_c_7259_n N_Z_c_9123_n 0.010348f $X=24.56 $Y=3.1 $X2=0 $Y2=0
cc_5706 N_VPWR_c_7262_n N_Z_c_9123_n 0.0274858f $X=25.5 $Y=3.1 $X2=0 $Y2=0
cc_5707 N_VPWR_c_7266_n N_Z_c_9123_n 0.0274858f $X=26.48 $Y=3.1 $X2=0 $Y2=0
cc_5708 N_VPWR_c_7269_n N_Z_c_9123_n 0.010348f $X=27.42 $Y=3.1 $X2=0 $Y2=0
cc_5709 N_VPWR_c_7272_n N_Z_c_9123_n 0.0106064f $X=28.36 $Y=3.1 $X2=0 $Y2=0
cc_5710 VPWR N_Z_c_9123_n 0.0762799f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5711 N_VPWR_M1016_d N_Z_c_9125_n 8.15553e-19 $X=31.21 $Y=1.625 $X2=0 $Y2=0
cc_5712 N_VPWR_M1095_d N_Z_c_9125_n 2.0504e-19 $X=32.13 $Y=1.625 $X2=0 $Y2=0
cc_5713 N_VPWR_M1022_s N_Z_c_9125_n 2.0504e-19 $X=32.92 $Y=1.625 $X2=0 $Y2=0
cc_5714 N_VPWR_M1256_s N_Z_c_9125_n 8.15553e-19 $X=33.84 $Y=1.625 $X2=0 $Y2=0
cc_5715 N_VPWR_c_7273_n N_Z_c_9125_n 0.0196216f $X=31.335 $Y=1.77 $X2=0 $Y2=0
cc_5716 N_VPWR_c_7275_n N_Z_c_9125_n 0.0222682f $X=32.275 $Y=1.77 $X2=0 $Y2=0
cc_5717 N_VPWR_c_7278_n N_Z_c_9125_n 0.0222682f $X=33.045 $Y=1.77 $X2=0 $Y2=0
cc_5718 N_VPWR_c_7280_n N_Z_c_9125_n 0.0196216f $X=33.985 $Y=1.77 $X2=0 $Y2=0
cc_5719 VPWR N_Z_c_9125_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5720 N_VPWR_M1120_d N_Z_c_9126_n 8.15553e-19 $X=31.21 $Y=2.995 $X2=0 $Y2=0
cc_5721 N_VPWR_M1201_d N_Z_c_9126_n 2.0504e-19 $X=32.13 $Y=2.995 $X2=0 $Y2=0
cc_5722 N_VPWR_M1034_d N_Z_c_9126_n 2.0504e-19 $X=32.92 $Y=2.995 $X2=0 $Y2=0
cc_5723 N_VPWR_M1130_d N_Z_c_9126_n 8.15553e-19 $X=33.84 $Y=2.995 $X2=0 $Y2=0
cc_5724 N_VPWR_c_7274_n N_Z_c_9126_n 0.0196216f $X=31.335 $Y=3.14 $X2=0 $Y2=0
cc_5725 N_VPWR_c_7276_n N_Z_c_9126_n 0.0222682f $X=32.275 $Y=3.14 $X2=0 $Y2=0
cc_5726 N_VPWR_c_7279_n N_Z_c_9126_n 0.0222682f $X=33.045 $Y=3.14 $X2=0 $Y2=0
cc_5727 N_VPWR_c_7281_n N_Z_c_9126_n 0.0196216f $X=33.985 $Y=3.14 $X2=0 $Y2=0
cc_5728 VPWR N_Z_c_9126_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5729 N_VPWR_M1088_d N_Z_c_9127_n 0.00213438f $X=36.835 $Y=1.485 $X2=0 $Y2=0
cc_5730 N_VPWR_M1183_d N_Z_c_9127_n 0.00236137f $X=37.755 $Y=1.485 $X2=0 $Y2=0
cc_5731 N_VPWR_M1255_d N_Z_c_9127_n 2.0504e-19 $X=38.695 $Y=1.485 $X2=0 $Y2=0
cc_5732 N_VPWR_M1099_d N_Z_c_9127_n 2.0504e-19 $X=39.235 $Y=1.485 $X2=0 $Y2=0
cc_5733 N_VPWR_M1176_d N_Z_c_9127_n 0.00236137f $X=40.155 $Y=1.485 $X2=0 $Y2=0
cc_5734 N_VPWR_M1282_d N_Z_c_9127_n 0.00213438f $X=41.095 $Y=1.485 $X2=0 $Y2=0
cc_5735 N_VPWR_c_7282_n N_Z_c_9127_n 0.0106064f $X=36.96 $Y=2 $X2=0 $Y2=0
cc_5736 N_VPWR_c_7284_n N_Z_c_9127_n 0.010348f $X=37.9 $Y=2 $X2=0 $Y2=0
cc_5737 N_VPWR_c_7286_n N_Z_c_9127_n 0.0276847f $X=38.84 $Y=1.66 $X2=0 $Y2=0
cc_5738 N_VPWR_c_7289_n N_Z_c_9127_n 0.0276847f $X=39.36 $Y=1.66 $X2=0 $Y2=0
cc_5739 N_VPWR_c_7291_n N_Z_c_9127_n 0.010348f $X=40.3 $Y=2 $X2=0 $Y2=0
cc_5740 N_VPWR_c_7294_n N_Z_c_9127_n 0.0106064f $X=41.24 $Y=2 $X2=0 $Y2=0
cc_5741 VPWR N_Z_c_9127_n 0.0537526f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5742 N_VPWR_M1102_d N_Z_c_9128_n 0.00213438f $X=36.835 $Y=2.955 $X2=0 $Y2=0
cc_5743 N_VPWR_M1186_d N_Z_c_9128_n 0.00236137f $X=37.755 $Y=2.955 $X2=0 $Y2=0
cc_5744 N_VPWR_M1264_d N_Z_c_9128_n 2.0504e-19 $X=38.695 $Y=2.955 $X2=0 $Y2=0
cc_5745 N_VPWR_M1109_d N_Z_c_9128_n 2.0504e-19 $X=39.235 $Y=2.955 $X2=0 $Y2=0
cc_5746 N_VPWR_M1184_d N_Z_c_9128_n 0.00236137f $X=40.155 $Y=2.955 $X2=0 $Y2=0
cc_5747 N_VPWR_M1293_d N_Z_c_9128_n 0.00213438f $X=41.095 $Y=2.955 $X2=0 $Y2=0
cc_5748 N_VPWR_c_7283_n N_Z_c_9128_n 0.0106064f $X=36.96 $Y=3.1 $X2=0 $Y2=0
cc_5749 N_VPWR_c_7285_n N_Z_c_9128_n 0.010348f $X=37.9 $Y=3.1 $X2=0 $Y2=0
cc_5750 N_VPWR_c_7287_n N_Z_c_9128_n 0.0276847f $X=38.84 $Y=3.1 $X2=0 $Y2=0
cc_5751 N_VPWR_c_7290_n N_Z_c_9128_n 0.0276847f $X=39.36 $Y=3.1 $X2=0 $Y2=0
cc_5752 N_VPWR_c_7292_n N_Z_c_9128_n 0.010348f $X=40.3 $Y=3.1 $X2=0 $Y2=0
cc_5753 N_VPWR_c_7295_n N_Z_c_9128_n 0.0106064f $X=41.24 $Y=3.1 $X2=0 $Y2=0
cc_5754 VPWR N_Z_c_9128_n 0.0537526f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5755 N_VPWR_M1015_d N_Z_c_9129_n 8.15553e-19 $X=44.09 $Y=1.625 $X2=0 $Y2=0
cc_5756 N_VPWR_M1063_d N_Z_c_9129_n 2.0504e-19 $X=45.01 $Y=1.625 $X2=0 $Y2=0
cc_5757 N_VPWR_M1142_d N_Z_c_9129_n 2.0504e-19 $X=45.8 $Y=1.625 $X2=0 $Y2=0
cc_5758 N_VPWR_M1185_d N_Z_c_9129_n 8.15553e-19 $X=46.72 $Y=1.625 $X2=0 $Y2=0
cc_5759 N_VPWR_c_7296_n N_Z_c_9129_n 0.0196216f $X=44.215 $Y=1.77 $X2=0 $Y2=0
cc_5760 N_VPWR_c_7298_n N_Z_c_9129_n 0.0222682f $X=45.155 $Y=1.77 $X2=0 $Y2=0
cc_5761 N_VPWR_c_7301_n N_Z_c_9129_n 0.0222682f $X=45.925 $Y=1.77 $X2=0 $Y2=0
cc_5762 N_VPWR_c_7303_n N_Z_c_9129_n 0.0196216f $X=46.865 $Y=1.77 $X2=0 $Y2=0
cc_5763 VPWR N_Z_c_9129_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5764 N_VPWR_M1124_d N_Z_c_9130_n 8.15553e-19 $X=44.09 $Y=2.995 $X2=0 $Y2=0
cc_5765 N_VPWR_M1170_d N_Z_c_9130_n 2.0504e-19 $X=45.01 $Y=2.995 $X2=0 $Y2=0
cc_5766 N_VPWR_M1233_d N_Z_c_9130_n 2.0504e-19 $X=45.8 $Y=2.995 $X2=0 $Y2=0
cc_5767 N_VPWR_M1279_d N_Z_c_9130_n 8.15553e-19 $X=46.72 $Y=2.995 $X2=0 $Y2=0
cc_5768 N_VPWR_c_7297_n N_Z_c_9130_n 0.0196216f $X=44.215 $Y=3.14 $X2=0 $Y2=0
cc_5769 N_VPWR_c_7299_n N_Z_c_9130_n 0.0222682f $X=45.155 $Y=3.14 $X2=0 $Y2=0
cc_5770 N_VPWR_c_7302_n N_Z_c_9130_n 0.0222682f $X=45.925 $Y=3.14 $X2=0 $Y2=0
cc_5771 N_VPWR_c_7304_n N_Z_c_9130_n 0.0196216f $X=46.865 $Y=3.14 $X2=0 $Y2=0
cc_5772 VPWR N_Z_c_9130_n 0.164379f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5773 VPWR N_Z_c_9131_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5774 N_VPWR_c_7351_n N_Z_c_9131_n 0.0123133f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_5775 N_VPWR_c_7311_n N_Z_c_9132_n 0.0123133f $X=4.95 $Y=2.72 $X2=0 $Y2=0
cc_5776 VPWR N_Z_c_9132_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5777 N_VPWR_c_7315_n N_Z_c_9133_n 0.0123133f $X=7.93 $Y=2.72 $X2=0 $Y2=0
cc_5778 VPWR N_Z_c_9133_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5779 N_VPWR_c_7318_n N_Z_c_9134_n 0.0123133f $X=10.605 $Y=2.72 $X2=0 $Y2=0
cc_5780 VPWR N_Z_c_9134_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5781 VPWR N_Z_c_9135_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5782 N_VPWR_c_7355_n N_Z_c_9135_n 0.0123133f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_5783 N_VPWR_c_7320_n N_Z_c_9136_n 0.0123133f $X=17.83 $Y=2.72 $X2=0 $Y2=0
cc_5784 VPWR N_Z_c_9136_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5785 N_VPWR_c_7324_n N_Z_c_9137_n 0.0123133f $X=20.81 $Y=2.72 $X2=0 $Y2=0
cc_5786 VPWR N_Z_c_9137_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5787 N_VPWR_c_7327_n N_Z_c_9138_n 0.0123133f $X=23.485 $Y=2.72 $X2=0 $Y2=0
cc_5788 VPWR N_Z_c_9138_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5789 VPWR N_Z_c_9139_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5790 N_VPWR_c_7362_n N_Z_c_9139_n 0.0123133f $X=28.75 $Y=2.72 $X2=0 $Y2=0
cc_5791 N_VPWR_c_7329_n N_Z_c_9140_n 0.0123133f $X=31.17 $Y=2.72 $X2=0 $Y2=0
cc_5792 VPWR N_Z_c_9140_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5793 N_VPWR_c_7333_n N_Z_c_9141_n 0.0123133f $X=34.15 $Y=2.72 $X2=0 $Y2=0
cc_5794 VPWR N_Z_c_9141_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5795 N_VPWR_c_7336_n N_Z_c_9142_n 0.0123133f $X=36.825 $Y=2.72 $X2=0 $Y2=0
cc_5796 VPWR N_Z_c_9142_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5797 VPWR N_Z_c_9143_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5798 N_VPWR_c_7366_n N_Z_c_9143_n 0.0123133f $X=41.63 $Y=2.72 $X2=0 $Y2=0
cc_5799 N_VPWR_c_7338_n N_Z_c_9144_n 0.0123133f $X=44.05 $Y=2.72 $X2=0 $Y2=0
cc_5800 VPWR N_Z_c_9144_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5801 N_VPWR_c_7342_n N_Z_c_9145_n 0.0123133f $X=47.03 $Y=2.72 $X2=0 $Y2=0
cc_5802 VPWR N_Z_c_9145_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5803 N_VPWR_c_7345_n N_Z_c_9146_n 0.0123133f $X=49.705 $Y=2.72 $X2=0 $Y2=0
cc_5804 VPWR N_Z_c_9146_n 0.0498209f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5805 VPWR N_A_1643_311#_M1002_d 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5806 VPWR N_A_1643_311#_M1134_d 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5807 N_VPWR_M1002_s N_A_1643_311#_c_10897_n 0.00715085f $X=10.615 $Y=1.485
+ $X2=0 $Y2=0
cc_5808 N_VPWR_c_7233_n N_A_1643_311#_c_10897_n 0.0152464f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5809 N_VPWR_M1038_s N_A_1643_311#_c_10919_n 0.00331615f $X=11.535 $Y=1.485
+ $X2=0 $Y2=0
cc_5810 N_VPWR_c_7235_n N_A_1643_311#_c_10919_n 0.0130979f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_5811 VPWR N_A_1643_311#_c_10906_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5812 N_VPWR_c_7231_n N_A_1643_311#_c_10948_n 0.00167067f $X=7.765 $Y=1.77
+ $X2=25.99 $Y2=1.87
cc_5813 VPWR N_A_1643_311#_c_10948_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5814 VPWR N_A_1643_311#_c_10908_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5815 VPWR N_A_1643_311#_c_10951_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5816 N_VPWR_c_7233_n N_A_1643_311#_c_10899_n 0.0156478f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5817 N_VPWR_c_7318_n N_A_1643_311#_c_10899_n 0.00115812f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_5818 VPWR N_A_1643_311#_c_10899_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5819 N_VPWR_c_7352_n N_A_1643_311#_c_10899_n 8.30334e-19 $X=11.545 $Y=2.72
+ $X2=0 $Y2=0
cc_5820 N_VPWR_c_7233_n N_A_1643_311#_c_10956_n 6.69936e-19 $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5821 VPWR N_A_1643_311#_c_10956_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5822 N_VPWR_c_7235_n N_A_1643_311#_c_10932_n 0.0153177f $X=11.68 $Y=2
+ $X2=25.99 $Y2=3.23
cc_5823 VPWR N_A_1643_311#_c_10932_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5824 N_VPWR_c_7352_n N_A_1643_311#_c_10932_n 8.30334e-19 $X=11.545 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5825 N_VPWR_c_7353_n N_A_1643_311#_c_10932_n 8.30334e-19 $X=12.485 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5826 N_VPWR_c_7233_n N_A_1643_311#_c_10962_n 6.68271e-19 $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5827 N_VPWR_c_7235_n N_A_1643_311#_c_10962_n 6.68271e-19 $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_5828 VPWR N_A_1643_311#_c_10962_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5829 N_VPWR_c_7233_n N_A_1643_311#_c_10934_n 0.0268237f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5830 N_VPWR_c_7235_n N_A_1643_311#_c_10934_n 0.0268237f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_5831 VPWR N_A_1643_311#_c_10934_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5832 N_VPWR_c_7352_n N_A_1643_311#_c_10934_n 0.0189467f $X=11.545 $Y=2.72
+ $X2=0 $Y2=0
cc_5833 N_VPWR_c_7235_n N_A_1643_311#_c_10969_n 6.68271e-19 $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_5834 N_VPWR_c_7237_n N_A_1643_311#_c_10969_n 0.00167228f $X=12.62 $Y=1.66
+ $X2=0 $Y2=0
cc_5835 VPWR N_A_1643_311#_c_10969_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5836 N_VPWR_c_7235_n N_A_1643_311#_c_10937_n 0.0268237f $X=11.68 $Y=2 $X2=0
+ $Y2=0
cc_5837 N_VPWR_c_7237_n N_A_1643_311#_c_10937_n 0.0318001f $X=12.62 $Y=1.66
+ $X2=0 $Y2=0
cc_5838 VPWR N_A_1643_311#_c_10937_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5839 N_VPWR_c_7353_n N_A_1643_311#_c_10937_n 0.0189467f $X=12.485 $Y=2.72
+ $X2=0 $Y2=0
cc_5840 N_VPWR_c_7231_n N_A_1643_311#_c_10900_n 0.0505494f $X=7.765 $Y=1.77
+ $X2=0 $Y2=0
cc_5841 N_VPWR_c_7315_n N_A_1643_311#_c_10900_n 0.0213652f $X=7.93 $Y=2.72 $X2=0
+ $Y2=0
cc_5842 VPWR N_A_1643_311#_c_10900_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5843 VPWR N_A_1643_311#_c_10901_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5844 N_VPWR_c_7233_n N_A_1643_311#_c_10902_n 0.0390576f $X=10.74 $Y=2 $X2=0
+ $Y2=0
cc_5845 N_VPWR_c_7318_n N_A_1643_311#_c_10902_n 0.0213652f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_5846 VPWR N_A_1643_311#_c_10902_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5847 VPWR N_A_1643_613#_M1011_d 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5848 VPWR N_A_1643_613#_M1148_d 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5849 N_VPWR_M1011_s N_A_1643_613#_c_11028_n 0.00715085f $X=10.615 $Y=2.955
+ $X2=0 $Y2=0
cc_5850 N_VPWR_c_7234_n N_A_1643_613#_c_11028_n 0.0152464f $X=10.74 $Y=3.1 $X2=0
+ $Y2=0
cc_5851 N_VPWR_M1051_s N_A_1643_613#_c_11050_n 0.00331615f $X=11.535 $Y=2.955
+ $X2=0 $Y2=0
cc_5852 N_VPWR_c_7236_n N_A_1643_613#_c_11050_n 0.0130979f $X=11.68 $Y=3.1 $X2=0
+ $Y2=0
cc_5853 VPWR N_A_1643_613#_c_11037_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5854 N_VPWR_c_7232_n N_A_1643_613#_c_11079_n 0.00167067f $X=7.765 $Y=3.14
+ $X2=25.99 $Y2=1.87
cc_5855 VPWR N_A_1643_613#_c_11079_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5856 VPWR N_A_1643_613#_c_11039_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5857 VPWR N_A_1643_613#_c_11082_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5858 N_VPWR_c_7234_n N_A_1643_613#_c_11030_n 0.0156478f $X=10.74 $Y=3.1 $X2=0
+ $Y2=0
cc_5859 N_VPWR_c_7318_n N_A_1643_613#_c_11030_n 0.00115812f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_5860 VPWR N_A_1643_613#_c_11030_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5861 N_VPWR_c_7352_n N_A_1643_613#_c_11030_n 8.30334e-19 $X=11.545 $Y=2.72
+ $X2=0 $Y2=0
cc_5862 N_VPWR_c_7234_n N_A_1643_613#_c_11087_n 6.69936e-19 $X=10.74 $Y=3.1
+ $X2=0 $Y2=0
cc_5863 VPWR N_A_1643_613#_c_11087_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5864 N_VPWR_c_7236_n N_A_1643_613#_c_11063_n 0.0153177f $X=11.68 $Y=3.1
+ $X2=25.99 $Y2=3.23
cc_5865 VPWR N_A_1643_613#_c_11063_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5866 N_VPWR_c_7352_n N_A_1643_613#_c_11063_n 8.30334e-19 $X=11.545 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5867 N_VPWR_c_7353_n N_A_1643_613#_c_11063_n 8.30334e-19 $X=12.485 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5868 N_VPWR_c_7234_n N_A_1643_613#_c_11093_n 6.68271e-19 $X=10.74 $Y=3.1
+ $X2=0 $Y2=0
cc_5869 N_VPWR_c_7236_n N_A_1643_613#_c_11093_n 6.68271e-19 $X=11.68 $Y=3.1
+ $X2=0 $Y2=0
cc_5870 VPWR N_A_1643_613#_c_11093_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5871 N_VPWR_c_7236_n N_A_1643_613#_c_11096_n 6.68271e-19 $X=11.68 $Y=3.1
+ $X2=0 $Y2=0
cc_5872 N_VPWR_c_7238_n N_A_1643_613#_c_11096_n 0.00167228f $X=12.62 $Y=3.1
+ $X2=0 $Y2=0
cc_5873 VPWR N_A_1643_613#_c_11096_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5874 N_VPWR_c_7232_n N_A_1643_613#_c_11031_n 0.0505494f $X=7.765 $Y=3.14
+ $X2=0 $Y2=0
cc_5875 N_VPWR_c_7315_n N_A_1643_613#_c_11031_n 0.0213652f $X=7.93 $Y=2.72 $X2=0
+ $Y2=0
cc_5876 VPWR N_A_1643_613#_c_11031_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5877 VPWR N_A_1643_613#_c_11032_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5878 N_VPWR_c_7234_n N_A_1643_613#_c_11033_n 0.0390576f $X=10.74 $Y=3.1 $X2=0
+ $Y2=0
cc_5879 N_VPWR_c_7318_n N_A_1643_613#_c_11033_n 0.0213652f $X=10.605 $Y=2.72
+ $X2=0 $Y2=0
cc_5880 VPWR N_A_1643_613#_c_11033_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5881 N_VPWR_c_7234_n N_A_1643_613#_c_11066_n 0.0268237f $X=10.74 $Y=3.1 $X2=0
+ $Y2=0
cc_5882 N_VPWR_c_7236_n N_A_1643_613#_c_11066_n 0.0268237f $X=11.68 $Y=3.1 $X2=0
+ $Y2=0
cc_5883 VPWR N_A_1643_613#_c_11066_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5884 N_VPWR_c_7352_n N_A_1643_613#_c_11066_n 0.0189467f $X=11.545 $Y=2.72
+ $X2=0 $Y2=0
cc_5885 N_VPWR_c_7236_n N_A_1643_613#_c_11069_n 0.0268237f $X=11.68 $Y=3.1 $X2=0
+ $Y2=0
cc_5886 N_VPWR_c_7238_n N_A_1643_613#_c_11069_n 0.0318001f $X=12.62 $Y=3.1 $X2=0
+ $Y2=0
cc_5887 VPWR N_A_1643_613#_c_11069_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5888 N_VPWR_c_7353_n N_A_1643_613#_c_11069_n 0.0189467f $X=12.485 $Y=2.72
+ $X2=0 $Y2=0
cc_5889 VPWR N_A_2693_297#_M1020_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_5890 VPWR N_A_2693_297#_M1157_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_5891 N_VPWR_M1067_s N_A_2693_297#_c_11164_n 0.00331615f $X=13.935 $Y=1.485
+ $X2=0 $Y2=0
cc_5892 N_VPWR_c_7242_n N_A_2693_297#_c_11164_n 0.0130979f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_5893 N_VPWR_M1301_s N_A_2693_297#_c_11159_n 0.00715085f $X=14.875 $Y=1.485
+ $X2=0 $Y2=0
cc_5894 N_VPWR_c_7245_n N_A_2693_297#_c_11159_n 0.0152464f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_5895 N_VPWR_c_7242_n N_A_2693_297#_c_11177_n 0.0153177f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_5896 N_VPWR_c_7244_n N_A_2693_297#_c_11177_n 8.30334e-19 $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5897 VPWR N_A_2693_297#_c_11177_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5898 N_VPWR_c_7354_n N_A_2693_297#_c_11177_n 8.30334e-19 $X=13.945 $Y=2.72
+ $X2=0 $Y2=0
cc_5899 N_VPWR_c_7240_n N_A_2693_297#_c_11212_n 0.00167228f $X=13.14 $Y=1.66
+ $X2=25.99 $Y2=1.87
cc_5900 N_VPWR_c_7242_n N_A_2693_297#_c_11212_n 6.68271e-19 $X=14.08 $Y=2
+ $X2=25.99 $Y2=1.87
cc_5901 VPWR N_A_2693_297#_c_11212_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5902 N_VPWR_c_7244_n N_A_2693_297#_c_11160_n 8.30334e-19 $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5903 N_VPWR_c_7245_n N_A_2693_297#_c_11160_n 0.0156478f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_5904 VPWR N_A_2693_297#_c_11160_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5905 N_VPWR_c_7355_n N_A_2693_297#_c_11160_n 0.00115812f $X=15.41 $Y=2.72
+ $X2=0 $Y2=0
cc_5906 N_VPWR_c_7242_n N_A_2693_297#_c_11219_n 6.68271e-19 $X=14.08 $Y=2
+ $X2=25.99 $Y2=2.21
cc_5907 N_VPWR_c_7245_n N_A_2693_297#_c_11219_n 6.68271e-19 $X=15.02 $Y=2
+ $X2=25.99 $Y2=2.21
cc_5908 VPWR N_A_2693_297#_c_11219_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5909 VPWR N_A_2693_297#_c_11188_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5910 N_VPWR_c_7245_n N_A_2693_297#_c_11223_n 6.69936e-19 $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_5911 VPWR N_A_2693_297#_c_11223_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5912 VPWR N_A_2693_297#_c_11190_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5913 VPWR N_A_2693_297#_c_11226_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5914 N_VPWR_c_7240_n N_A_2693_297#_c_11180_n 0.0318001f $X=13.14 $Y=1.66
+ $X2=25.99 $Y2=3.57
cc_5915 N_VPWR_c_7242_n N_A_2693_297#_c_11180_n 0.0268237f $X=14.08 $Y=2
+ $X2=25.99 $Y2=3.57
cc_5916 VPWR N_A_2693_297#_c_11180_n 0.00313104f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.57
cc_5917 N_VPWR_c_7354_n N_A_2693_297#_c_11180_n 0.0189467f $X=13.945 $Y=2.72
+ $X2=25.99 $Y2=3.57
cc_5918 N_VPWR_c_7242_n N_A_2693_297#_c_11183_n 0.0268237f $X=14.08 $Y=2 $X2=0
+ $Y2=0
cc_5919 N_VPWR_c_7244_n N_A_2693_297#_c_11183_n 0.0189467f $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5920 N_VPWR_c_7245_n N_A_2693_297#_c_11183_n 0.0268237f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_5921 VPWR N_A_2693_297#_c_11183_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5922 N_VPWR_c_7247_n N_A_2693_297#_c_11235_n 0.00167067f $X=17.995 $Y=1.77
+ $X2=0 $Y2=0
cc_5923 VPWR N_A_2693_297#_c_11235_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5924 N_VPWR_c_7245_n N_A_2693_297#_c_11161_n 0.0390576f $X=15.02 $Y=2 $X2=0
+ $Y2=0
cc_5925 VPWR N_A_2693_297#_c_11161_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5926 N_VPWR_c_7355_n N_A_2693_297#_c_11161_n 0.0213652f $X=15.41 $Y=2.72
+ $X2=0 $Y2=0
cc_5927 VPWR N_A_2693_297#_c_11162_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5928 N_VPWR_c_7247_n N_A_2693_297#_c_11163_n 0.0505494f $X=17.995 $Y=1.77
+ $X2=0 $Y2=0
cc_5929 N_VPWR_c_7320_n N_A_2693_297#_c_11163_n 0.0213652f $X=17.83 $Y=2.72
+ $X2=0 $Y2=0
cc_5930 VPWR N_A_2693_297#_c_11163_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5931 VPWR N_A_2693_591#_M1024_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_5932 VPWR N_A_2693_591#_M1164_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_5933 N_VPWR_M1076_s N_A_2693_591#_c_11292_n 0.00331615f $X=13.935 $Y=2.955
+ $X2=0 $Y2=0
cc_5934 N_VPWR_c_7243_n N_A_2693_591#_c_11292_n 0.0130979f $X=14.08 $Y=3.1 $X2=0
+ $Y2=0
cc_5935 N_VPWR_M1309_s N_A_2693_591#_c_11287_n 0.00715085f $X=14.875 $Y=2.955
+ $X2=0 $Y2=0
cc_5936 N_VPWR_c_7246_n N_A_2693_591#_c_11287_n 0.0152464f $X=15.02 $Y=3.1 $X2=0
+ $Y2=0
cc_5937 N_VPWR_c_7243_n N_A_2693_591#_c_11305_n 0.0153177f $X=14.08 $Y=3.1 $X2=0
+ $Y2=0
cc_5938 N_VPWR_c_7244_n N_A_2693_591#_c_11305_n 8.30334e-19 $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5939 VPWR N_A_2693_591#_c_11305_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5940 N_VPWR_c_7354_n N_A_2693_591#_c_11305_n 8.30334e-19 $X=13.945 $Y=2.72
+ $X2=0 $Y2=0
cc_5941 N_VPWR_c_7241_n N_A_2693_591#_c_11340_n 0.00167228f $X=13.14 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_5942 N_VPWR_c_7243_n N_A_2693_591#_c_11340_n 6.68271e-19 $X=14.08 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_5943 VPWR N_A_2693_591#_c_11340_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5944 N_VPWR_c_7244_n N_A_2693_591#_c_11288_n 8.30334e-19 $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5945 N_VPWR_c_7246_n N_A_2693_591#_c_11288_n 0.0156478f $X=15.02 $Y=3.1 $X2=0
+ $Y2=0
cc_5946 VPWR N_A_2693_591#_c_11288_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5947 N_VPWR_c_7355_n N_A_2693_591#_c_11288_n 0.00115812f $X=15.41 $Y=2.72
+ $X2=0 $Y2=0
cc_5948 N_VPWR_c_7243_n N_A_2693_591#_c_11347_n 6.68271e-19 $X=14.08 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_5949 N_VPWR_c_7246_n N_A_2693_591#_c_11347_n 6.68271e-19 $X=15.02 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_5950 VPWR N_A_2693_591#_c_11347_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5951 VPWR N_A_2693_591#_c_11316_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5952 N_VPWR_c_7246_n N_A_2693_591#_c_11351_n 6.69936e-19 $X=15.02 $Y=3.1
+ $X2=0 $Y2=0
cc_5953 VPWR N_A_2693_591#_c_11351_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5954 VPWR N_A_2693_591#_c_11318_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5955 VPWR N_A_2693_591#_c_11354_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5956 N_VPWR_c_7248_n N_A_2693_591#_c_11355_n 0.00167067f $X=17.995 $Y=3.14
+ $X2=0 $Y2=0
cc_5957 VPWR N_A_2693_591#_c_11355_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5958 N_VPWR_c_7241_n N_A_2693_591#_c_11308_n 0.0318001f $X=13.14 $Y=3.1 $X2=0
+ $Y2=0
cc_5959 N_VPWR_c_7243_n N_A_2693_591#_c_11308_n 0.0268237f $X=14.08 $Y=3.1 $X2=0
+ $Y2=0
cc_5960 VPWR N_A_2693_591#_c_11308_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5961 N_VPWR_c_7354_n N_A_2693_591#_c_11308_n 0.0189467f $X=13.945 $Y=2.72
+ $X2=0 $Y2=0
cc_5962 N_VPWR_c_7243_n N_A_2693_591#_c_11311_n 0.0268237f $X=14.08 $Y=3.1 $X2=0
+ $Y2=0
cc_5963 N_VPWR_c_7244_n N_A_2693_591#_c_11311_n 0.0189467f $X=14.885 $Y=2.72
+ $X2=0 $Y2=0
cc_5964 N_VPWR_c_7246_n N_A_2693_591#_c_11311_n 0.0268237f $X=15.02 $Y=3.1 $X2=0
+ $Y2=0
cc_5965 VPWR N_A_2693_591#_c_11311_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5966 N_VPWR_c_7246_n N_A_2693_591#_c_11289_n 0.0390576f $X=15.02 $Y=3.1 $X2=0
+ $Y2=0
cc_5967 VPWR N_A_2693_591#_c_11289_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5968 N_VPWR_c_7355_n N_A_2693_591#_c_11289_n 0.0213652f $X=15.41 $Y=2.72
+ $X2=0 $Y2=0
cc_5969 VPWR N_A_2693_591#_c_11290_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5970 N_VPWR_c_7248_n N_A_2693_591#_c_11291_n 0.0505494f $X=17.995 $Y=3.14
+ $X2=0 $Y2=0
cc_5971 N_VPWR_c_7320_n N_A_2693_591#_c_11291_n 0.0213652f $X=17.83 $Y=2.72
+ $X2=0 $Y2=0
cc_5972 VPWR N_A_2693_591#_c_11291_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5973 VPWR N_A_4219_311#_M1042_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5974 VPWR N_A_4219_311#_M1116_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5975 N_VPWR_M1042_d N_A_4219_311#_c_11415_n 0.00715085f $X=23.495 $Y=1.485
+ $X2=0 $Y2=0
cc_5976 N_VPWR_c_7256_n N_A_4219_311#_c_11415_n 0.0152464f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_5977 N_VPWR_M1089_d N_A_4219_311#_c_11437_n 0.00331615f $X=24.415 $Y=1.485
+ $X2=0 $Y2=0
cc_5978 N_VPWR_c_7258_n N_A_4219_311#_c_11437_n 0.0130979f $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_5979 VPWR N_A_4219_311#_c_11424_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5980 N_VPWR_c_7254_n N_A_4219_311#_c_11466_n 0.00167067f $X=20.645 $Y=1.77
+ $X2=25.99 $Y2=1.87
cc_5981 VPWR N_A_4219_311#_c_11466_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_5982 VPWR N_A_4219_311#_c_11426_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5983 VPWR N_A_4219_311#_c_11469_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_5984 N_VPWR_c_7256_n N_A_4219_311#_c_11417_n 0.0156478f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_5985 N_VPWR_c_7327_n N_A_4219_311#_c_11417_n 0.00115812f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_5986 VPWR N_A_4219_311#_c_11417_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5987 N_VPWR_c_7356_n N_A_4219_311#_c_11417_n 8.30334e-19 $X=24.425 $Y=2.72
+ $X2=0 $Y2=0
cc_5988 N_VPWR_c_7256_n N_A_4219_311#_c_11474_n 6.69936e-19 $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_5989 VPWR N_A_4219_311#_c_11474_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5990 N_VPWR_c_7258_n N_A_4219_311#_c_11450_n 0.0153177f $X=24.56 $Y=2
+ $X2=25.99 $Y2=3.23
cc_5991 VPWR N_A_4219_311#_c_11450_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_5992 N_VPWR_c_7356_n N_A_4219_311#_c_11450_n 8.30334e-19 $X=24.425 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5993 N_VPWR_c_7357_n N_A_4219_311#_c_11450_n 8.30334e-19 $X=25.365 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_5994 N_VPWR_c_7256_n N_A_4219_311#_c_11480_n 6.68271e-19 $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_5995 N_VPWR_c_7258_n N_A_4219_311#_c_11480_n 6.68271e-19 $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_5996 VPWR N_A_4219_311#_c_11480_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_5997 N_VPWR_c_7256_n N_A_4219_311#_c_11452_n 0.0268237f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_5998 N_VPWR_c_7258_n N_A_4219_311#_c_11452_n 0.0268237f $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_5999 VPWR N_A_4219_311#_c_11452_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6000 N_VPWR_c_7356_n N_A_4219_311#_c_11452_n 0.0189467f $X=24.425 $Y=2.72
+ $X2=0 $Y2=0
cc_6001 N_VPWR_c_7258_n N_A_4219_311#_c_11487_n 6.68271e-19 $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_6002 N_VPWR_c_7260_n N_A_4219_311#_c_11487_n 0.00167228f $X=25.5 $Y=1.66
+ $X2=0 $Y2=0
cc_6003 VPWR N_A_4219_311#_c_11487_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6004 N_VPWR_c_7258_n N_A_4219_311#_c_11455_n 0.0268237f $X=24.56 $Y=2 $X2=0
+ $Y2=0
cc_6005 N_VPWR_c_7260_n N_A_4219_311#_c_11455_n 0.0318001f $X=25.5 $Y=1.66 $X2=0
+ $Y2=0
cc_6006 VPWR N_A_4219_311#_c_11455_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6007 N_VPWR_c_7357_n N_A_4219_311#_c_11455_n 0.0189467f $X=25.365 $Y=2.72
+ $X2=0 $Y2=0
cc_6008 N_VPWR_c_7254_n N_A_4219_311#_c_11418_n 0.0505494f $X=20.645 $Y=1.77
+ $X2=0 $Y2=0
cc_6009 N_VPWR_c_7324_n N_A_4219_311#_c_11418_n 0.0213652f $X=20.81 $Y=2.72
+ $X2=0 $Y2=0
cc_6010 VPWR N_A_4219_311#_c_11418_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6011 VPWR N_A_4219_311#_c_11419_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6012 N_VPWR_c_7256_n N_A_4219_311#_c_11420_n 0.0390576f $X=23.62 $Y=2 $X2=0
+ $Y2=0
cc_6013 N_VPWR_c_7327_n N_A_4219_311#_c_11420_n 0.0213652f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_6014 VPWR N_A_4219_311#_c_11420_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6015 VPWR N_A_4219_613#_M1052_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6016 VPWR N_A_4219_613#_M1129_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6017 N_VPWR_M1052_d N_A_4219_613#_c_11546_n 0.00715085f $X=23.495 $Y=2.955
+ $X2=0 $Y2=0
cc_6018 N_VPWR_c_7257_n N_A_4219_613#_c_11546_n 0.0152464f $X=23.62 $Y=3.1 $X2=0
+ $Y2=0
cc_6019 N_VPWR_M1101_d N_A_4219_613#_c_11568_n 0.00331615f $X=24.415 $Y=2.955
+ $X2=0 $Y2=0
cc_6020 N_VPWR_c_7259_n N_A_4219_613#_c_11568_n 0.0130979f $X=24.56 $Y=3.1 $X2=0
+ $Y2=0
cc_6021 VPWR N_A_4219_613#_c_11555_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6022 N_VPWR_c_7255_n N_A_4219_613#_c_11597_n 0.00167067f $X=20.645 $Y=3.14
+ $X2=25.99 $Y2=1.87
cc_6023 VPWR N_A_4219_613#_c_11597_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6024 VPWR N_A_4219_613#_c_11557_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6025 VPWR N_A_4219_613#_c_11600_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6026 N_VPWR_c_7257_n N_A_4219_613#_c_11548_n 0.0156478f $X=23.62 $Y=3.1 $X2=0
+ $Y2=0
cc_6027 N_VPWR_c_7327_n N_A_4219_613#_c_11548_n 0.00115812f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_6028 VPWR N_A_4219_613#_c_11548_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6029 N_VPWR_c_7356_n N_A_4219_613#_c_11548_n 8.30334e-19 $X=24.425 $Y=2.72
+ $X2=0 $Y2=0
cc_6030 N_VPWR_c_7257_n N_A_4219_613#_c_11605_n 6.69936e-19 $X=23.62 $Y=3.1
+ $X2=0 $Y2=0
cc_6031 VPWR N_A_4219_613#_c_11605_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6032 N_VPWR_c_7259_n N_A_4219_613#_c_11581_n 0.0153177f $X=24.56 $Y=3.1
+ $X2=25.99 $Y2=3.23
cc_6033 VPWR N_A_4219_613#_c_11581_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6034 N_VPWR_c_7356_n N_A_4219_613#_c_11581_n 8.30334e-19 $X=24.425 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6035 N_VPWR_c_7357_n N_A_4219_613#_c_11581_n 8.30334e-19 $X=25.365 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6036 N_VPWR_c_7257_n N_A_4219_613#_c_11611_n 6.68271e-19 $X=23.62 $Y=3.1
+ $X2=0 $Y2=0
cc_6037 N_VPWR_c_7259_n N_A_4219_613#_c_11611_n 6.68271e-19 $X=24.56 $Y=3.1
+ $X2=0 $Y2=0
cc_6038 VPWR N_A_4219_613#_c_11611_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6039 N_VPWR_c_7259_n N_A_4219_613#_c_11614_n 6.68271e-19 $X=24.56 $Y=3.1
+ $X2=0 $Y2=0
cc_6040 N_VPWR_c_7262_n N_A_4219_613#_c_11614_n 0.00167228f $X=25.5 $Y=3.1 $X2=0
+ $Y2=0
cc_6041 VPWR N_A_4219_613#_c_11614_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6042 N_VPWR_c_7255_n N_A_4219_613#_c_11549_n 0.0505494f $X=20.645 $Y=3.14
+ $X2=0 $Y2=0
cc_6043 N_VPWR_c_7324_n N_A_4219_613#_c_11549_n 0.0213652f $X=20.81 $Y=2.72
+ $X2=0 $Y2=0
cc_6044 VPWR N_A_4219_613#_c_11549_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6045 VPWR N_A_4219_613#_c_11550_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6046 N_VPWR_c_7257_n N_A_4219_613#_c_11551_n 0.0390576f $X=23.62 $Y=3.1 $X2=0
+ $Y2=0
cc_6047 N_VPWR_c_7327_n N_A_4219_613#_c_11551_n 0.0213652f $X=23.485 $Y=2.72
+ $X2=0 $Y2=0
cc_6048 VPWR N_A_4219_613#_c_11551_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6049 N_VPWR_c_7257_n N_A_4219_613#_c_11584_n 0.0268237f $X=23.62 $Y=3.1 $X2=0
+ $Y2=0
cc_6050 N_VPWR_c_7259_n N_A_4219_613#_c_11584_n 0.0268237f $X=24.56 $Y=3.1 $X2=0
+ $Y2=0
cc_6051 VPWR N_A_4219_613#_c_11584_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6052 N_VPWR_c_7356_n N_A_4219_613#_c_11584_n 0.0189467f $X=24.425 $Y=2.72
+ $X2=0 $Y2=0
cc_6053 N_VPWR_c_7259_n N_A_4219_613#_c_11587_n 0.0268237f $X=24.56 $Y=3.1 $X2=0
+ $Y2=0
cc_6054 N_VPWR_c_7262_n N_A_4219_613#_c_11587_n 0.0318001f $X=25.5 $Y=3.1 $X2=0
+ $Y2=0
cc_6055 VPWR N_A_4219_613#_c_11587_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6056 N_VPWR_c_7357_n N_A_4219_613#_c_11587_n 0.0189467f $X=25.365 $Y=2.72
+ $X2=0 $Y2=0
cc_6057 VPWR N_A_5361_297#_M1158_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_6058 VPWR N_A_5361_297#_M1265_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_6059 N_VPWR_M1194_d N_A_5361_297#_c_11682_n 0.00331615f $X=27.275 $Y=1.485
+ $X2=0 $Y2=0
cc_6060 N_VPWR_c_7268_n N_A_5361_297#_c_11682_n 0.0130979f $X=27.42 $Y=2 $X2=0
+ $Y2=0
cc_6061 N_VPWR_M1319_d N_A_5361_297#_c_11677_n 0.00715085f $X=28.215 $Y=1.485
+ $X2=0 $Y2=0
cc_6062 N_VPWR_c_7271_n N_A_5361_297#_c_11677_n 0.0152464f $X=28.36 $Y=2 $X2=0
+ $Y2=0
cc_6063 N_VPWR_c_7268_n N_A_5361_297#_c_11695_n 0.0153177f $X=27.42 $Y=2 $X2=0
+ $Y2=0
cc_6064 N_VPWR_c_7270_n N_A_5361_297#_c_11695_n 8.30334e-19 $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6065 VPWR N_A_5361_297#_c_11695_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6066 N_VPWR_c_7361_n N_A_5361_297#_c_11695_n 8.30334e-19 $X=27.285 $Y=2.72
+ $X2=0 $Y2=0
cc_6067 N_VPWR_c_7264_n N_A_5361_297#_c_11730_n 0.00167228f $X=26.48 $Y=1.66
+ $X2=25.99 $Y2=1.87
cc_6068 N_VPWR_c_7268_n N_A_5361_297#_c_11730_n 6.68271e-19 $X=27.42 $Y=2
+ $X2=25.99 $Y2=1.87
cc_6069 VPWR N_A_5361_297#_c_11730_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6070 N_VPWR_c_7270_n N_A_5361_297#_c_11678_n 8.30334e-19 $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6071 N_VPWR_c_7271_n N_A_5361_297#_c_11678_n 0.0156478f $X=28.36 $Y=2 $X2=0
+ $Y2=0
cc_6072 VPWR N_A_5361_297#_c_11678_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6073 N_VPWR_c_7362_n N_A_5361_297#_c_11678_n 0.00115812f $X=28.75 $Y=2.72
+ $X2=0 $Y2=0
cc_6074 N_VPWR_c_7268_n N_A_5361_297#_c_11737_n 6.68271e-19 $X=27.42 $Y=2
+ $X2=25.99 $Y2=2.21
cc_6075 N_VPWR_c_7271_n N_A_5361_297#_c_11737_n 6.68271e-19 $X=28.36 $Y=2
+ $X2=25.99 $Y2=2.21
cc_6076 VPWR N_A_5361_297#_c_11737_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6077 VPWR N_A_5361_297#_c_11706_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6078 N_VPWR_c_7271_n N_A_5361_297#_c_11741_n 6.69936e-19 $X=28.36 $Y=2 $X2=0
+ $Y2=0
cc_6079 VPWR N_A_5361_297#_c_11741_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6080 VPWR N_A_5361_297#_c_11708_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6081 VPWR N_A_5361_297#_c_11744_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6082 N_VPWR_c_7264_n N_A_5361_297#_c_11698_n 0.0318001f $X=26.48 $Y=1.66
+ $X2=25.99 $Y2=3.57
cc_6083 N_VPWR_c_7268_n N_A_5361_297#_c_11698_n 0.0268237f $X=27.42 $Y=2
+ $X2=25.99 $Y2=3.57
cc_6084 VPWR N_A_5361_297#_c_11698_n 0.00313104f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.57
cc_6085 N_VPWR_c_7361_n N_A_5361_297#_c_11698_n 0.0189467f $X=27.285 $Y=2.72
+ $X2=25.99 $Y2=3.57
cc_6086 N_VPWR_c_7268_n N_A_5361_297#_c_11701_n 0.0268237f $X=27.42 $Y=2 $X2=0
+ $Y2=0
cc_6087 N_VPWR_c_7270_n N_A_5361_297#_c_11701_n 0.0189467f $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6088 N_VPWR_c_7271_n N_A_5361_297#_c_11701_n 0.0268237f $X=28.36 $Y=2 $X2=0
+ $Y2=0
cc_6089 VPWR N_A_5361_297#_c_11701_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6090 N_VPWR_c_7273_n N_A_5361_297#_c_11753_n 0.00167067f $X=31.335 $Y=1.77
+ $X2=0 $Y2=0
cc_6091 VPWR N_A_5361_297#_c_11753_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6092 N_VPWR_c_7271_n N_A_5361_297#_c_11679_n 0.0390576f $X=28.36 $Y=2 $X2=0
+ $Y2=0
cc_6093 VPWR N_A_5361_297#_c_11679_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6094 N_VPWR_c_7362_n N_A_5361_297#_c_11679_n 0.0213652f $X=28.75 $Y=2.72
+ $X2=0 $Y2=0
cc_6095 VPWR N_A_5361_297#_c_11680_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6096 N_VPWR_c_7273_n N_A_5361_297#_c_11681_n 0.0505494f $X=31.335 $Y=1.77
+ $X2=0 $Y2=0
cc_6097 N_VPWR_c_7329_n N_A_5361_297#_c_11681_n 0.0213652f $X=31.17 $Y=2.72
+ $X2=0 $Y2=0
cc_6098 VPWR N_A_5361_297#_c_11681_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6099 VPWR N_A_5361_591#_M1006_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_6100 VPWR N_A_5361_591#_M1203_d 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_6101 N_VPWR_M1165_s N_A_5361_591#_c_11810_n 0.00331615f $X=27.275 $Y=2.955
+ $X2=0 $Y2=0
cc_6102 N_VPWR_c_7269_n N_A_5361_591#_c_11810_n 0.0130979f $X=27.42 $Y=3.1 $X2=0
+ $Y2=0
cc_6103 N_VPWR_M1277_s N_A_5361_591#_c_11805_n 0.00715085f $X=28.215 $Y=2.955
+ $X2=0 $Y2=0
cc_6104 N_VPWR_c_7272_n N_A_5361_591#_c_11805_n 0.0152464f $X=28.36 $Y=3.1 $X2=0
+ $Y2=0
cc_6105 N_VPWR_c_7269_n N_A_5361_591#_c_11823_n 0.0153177f $X=27.42 $Y=3.1 $X2=0
+ $Y2=0
cc_6106 N_VPWR_c_7270_n N_A_5361_591#_c_11823_n 8.30334e-19 $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6107 VPWR N_A_5361_591#_c_11823_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6108 N_VPWR_c_7361_n N_A_5361_591#_c_11823_n 8.30334e-19 $X=27.285 $Y=2.72
+ $X2=0 $Y2=0
cc_6109 N_VPWR_c_7266_n N_A_5361_591#_c_11858_n 0.00167228f $X=26.48 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_6110 N_VPWR_c_7269_n N_A_5361_591#_c_11858_n 6.68271e-19 $X=27.42 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_6111 VPWR N_A_5361_591#_c_11858_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6112 N_VPWR_c_7270_n N_A_5361_591#_c_11806_n 8.30334e-19 $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6113 N_VPWR_c_7272_n N_A_5361_591#_c_11806_n 0.0156478f $X=28.36 $Y=3.1 $X2=0
+ $Y2=0
cc_6114 VPWR N_A_5361_591#_c_11806_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6115 N_VPWR_c_7362_n N_A_5361_591#_c_11806_n 0.00115812f $X=28.75 $Y=2.72
+ $X2=0 $Y2=0
cc_6116 N_VPWR_c_7269_n N_A_5361_591#_c_11865_n 6.68271e-19 $X=27.42 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_6117 N_VPWR_c_7272_n N_A_5361_591#_c_11865_n 6.68271e-19 $X=28.36 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_6118 VPWR N_A_5361_591#_c_11865_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6119 VPWR N_A_5361_591#_c_11834_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6120 N_VPWR_c_7272_n N_A_5361_591#_c_11869_n 6.69936e-19 $X=28.36 $Y=3.1
+ $X2=0 $Y2=0
cc_6121 VPWR N_A_5361_591#_c_11869_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6122 VPWR N_A_5361_591#_c_11836_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6123 VPWR N_A_5361_591#_c_11872_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6124 N_VPWR_c_7274_n N_A_5361_591#_c_11873_n 0.00167067f $X=31.335 $Y=3.14
+ $X2=0 $Y2=0
cc_6125 VPWR N_A_5361_591#_c_11873_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6126 N_VPWR_c_7266_n N_A_5361_591#_c_11826_n 0.0318001f $X=26.48 $Y=3.1 $X2=0
+ $Y2=0
cc_6127 N_VPWR_c_7269_n N_A_5361_591#_c_11826_n 0.0268237f $X=27.42 $Y=3.1 $X2=0
+ $Y2=0
cc_6128 VPWR N_A_5361_591#_c_11826_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6129 N_VPWR_c_7361_n N_A_5361_591#_c_11826_n 0.0189467f $X=27.285 $Y=2.72
+ $X2=0 $Y2=0
cc_6130 N_VPWR_c_7269_n N_A_5361_591#_c_11829_n 0.0268237f $X=27.42 $Y=3.1 $X2=0
+ $Y2=0
cc_6131 N_VPWR_c_7270_n N_A_5361_591#_c_11829_n 0.0189467f $X=28.225 $Y=2.72
+ $X2=0 $Y2=0
cc_6132 N_VPWR_c_7272_n N_A_5361_591#_c_11829_n 0.0268237f $X=28.36 $Y=3.1 $X2=0
+ $Y2=0
cc_6133 VPWR N_A_5361_591#_c_11829_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6134 N_VPWR_c_7272_n N_A_5361_591#_c_11807_n 0.0390576f $X=28.36 $Y=3.1 $X2=0
+ $Y2=0
cc_6135 VPWR N_A_5361_591#_c_11807_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6136 N_VPWR_c_7362_n N_A_5361_591#_c_11807_n 0.0213652f $X=28.75 $Y=2.72
+ $X2=0 $Y2=0
cc_6137 VPWR N_A_5361_591#_c_11808_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6138 N_VPWR_c_7274_n N_A_5361_591#_c_11809_n 0.0505494f $X=31.335 $Y=3.14
+ $X2=0 $Y2=0
cc_6139 N_VPWR_c_7329_n N_A_5361_591#_c_11809_n 0.0213652f $X=31.17 $Y=2.72
+ $X2=0 $Y2=0
cc_6140 VPWR N_A_5361_591#_c_11809_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6141 VPWR N_A_6887_311#_M1088_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6142 VPWR N_A_6887_311#_M1217_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6143 N_VPWR_M1088_d N_A_6887_311#_c_11933_n 0.00715085f $X=36.835 $Y=1.485
+ $X2=0 $Y2=0
cc_6144 N_VPWR_c_7282_n N_A_6887_311#_c_11933_n 0.0152464f $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6145 N_VPWR_M1183_d N_A_6887_311#_c_11955_n 0.00331615f $X=37.755 $Y=1.485
+ $X2=0 $Y2=0
cc_6146 N_VPWR_c_7284_n N_A_6887_311#_c_11955_n 0.0130979f $X=37.9 $Y=2 $X2=0
+ $Y2=0
cc_6147 VPWR N_A_6887_311#_c_11942_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6148 N_VPWR_c_7280_n N_A_6887_311#_c_11984_n 0.00167067f $X=33.985 $Y=1.77
+ $X2=25.99 $Y2=1.87
cc_6149 VPWR N_A_6887_311#_c_11984_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6150 VPWR N_A_6887_311#_c_11944_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6151 VPWR N_A_6887_311#_c_11987_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6152 N_VPWR_c_7282_n N_A_6887_311#_c_11935_n 0.0156478f $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6153 N_VPWR_c_7336_n N_A_6887_311#_c_11935_n 0.00115812f $X=36.825 $Y=2.72
+ $X2=0 $Y2=0
cc_6154 VPWR N_A_6887_311#_c_11935_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6155 N_VPWR_c_7363_n N_A_6887_311#_c_11935_n 8.30334e-19 $X=37.765 $Y=2.72
+ $X2=0 $Y2=0
cc_6156 N_VPWR_c_7282_n N_A_6887_311#_c_11992_n 6.69936e-19 $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6157 VPWR N_A_6887_311#_c_11992_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6158 N_VPWR_c_7284_n N_A_6887_311#_c_11968_n 0.0153177f $X=37.9 $Y=2
+ $X2=25.99 $Y2=3.23
cc_6159 VPWR N_A_6887_311#_c_11968_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6160 N_VPWR_c_7363_n N_A_6887_311#_c_11968_n 8.30334e-19 $X=37.765 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6161 N_VPWR_c_7364_n N_A_6887_311#_c_11968_n 8.30334e-19 $X=38.705 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6162 N_VPWR_c_7282_n N_A_6887_311#_c_11998_n 6.68271e-19 $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6163 N_VPWR_c_7284_n N_A_6887_311#_c_11998_n 6.68271e-19 $X=37.9 $Y=2 $X2=0
+ $Y2=0
cc_6164 VPWR N_A_6887_311#_c_11998_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6165 N_VPWR_c_7282_n N_A_6887_311#_c_11970_n 0.0268237f $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6166 N_VPWR_c_7284_n N_A_6887_311#_c_11970_n 0.0268237f $X=37.9 $Y=2 $X2=0
+ $Y2=0
cc_6167 VPWR N_A_6887_311#_c_11970_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6168 N_VPWR_c_7363_n N_A_6887_311#_c_11970_n 0.0189467f $X=37.765 $Y=2.72
+ $X2=0 $Y2=0
cc_6169 N_VPWR_c_7284_n N_A_6887_311#_c_12005_n 6.68271e-19 $X=37.9 $Y=2 $X2=0
+ $Y2=0
cc_6170 N_VPWR_c_7286_n N_A_6887_311#_c_12005_n 0.00167228f $X=38.84 $Y=1.66
+ $X2=0 $Y2=0
cc_6171 VPWR N_A_6887_311#_c_12005_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6172 N_VPWR_c_7284_n N_A_6887_311#_c_11973_n 0.0268237f $X=37.9 $Y=2 $X2=0
+ $Y2=0
cc_6173 N_VPWR_c_7286_n N_A_6887_311#_c_11973_n 0.0318001f $X=38.84 $Y=1.66
+ $X2=0 $Y2=0
cc_6174 VPWR N_A_6887_311#_c_11973_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6175 N_VPWR_c_7364_n N_A_6887_311#_c_11973_n 0.0189467f $X=38.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6176 N_VPWR_c_7280_n N_A_6887_311#_c_11936_n 0.0505494f $X=33.985 $Y=1.77
+ $X2=0 $Y2=0
cc_6177 N_VPWR_c_7333_n N_A_6887_311#_c_11936_n 0.0213652f $X=34.15 $Y=2.72
+ $X2=0 $Y2=0
cc_6178 VPWR N_A_6887_311#_c_11936_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6179 VPWR N_A_6887_311#_c_11937_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6180 N_VPWR_c_7282_n N_A_6887_311#_c_11938_n 0.0390576f $X=36.96 $Y=2 $X2=0
+ $Y2=0
cc_6181 N_VPWR_c_7336_n N_A_6887_311#_c_11938_n 0.0213652f $X=36.825 $Y=2.72
+ $X2=0 $Y2=0
cc_6182 VPWR N_A_6887_311#_c_11938_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6183 VPWR N_A_6887_613#_M1102_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6184 VPWR N_A_6887_613#_M1224_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6185 N_VPWR_M1102_d N_A_6887_613#_c_12064_n 0.00715085f $X=36.835 $Y=2.955
+ $X2=0 $Y2=0
cc_6186 N_VPWR_c_7283_n N_A_6887_613#_c_12064_n 0.0152464f $X=36.96 $Y=3.1 $X2=0
+ $Y2=0
cc_6187 N_VPWR_M1186_d N_A_6887_613#_c_12086_n 0.00331615f $X=37.755 $Y=2.955
+ $X2=0 $Y2=0
cc_6188 N_VPWR_c_7285_n N_A_6887_613#_c_12086_n 0.0130979f $X=37.9 $Y=3.1 $X2=0
+ $Y2=0
cc_6189 VPWR N_A_6887_613#_c_12073_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6190 N_VPWR_c_7281_n N_A_6887_613#_c_12115_n 0.00167067f $X=33.985 $Y=3.14
+ $X2=25.99 $Y2=1.87
cc_6191 VPWR N_A_6887_613#_c_12115_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6192 VPWR N_A_6887_613#_c_12075_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6193 VPWR N_A_6887_613#_c_12118_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6194 N_VPWR_c_7283_n N_A_6887_613#_c_12066_n 0.0156478f $X=36.96 $Y=3.1 $X2=0
+ $Y2=0
cc_6195 N_VPWR_c_7336_n N_A_6887_613#_c_12066_n 0.00115812f $X=36.825 $Y=2.72
+ $X2=0 $Y2=0
cc_6196 VPWR N_A_6887_613#_c_12066_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6197 N_VPWR_c_7363_n N_A_6887_613#_c_12066_n 8.30334e-19 $X=37.765 $Y=2.72
+ $X2=0 $Y2=0
cc_6198 N_VPWR_c_7283_n N_A_6887_613#_c_12123_n 6.69936e-19 $X=36.96 $Y=3.1
+ $X2=0 $Y2=0
cc_6199 VPWR N_A_6887_613#_c_12123_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6200 N_VPWR_c_7285_n N_A_6887_613#_c_12099_n 0.0153177f $X=37.9 $Y=3.1
+ $X2=25.99 $Y2=3.23
cc_6201 VPWR N_A_6887_613#_c_12099_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6202 N_VPWR_c_7363_n N_A_6887_613#_c_12099_n 8.30334e-19 $X=37.765 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6203 N_VPWR_c_7364_n N_A_6887_613#_c_12099_n 8.30334e-19 $X=38.705 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6204 N_VPWR_c_7283_n N_A_6887_613#_c_12129_n 6.68271e-19 $X=36.96 $Y=3.1
+ $X2=0 $Y2=0
cc_6205 N_VPWR_c_7285_n N_A_6887_613#_c_12129_n 6.68271e-19 $X=37.9 $Y=3.1 $X2=0
+ $Y2=0
cc_6206 VPWR N_A_6887_613#_c_12129_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6207 N_VPWR_c_7285_n N_A_6887_613#_c_12132_n 6.68271e-19 $X=37.9 $Y=3.1 $X2=0
+ $Y2=0
cc_6208 N_VPWR_c_7287_n N_A_6887_613#_c_12132_n 0.00167228f $X=38.84 $Y=3.1
+ $X2=0 $Y2=0
cc_6209 VPWR N_A_6887_613#_c_12132_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6210 N_VPWR_c_7281_n N_A_6887_613#_c_12067_n 0.0505494f $X=33.985 $Y=3.14
+ $X2=0 $Y2=0
cc_6211 N_VPWR_c_7333_n N_A_6887_613#_c_12067_n 0.0213652f $X=34.15 $Y=2.72
+ $X2=0 $Y2=0
cc_6212 VPWR N_A_6887_613#_c_12067_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6213 VPWR N_A_6887_613#_c_12068_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6214 N_VPWR_c_7283_n N_A_6887_613#_c_12069_n 0.0390576f $X=36.96 $Y=3.1 $X2=0
+ $Y2=0
cc_6215 N_VPWR_c_7336_n N_A_6887_613#_c_12069_n 0.0213652f $X=36.825 $Y=2.72
+ $X2=0 $Y2=0
cc_6216 VPWR N_A_6887_613#_c_12069_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6217 N_VPWR_c_7283_n N_A_6887_613#_c_12102_n 0.0268237f $X=36.96 $Y=3.1 $X2=0
+ $Y2=0
cc_6218 N_VPWR_c_7285_n N_A_6887_613#_c_12102_n 0.0268237f $X=37.9 $Y=3.1 $X2=0
+ $Y2=0
cc_6219 VPWR N_A_6887_613#_c_12102_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6220 N_VPWR_c_7363_n N_A_6887_613#_c_12102_n 0.0189467f $X=37.765 $Y=2.72
+ $X2=0 $Y2=0
cc_6221 N_VPWR_c_7285_n N_A_6887_613#_c_12105_n 0.0268237f $X=37.9 $Y=3.1 $X2=0
+ $Y2=0
cc_6222 N_VPWR_c_7287_n N_A_6887_613#_c_12105_n 0.0318001f $X=38.84 $Y=3.1 $X2=0
+ $Y2=0
cc_6223 VPWR N_A_6887_613#_c_12105_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6224 N_VPWR_c_7364_n N_A_6887_613#_c_12105_n 0.0189467f $X=38.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6225 VPWR N_A_7937_297#_M1099_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_6226 VPWR N_A_7937_297#_M1246_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_6227 N_VPWR_M1176_d N_A_7937_297#_c_12200_n 0.00331615f $X=40.155 $Y=1.485
+ $X2=0 $Y2=0
cc_6228 N_VPWR_c_7291_n N_A_7937_297#_c_12200_n 0.0130979f $X=40.3 $Y=2 $X2=0
+ $Y2=0
cc_6229 N_VPWR_M1282_d N_A_7937_297#_c_12195_n 0.00715085f $X=41.095 $Y=1.485
+ $X2=0 $Y2=0
cc_6230 N_VPWR_c_7294_n N_A_7937_297#_c_12195_n 0.0152464f $X=41.24 $Y=2 $X2=0
+ $Y2=0
cc_6231 N_VPWR_c_7291_n N_A_7937_297#_c_12213_n 0.0153177f $X=40.3 $Y=2 $X2=0
+ $Y2=0
cc_6232 N_VPWR_c_7293_n N_A_7937_297#_c_12213_n 8.30334e-19 $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6233 VPWR N_A_7937_297#_c_12213_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6234 N_VPWR_c_7365_n N_A_7937_297#_c_12213_n 8.30334e-19 $X=40.165 $Y=2.72
+ $X2=0 $Y2=0
cc_6235 N_VPWR_c_7289_n N_A_7937_297#_c_12248_n 0.00167228f $X=39.36 $Y=1.66
+ $X2=25.99 $Y2=1.87
cc_6236 N_VPWR_c_7291_n N_A_7937_297#_c_12248_n 6.68271e-19 $X=40.3 $Y=2
+ $X2=25.99 $Y2=1.87
cc_6237 VPWR N_A_7937_297#_c_12248_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6238 N_VPWR_c_7293_n N_A_7937_297#_c_12196_n 8.30334e-19 $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6239 N_VPWR_c_7294_n N_A_7937_297#_c_12196_n 0.0156478f $X=41.24 $Y=2 $X2=0
+ $Y2=0
cc_6240 VPWR N_A_7937_297#_c_12196_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6241 N_VPWR_c_7366_n N_A_7937_297#_c_12196_n 0.00115812f $X=41.63 $Y=2.72
+ $X2=0 $Y2=0
cc_6242 N_VPWR_c_7291_n N_A_7937_297#_c_12255_n 6.68271e-19 $X=40.3 $Y=2
+ $X2=25.99 $Y2=2.21
cc_6243 N_VPWR_c_7294_n N_A_7937_297#_c_12255_n 6.68271e-19 $X=41.24 $Y=2
+ $X2=25.99 $Y2=2.21
cc_6244 VPWR N_A_7937_297#_c_12255_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6245 VPWR N_A_7937_297#_c_12224_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6246 N_VPWR_c_7294_n N_A_7937_297#_c_12259_n 6.69936e-19 $X=41.24 $Y=2 $X2=0
+ $Y2=0
cc_6247 VPWR N_A_7937_297#_c_12259_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6248 VPWR N_A_7937_297#_c_12226_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6249 VPWR N_A_7937_297#_c_12262_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6250 N_VPWR_c_7289_n N_A_7937_297#_c_12216_n 0.0318001f $X=39.36 $Y=1.66
+ $X2=25.99 $Y2=3.57
cc_6251 N_VPWR_c_7291_n N_A_7937_297#_c_12216_n 0.0268237f $X=40.3 $Y=2
+ $X2=25.99 $Y2=3.57
cc_6252 VPWR N_A_7937_297#_c_12216_n 0.00313104f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.57
cc_6253 N_VPWR_c_7365_n N_A_7937_297#_c_12216_n 0.0189467f $X=40.165 $Y=2.72
+ $X2=25.99 $Y2=3.57
cc_6254 N_VPWR_c_7291_n N_A_7937_297#_c_12219_n 0.0268237f $X=40.3 $Y=2 $X2=0
+ $Y2=0
cc_6255 N_VPWR_c_7293_n N_A_7937_297#_c_12219_n 0.0189467f $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6256 N_VPWR_c_7294_n N_A_7937_297#_c_12219_n 0.0268237f $X=41.24 $Y=2 $X2=0
+ $Y2=0
cc_6257 VPWR N_A_7937_297#_c_12219_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6258 N_VPWR_c_7296_n N_A_7937_297#_c_12271_n 0.00167067f $X=44.215 $Y=1.77
+ $X2=0 $Y2=0
cc_6259 VPWR N_A_7937_297#_c_12271_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6260 N_VPWR_c_7294_n N_A_7937_297#_c_12197_n 0.0390576f $X=41.24 $Y=2 $X2=0
+ $Y2=0
cc_6261 VPWR N_A_7937_297#_c_12197_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6262 N_VPWR_c_7366_n N_A_7937_297#_c_12197_n 0.0213652f $X=41.63 $Y=2.72
+ $X2=0 $Y2=0
cc_6263 VPWR N_A_7937_297#_c_12198_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6264 N_VPWR_c_7296_n N_A_7937_297#_c_12199_n 0.0505494f $X=44.215 $Y=1.77
+ $X2=0 $Y2=0
cc_6265 N_VPWR_c_7338_n N_A_7937_297#_c_12199_n 0.0213652f $X=44.05 $Y=2.72
+ $X2=0 $Y2=0
cc_6266 VPWR N_A_7937_297#_c_12199_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6267 VPWR N_A_7937_591#_M1109_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=1.525
cc_6268 VPWR N_A_7937_591#_M1251_s 0.0011753f $X=51.665 $Y=2.635 $X2=25.905
+ $Y2=3.04
cc_6269 N_VPWR_M1184_d N_A_7937_591#_c_12328_n 0.00331615f $X=40.155 $Y=2.955
+ $X2=0 $Y2=0
cc_6270 N_VPWR_c_7292_n N_A_7937_591#_c_12328_n 0.0130979f $X=40.3 $Y=3.1 $X2=0
+ $Y2=0
cc_6271 N_VPWR_M1293_d N_A_7937_591#_c_12323_n 0.00715085f $X=41.095 $Y=2.955
+ $X2=0 $Y2=0
cc_6272 N_VPWR_c_7295_n N_A_7937_591#_c_12323_n 0.0152464f $X=41.24 $Y=3.1 $X2=0
+ $Y2=0
cc_6273 N_VPWR_c_7292_n N_A_7937_591#_c_12341_n 0.0153177f $X=40.3 $Y=3.1 $X2=0
+ $Y2=0
cc_6274 N_VPWR_c_7293_n N_A_7937_591#_c_12341_n 8.30334e-19 $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6275 VPWR N_A_7937_591#_c_12341_n 0.0558368f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6276 N_VPWR_c_7365_n N_A_7937_591#_c_12341_n 8.30334e-19 $X=40.165 $Y=2.72
+ $X2=0 $Y2=0
cc_6277 N_VPWR_c_7290_n N_A_7937_591#_c_12376_n 0.00167228f $X=39.36 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_6278 N_VPWR_c_7292_n N_A_7937_591#_c_12376_n 6.68271e-19 $X=40.3 $Y=3.1
+ $X2=25.99 $Y2=1.87
cc_6279 VPWR N_A_7937_591#_c_12376_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6280 N_VPWR_c_7293_n N_A_7937_591#_c_12324_n 8.30334e-19 $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6281 N_VPWR_c_7295_n N_A_7937_591#_c_12324_n 0.0156478f $X=41.24 $Y=3.1 $X2=0
+ $Y2=0
cc_6282 VPWR N_A_7937_591#_c_12324_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6283 N_VPWR_c_7366_n N_A_7937_591#_c_12324_n 0.00115812f $X=41.63 $Y=2.72
+ $X2=0 $Y2=0
cc_6284 N_VPWR_c_7292_n N_A_7937_591#_c_12383_n 6.68271e-19 $X=40.3 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_6285 N_VPWR_c_7295_n N_A_7937_591#_c_12383_n 6.68271e-19 $X=41.24 $Y=3.1
+ $X2=25.99 $Y2=2.21
cc_6286 VPWR N_A_7937_591#_c_12383_n 0.0295747f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6287 VPWR N_A_7937_591#_c_12352_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6288 N_VPWR_c_7295_n N_A_7937_591#_c_12387_n 6.69936e-19 $X=41.24 $Y=3.1
+ $X2=0 $Y2=0
cc_6289 VPWR N_A_7937_591#_c_12387_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6290 VPWR N_A_7937_591#_c_12354_n 0.0571367f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6291 VPWR N_A_7937_591#_c_12390_n 0.0296491f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6292 N_VPWR_c_7297_n N_A_7937_591#_c_12391_n 0.00167067f $X=44.215 $Y=3.14
+ $X2=0 $Y2=0
cc_6293 VPWR N_A_7937_591#_c_12391_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6294 N_VPWR_c_7290_n N_A_7937_591#_c_12344_n 0.0318001f $X=39.36 $Y=3.1 $X2=0
+ $Y2=0
cc_6295 N_VPWR_c_7292_n N_A_7937_591#_c_12344_n 0.0268237f $X=40.3 $Y=3.1 $X2=0
+ $Y2=0
cc_6296 VPWR N_A_7937_591#_c_12344_n 0.00313104f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6297 N_VPWR_c_7365_n N_A_7937_591#_c_12344_n 0.0189467f $X=40.165 $Y=2.72
+ $X2=0 $Y2=0
cc_6298 N_VPWR_c_7292_n N_A_7937_591#_c_12347_n 0.0268237f $X=40.3 $Y=3.1 $X2=0
+ $Y2=0
cc_6299 N_VPWR_c_7293_n N_A_7937_591#_c_12347_n 0.0189467f $X=41.105 $Y=2.72
+ $X2=0 $Y2=0
cc_6300 N_VPWR_c_7295_n N_A_7937_591#_c_12347_n 0.0268237f $X=41.24 $Y=3.1 $X2=0
+ $Y2=0
cc_6301 VPWR N_A_7937_591#_c_12347_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6302 N_VPWR_c_7295_n N_A_7937_591#_c_12325_n 0.0390576f $X=41.24 $Y=3.1 $X2=0
+ $Y2=0
cc_6303 VPWR N_A_7937_591#_c_12325_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6304 N_VPWR_c_7366_n N_A_7937_591#_c_12325_n 0.0213652f $X=41.63 $Y=2.72
+ $X2=0 $Y2=0
cc_6305 VPWR N_A_7937_591#_c_12326_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6306 N_VPWR_c_7297_n N_A_7937_591#_c_12327_n 0.0505494f $X=44.215 $Y=3.14
+ $X2=0 $Y2=0
cc_6307 N_VPWR_c_7338_n N_A_7937_591#_c_12327_n 0.0213652f $X=44.05 $Y=2.72
+ $X2=0 $Y2=0
cc_6308 VPWR N_A_7937_591#_c_12327_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6309 VPWR N_A_9463_311#_M1040_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6310 VPWR N_A_9463_311#_M1131_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6311 N_VPWR_M1040_d N_A_9463_311#_c_12451_n 0.00732532f $X=49.715 $Y=1.485
+ $X2=0 $Y2=0
cc_6312 N_VPWR_c_7305_n N_A_9463_311#_c_12451_n 0.0175034f $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6313 N_VPWR_M1087_d N_A_9463_311#_c_12473_n 0.00346031f $X=50.635 $Y=1.485
+ $X2=0 $Y2=0
cc_6314 N_VPWR_c_7307_n N_A_9463_311#_c_12473_n 0.0138552f $X=50.78 $Y=2 $X2=0
+ $Y2=0
cc_6315 VPWR N_A_9463_311#_c_12460_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6316 N_VPWR_c_7303_n N_A_9463_311#_c_12502_n 0.00167067f $X=46.865 $Y=1.77
+ $X2=25.99 $Y2=1.87
cc_6317 VPWR N_A_9463_311#_c_12502_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6318 VPWR N_A_9463_311#_c_12462_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6319 VPWR N_A_9463_311#_c_12505_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6320 N_VPWR_c_7305_n N_A_9463_311#_c_12453_n 0.0160196f $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6321 N_VPWR_c_7345_n N_A_9463_311#_c_12453_n 0.00115812f $X=49.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6322 VPWR N_A_9463_311#_c_12453_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6323 N_VPWR_c_7367_n N_A_9463_311#_c_12453_n 8.30334e-19 $X=50.645 $Y=2.72
+ $X2=0 $Y2=0
cc_6324 N_VPWR_c_7305_n N_A_9463_311#_c_12510_n 6.69936e-19 $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6325 VPWR N_A_9463_311#_c_12510_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6326 N_VPWR_M1087_d N_A_9463_311#_c_12486_n 2.7385e-19 $X=50.635 $Y=1.485
+ $X2=25.99 $Y2=3.23
cc_6327 N_VPWR_c_7307_n N_A_9463_311#_c_12486_n 0.0156895f $X=50.78 $Y=2
+ $X2=25.99 $Y2=3.23
cc_6328 VPWR N_A_9463_311#_c_12486_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6329 N_VPWR_c_7367_n N_A_9463_311#_c_12486_n 8.30334e-19 $X=50.645 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6330 N_VPWR_c_7368_n N_A_9463_311#_c_12486_n 8.30334e-19 $X=51.585 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6331 N_VPWR_c_7305_n N_A_9463_311#_c_12517_n 6.68271e-19 $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6332 N_VPWR_c_7307_n N_A_9463_311#_c_12517_n 6.68271e-19 $X=50.78 $Y=2 $X2=0
+ $Y2=0
cc_6333 VPWR N_A_9463_311#_c_12517_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6334 N_VPWR_c_7305_n N_A_9463_311#_c_12488_n 0.0254588f $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6335 N_VPWR_c_7307_n N_A_9463_311#_c_12488_n 0.0254588f $X=50.78 $Y=2 $X2=0
+ $Y2=0
cc_6336 VPWR N_A_9463_311#_c_12488_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6337 N_VPWR_c_7367_n N_A_9463_311#_c_12488_n 0.0189467f $X=50.645 $Y=2.72
+ $X2=0 $Y2=0
cc_6338 N_VPWR_c_7307_n N_A_9463_311#_c_12524_n 6.68271e-19 $X=50.78 $Y=2 $X2=0
+ $Y2=0
cc_6339 N_VPWR_c_7309_n N_A_9463_311#_c_12524_n 0.00167228f $X=51.72 $Y=1.66
+ $X2=0 $Y2=0
cc_6340 VPWR N_A_9463_311#_c_12524_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6341 N_VPWR_c_7307_n N_A_9463_311#_c_12491_n 0.0254588f $X=50.78 $Y=2 $X2=0
+ $Y2=0
cc_6342 VPWR N_A_9463_311#_c_12491_n 0.00345059f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6343 N_VPWR_c_7368_n N_A_9463_311#_c_12491_n 0.0189467f $X=51.585 $Y=2.72
+ $X2=0 $Y2=0
cc_6344 N_VPWR_c_7303_n N_A_9463_311#_c_12454_n 0.0505494f $X=46.865 $Y=1.77
+ $X2=0 $Y2=0
cc_6345 N_VPWR_c_7342_n N_A_9463_311#_c_12454_n 0.0213652f $X=47.03 $Y=2.72
+ $X2=0 $Y2=0
cc_6346 VPWR N_A_9463_311#_c_12454_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6347 VPWR N_A_9463_311#_c_12455_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6348 N_VPWR_c_7305_n N_A_9463_311#_c_12456_n 0.0403522f $X=49.84 $Y=2 $X2=0
+ $Y2=0
cc_6349 N_VPWR_c_7345_n N_A_9463_311#_c_12456_n 0.0213652f $X=49.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6350 VPWR N_A_9463_311#_c_12456_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6351 VPWR N_A_9463_613#_M1056_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6352 VPWR N_A_9463_613#_M1145_s 0.0011753f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6353 N_VPWR_M1056_d N_A_9463_613#_c_12570_n 0.00732532f $X=49.715 $Y=2.955
+ $X2=0 $Y2=0
cc_6354 N_VPWR_c_7306_n N_A_9463_613#_c_12570_n 0.0175034f $X=49.84 $Y=3.1 $X2=0
+ $Y2=0
cc_6355 N_VPWR_M1103_d N_A_9463_613#_c_12592_n 0.00346031f $X=50.635 $Y=2.955
+ $X2=0 $Y2=0
cc_6356 N_VPWR_c_7308_n N_A_9463_613#_c_12592_n 0.0138552f $X=50.78 $Y=3.1 $X2=0
+ $Y2=0
cc_6357 VPWR N_A_9463_613#_c_12579_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6358 N_VPWR_c_7304_n N_A_9463_613#_c_12621_n 0.00167067f $X=46.865 $Y=3.14
+ $X2=25.99 $Y2=1.87
cc_6359 VPWR N_A_9463_613#_c_12621_n 0.0297857f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=1.87
cc_6360 VPWR N_A_9463_613#_c_12581_n 0.0571367f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6361 VPWR N_A_9463_613#_c_12624_n 0.0296491f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=2.21
cc_6362 N_VPWR_c_7306_n N_A_9463_613#_c_12572_n 0.0160196f $X=49.84 $Y=3.1 $X2=0
+ $Y2=0
cc_6363 N_VPWR_c_7345_n N_A_9463_613#_c_12572_n 0.00115812f $X=49.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6364 VPWR N_A_9463_613#_c_12572_n 0.0605692f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6365 N_VPWR_c_7367_n N_A_9463_613#_c_12572_n 8.30334e-19 $X=50.645 $Y=2.72
+ $X2=0 $Y2=0
cc_6366 N_VPWR_c_7306_n N_A_9463_613#_c_12629_n 6.69936e-19 $X=49.84 $Y=3.1
+ $X2=0 $Y2=0
cc_6367 VPWR N_A_9463_613#_c_12629_n 0.0297857f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6368 N_VPWR_M1103_d N_A_9463_613#_c_12605_n 2.7385e-19 $X=50.635 $Y=2.955
+ $X2=25.99 $Y2=3.23
cc_6369 N_VPWR_c_7308_n N_A_9463_613#_c_12605_n 0.0156895f $X=50.78 $Y=3.1
+ $X2=25.99 $Y2=3.23
cc_6370 VPWR N_A_9463_613#_c_12605_n 0.0558368f $X=51.665 $Y=2.635 $X2=25.99
+ $Y2=3.23
cc_6371 N_VPWR_c_7367_n N_A_9463_613#_c_12605_n 8.30334e-19 $X=50.645 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6372 N_VPWR_c_7368_n N_A_9463_613#_c_12605_n 8.30334e-19 $X=51.585 $Y=2.72
+ $X2=25.99 $Y2=3.23
cc_6373 N_VPWR_c_7306_n N_A_9463_613#_c_12636_n 6.68271e-19 $X=49.84 $Y=3.1
+ $X2=0 $Y2=0
cc_6374 N_VPWR_c_7308_n N_A_9463_613#_c_12636_n 6.68271e-19 $X=50.78 $Y=3.1
+ $X2=0 $Y2=0
cc_6375 VPWR N_A_9463_613#_c_12636_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6376 N_VPWR_c_7308_n N_A_9463_613#_c_12639_n 6.68271e-19 $X=50.78 $Y=3.1
+ $X2=0 $Y2=0
cc_6377 N_VPWR_c_7310_n N_A_9463_613#_c_12639_n 0.00167228f $X=51.72 $Y=3.1
+ $X2=0 $Y2=0
cc_6378 VPWR N_A_9463_613#_c_12639_n 0.0295747f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6379 N_VPWR_c_7304_n N_A_9463_613#_c_12573_n 0.0505494f $X=46.865 $Y=3.14
+ $X2=0 $Y2=0
cc_6380 N_VPWR_c_7342_n N_A_9463_613#_c_12573_n 0.0213652f $X=47.03 $Y=2.72
+ $X2=0 $Y2=0
cc_6381 VPWR N_A_9463_613#_c_12573_n 0.00284741f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6382 VPWR N_A_9463_613#_c_12574_n 0.00468575f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6383 N_VPWR_c_7306_n N_A_9463_613#_c_12575_n 0.0403522f $X=49.84 $Y=3.1 $X2=0
+ $Y2=0
cc_6384 N_VPWR_c_7345_n N_A_9463_613#_c_12575_n 0.0213652f $X=49.705 $Y=2.72
+ $X2=0 $Y2=0
cc_6385 VPWR N_A_9463_613#_c_12575_n 0.0027766f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6386 N_VPWR_c_7306_n N_A_9463_613#_c_12608_n 0.0254588f $X=49.84 $Y=3.1 $X2=0
+ $Y2=0
cc_6387 N_VPWR_c_7308_n N_A_9463_613#_c_12608_n 0.0254588f $X=50.78 $Y=3.1 $X2=0
+ $Y2=0
cc_6388 VPWR N_A_9463_613#_c_12608_n 0.00300637f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6389 N_VPWR_c_7367_n N_A_9463_613#_c_12608_n 0.0189467f $X=50.645 $Y=2.72
+ $X2=0 $Y2=0
cc_6390 N_VPWR_c_7308_n N_A_9463_613#_c_12611_n 0.0254588f $X=50.78 $Y=3.1 $X2=0
+ $Y2=0
cc_6391 VPWR N_A_9463_613#_c_12611_n 0.00345059f $X=51.665 $Y=2.635 $X2=0 $Y2=0
cc_6392 N_VPWR_c_7368_n N_A_9463_613#_c_12611_n 0.0189467f $X=51.585 $Y=2.72
+ $X2=0 $Y2=0
cc_6393 N_VPWR_c_7217_n N_VGND_c_12690_n 0.00764703f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_6394 N_VPWR_c_7218_n N_VGND_c_12692_n 0.00764703f $X=0.26 $Y=3.1 $X2=0 $Y2=0
cc_6395 N_VPWR_c_7237_n N_VGND_c_12711_n 0.00764703f $X=12.62 $Y=1.66 $X2=0
+ $Y2=0
cc_6396 N_VPWR_c_7238_n N_VGND_c_12712_n 0.00764703f $X=12.62 $Y=3.1 $X2=0 $Y2=0
cc_6397 N_VPWR_c_7240_n N_VGND_c_12715_n 0.00764703f $X=13.14 $Y=1.66 $X2=0
+ $Y2=0
cc_6398 N_VPWR_c_7241_n N_VGND_c_12716_n 0.00764703f $X=13.14 $Y=3.1 $X2=0 $Y2=0
cc_6399 N_VPWR_c_7260_n N_VGND_c_12735_n 0.00764703f $X=25.5 $Y=1.66 $X2=0 $Y2=0
cc_6400 N_VPWR_c_7262_n N_VGND_c_12737_n 0.00764703f $X=25.5 $Y=3.1 $X2=0 $Y2=0
cc_6401 N_VPWR_c_7264_n N_VGND_c_12738_n 0.00764703f $X=26.48 $Y=1.66 $X2=0
+ $Y2=0
cc_6402 N_VPWR_c_7266_n N_VGND_c_12740_n 0.00764703f $X=26.48 $Y=3.1 $X2=0 $Y2=0
cc_6403 N_VPWR_c_7286_n N_VGND_c_12759_n 0.00764703f $X=38.84 $Y=1.66 $X2=0
+ $Y2=0
cc_6404 N_VPWR_c_7287_n N_VGND_c_12760_n 0.00764703f $X=38.84 $Y=3.1 $X2=0 $Y2=0
cc_6405 N_VPWR_c_7289_n N_VGND_c_12763_n 0.00764703f $X=39.36 $Y=1.66 $X2=0
+ $Y2=0
cc_6406 N_VPWR_c_7290_n N_VGND_c_12764_n 0.00764703f $X=39.36 $Y=3.1 $X2=0 $Y2=0
cc_6407 N_VPWR_c_7309_n N_VGND_c_12784_n 0.00764703f $X=51.72 $Y=1.66 $X2=0
+ $Y2=0
cc_6408 N_VPWR_c_7310_n N_VGND_c_12786_n 0.00764703f $X=51.72 $Y=3.1 $X2=0 $Y2=0
cc_6409 N_A_117_297#_c_8774_n N_A_117_591#_c_8890_n 0.00460759f $X=3.6 $Y=1.7
+ $X2=0 $Y2=0
cc_6410 N_A_117_297#_c_8774_n N_Z_c_9004_n 0.0192125f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_6411 N_A_117_297#_c_8774_n N_Z_c_9048_n 0.0024794f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_6412 N_A_117_297#_M1299_d N_Z_c_9115_n 2.15519e-19 $X=4.395 $Y=1.555 $X2=0
+ $Y2=0
cc_6413 N_A_117_297#_c_8802_n N_Z_c_9115_n 0.0146113f $X=4.405 $Y=2.225 $X2=0
+ $Y2=0
cc_6414 N_A_117_297#_c_8847_n N_Z_c_9115_n 0.0238046f $X=4.55 $Y=2.225 $X2=0
+ $Y2=0
cc_6415 N_A_117_297#_c_8775_n N_Z_c_9115_n 0.0169532f $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_6416 N_A_117_297#_c_8802_n N_Z_c_10135_n 0.0238869f $X=4.405 $Y=2.225 $X2=0
+ $Y2=0
cc_6417 N_A_117_297#_c_8774_n N_Z_c_10135_n 6.68271e-19 $X=3.6 $Y=1.7 $X2=0
+ $Y2=0
cc_6418 N_A_117_297#_c_8775_n N_Z_c_10135_n 6.74054e-19 $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_6419 N_A_117_297#_M1207_d Z 3.28377e-19 $X=3.455 $Y=1.555 $X2=0 $Y2=0
cc_6420 N_A_117_297#_c_8800_n Z 0.0139315f $X=3.455 $Y=2.225 $X2=0 $Y2=0
cc_6421 N_A_117_297#_c_8802_n Z 0.0139315f $X=4.405 $Y=2.225 $X2=0 $Y2=0
cc_6422 N_A_117_297#_c_8839_n Z 0.0236317f $X=3.745 $Y=2.225 $X2=0 $Y2=0
cc_6423 N_A_117_297#_c_8774_n Z 0.0151604f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_6424 N_A_117_297#_c_8771_n N_Z_c_9131_n 0.00915958f $X=2.495 $Y=1.58 $X2=0
+ $Y2=0
cc_6425 N_A_117_297#_c_8800_n N_Z_c_9131_n 0.0181912f $X=3.455 $Y=2.225 $X2=0
+ $Y2=0
cc_6426 N_A_117_297#_c_8836_n N_Z_c_9131_n 0.0025679f $X=2.795 $Y=2.225 $X2=0
+ $Y2=0
cc_6427 N_A_117_297#_c_8839_n N_Z_c_9131_n 0.00259673f $X=3.745 $Y=2.225 $X2=0
+ $Y2=0
cc_6428 N_A_117_297#_c_8773_n N_Z_c_9131_n 0.0364724f $X=2.66 $Y=1.7 $X2=0 $Y2=0
cc_6429 N_A_117_297#_c_8774_n N_Z_c_9131_n 0.0438531f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_6430 N_A_117_297#_c_8802_n N_Z_c_9132_n 0.0174871f $X=4.405 $Y=2.225 $X2=0
+ $Y2=0
cc_6431 N_A_117_297#_c_8839_n N_Z_c_9132_n 0.00259673f $X=3.745 $Y=2.225 $X2=0
+ $Y2=0
cc_6432 N_A_117_297#_c_8847_n N_Z_c_9132_n 0.0025679f $X=4.55 $Y=2.225 $X2=0
+ $Y2=0
cc_6433 N_A_117_297#_c_8774_n N_Z_c_9132_n 0.0438531f $X=3.6 $Y=1.7 $X2=0 $Y2=0
cc_6434 N_A_117_297#_c_8775_n N_Z_c_9132_n 0.0420527f $X=4.54 $Y=1.73 $X2=0
+ $Y2=0
cc_6435 N_A_117_297#_c_8800_n N_Z_c_10154_n 0.0238869f $X=3.455 $Y=2.225 $X2=0
+ $Y2=0
cc_6436 N_A_117_297#_c_8773_n N_Z_c_10154_n 0.00168706f $X=2.66 $Y=1.7 $X2=0
+ $Y2=0
cc_6437 N_A_117_297#_c_8774_n N_Z_c_10154_n 6.68271e-19 $X=3.6 $Y=1.7 $X2=0
+ $Y2=0
cc_6438 N_A_117_297#_c_8771_n N_A_119_47#_c_14050_n 0.0247972f $X=2.495 $Y=1.58
+ $X2=25.99 $Y2=1.73
cc_6439 N_A_117_297#_c_8785_n N_A_119_47#_c_14056_n 6.95815e-19 $X=1.67 $Y=1.66
+ $X2=0 $Y2=0
cc_6440 N_A_117_591#_c_8890_n N_Z_c_9005_n 0.0192125f $X=3.6 $Y=3.21 $X2=0 $Y2=0
cc_6441 N_A_117_591#_c_8890_n N_Z_c_9049_n 0.0024794f $X=3.6 $Y=3.21 $X2=0 $Y2=0
cc_6442 N_A_117_591#_M1269_s N_Z_c_9116_n 2.15519e-19 $X=4.395 $Y=3.065 $X2=0
+ $Y2=0
cc_6443 N_A_117_591#_c_8918_n N_Z_c_9116_n 0.0146113f $X=4.405 $Y=3.215 $X2=0
+ $Y2=0
cc_6444 N_A_117_591#_c_8956_n N_Z_c_9116_n 0.0238046f $X=4.55 $Y=3.215 $X2=0
+ $Y2=0
cc_6445 N_A_117_591#_c_8891_n N_Z_c_9116_n 0.0169532f $X=4.54 $Y=3.21 $X2=0
+ $Y2=0
cc_6446 N_A_117_591#_c_8918_n N_Z_c_10163_n 0.0238869f $X=4.405 $Y=3.215 $X2=0
+ $Y2=0
cc_6447 N_A_117_591#_c_8890_n N_Z_c_10163_n 6.68271e-19 $X=3.6 $Y=3.21 $X2=0
+ $Y2=0
cc_6448 N_A_117_591#_c_8891_n N_Z_c_10163_n 6.74054e-19 $X=4.54 $Y=3.21 $X2=0
+ $Y2=0
cc_6449 N_A_117_591#_M1079_s Z 3.28377e-19 $X=3.455 $Y=3.065 $X2=0 $Y2=0
cc_6450 N_A_117_591#_c_8916_n Z 0.0139315f $X=3.455 $Y=3.215 $X2=0 $Y2=0
cc_6451 N_A_117_591#_c_8918_n Z 0.0139315f $X=4.405 $Y=3.215 $X2=0 $Y2=0
cc_6452 N_A_117_591#_c_8955_n Z 0.0236317f $X=3.745 $Y=3.215 $X2=0 $Y2=0
cc_6453 N_A_117_591#_c_8890_n Z 0.0151604f $X=3.6 $Y=3.21 $X2=0 $Y2=0
cc_6454 N_A_117_591#_c_8887_n N_Z_c_9131_n 0.00915958f $X=2.495 $Y=3.86 $X2=0
+ $Y2=0
cc_6455 N_A_117_591#_c_8916_n N_Z_c_9131_n 0.0181912f $X=3.455 $Y=3.215 $X2=0
+ $Y2=0
cc_6456 N_A_117_591#_c_8952_n N_Z_c_9131_n 0.0025679f $X=2.795 $Y=3.215 $X2=0
+ $Y2=0
cc_6457 N_A_117_591#_c_8955_n N_Z_c_9131_n 0.00259673f $X=3.745 $Y=3.215 $X2=0
+ $Y2=0
cc_6458 N_A_117_591#_c_8889_n N_Z_c_9131_n 0.0364724f $X=2.66 $Y=3.21 $X2=0
+ $Y2=0
cc_6459 N_A_117_591#_c_8890_n N_Z_c_9131_n 0.0438531f $X=3.6 $Y=3.21 $X2=0 $Y2=0
cc_6460 N_A_117_591#_c_8918_n N_Z_c_9132_n 0.0174871f $X=4.405 $Y=3.215 $X2=0
+ $Y2=0
cc_6461 N_A_117_591#_c_8955_n N_Z_c_9132_n 0.00259673f $X=3.745 $Y=3.215 $X2=0
+ $Y2=0
cc_6462 N_A_117_591#_c_8956_n N_Z_c_9132_n 0.0025679f $X=4.55 $Y=3.215 $X2=0
+ $Y2=0
cc_6463 N_A_117_591#_c_8890_n N_Z_c_9132_n 0.0438531f $X=3.6 $Y=3.21 $X2=0 $Y2=0
cc_6464 N_A_117_591#_c_8891_n N_Z_c_9132_n 0.0420527f $X=4.54 $Y=3.21 $X2=0
+ $Y2=0
cc_6465 N_A_117_591#_c_8916_n N_Z_c_10182_n 0.0238869f $X=3.455 $Y=3.215 $X2=0
+ $Y2=0
cc_6466 N_A_117_591#_c_8889_n N_Z_c_10182_n 0.00168706f $X=2.66 $Y=3.21 $X2=0
+ $Y2=0
cc_6467 N_A_117_591#_c_8890_n N_Z_c_10182_n 6.68271e-19 $X=3.6 $Y=3.21 $X2=0
+ $Y2=0
cc_6468 N_A_117_591#_c_8887_n N_A_119_911#_c_14132_n 0.0247972f $X=2.495 $Y=3.86
+ $X2=0 $Y2=0
cc_6469 N_A_117_591#_c_8901_n N_A_119_911#_c_14139_n 6.95815e-19 $X=1.67 $Y=3.78
+ $X2=0 $Y2=0
cc_6470 N_Z_c_9115_n N_A_1643_311#_M1007_s 2.15519e-19 $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_6471 N_Z_c_9288_n N_A_1643_311#_M1048_s 3.28377e-19 $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_6472 N_Z_c_9117_n N_A_1643_311#_M1284_s 2.15519e-19 $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6473 N_Z_c_9117_n N_A_1643_311#_c_10897_n 0.0242319f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6474 N_Z_c_9134_n N_A_1643_311#_c_10898_n 0.00915958f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6475 N_Z_c_9117_n N_A_1643_311#_c_10919_n 0.020688f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6476 N_Z_c_9115_n N_A_1643_311#_c_10906_n 0.0146113f $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_6477 N_Z_c_9288_n N_A_1643_311#_c_10906_n 0.0139315f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_6478 Z N_A_1643_311#_c_10906_n 0.0238869f $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_6479 N_Z_c_9133_n N_A_1643_311#_c_10906_n 0.0174871f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6480 N_Z_c_9115_n N_A_1643_311#_c_10948_n 0.0238046f $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_6481 N_Z_c_9133_n N_A_1643_311#_c_10948_n 0.0025679f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6482 N_Z_c_9117_n N_A_1643_311#_c_10908_n 0.0146113f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6483 N_Z_c_10198_p N_A_1643_311#_c_10908_n 0.0238869f $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_6484 N_Z_c_9288_n N_A_1643_311#_c_10908_n 0.0139315f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_6485 N_Z_c_9134_n N_A_1643_311#_c_10908_n 0.0174871f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6486 N_Z_c_9288_n N_A_1643_311#_c_10951_n 0.0236317f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_6487 N_Z_c_9133_n N_A_1643_311#_c_10951_n 0.00259673f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6488 N_Z_c_9134_n N_A_1643_311#_c_10951_n 0.00259673f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6489 N_Z_c_9117_n N_A_1643_311#_c_10899_n 0.0521734f $X=15.865 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6490 N_Z_c_9117_n N_A_1643_311#_c_10956_n 0.0238046f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6491 N_Z_c_9134_n N_A_1643_311#_c_10956_n 0.0025679f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6492 N_Z_c_9117_n N_A_1643_311#_c_10932_n 0.0481433f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6493 N_Z_c_9117_n N_A_1643_311#_c_10962_n 0.0238869f $X=15.865 $Y=1.87
+ $X2=25.99 $Y2=0.64
cc_6494 N_Z_c_9117_n N_A_1643_311#_c_10934_n 0.0205035f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6495 N_Z_c_9117_n N_A_1643_311#_c_10969_n 0.0238869f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6496 N_Z_c_9117_n N_A_1643_311#_c_10937_n 0.0187608f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6497 N_Z_c_9115_n N_A_1643_311#_c_10900_n 0.0169532f $X=8.665 $Y=1.87 $X2=0
+ $Y2=0
cc_6498 Z N_A_1643_311#_c_10900_n 6.74054e-19 $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_6499 N_Z_c_9133_n N_A_1643_311#_c_10900_n 0.0420527f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6500 N_Z_c_9010_n N_A_1643_311#_c_10901_n 0.0192125f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_6501 N_Z_c_9050_n N_A_1643_311#_c_10901_n 0.0024794f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_6502 N_Z_c_10198_p N_A_1643_311#_c_10901_n 6.68271e-19 $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_6503 N_Z_c_9288_n N_A_1643_311#_c_10901_n 0.0151604f $X=9.605 $Y=1.87 $X2=0
+ $Y2=0
cc_6504 Z N_A_1643_311#_c_10901_n 6.68271e-19 $X=8.785 $Y=1.785 $X2=0 $Y2=0
cc_6505 N_Z_c_9133_n N_A_1643_311#_c_10901_n 0.0438531f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6506 N_Z_c_9134_n N_A_1643_311#_c_10901_n 0.0438531f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6507 N_Z_c_9117_n N_A_1643_311#_c_10902_n 0.026602f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6508 N_Z_c_10198_p N_A_1643_311#_c_10902_n 6.74054e-19 $X=9.895 $Y=1.87 $X2=0
+ $Y2=0
cc_6509 N_Z_c_9134_n N_A_1643_311#_c_10902_n 0.0383005f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6510 N_Z_c_9116_n N_A_1643_613#_M1112_d 2.15519e-19 $X=8.665 $Y=3.57 $X2=0
+ $Y2=0
cc_6511 N_Z_c_9317_n N_A_1643_613#_M1161_d 3.28377e-19 $X=9.605 $Y=3.57 $X2=0
+ $Y2=0
cc_6512 N_Z_c_9118_n N_A_1643_613#_M1273_d 2.15519e-19 $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6513 N_Z_c_9118_n N_A_1643_613#_c_11028_n 0.0242319f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6514 N_Z_c_9134_n N_A_1643_613#_c_11029_n 0.00915958f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6515 N_Z_c_9118_n N_A_1643_613#_c_11050_n 0.020688f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6516 N_Z_c_9116_n N_A_1643_613#_c_11037_n 0.0146113f $X=8.665 $Y=3.57 $X2=0
+ $Y2=0
cc_6517 N_Z_c_9317_n N_A_1643_613#_c_11037_n 0.0139315f $X=9.605 $Y=3.57 $X2=0
+ $Y2=0
cc_6518 Z N_A_1643_613#_c_11037_n 0.0238869f $X=8.785 $Y=3.485 $X2=0 $Y2=0
cc_6519 N_Z_c_9133_n N_A_1643_613#_c_11037_n 0.0174871f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6520 N_Z_c_9116_n N_A_1643_613#_c_11079_n 0.0238046f $X=8.665 $Y=3.57 $X2=0
+ $Y2=0
cc_6521 N_Z_c_9133_n N_A_1643_613#_c_11079_n 0.0025679f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6522 N_Z_c_9118_n N_A_1643_613#_c_11039_n 0.0146113f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6523 N_Z_c_10238_p N_A_1643_613#_c_11039_n 0.0238869f $X=9.895 $Y=3.57 $X2=0
+ $Y2=0
cc_6524 N_Z_c_9317_n N_A_1643_613#_c_11039_n 0.0139315f $X=9.605 $Y=3.57 $X2=0
+ $Y2=0
cc_6525 N_Z_c_9134_n N_A_1643_613#_c_11039_n 0.0174871f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6526 N_Z_c_9317_n N_A_1643_613#_c_11082_n 0.0236317f $X=9.605 $Y=3.57 $X2=0
+ $Y2=0
cc_6527 N_Z_c_9133_n N_A_1643_613#_c_11082_n 0.00259673f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6528 N_Z_c_9134_n N_A_1643_613#_c_11082_n 0.00259673f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6529 N_Z_c_9118_n N_A_1643_613#_c_11030_n 0.0521734f $X=15.865 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6530 N_Z_c_9118_n N_A_1643_613#_c_11087_n 0.0238046f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6531 N_Z_c_9134_n N_A_1643_613#_c_11087_n 0.0025679f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6532 N_Z_c_9118_n N_A_1643_613#_c_11063_n 0.0481433f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6533 N_Z_c_9118_n N_A_1643_613#_c_11093_n 0.0238869f $X=15.865 $Y=3.57
+ $X2=25.99 $Y2=0.64
cc_6534 N_Z_c_9118_n N_A_1643_613#_c_11096_n 0.0238869f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6535 N_Z_c_9116_n N_A_1643_613#_c_11031_n 0.0169532f $X=8.665 $Y=3.57 $X2=0
+ $Y2=0
cc_6536 Z N_A_1643_613#_c_11031_n 6.74054e-19 $X=8.785 $Y=3.485 $X2=0 $Y2=0
cc_6537 N_Z_c_9133_n N_A_1643_613#_c_11031_n 0.0420527f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6538 N_Z_c_9011_n N_A_1643_613#_c_11032_n 0.0192125f $X=9.585 $Y=4.225 $X2=0
+ $Y2=0
cc_6539 N_Z_c_9051_n N_A_1643_613#_c_11032_n 0.0024794f $X=8.91 $Y=4.225 $X2=0
+ $Y2=0
cc_6540 N_Z_c_10238_p N_A_1643_613#_c_11032_n 6.68271e-19 $X=9.895 $Y=3.57 $X2=0
+ $Y2=0
cc_6541 N_Z_c_9317_n N_A_1643_613#_c_11032_n 0.0151604f $X=9.605 $Y=3.57 $X2=0
+ $Y2=0
cc_6542 Z N_A_1643_613#_c_11032_n 6.68271e-19 $X=8.785 $Y=3.485 $X2=0 $Y2=0
cc_6543 N_Z_c_9133_n N_A_1643_613#_c_11032_n 0.0438531f $X=8.81 $Y=1.7 $X2=0
+ $Y2=0
cc_6544 N_Z_c_9134_n N_A_1643_613#_c_11032_n 0.0438531f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6545 N_Z_c_9118_n N_A_1643_613#_c_11033_n 0.026602f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6546 N_Z_c_10238_p N_A_1643_613#_c_11033_n 6.74054e-19 $X=9.895 $Y=3.57 $X2=0
+ $Y2=0
cc_6547 N_Z_c_9134_n N_A_1643_613#_c_11033_n 0.0383005f $X=9.75 $Y=1.7 $X2=0
+ $Y2=0
cc_6548 N_Z_c_9118_n N_A_1643_613#_c_11066_n 0.0205035f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6549 N_Z_c_9118_n N_A_1643_613#_c_11069_n 0.0187608f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6550 N_Z_c_9117_n N_A_2693_297#_M1082_d 2.15519e-19 $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6551 Z N_A_2693_297#_M1138_d 3.28377e-19 $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_6552 N_Z_c_9119_n N_A_2693_297#_M1250_d 2.15519e-19 $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6553 N_Z_c_9117_n N_A_2693_297#_c_11164_n 0.020688f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6554 N_Z_c_9117_n N_A_2693_297#_c_11159_n 0.0242319f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6555 N_Z_c_9135_n N_A_2693_297#_c_11159_n 0.00915958f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6556 N_Z_c_9117_n N_A_2693_297#_c_11177_n 0.0481433f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6557 N_Z_c_9117_n N_A_2693_297#_c_11212_n 0.0238869f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6558 N_Z_c_9117_n N_A_2693_297#_c_11160_n 0.0521734f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6559 N_Z_c_9117_n N_A_2693_297#_c_11219_n 0.0238869f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6560 N_Z_c_9117_n N_A_2693_297#_c_11188_n 0.0146113f $X=15.865 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6561 N_Z_c_10276_p N_A_2693_297#_c_11188_n 0.0238869f $X=16.155 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6562 Z N_A_2693_297#_c_11188_n 0.0139315f $X=16.805 $Y=1.785 $X2=25.99
+ $Y2=0.51
cc_6563 N_Z_c_9135_n N_A_2693_297#_c_11188_n 0.0174871f $X=16.01 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6564 N_Z_c_9117_n N_A_2693_297#_c_11223_n 0.0238046f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6565 N_Z_c_9135_n N_A_2693_297#_c_11223_n 0.0025679f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6566 N_Z_c_9119_n N_A_2693_297#_c_11190_n 0.0146113f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6567 N_Z_c_10282_p N_A_2693_297#_c_11190_n 0.0238869f $X=17.095 $Y=1.87 $X2=0
+ $Y2=0
cc_6568 Z N_A_2693_297#_c_11190_n 0.0139315f $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_6569 N_Z_c_9136_n N_A_2693_297#_c_11190_n 0.0174871f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6570 Z N_A_2693_297#_c_11226_n 0.0236317f $X=16.805 $Y=1.785 $X2=25.99
+ $Y2=0.64
cc_6571 N_Z_c_9135_n N_A_2693_297#_c_11226_n 0.00259673f $X=16.01 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6572 N_Z_c_9136_n N_A_2693_297#_c_11226_n 0.00259673f $X=16.95 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6573 N_Z_c_9117_n N_A_2693_297#_c_11180_n 0.0187608f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6574 N_Z_c_9117_n N_A_2693_297#_c_11183_n 0.0205035f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6575 N_Z_c_9119_n N_A_2693_297#_c_11235_n 0.0238046f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6576 N_Z_c_9136_n N_A_2693_297#_c_11235_n 0.0025679f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6577 N_Z_c_9117_n N_A_2693_297#_c_11161_n 0.026602f $X=15.865 $Y=1.87 $X2=0
+ $Y2=0
cc_6578 N_Z_c_10276_p N_A_2693_297#_c_11161_n 6.74054e-19 $X=16.155 $Y=1.87
+ $X2=0 $Y2=0
cc_6579 N_Z_c_9135_n N_A_2693_297#_c_11161_n 0.0383005f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6580 N_Z_c_9014_n N_A_2693_297#_c_11162_n 0.0192125f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_6581 N_Z_c_9062_n N_A_2693_297#_c_11162_n 0.0024794f $X=16.85 $Y=1.215 $X2=0
+ $Y2=0
cc_6582 N_Z_c_10282_p N_A_2693_297#_c_11162_n 6.68271e-19 $X=17.095 $Y=1.87
+ $X2=0 $Y2=0
cc_6583 N_Z_c_10276_p N_A_2693_297#_c_11162_n 6.68271e-19 $X=16.155 $Y=1.87
+ $X2=0 $Y2=0
cc_6584 Z N_A_2693_297#_c_11162_n 0.0151604f $X=16.805 $Y=1.785 $X2=0 $Y2=0
cc_6585 N_Z_c_9135_n N_A_2693_297#_c_11162_n 0.0438531f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6586 N_Z_c_9136_n N_A_2693_297#_c_11162_n 0.0438531f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6587 N_Z_c_9119_n N_A_2693_297#_c_11163_n 0.0169532f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6588 N_Z_c_10282_p N_A_2693_297#_c_11163_n 6.74054e-19 $X=17.095 $Y=1.87
+ $X2=0 $Y2=0
cc_6589 N_Z_c_9136_n N_A_2693_297#_c_11163_n 0.0420527f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6590 N_Z_c_9118_n N_A_2693_591#_M1000_d 2.15519e-19 $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6591 Z N_A_2693_591#_M1080_d 3.28377e-19 $X=16.805 $Y=3.485 $X2=0 $Y2=0
cc_6592 N_Z_c_9120_n N_A_2693_591#_M1270_d 2.15519e-19 $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6593 N_Z_c_9118_n N_A_2693_591#_c_11292_n 0.020688f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6594 N_Z_c_9118_n N_A_2693_591#_c_11287_n 0.0242319f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6595 N_Z_c_9135_n N_A_2693_591#_c_11287_n 0.00915958f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6596 N_Z_c_9118_n N_A_2693_591#_c_11305_n 0.0481433f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6597 N_Z_c_9118_n N_A_2693_591#_c_11340_n 0.0238869f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6598 N_Z_c_9118_n N_A_2693_591#_c_11288_n 0.0521734f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6599 N_Z_c_9118_n N_A_2693_591#_c_11347_n 0.0238869f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6600 N_Z_c_9118_n N_A_2693_591#_c_11316_n 0.0146113f $X=15.865 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6601 N_Z_c_10316_p N_A_2693_591#_c_11316_n 0.0238869f $X=16.155 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6602 Z N_A_2693_591#_c_11316_n 0.0139315f $X=16.805 $Y=3.485 $X2=25.99
+ $Y2=0.51
cc_6603 N_Z_c_9135_n N_A_2693_591#_c_11316_n 0.0174871f $X=16.01 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6604 N_Z_c_9118_n N_A_2693_591#_c_11351_n 0.0238046f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6605 N_Z_c_9135_n N_A_2693_591#_c_11351_n 0.0025679f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6606 N_Z_c_9120_n N_A_2693_591#_c_11318_n 0.0146113f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6607 N_Z_c_10322_p N_A_2693_591#_c_11318_n 0.0238869f $X=17.095 $Y=3.57 $X2=0
+ $Y2=0
cc_6608 Z N_A_2693_591#_c_11318_n 0.0139315f $X=16.805 $Y=3.485 $X2=0 $Y2=0
cc_6609 N_Z_c_9136_n N_A_2693_591#_c_11318_n 0.0174871f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6610 Z N_A_2693_591#_c_11354_n 0.0236317f $X=16.805 $Y=3.485 $X2=25.99
+ $Y2=0.64
cc_6611 N_Z_c_9135_n N_A_2693_591#_c_11354_n 0.00259673f $X=16.01 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6612 N_Z_c_9136_n N_A_2693_591#_c_11354_n 0.00259673f $X=16.95 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6613 N_Z_c_9120_n N_A_2693_591#_c_11355_n 0.0238046f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6614 N_Z_c_9136_n N_A_2693_591#_c_11355_n 0.0025679f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6615 N_Z_c_9118_n N_A_2693_591#_c_11308_n 0.0187608f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6616 N_Z_c_9118_n N_A_2693_591#_c_11311_n 0.0205035f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6617 N_Z_c_9118_n N_A_2693_591#_c_11289_n 0.026602f $X=15.865 $Y=3.57 $X2=0
+ $Y2=0
cc_6618 N_Z_c_10316_p N_A_2693_591#_c_11289_n 6.74054e-19 $X=16.155 $Y=3.57
+ $X2=0 $Y2=0
cc_6619 N_Z_c_9135_n N_A_2693_591#_c_11289_n 0.0383005f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6620 N_Z_c_9015_n N_A_2693_591#_c_11290_n 0.0192125f $X=16.585 $Y=4.225 $X2=0
+ $Y2=0
cc_6621 N_Z_c_9063_n N_A_2693_591#_c_11290_n 0.0024794f $X=16.85 $Y=4.225 $X2=0
+ $Y2=0
cc_6622 N_Z_c_10322_p N_A_2693_591#_c_11290_n 6.68271e-19 $X=17.095 $Y=3.57
+ $X2=0 $Y2=0
cc_6623 N_Z_c_10316_p N_A_2693_591#_c_11290_n 6.68271e-19 $X=16.155 $Y=3.57
+ $X2=0 $Y2=0
cc_6624 Z N_A_2693_591#_c_11290_n 0.0151604f $X=16.805 $Y=3.485 $X2=0 $Y2=0
cc_6625 N_Z_c_9135_n N_A_2693_591#_c_11290_n 0.0438531f $X=16.01 $Y=1.7 $X2=0
+ $Y2=0
cc_6626 N_Z_c_9136_n N_A_2693_591#_c_11290_n 0.0438531f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6627 N_Z_c_9120_n N_A_2693_591#_c_11291_n 0.0169532f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6628 N_Z_c_10322_p N_A_2693_591#_c_11291_n 6.74054e-19 $X=17.095 $Y=3.57
+ $X2=0 $Y2=0
cc_6629 N_Z_c_9136_n N_A_2693_591#_c_11291_n 0.0420527f $X=16.95 $Y=1.7 $X2=0
+ $Y2=0
cc_6630 N_Z_c_9119_n N_A_4219_311#_M1121_d 2.15519e-19 $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6631 N_Z_c_9494_n N_A_4219_311#_M1171_d 3.28377e-19 $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_6632 N_Z_c_9121_n N_A_4219_311#_M1287_d 2.15519e-19 $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6633 N_Z_c_9121_n N_A_4219_311#_c_11415_n 0.0242319f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6634 N_Z_c_9138_n N_A_4219_311#_c_11416_n 0.00915958f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6635 N_Z_c_9121_n N_A_4219_311#_c_11437_n 0.020688f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6636 N_Z_c_9119_n N_A_4219_311#_c_11424_n 0.0146113f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6637 N_Z_c_9494_n N_A_4219_311#_c_11424_n 0.0139315f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_6638 Z N_A_4219_311#_c_11424_n 0.0238869f $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_6639 N_Z_c_9137_n N_A_4219_311#_c_11424_n 0.0174871f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6640 N_Z_c_9119_n N_A_4219_311#_c_11466_n 0.0238046f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6641 N_Z_c_9137_n N_A_4219_311#_c_11466_n 0.0025679f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6642 N_Z_c_9121_n N_A_4219_311#_c_11426_n 0.0146113f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6643 N_Z_c_10358_p N_A_4219_311#_c_11426_n 0.0238869f $X=22.775 $Y=1.87 $X2=0
+ $Y2=0
cc_6644 N_Z_c_9494_n N_A_4219_311#_c_11426_n 0.0139315f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_6645 N_Z_c_9138_n N_A_4219_311#_c_11426_n 0.0174871f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6646 N_Z_c_9494_n N_A_4219_311#_c_11469_n 0.0236317f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_6647 N_Z_c_9137_n N_A_4219_311#_c_11469_n 0.00259673f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6648 N_Z_c_9138_n N_A_4219_311#_c_11469_n 0.00259673f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6649 N_Z_c_9121_n N_A_4219_311#_c_11417_n 0.0521734f $X=29.205 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6650 N_Z_c_9121_n N_A_4219_311#_c_11474_n 0.0238046f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6651 N_Z_c_9138_n N_A_4219_311#_c_11474_n 0.0025679f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6652 N_Z_c_9121_n N_A_4219_311#_c_11450_n 0.0481433f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6653 N_Z_c_9121_n N_A_4219_311#_c_11480_n 0.0238869f $X=29.205 $Y=1.87
+ $X2=25.99 $Y2=0.64
cc_6654 N_Z_c_9121_n N_A_4219_311#_c_11452_n 0.0205035f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6655 N_Z_c_9121_n N_A_4219_311#_c_11487_n 0.0238869f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6656 N_Z_c_9121_n N_A_4219_311#_c_11455_n 0.0187608f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6657 N_Z_c_9119_n N_A_4219_311#_c_11418_n 0.0169532f $X=21.545 $Y=1.87 $X2=0
+ $Y2=0
cc_6658 Z N_A_4219_311#_c_11418_n 6.74054e-19 $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_6659 N_Z_c_9137_n N_A_4219_311#_c_11418_n 0.0420527f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6660 N_Z_c_9020_n N_A_4219_311#_c_11419_n 0.0192125f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_6661 N_Z_c_9064_n N_A_4219_311#_c_11419_n 0.0024794f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_6662 N_Z_c_10358_p N_A_4219_311#_c_11419_n 6.68271e-19 $X=22.775 $Y=1.87
+ $X2=0 $Y2=0
cc_6663 N_Z_c_9494_n N_A_4219_311#_c_11419_n 0.0151604f $X=22.485 $Y=1.87 $X2=0
+ $Y2=0
cc_6664 Z N_A_4219_311#_c_11419_n 6.68271e-19 $X=21.665 $Y=1.785 $X2=0 $Y2=0
cc_6665 N_Z_c_9137_n N_A_4219_311#_c_11419_n 0.0438531f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6666 N_Z_c_9138_n N_A_4219_311#_c_11419_n 0.0438531f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6667 N_Z_c_9121_n N_A_4219_311#_c_11420_n 0.026602f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6668 N_Z_c_10358_p N_A_4219_311#_c_11420_n 6.74054e-19 $X=22.775 $Y=1.87
+ $X2=0 $Y2=0
cc_6669 N_Z_c_9138_n N_A_4219_311#_c_11420_n 0.0383005f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6670 N_Z_c_9120_n N_A_4219_613#_M1071_d 2.15519e-19 $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6671 N_Z_c_9523_n N_A_4219_613#_M1114_d 3.28377e-19 $X=22.485 $Y=3.57 $X2=0
+ $Y2=0
cc_6672 N_Z_c_9123_n N_A_4219_613#_M1313_d 2.15519e-19 $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6673 N_Z_c_9123_n N_A_4219_613#_c_11546_n 0.0242319f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6674 N_Z_c_9138_n N_A_4219_613#_c_11547_n 0.00915958f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6675 N_Z_c_9123_n N_A_4219_613#_c_11568_n 0.020688f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6676 N_Z_c_9120_n N_A_4219_613#_c_11555_n 0.0146113f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6677 N_Z_c_9523_n N_A_4219_613#_c_11555_n 0.0139315f $X=22.485 $Y=3.57 $X2=0
+ $Y2=0
cc_6678 Z N_A_4219_613#_c_11555_n 0.0238869f $X=21.665 $Y=3.485 $X2=0 $Y2=0
cc_6679 N_Z_c_9137_n N_A_4219_613#_c_11555_n 0.0174871f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6680 N_Z_c_9120_n N_A_4219_613#_c_11597_n 0.0238046f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6681 N_Z_c_9137_n N_A_4219_613#_c_11597_n 0.0025679f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6682 N_Z_c_9123_n N_A_4219_613#_c_11557_n 0.0146113f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6683 N_Z_c_10398_p N_A_4219_613#_c_11557_n 0.0238869f $X=22.775 $Y=3.57 $X2=0
+ $Y2=0
cc_6684 N_Z_c_9523_n N_A_4219_613#_c_11557_n 0.0139315f $X=22.485 $Y=3.57 $X2=0
+ $Y2=0
cc_6685 N_Z_c_9138_n N_A_4219_613#_c_11557_n 0.0174871f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6686 N_Z_c_9523_n N_A_4219_613#_c_11600_n 0.0236317f $X=22.485 $Y=3.57 $X2=0
+ $Y2=0
cc_6687 N_Z_c_9137_n N_A_4219_613#_c_11600_n 0.00259673f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6688 N_Z_c_9138_n N_A_4219_613#_c_11600_n 0.00259673f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6689 N_Z_c_9123_n N_A_4219_613#_c_11548_n 0.0521734f $X=29.205 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6690 N_Z_c_9123_n N_A_4219_613#_c_11605_n 0.0238046f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6691 N_Z_c_9138_n N_A_4219_613#_c_11605_n 0.0025679f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6692 N_Z_c_9123_n N_A_4219_613#_c_11581_n 0.0481433f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6693 N_Z_c_9123_n N_A_4219_613#_c_11611_n 0.0238869f $X=29.205 $Y=3.57
+ $X2=25.99 $Y2=0.64
cc_6694 N_Z_c_9123_n N_A_4219_613#_c_11614_n 0.0238869f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6695 N_Z_c_9120_n N_A_4219_613#_c_11549_n 0.0169532f $X=21.545 $Y=3.57 $X2=0
+ $Y2=0
cc_6696 Z N_A_4219_613#_c_11549_n 6.74054e-19 $X=21.665 $Y=3.485 $X2=0 $Y2=0
cc_6697 N_Z_c_9137_n N_A_4219_613#_c_11549_n 0.0420527f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6698 N_Z_c_9021_n N_A_4219_613#_c_11550_n 0.0192125f $X=22.465 $Y=4.225 $X2=0
+ $Y2=0
cc_6699 N_Z_c_9065_n N_A_4219_613#_c_11550_n 0.0024794f $X=21.79 $Y=4.225 $X2=0
+ $Y2=0
cc_6700 N_Z_c_10398_p N_A_4219_613#_c_11550_n 6.68271e-19 $X=22.775 $Y=3.57
+ $X2=0 $Y2=0
cc_6701 N_Z_c_9523_n N_A_4219_613#_c_11550_n 0.0151604f $X=22.485 $Y=3.57 $X2=0
+ $Y2=0
cc_6702 Z N_A_4219_613#_c_11550_n 6.68271e-19 $X=21.665 $Y=3.485 $X2=0 $Y2=0
cc_6703 N_Z_c_9137_n N_A_4219_613#_c_11550_n 0.0438531f $X=21.69 $Y=1.7 $X2=0
+ $Y2=0
cc_6704 N_Z_c_9138_n N_A_4219_613#_c_11550_n 0.0438531f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6705 N_Z_c_9123_n N_A_4219_613#_c_11551_n 0.026602f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6706 N_Z_c_10398_p N_A_4219_613#_c_11551_n 6.74054e-19 $X=22.775 $Y=3.57
+ $X2=0 $Y2=0
cc_6707 N_Z_c_9138_n N_A_4219_613#_c_11551_n 0.0383005f $X=22.63 $Y=1.7 $X2=0
+ $Y2=0
cc_6708 N_Z_c_9123_n N_A_4219_613#_c_11584_n 0.0205035f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6709 N_Z_c_9123_n N_A_4219_613#_c_11587_n 0.0187608f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6710 N_Z_c_9121_n N_A_5361_297#_M1050_d 2.15519e-19 $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6711 Z N_A_5361_297#_M1118_d 3.28377e-19 $X=30.145 $Y=1.785 $X2=0 $Y2=0
cc_6712 N_Z_c_9125_n N_A_5361_297#_M1295_d 2.15519e-19 $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6713 N_Z_c_9121_n N_A_5361_297#_c_11682_n 0.020688f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6714 N_Z_c_9121_n N_A_5361_297#_c_11677_n 0.0242319f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6715 N_Z_c_9139_n N_A_5361_297#_c_11677_n 0.00915958f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6716 N_Z_c_9121_n N_A_5361_297#_c_11695_n 0.0481433f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6717 N_Z_c_9121_n N_A_5361_297#_c_11730_n 0.0238869f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6718 N_Z_c_9121_n N_A_5361_297#_c_11678_n 0.0521734f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6719 N_Z_c_9121_n N_A_5361_297#_c_11737_n 0.0238869f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6720 N_Z_c_9121_n N_A_5361_297#_c_11706_n 0.0146113f $X=29.205 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6721 N_Z_c_10436_p N_A_5361_297#_c_11706_n 0.0238869f $X=29.495 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6722 Z N_A_5361_297#_c_11706_n 0.0139315f $X=30.145 $Y=1.785 $X2=25.99
+ $Y2=0.51
cc_6723 N_Z_c_9139_n N_A_5361_297#_c_11706_n 0.0174871f $X=29.35 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6724 N_Z_c_9121_n N_A_5361_297#_c_11741_n 0.0238046f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6725 N_Z_c_9139_n N_A_5361_297#_c_11741_n 0.0025679f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6726 N_Z_c_9125_n N_A_5361_297#_c_11708_n 0.0146113f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6727 N_Z_c_10442_p N_A_5361_297#_c_11708_n 0.0238869f $X=30.435 $Y=1.87 $X2=0
+ $Y2=0
cc_6728 Z N_A_5361_297#_c_11708_n 0.0139315f $X=30.145 $Y=1.785 $X2=0 $Y2=0
cc_6729 N_Z_c_9140_n N_A_5361_297#_c_11708_n 0.0174871f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6730 Z N_A_5361_297#_c_11744_n 0.0236317f $X=30.145 $Y=1.785 $X2=25.99
+ $Y2=0.64
cc_6731 N_Z_c_9139_n N_A_5361_297#_c_11744_n 0.00259673f $X=29.35 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6732 N_Z_c_9140_n N_A_5361_297#_c_11744_n 0.00259673f $X=30.29 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6733 N_Z_c_9121_n N_A_5361_297#_c_11698_n 0.0187608f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6734 N_Z_c_9121_n N_A_5361_297#_c_11701_n 0.0205035f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6735 N_Z_c_9125_n N_A_5361_297#_c_11753_n 0.0238046f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6736 N_Z_c_9140_n N_A_5361_297#_c_11753_n 0.0025679f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6737 N_Z_c_9121_n N_A_5361_297#_c_11679_n 0.026602f $X=29.205 $Y=1.87 $X2=0
+ $Y2=0
cc_6738 N_Z_c_10436_p N_A_5361_297#_c_11679_n 6.74054e-19 $X=29.495 $Y=1.87
+ $X2=0 $Y2=0
cc_6739 N_Z_c_9139_n N_A_5361_297#_c_11679_n 0.0383005f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6740 N_Z_c_9024_n N_A_5361_297#_c_11680_n 0.0192125f $X=29.925 $Y=1.215 $X2=0
+ $Y2=0
cc_6741 N_Z_c_9076_n N_A_5361_297#_c_11680_n 0.0024794f $X=30.19 $Y=1.215 $X2=0
+ $Y2=0
cc_6742 N_Z_c_10442_p N_A_5361_297#_c_11680_n 6.68271e-19 $X=30.435 $Y=1.87
+ $X2=0 $Y2=0
cc_6743 N_Z_c_10436_p N_A_5361_297#_c_11680_n 6.68271e-19 $X=29.495 $Y=1.87
+ $X2=0 $Y2=0
cc_6744 Z N_A_5361_297#_c_11680_n 0.0151604f $X=30.145 $Y=1.785 $X2=0 $Y2=0
cc_6745 N_Z_c_9139_n N_A_5361_297#_c_11680_n 0.0438531f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6746 N_Z_c_9140_n N_A_5361_297#_c_11680_n 0.0438531f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6747 N_Z_c_9125_n N_A_5361_297#_c_11681_n 0.0169532f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6748 N_Z_c_10442_p N_A_5361_297#_c_11681_n 6.74054e-19 $X=30.435 $Y=1.87
+ $X2=0 $Y2=0
cc_6749 N_Z_c_9140_n N_A_5361_297#_c_11681_n 0.0420527f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6750 N_Z_c_9123_n N_A_5361_591#_M1055_s 2.15519e-19 $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6751 Z N_A_5361_591#_M1119_s 3.28377e-19 $X=30.145 $Y=3.485 $X2=0 $Y2=0
cc_6752 N_Z_c_9126_n N_A_5361_591#_M1257_s 2.15519e-19 $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6753 N_Z_c_9123_n N_A_5361_591#_c_11810_n 0.020688f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6754 N_Z_c_9123_n N_A_5361_591#_c_11805_n 0.0242319f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6755 N_Z_c_9139_n N_A_5361_591#_c_11805_n 0.00915958f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6756 N_Z_c_9123_n N_A_5361_591#_c_11823_n 0.0481433f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6757 N_Z_c_9123_n N_A_5361_591#_c_11858_n 0.0238869f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6758 N_Z_c_9123_n N_A_5361_591#_c_11806_n 0.0521734f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6759 N_Z_c_9123_n N_A_5361_591#_c_11865_n 0.0238869f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6760 N_Z_c_9123_n N_A_5361_591#_c_11834_n 0.0146113f $X=29.205 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6761 N_Z_c_10476_p N_A_5361_591#_c_11834_n 0.0238869f $X=29.495 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6762 Z N_A_5361_591#_c_11834_n 0.0139315f $X=30.145 $Y=3.485 $X2=25.99
+ $Y2=0.51
cc_6763 N_Z_c_9139_n N_A_5361_591#_c_11834_n 0.0174871f $X=29.35 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6764 N_Z_c_9123_n N_A_5361_591#_c_11869_n 0.0238046f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6765 N_Z_c_9139_n N_A_5361_591#_c_11869_n 0.0025679f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6766 N_Z_c_9126_n N_A_5361_591#_c_11836_n 0.0146113f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6767 N_Z_c_10482_p N_A_5361_591#_c_11836_n 0.0238869f $X=30.435 $Y=3.57 $X2=0
+ $Y2=0
cc_6768 Z N_A_5361_591#_c_11836_n 0.0139315f $X=30.145 $Y=3.485 $X2=0 $Y2=0
cc_6769 N_Z_c_9140_n N_A_5361_591#_c_11836_n 0.0174871f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6770 Z N_A_5361_591#_c_11872_n 0.0236317f $X=30.145 $Y=3.485 $X2=25.99
+ $Y2=0.64
cc_6771 N_Z_c_9139_n N_A_5361_591#_c_11872_n 0.00259673f $X=29.35 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6772 N_Z_c_9140_n N_A_5361_591#_c_11872_n 0.00259673f $X=30.29 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6773 N_Z_c_9126_n N_A_5361_591#_c_11873_n 0.0238046f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6774 N_Z_c_9140_n N_A_5361_591#_c_11873_n 0.0025679f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6775 N_Z_c_9123_n N_A_5361_591#_c_11826_n 0.0187608f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6776 N_Z_c_9123_n N_A_5361_591#_c_11829_n 0.0205035f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6777 N_Z_c_9123_n N_A_5361_591#_c_11807_n 0.026602f $X=29.205 $Y=3.57 $X2=0
+ $Y2=0
cc_6778 N_Z_c_10476_p N_A_5361_591#_c_11807_n 6.74054e-19 $X=29.495 $Y=3.57
+ $X2=0 $Y2=0
cc_6779 N_Z_c_9139_n N_A_5361_591#_c_11807_n 0.0383005f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6780 N_Z_c_9025_n N_A_5361_591#_c_11808_n 0.0192125f $X=29.925 $Y=4.225 $X2=0
+ $Y2=0
cc_6781 N_Z_c_9077_n N_A_5361_591#_c_11808_n 0.0024794f $X=30.19 $Y=4.225 $X2=0
+ $Y2=0
cc_6782 N_Z_c_10482_p N_A_5361_591#_c_11808_n 6.68271e-19 $X=30.435 $Y=3.57
+ $X2=0 $Y2=0
cc_6783 N_Z_c_10476_p N_A_5361_591#_c_11808_n 6.68271e-19 $X=29.495 $Y=3.57
+ $X2=0 $Y2=0
cc_6784 Z N_A_5361_591#_c_11808_n 0.0151604f $X=30.145 $Y=3.485 $X2=0 $Y2=0
cc_6785 N_Z_c_9139_n N_A_5361_591#_c_11808_n 0.0438531f $X=29.35 $Y=1.7 $X2=0
+ $Y2=0
cc_6786 N_Z_c_9140_n N_A_5361_591#_c_11808_n 0.0438531f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6787 N_Z_c_9126_n N_A_5361_591#_c_11809_n 0.0169532f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6788 N_Z_c_10482_p N_A_5361_591#_c_11809_n 6.74054e-19 $X=30.435 $Y=3.57
+ $X2=0 $Y2=0
cc_6789 N_Z_c_9140_n N_A_5361_591#_c_11809_n 0.0420527f $X=30.29 $Y=1.7 $X2=0
+ $Y2=0
cc_6790 N_Z_c_9125_n N_A_6887_311#_M1046_s 2.15519e-19 $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6791 N_Z_c_9700_n N_A_6887_311#_M1094_s 3.28377e-19 $X=35.825 $Y=1.87 $X2=0
+ $Y2=0
cc_6792 N_Z_c_9127_n N_A_6887_311#_M1292_s 2.15519e-19 $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6793 N_Z_c_9127_n N_A_6887_311#_c_11933_n 0.0242319f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6794 N_Z_c_9142_n N_A_6887_311#_c_11934_n 0.00915958f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6795 N_Z_c_9127_n N_A_6887_311#_c_11955_n 0.020688f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6796 N_Z_c_9125_n N_A_6887_311#_c_11942_n 0.0146113f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6797 N_Z_c_9700_n N_A_6887_311#_c_11942_n 0.0139315f $X=35.825 $Y=1.87 $X2=0
+ $Y2=0
cc_6798 Z N_A_6887_311#_c_11942_n 0.0238869f $X=35.005 $Y=1.785 $X2=0 $Y2=0
cc_6799 N_Z_c_9141_n N_A_6887_311#_c_11942_n 0.0174871f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6800 N_Z_c_9125_n N_A_6887_311#_c_11984_n 0.0238046f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6801 N_Z_c_9141_n N_A_6887_311#_c_11984_n 0.0025679f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6802 N_Z_c_9127_n N_A_6887_311#_c_11944_n 0.0146113f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6803 N_Z_c_10518_p N_A_6887_311#_c_11944_n 0.0238869f $X=36.115 $Y=1.87 $X2=0
+ $Y2=0
cc_6804 N_Z_c_9700_n N_A_6887_311#_c_11944_n 0.0139315f $X=35.825 $Y=1.87 $X2=0
+ $Y2=0
cc_6805 N_Z_c_9142_n N_A_6887_311#_c_11944_n 0.0174871f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6806 N_Z_c_9700_n N_A_6887_311#_c_11987_n 0.0236317f $X=35.825 $Y=1.87 $X2=0
+ $Y2=0
cc_6807 N_Z_c_9141_n N_A_6887_311#_c_11987_n 0.00259673f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6808 N_Z_c_9142_n N_A_6887_311#_c_11987_n 0.00259673f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6809 N_Z_c_9127_n N_A_6887_311#_c_11935_n 0.0521734f $X=42.085 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6810 N_Z_c_9127_n N_A_6887_311#_c_11992_n 0.0238046f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6811 N_Z_c_9142_n N_A_6887_311#_c_11992_n 0.0025679f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6812 N_Z_c_9127_n N_A_6887_311#_c_11968_n 0.0481433f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6813 N_Z_c_9127_n N_A_6887_311#_c_11998_n 0.0238869f $X=42.085 $Y=1.87
+ $X2=25.99 $Y2=0.64
cc_6814 N_Z_c_9127_n N_A_6887_311#_c_11970_n 0.0205035f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6815 N_Z_c_9127_n N_A_6887_311#_c_12005_n 0.0238869f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6816 N_Z_c_9127_n N_A_6887_311#_c_11973_n 0.0187608f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6817 N_Z_c_9125_n N_A_6887_311#_c_11936_n 0.0169532f $X=34.885 $Y=1.87 $X2=0
+ $Y2=0
cc_6818 Z N_A_6887_311#_c_11936_n 6.74054e-19 $X=35.005 $Y=1.785 $X2=0 $Y2=0
cc_6819 N_Z_c_9141_n N_A_6887_311#_c_11936_n 0.0420527f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6820 N_Z_c_9030_n N_A_6887_311#_c_11937_n 0.0192125f $X=35.805 $Y=1.215 $X2=0
+ $Y2=0
cc_6821 N_Z_c_9078_n N_A_6887_311#_c_11937_n 0.0024794f $X=35.13 $Y=1.215 $X2=0
+ $Y2=0
cc_6822 N_Z_c_10518_p N_A_6887_311#_c_11937_n 6.68271e-19 $X=36.115 $Y=1.87
+ $X2=0 $Y2=0
cc_6823 N_Z_c_9700_n N_A_6887_311#_c_11937_n 0.0151604f $X=35.825 $Y=1.87 $X2=0
+ $Y2=0
cc_6824 Z N_A_6887_311#_c_11937_n 6.68271e-19 $X=35.005 $Y=1.785 $X2=0 $Y2=0
cc_6825 N_Z_c_9141_n N_A_6887_311#_c_11937_n 0.0438531f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6826 N_Z_c_9142_n N_A_6887_311#_c_11937_n 0.0438531f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6827 N_Z_c_9127_n N_A_6887_311#_c_11938_n 0.026602f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6828 N_Z_c_10518_p N_A_6887_311#_c_11938_n 6.74054e-19 $X=36.115 $Y=1.87
+ $X2=0 $Y2=0
cc_6829 N_Z_c_9142_n N_A_6887_311#_c_11938_n 0.0383005f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6830 N_Z_c_9126_n N_A_6887_613#_M1092_s 2.15519e-19 $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6831 N_Z_c_9729_n N_A_6887_613#_M1117_s 3.28377e-19 $X=35.825 $Y=3.57 $X2=0
+ $Y2=0
cc_6832 N_Z_c_9128_n N_A_6887_613#_M1238_s 2.15519e-19 $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6833 N_Z_c_9128_n N_A_6887_613#_c_12064_n 0.0242319f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6834 N_Z_c_9142_n N_A_6887_613#_c_12065_n 0.00915958f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6835 N_Z_c_9128_n N_A_6887_613#_c_12086_n 0.020688f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6836 N_Z_c_9126_n N_A_6887_613#_c_12073_n 0.0146113f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6837 N_Z_c_9729_n N_A_6887_613#_c_12073_n 0.0139315f $X=35.825 $Y=3.57 $X2=0
+ $Y2=0
cc_6838 Z N_A_6887_613#_c_12073_n 0.0238869f $X=35.005 $Y=3.485 $X2=0 $Y2=0
cc_6839 N_Z_c_9141_n N_A_6887_613#_c_12073_n 0.0174871f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6840 N_Z_c_9126_n N_A_6887_613#_c_12115_n 0.0238046f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6841 N_Z_c_9141_n N_A_6887_613#_c_12115_n 0.0025679f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6842 N_Z_c_9128_n N_A_6887_613#_c_12075_n 0.0146113f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6843 N_Z_c_10558_p N_A_6887_613#_c_12075_n 0.0238869f $X=36.115 $Y=3.57 $X2=0
+ $Y2=0
cc_6844 N_Z_c_9729_n N_A_6887_613#_c_12075_n 0.0139315f $X=35.825 $Y=3.57 $X2=0
+ $Y2=0
cc_6845 N_Z_c_9142_n N_A_6887_613#_c_12075_n 0.0174871f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6846 N_Z_c_9729_n N_A_6887_613#_c_12118_n 0.0236317f $X=35.825 $Y=3.57 $X2=0
+ $Y2=0
cc_6847 N_Z_c_9141_n N_A_6887_613#_c_12118_n 0.00259673f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6848 N_Z_c_9142_n N_A_6887_613#_c_12118_n 0.00259673f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6849 N_Z_c_9128_n N_A_6887_613#_c_12066_n 0.0521734f $X=42.085 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6850 N_Z_c_9128_n N_A_6887_613#_c_12123_n 0.0238046f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6851 N_Z_c_9142_n N_A_6887_613#_c_12123_n 0.0025679f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6852 N_Z_c_9128_n N_A_6887_613#_c_12099_n 0.0481433f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6853 N_Z_c_9128_n N_A_6887_613#_c_12129_n 0.0238869f $X=42.085 $Y=3.57
+ $X2=25.99 $Y2=0.64
cc_6854 N_Z_c_9128_n N_A_6887_613#_c_12132_n 0.0238869f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6855 N_Z_c_9126_n N_A_6887_613#_c_12067_n 0.0169532f $X=34.885 $Y=3.57 $X2=0
+ $Y2=0
cc_6856 Z N_A_6887_613#_c_12067_n 6.74054e-19 $X=35.005 $Y=3.485 $X2=0 $Y2=0
cc_6857 N_Z_c_9141_n N_A_6887_613#_c_12067_n 0.0420527f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6858 N_Z_c_9031_n N_A_6887_613#_c_12068_n 0.0192125f $X=35.805 $Y=4.225 $X2=0
+ $Y2=0
cc_6859 N_Z_c_9079_n N_A_6887_613#_c_12068_n 0.0024794f $X=35.13 $Y=4.225 $X2=0
+ $Y2=0
cc_6860 N_Z_c_10558_p N_A_6887_613#_c_12068_n 6.68271e-19 $X=36.115 $Y=3.57
+ $X2=0 $Y2=0
cc_6861 N_Z_c_9729_n N_A_6887_613#_c_12068_n 0.0151604f $X=35.825 $Y=3.57 $X2=0
+ $Y2=0
cc_6862 Z N_A_6887_613#_c_12068_n 6.68271e-19 $X=35.005 $Y=3.485 $X2=0 $Y2=0
cc_6863 N_Z_c_9141_n N_A_6887_613#_c_12068_n 0.0438531f $X=35.03 $Y=1.7 $X2=0
+ $Y2=0
cc_6864 N_Z_c_9142_n N_A_6887_613#_c_12068_n 0.0438531f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6865 N_Z_c_9128_n N_A_6887_613#_c_12069_n 0.026602f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6866 N_Z_c_10558_p N_A_6887_613#_c_12069_n 6.74054e-19 $X=36.115 $Y=3.57
+ $X2=0 $Y2=0
cc_6867 N_Z_c_9142_n N_A_6887_613#_c_12069_n 0.0383005f $X=35.97 $Y=1.7 $X2=0
+ $Y2=0
cc_6868 N_Z_c_9128_n N_A_6887_613#_c_12102_n 0.0205035f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6869 N_Z_c_9128_n N_A_6887_613#_c_12105_n 0.0187608f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6870 N_Z_c_9127_n N_A_7937_297#_M1081_d 2.15519e-19 $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6871 Z N_A_7937_297#_M1168_d 3.28377e-19 $X=43.025 $Y=1.785 $X2=0 $Y2=0
cc_6872 N_Z_c_9129_n N_A_7937_297#_M1248_d 2.15519e-19 $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6873 N_Z_c_9127_n N_A_7937_297#_c_12200_n 0.020688f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6874 N_Z_c_9127_n N_A_7937_297#_c_12195_n 0.0242319f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6875 N_Z_c_9143_n N_A_7937_297#_c_12195_n 0.00915958f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6876 N_Z_c_9127_n N_A_7937_297#_c_12213_n 0.0481433f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6877 N_Z_c_9127_n N_A_7937_297#_c_12248_n 0.0238869f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6878 N_Z_c_9127_n N_A_7937_297#_c_12196_n 0.0521734f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6879 N_Z_c_9127_n N_A_7937_297#_c_12255_n 0.0238869f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6880 N_Z_c_9127_n N_A_7937_297#_c_12224_n 0.0146113f $X=42.085 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6881 N_Z_c_10596_p N_A_7937_297#_c_12224_n 0.0238869f $X=42.375 $Y=1.87
+ $X2=25.99 $Y2=0.51
cc_6882 Z N_A_7937_297#_c_12224_n 0.0139315f $X=43.025 $Y=1.785 $X2=25.99
+ $Y2=0.51
cc_6883 N_Z_c_9143_n N_A_7937_297#_c_12224_n 0.0174871f $X=42.23 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6884 N_Z_c_9127_n N_A_7937_297#_c_12259_n 0.0238046f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6885 N_Z_c_9143_n N_A_7937_297#_c_12259_n 0.0025679f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6886 N_Z_c_9129_n N_A_7937_297#_c_12226_n 0.0146113f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6887 N_Z_c_10602_p N_A_7937_297#_c_12226_n 0.0238869f $X=43.315 $Y=1.87 $X2=0
+ $Y2=0
cc_6888 Z N_A_7937_297#_c_12226_n 0.0139315f $X=43.025 $Y=1.785 $X2=0 $Y2=0
cc_6889 N_Z_c_9144_n N_A_7937_297#_c_12226_n 0.0174871f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6890 Z N_A_7937_297#_c_12262_n 0.0236317f $X=43.025 $Y=1.785 $X2=25.99
+ $Y2=0.64
cc_6891 N_Z_c_9143_n N_A_7937_297#_c_12262_n 0.00259673f $X=42.23 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6892 N_Z_c_9144_n N_A_7937_297#_c_12262_n 0.00259673f $X=43.17 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6893 N_Z_c_9127_n N_A_7937_297#_c_12216_n 0.0187608f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6894 N_Z_c_9127_n N_A_7937_297#_c_12219_n 0.0205035f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6895 N_Z_c_9129_n N_A_7937_297#_c_12271_n 0.0238046f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6896 N_Z_c_9144_n N_A_7937_297#_c_12271_n 0.0025679f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6897 N_Z_c_9127_n N_A_7937_297#_c_12197_n 0.026602f $X=42.085 $Y=1.87 $X2=0
+ $Y2=0
cc_6898 N_Z_c_10596_p N_A_7937_297#_c_12197_n 6.74054e-19 $X=42.375 $Y=1.87
+ $X2=0 $Y2=0
cc_6899 N_Z_c_9143_n N_A_7937_297#_c_12197_n 0.0383005f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6900 N_Z_c_9034_n N_A_7937_297#_c_12198_n 0.0192125f $X=42.805 $Y=1.215 $X2=0
+ $Y2=0
cc_6901 N_Z_c_9090_n N_A_7937_297#_c_12198_n 0.0024794f $X=43.07 $Y=1.215 $X2=0
+ $Y2=0
cc_6902 N_Z_c_10602_p N_A_7937_297#_c_12198_n 6.68271e-19 $X=43.315 $Y=1.87
+ $X2=0 $Y2=0
cc_6903 N_Z_c_10596_p N_A_7937_297#_c_12198_n 6.68271e-19 $X=42.375 $Y=1.87
+ $X2=0 $Y2=0
cc_6904 Z N_A_7937_297#_c_12198_n 0.0151604f $X=43.025 $Y=1.785 $X2=0 $Y2=0
cc_6905 N_Z_c_9143_n N_A_7937_297#_c_12198_n 0.0438531f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6906 N_Z_c_9144_n N_A_7937_297#_c_12198_n 0.0438531f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6907 N_Z_c_9129_n N_A_7937_297#_c_12199_n 0.0169532f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6908 N_Z_c_10602_p N_A_7937_297#_c_12199_n 6.74054e-19 $X=43.315 $Y=1.87
+ $X2=0 $Y2=0
cc_6909 N_Z_c_9144_n N_A_7937_297#_c_12199_n 0.0420527f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6910 N_Z_c_9128_n N_A_7937_591#_M1025_d 2.15519e-19 $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6911 Z N_A_7937_591#_M1077_d 3.28377e-19 $X=43.025 $Y=3.485 $X2=0 $Y2=0
cc_6912 N_Z_c_9130_n N_A_7937_591#_M1314_d 2.15519e-19 $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6913 N_Z_c_9128_n N_A_7937_591#_c_12328_n 0.020688f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6914 N_Z_c_9128_n N_A_7937_591#_c_12323_n 0.0242319f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6915 N_Z_c_9143_n N_A_7937_591#_c_12323_n 0.00915958f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6916 N_Z_c_9128_n N_A_7937_591#_c_12341_n 0.0481433f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6917 N_Z_c_9128_n N_A_7937_591#_c_12376_n 0.0238869f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6918 N_Z_c_9128_n N_A_7937_591#_c_12324_n 0.0521734f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6919 N_Z_c_9128_n N_A_7937_591#_c_12383_n 0.0238869f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6920 N_Z_c_9128_n N_A_7937_591#_c_12352_n 0.0146113f $X=42.085 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6921 N_Z_c_10636_p N_A_7937_591#_c_12352_n 0.0238869f $X=42.375 $Y=3.57
+ $X2=25.99 $Y2=0.51
cc_6922 Z N_A_7937_591#_c_12352_n 0.0139315f $X=43.025 $Y=3.485 $X2=25.99
+ $Y2=0.51
cc_6923 N_Z_c_9143_n N_A_7937_591#_c_12352_n 0.0174871f $X=42.23 $Y=1.7
+ $X2=25.99 $Y2=0.51
cc_6924 N_Z_c_9128_n N_A_7937_591#_c_12387_n 0.0238046f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6925 N_Z_c_9143_n N_A_7937_591#_c_12387_n 0.0025679f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6926 N_Z_c_9130_n N_A_7937_591#_c_12354_n 0.0146113f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6927 N_Z_c_10642_p N_A_7937_591#_c_12354_n 0.0238869f $X=43.315 $Y=3.57 $X2=0
+ $Y2=0
cc_6928 Z N_A_7937_591#_c_12354_n 0.0139315f $X=43.025 $Y=3.485 $X2=0 $Y2=0
cc_6929 N_Z_c_9144_n N_A_7937_591#_c_12354_n 0.0174871f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6930 Z N_A_7937_591#_c_12390_n 0.0236317f $X=43.025 $Y=3.485 $X2=25.99
+ $Y2=0.64
cc_6931 N_Z_c_9143_n N_A_7937_591#_c_12390_n 0.00259673f $X=42.23 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6932 N_Z_c_9144_n N_A_7937_591#_c_12390_n 0.00259673f $X=43.17 $Y=1.7
+ $X2=25.99 $Y2=0.64
cc_6933 N_Z_c_9130_n N_A_7937_591#_c_12391_n 0.0238046f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6934 N_Z_c_9144_n N_A_7937_591#_c_12391_n 0.0025679f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6935 N_Z_c_9128_n N_A_7937_591#_c_12344_n 0.0187608f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6936 N_Z_c_9128_n N_A_7937_591#_c_12347_n 0.0205035f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6937 N_Z_c_9128_n N_A_7937_591#_c_12325_n 0.026602f $X=42.085 $Y=3.57 $X2=0
+ $Y2=0
cc_6938 N_Z_c_10636_p N_A_7937_591#_c_12325_n 6.74054e-19 $X=42.375 $Y=3.57
+ $X2=0 $Y2=0
cc_6939 N_Z_c_9143_n N_A_7937_591#_c_12325_n 0.0383005f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6940 N_Z_c_9035_n N_A_7937_591#_c_12326_n 0.0192125f $X=42.805 $Y=4.225 $X2=0
+ $Y2=0
cc_6941 N_Z_c_9091_n N_A_7937_591#_c_12326_n 0.0024794f $X=43.07 $Y=4.225 $X2=0
+ $Y2=0
cc_6942 N_Z_c_10642_p N_A_7937_591#_c_12326_n 6.68271e-19 $X=43.315 $Y=3.57
+ $X2=0 $Y2=0
cc_6943 N_Z_c_10636_p N_A_7937_591#_c_12326_n 6.68271e-19 $X=42.375 $Y=3.57
+ $X2=0 $Y2=0
cc_6944 Z N_A_7937_591#_c_12326_n 0.0151604f $X=43.025 $Y=3.485 $X2=0 $Y2=0
cc_6945 N_Z_c_9143_n N_A_7937_591#_c_12326_n 0.0438531f $X=42.23 $Y=1.7 $X2=0
+ $Y2=0
cc_6946 N_Z_c_9144_n N_A_7937_591#_c_12326_n 0.0438531f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6947 N_Z_c_9130_n N_A_7937_591#_c_12327_n 0.0169532f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6948 N_Z_c_10642_p N_A_7937_591#_c_12327_n 6.74054e-19 $X=43.315 $Y=3.57
+ $X2=0 $Y2=0
cc_6949 N_Z_c_9144_n N_A_7937_591#_c_12327_n 0.0420527f $X=43.17 $Y=1.7 $X2=0
+ $Y2=0
cc_6950 N_Z_c_9129_n N_A_9463_311#_M1013_s 2.15519e-19 $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6951 N_Z_c_9905_n N_A_9463_311#_M1058_s 3.28377e-19 $X=48.705 $Y=1.87 $X2=0
+ $Y2=0
cc_6952 N_Z_c_9146_n N_A_9463_311#_c_12452_n 0.00915958f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6953 N_Z_c_9129_n N_A_9463_311#_c_12460_n 0.0146113f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6954 N_Z_c_9905_n N_A_9463_311#_c_12460_n 0.0139315f $X=48.705 $Y=1.87 $X2=0
+ $Y2=0
cc_6955 Z N_A_9463_311#_c_12460_n 0.0238869f $X=47.885 $Y=1.785 $X2=0 $Y2=0
cc_6956 N_Z_c_9145_n N_A_9463_311#_c_12460_n 0.0174871f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6957 N_Z_c_9129_n N_A_9463_311#_c_12502_n 0.0238046f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6958 N_Z_c_9145_n N_A_9463_311#_c_12502_n 0.0025679f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6959 N_Z_c_9905_n N_A_9463_311#_c_12462_n 0.0139315f $X=48.705 $Y=1.87 $X2=0
+ $Y2=0
cc_6960 N_Z_c_10675_p N_A_9463_311#_c_12462_n 0.0238869f $X=48.85 $Y=1.87 $X2=0
+ $Y2=0
cc_6961 N_Z_c_9146_n N_A_9463_311#_c_12462_n 0.0181912f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6962 N_Z_c_9905_n N_A_9463_311#_c_12505_n 0.0236317f $X=48.705 $Y=1.87 $X2=0
+ $Y2=0
cc_6963 N_Z_c_9145_n N_A_9463_311#_c_12505_n 0.00259673f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6964 N_Z_c_9146_n N_A_9463_311#_c_12505_n 0.00259673f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6965 N_Z_c_9146_n N_A_9463_311#_c_12510_n 0.0025679f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6966 N_Z_c_9129_n N_A_9463_311#_c_12454_n 0.0169532f $X=47.765 $Y=1.87 $X2=0
+ $Y2=0
cc_6967 Z N_A_9463_311#_c_12454_n 6.74054e-19 $X=47.885 $Y=1.785 $X2=0 $Y2=0
cc_6968 N_Z_c_9145_n N_A_9463_311#_c_12454_n 0.0420527f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6969 N_Z_c_9040_n N_A_9463_311#_c_12455_n 0.0192125f $X=48.685 $Y=1.215 $X2=0
+ $Y2=0
cc_6970 N_Z_c_9092_n N_A_9463_311#_c_12455_n 0.0024794f $X=48.01 $Y=1.215 $X2=0
+ $Y2=0
cc_6971 N_Z_c_9905_n N_A_9463_311#_c_12455_n 0.0151604f $X=48.705 $Y=1.87 $X2=0
+ $Y2=0
cc_6972 N_Z_c_10675_p N_A_9463_311#_c_12455_n 6.68271e-19 $X=48.85 $Y=1.87 $X2=0
+ $Y2=0
cc_6973 Z N_A_9463_311#_c_12455_n 6.68271e-19 $X=47.885 $Y=1.785 $X2=0 $Y2=0
cc_6974 N_Z_c_9145_n N_A_9463_311#_c_12455_n 0.0438531f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6975 N_Z_c_9146_n N_A_9463_311#_c_12455_n 0.0438531f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6976 N_Z_c_10675_p N_A_9463_311#_c_12456_n 0.00168706f $X=48.85 $Y=1.87 $X2=0
+ $Y2=0
cc_6977 N_Z_c_9146_n N_A_9463_311#_c_12456_n 0.0364724f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6978 N_Z_c_9130_n N_A_9463_613#_M1166_s 2.15519e-19 $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6979 N_Z_c_9933_n N_A_9463_613#_M1204_s 3.28377e-19 $X=48.705 $Y=3.57 $X2=0
+ $Y2=0
cc_6980 N_Z_c_9146_n N_A_9463_613#_c_12571_n 0.00915958f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6981 N_Z_c_9130_n N_A_9463_613#_c_12579_n 0.0146113f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6982 N_Z_c_9933_n N_A_9463_613#_c_12579_n 0.0139315f $X=48.705 $Y=3.57 $X2=0
+ $Y2=0
cc_6983 Z N_A_9463_613#_c_12579_n 0.0238869f $X=47.885 $Y=3.485 $X2=0 $Y2=0
cc_6984 N_Z_c_9145_n N_A_9463_613#_c_12579_n 0.0174871f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6985 N_Z_c_9130_n N_A_9463_613#_c_12621_n 0.0238046f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6986 N_Z_c_9145_n N_A_9463_613#_c_12621_n 0.0025679f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6987 N_Z_c_9933_n N_A_9463_613#_c_12581_n 0.0139315f $X=48.705 $Y=3.57 $X2=0
+ $Y2=0
cc_6988 N_Z_c_10703_p N_A_9463_613#_c_12581_n 0.0238869f $X=48.85 $Y=3.57 $X2=0
+ $Y2=0
cc_6989 N_Z_c_9146_n N_A_9463_613#_c_12581_n 0.0181912f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6990 N_Z_c_9933_n N_A_9463_613#_c_12624_n 0.0236317f $X=48.705 $Y=3.57 $X2=0
+ $Y2=0
cc_6991 N_Z_c_9145_n N_A_9463_613#_c_12624_n 0.00259673f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6992 N_Z_c_9146_n N_A_9463_613#_c_12624_n 0.00259673f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6993 N_Z_c_9146_n N_A_9463_613#_c_12629_n 0.0025679f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_6994 N_Z_c_9130_n N_A_9463_613#_c_12573_n 0.0169532f $X=47.765 $Y=3.57 $X2=0
+ $Y2=0
cc_6995 Z N_A_9463_613#_c_12573_n 6.74054e-19 $X=47.885 $Y=3.485 $X2=0 $Y2=0
cc_6996 N_Z_c_9145_n N_A_9463_613#_c_12573_n 0.0420527f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_6997 N_Z_c_9041_n N_A_9463_613#_c_12574_n 0.0192125f $X=48.685 $Y=4.225 $X2=0
+ $Y2=0
cc_6998 N_Z_c_9093_n N_A_9463_613#_c_12574_n 0.0024794f $X=48.01 $Y=4.225 $X2=0
+ $Y2=0
cc_6999 N_Z_c_9933_n N_A_9463_613#_c_12574_n 0.0151604f $X=48.705 $Y=3.57 $X2=0
+ $Y2=0
cc_7000 N_Z_c_10703_p N_A_9463_613#_c_12574_n 6.68271e-19 $X=48.85 $Y=3.57 $X2=0
+ $Y2=0
cc_7001 Z N_A_9463_613#_c_12574_n 6.68271e-19 $X=47.885 $Y=3.485 $X2=0 $Y2=0
cc_7002 N_Z_c_9145_n N_A_9463_613#_c_12574_n 0.0438531f $X=47.91 $Y=1.7 $X2=0
+ $Y2=0
cc_7003 N_Z_c_9146_n N_A_9463_613#_c_12574_n 0.0438531f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_7004 N_Z_c_10703_p N_A_9463_613#_c_12575_n 0.00168706f $X=48.85 $Y=3.57 $X2=0
+ $Y2=0
cc_7005 N_Z_c_9146_n N_A_9463_613#_c_12575_n 0.0364724f $X=48.85 $Y=1.7 $X2=0
+ $Y2=0
cc_7006 N_Z_c_9043_n N_A_119_47#_c_14050_n 0.00799417f $X=3.03 $Y=0.68 $X2=0
+ $Y2=0
cc_7007 N_Z_M1053_s N_A_119_47#_c_14052_n 0.00165831f $X=2.895 $Y=0.33 $X2=0
+ $Y2=0
cc_7008 N_Z_c_9004_n N_A_119_47#_c_14052_n 0.00133192f $X=3.705 $Y=1.215 $X2=0
+ $Y2=0
cc_7009 N_Z_c_9043_n N_A_119_47#_c_14052_n 0.0157607f $X=3.03 $Y=0.68 $X2=0
+ $Y2=0
cc_7010 N_Z_c_9046_n N_A_119_47#_c_14052_n 0.00293855f $X=3.13 $Y=1.215 $X2=0
+ $Y2=0
cc_7011 N_Z_c_9004_n N_A_119_47#_c_14077_n 0.00918654f $X=3.705 $Y=1.215 $X2=0
+ $Y2=0
cc_7012 N_Z_M1105_s N_A_119_47#_c_14054_n 0.00165831f $X=3.735 $Y=0.33 $X2=25.99
+ $Y2=4.8
cc_7013 N_Z_c_9004_n N_A_119_47#_c_14054_n 0.00405549f $X=3.705 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7014 N_Z_c_9006_n N_A_119_47#_c_14054_n 0.015949f $X=3.87 $Y=0.68 $X2=25.99
+ $Y2=4.8
cc_7015 N_Z_c_9048_n N_A_119_47#_c_14054_n 0.00443806f $X=3.97 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7016 N_Z_c_9048_n N_A_119_47#_c_14055_n 0.00158445f $X=3.97 $Y=1.215
+ $X2=25.99 $Y2=4.93
cc_7017 N_Z_c_9044_n N_A_119_911#_c_14132_n 0.00799417f $X=3.03 $Y=4.76 $X2=0
+ $Y2=0
cc_7018 N_Z_M1070_d N_A_119_911#_c_14134_n 0.00165831f $X=2.895 $Y=4.59 $X2=0
+ $Y2=0
cc_7019 N_Z_c_9005_n N_A_119_911#_c_14134_n 0.00133192f $X=3.705 $Y=4.225 $X2=0
+ $Y2=0
cc_7020 N_Z_c_9044_n N_A_119_911#_c_14134_n 0.0157607f $X=3.03 $Y=4.76 $X2=0
+ $Y2=0
cc_7021 N_Z_c_9047_n N_A_119_911#_c_14134_n 0.00293855f $X=3.13 $Y=4.225 $X2=0
+ $Y2=0
cc_7022 N_Z_c_9005_n N_A_119_911#_c_14156_n 0.00918654f $X=3.705 $Y=4.225 $X2=0
+ $Y2=0
cc_7023 N_Z_M1236_d N_A_119_911#_c_14136_n 0.00165831f $X=3.735 $Y=4.59
+ $X2=25.99 $Y2=0.64
cc_7024 N_Z_c_9005_n N_A_119_911#_c_14136_n 0.00405549f $X=3.705 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7025 N_Z_c_9007_n N_A_119_911#_c_14136_n 0.015949f $X=3.87 $Y=4.76 $X2=25.99
+ $Y2=0.64
cc_7026 N_Z_c_9049_n N_A_119_911#_c_14136_n 0.00443806f $X=3.97 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7027 N_Z_c_9049_n N_A_119_911#_c_14137_n 0.00158445f $X=3.97 $Y=4.225
+ $X2=25.99 $Y2=4.8
cc_7028 N_Z_c_9050_n N_A_1693_66#_c_14211_n 0.00158445f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_7029 N_Z_M1039_d N_A_1693_66#_c_14212_n 0.00165831f $X=8.875 $Y=0.33 $X2=0
+ $Y2=0
cc_7030 N_Z_c_9008_n N_A_1693_66#_c_14212_n 0.015949f $X=9.01 $Y=0.68 $X2=0
+ $Y2=0
cc_7031 N_Z_c_9010_n N_A_1693_66#_c_14212_n 0.00405549f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_7032 N_Z_c_9050_n N_A_1693_66#_c_14212_n 0.00443806f $X=8.91 $Y=1.215 $X2=0
+ $Y2=0
cc_7033 N_Z_c_9010_n N_A_1693_66#_c_14233_n 0.00918654f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_7034 N_Z_M1093_d N_A_1693_66#_c_14214_n 0.00165831f $X=9.715 $Y=0.33 $X2=0
+ $Y2=0
cc_7035 N_Z_c_9010_n N_A_1693_66#_c_14214_n 0.00133192f $X=9.585 $Y=1.215 $X2=0
+ $Y2=0
cc_7036 N_Z_c_9052_n N_A_1693_66#_c_14214_n 0.00293855f $X=9.75 $Y=1.215 $X2=0
+ $Y2=0
cc_7037 N_Z_c_9054_n N_A_1693_66#_c_14214_n 0.0157607f $X=9.85 $Y=0.68 $X2=0
+ $Y2=0
cc_7038 N_Z_c_9054_n N_A_1693_66#_c_14217_n 0.00799417f $X=9.85 $Y=0.68 $X2=0
+ $Y2=0
cc_7039 N_Z_c_9051_n N_A_1693_918#_c_14295_n 0.00158445f $X=8.91 $Y=4.225 $X2=0
+ $Y2=0
cc_7040 N_Z_M1027_d N_A_1693_918#_c_14296_n 0.00165831f $X=8.875 $Y=4.59 $X2=0
+ $Y2=0
cc_7041 N_Z_c_9009_n N_A_1693_918#_c_14296_n 0.015949f $X=9.01 $Y=4.76 $X2=0
+ $Y2=0
cc_7042 N_Z_c_9011_n N_A_1693_918#_c_14296_n 0.00405549f $X=9.585 $Y=4.225 $X2=0
+ $Y2=0
cc_7043 N_Z_c_9051_n N_A_1693_918#_c_14296_n 0.00443806f $X=8.91 $Y=4.225 $X2=0
+ $Y2=0
cc_7044 N_Z_c_9011_n N_A_1693_918#_c_14317_n 0.00918654f $X=9.585 $Y=4.225 $X2=0
+ $Y2=0
cc_7045 N_Z_M1096_d N_A_1693_918#_c_14298_n 0.00165831f $X=9.715 $Y=4.59 $X2=0
+ $Y2=0
cc_7046 N_Z_c_9011_n N_A_1693_918#_c_14298_n 0.00133192f $X=9.585 $Y=4.225 $X2=0
+ $Y2=0
cc_7047 N_Z_c_9053_n N_A_1693_918#_c_14298_n 0.00293855f $X=9.75 $Y=4.225 $X2=0
+ $Y2=0
cc_7048 N_Z_c_9055_n N_A_1693_918#_c_14298_n 0.0157607f $X=9.85 $Y=4.76 $X2=0
+ $Y2=0
cc_7049 N_Z_c_9055_n N_A_1693_918#_c_14301_n 0.00799417f $X=9.85 $Y=4.76 $X2=0
+ $Y2=0
cc_7050 N_Z_c_9057_n N_A_2695_47#_c_14378_n 0.00799417f $X=15.91 $Y=0.68 $X2=0
+ $Y2=0
cc_7051 N_Z_M1035_d N_A_2695_47#_c_14380_n 0.00165831f $X=15.775 $Y=0.33 $X2=0
+ $Y2=0
cc_7052 N_Z_c_9014_n N_A_2695_47#_c_14380_n 0.00133192f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_7053 N_Z_c_9057_n N_A_2695_47#_c_14380_n 0.0157607f $X=15.91 $Y=0.68 $X2=0
+ $Y2=0
cc_7054 N_Z_c_9060_n N_A_2695_47#_c_14380_n 0.00293855f $X=16.01 $Y=1.215 $X2=0
+ $Y2=0
cc_7055 N_Z_c_9014_n N_A_2695_47#_c_14405_n 0.00918654f $X=16.585 $Y=1.215 $X2=0
+ $Y2=0
cc_7056 N_Z_M1108_d N_A_2695_47#_c_14382_n 0.00165831f $X=16.615 $Y=0.33
+ $X2=25.99 $Y2=4.8
cc_7057 N_Z_c_9014_n N_A_2695_47#_c_14382_n 0.00405549f $X=16.585 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7058 N_Z_c_9016_n N_A_2695_47#_c_14382_n 0.015949f $X=16.75 $Y=0.68 $X2=25.99
+ $Y2=4.8
cc_7059 N_Z_c_9062_n N_A_2695_47#_c_14382_n 0.00443806f $X=16.85 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7060 N_Z_c_9062_n N_A_2695_47#_c_14383_n 0.00158445f $X=16.85 $Y=1.215
+ $X2=25.99 $Y2=4.93
cc_7061 N_Z_c_9058_n N_A_2695_911#_c_14460_n 0.00799417f $X=15.91 $Y=4.76 $X2=0
+ $Y2=0
cc_7062 N_Z_M1010_s N_A_2695_911#_c_14462_n 0.00165831f $X=15.775 $Y=4.59 $X2=0
+ $Y2=0
cc_7063 N_Z_c_9015_n N_A_2695_911#_c_14462_n 0.00133192f $X=16.585 $Y=4.225
+ $X2=0 $Y2=0
cc_7064 N_Z_c_9058_n N_A_2695_911#_c_14462_n 0.0157607f $X=15.91 $Y=4.76 $X2=0
+ $Y2=0
cc_7065 N_Z_c_9061_n N_A_2695_911#_c_14462_n 0.00293855f $X=16.01 $Y=4.225 $X2=0
+ $Y2=0
cc_7066 N_Z_c_9015_n N_A_2695_911#_c_14484_n 0.00918654f $X=16.585 $Y=4.225
+ $X2=0 $Y2=0
cc_7067 N_Z_M1263_s N_A_2695_911#_c_14464_n 0.00165831f $X=16.615 $Y=4.59
+ $X2=25.99 $Y2=0.64
cc_7068 N_Z_c_9015_n N_A_2695_911#_c_14464_n 0.00405549f $X=16.585 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7069 N_Z_c_9017_n N_A_2695_911#_c_14464_n 0.015949f $X=16.75 $Y=4.76
+ $X2=25.99 $Y2=0.64
cc_7070 N_Z_c_9063_n N_A_2695_911#_c_14464_n 0.00443806f $X=16.85 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7071 N_Z_c_9063_n N_A_2695_911#_c_14465_n 0.00158445f $X=16.85 $Y=4.225
+ $X2=25.99 $Y2=4.8
cc_7072 N_Z_c_9064_n N_A_4269_66#_c_14539_n 0.00158445f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_7073 N_Z_M1030_s N_A_4269_66#_c_14540_n 0.00165831f $X=21.755 $Y=0.33 $X2=0
+ $Y2=0
cc_7074 N_Z_c_9018_n N_A_4269_66#_c_14540_n 0.015949f $X=21.89 $Y=0.68 $X2=0
+ $Y2=0
cc_7075 N_Z_c_9020_n N_A_4269_66#_c_14540_n 0.00405549f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_7076 N_Z_c_9064_n N_A_4269_66#_c_14540_n 0.00443806f $X=21.79 $Y=1.215 $X2=0
+ $Y2=0
cc_7077 N_Z_c_9020_n N_A_4269_66#_c_14561_n 0.00918654f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_7078 N_Z_M1059_s N_A_4269_66#_c_14542_n 0.00165831f $X=22.595 $Y=0.33 $X2=0
+ $Y2=0
cc_7079 N_Z_c_9020_n N_A_4269_66#_c_14542_n 0.00133192f $X=22.465 $Y=1.215 $X2=0
+ $Y2=0
cc_7080 N_Z_c_9066_n N_A_4269_66#_c_14542_n 0.00293855f $X=22.63 $Y=1.215 $X2=0
+ $Y2=0
cc_7081 N_Z_c_9068_n N_A_4269_66#_c_14542_n 0.0157607f $X=22.73 $Y=0.68 $X2=0
+ $Y2=0
cc_7082 N_Z_c_9068_n N_A_4269_66#_c_14545_n 0.00799417f $X=22.73 $Y=0.68 $X2=0
+ $Y2=0
cc_7083 N_Z_c_9065_n N_A_4269_918#_c_14623_n 0.00158445f $X=21.79 $Y=4.225 $X2=0
+ $Y2=0
cc_7084 N_Z_M1047_s N_A_4269_918#_c_14624_n 0.00165831f $X=21.755 $Y=4.59 $X2=0
+ $Y2=0
cc_7085 N_Z_c_9019_n N_A_4269_918#_c_14624_n 0.015949f $X=21.89 $Y=4.76 $X2=0
+ $Y2=0
cc_7086 N_Z_c_9021_n N_A_4269_918#_c_14624_n 0.00405549f $X=22.465 $Y=4.225
+ $X2=0 $Y2=0
cc_7087 N_Z_c_9065_n N_A_4269_918#_c_14624_n 0.00443806f $X=21.79 $Y=4.225 $X2=0
+ $Y2=0
cc_7088 N_Z_c_9021_n N_A_4269_918#_c_14645_n 0.00918654f $X=22.465 $Y=4.225
+ $X2=0 $Y2=0
cc_7089 N_Z_M1316_s N_A_4269_918#_c_14626_n 0.00165831f $X=22.595 $Y=4.59 $X2=0
+ $Y2=0
cc_7090 N_Z_c_9021_n N_A_4269_918#_c_14626_n 0.00133192f $X=22.465 $Y=4.225
+ $X2=0 $Y2=0
cc_7091 N_Z_c_9067_n N_A_4269_918#_c_14626_n 0.00293855f $X=22.63 $Y=4.225 $X2=0
+ $Y2=0
cc_7092 N_Z_c_9069_n N_A_4269_918#_c_14626_n 0.0157607f $X=22.73 $Y=4.76 $X2=0
+ $Y2=0
cc_7093 N_Z_c_9069_n N_A_4269_918#_c_14629_n 0.00799417f $X=22.73 $Y=4.76 $X2=0
+ $Y2=0
cc_7094 N_Z_c_9071_n N_A_5363_47#_c_14706_n 0.00799417f $X=29.25 $Y=0.68 $X2=0
+ $Y2=0
cc_7095 N_Z_M1154_d N_A_5363_47#_c_14708_n 0.00165831f $X=29.115 $Y=0.33 $X2=0
+ $Y2=0
cc_7096 N_Z_c_9024_n N_A_5363_47#_c_14708_n 0.00133192f $X=29.925 $Y=1.215 $X2=0
+ $Y2=0
cc_7097 N_Z_c_9071_n N_A_5363_47#_c_14708_n 0.0157607f $X=29.25 $Y=0.68 $X2=0
+ $Y2=0
cc_7098 N_Z_c_9074_n N_A_5363_47#_c_14708_n 0.00293855f $X=29.35 $Y=1.215 $X2=0
+ $Y2=0
cc_7099 N_Z_c_9024_n N_A_5363_47#_c_14733_n 0.00918654f $X=29.925 $Y=1.215 $X2=0
+ $Y2=0
cc_7100 N_Z_M1205_d N_A_5363_47#_c_14710_n 0.00165831f $X=29.955 $Y=0.33
+ $X2=25.99 $Y2=4.8
cc_7101 N_Z_c_9024_n N_A_5363_47#_c_14710_n 0.00405549f $X=29.925 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7102 N_Z_c_9026_n N_A_5363_47#_c_14710_n 0.015949f $X=30.09 $Y=0.68 $X2=25.99
+ $Y2=4.8
cc_7103 N_Z_c_9076_n N_A_5363_47#_c_14710_n 0.00443806f $X=30.19 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7104 N_Z_c_9076_n N_A_5363_47#_c_14711_n 0.00158445f $X=30.19 $Y=1.215
+ $X2=25.99 $Y2=4.93
cc_7105 N_Z_c_9072_n N_A_5363_911#_c_14788_n 0.00799417f $X=29.25 $Y=4.76 $X2=0
+ $Y2=0
cc_7106 N_Z_M1044_s N_A_5363_911#_c_14790_n 0.00165831f $X=29.115 $Y=4.59 $X2=0
+ $Y2=0
cc_7107 N_Z_c_9025_n N_A_5363_911#_c_14790_n 0.00133192f $X=29.925 $Y=4.225
+ $X2=0 $Y2=0
cc_7108 N_Z_c_9072_n N_A_5363_911#_c_14790_n 0.0157607f $X=29.25 $Y=4.76 $X2=0
+ $Y2=0
cc_7109 N_Z_c_9075_n N_A_5363_911#_c_14790_n 0.00293855f $X=29.35 $Y=4.225 $X2=0
+ $Y2=0
cc_7110 N_Z_c_9025_n N_A_5363_911#_c_14812_n 0.00918654f $X=29.925 $Y=4.225
+ $X2=0 $Y2=0
cc_7111 N_Z_M1218_s N_A_5363_911#_c_14792_n 0.00165831f $X=29.955 $Y=4.59
+ $X2=25.99 $Y2=0.64
cc_7112 N_Z_c_9025_n N_A_5363_911#_c_14792_n 0.00405549f $X=29.925 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7113 N_Z_c_9027_n N_A_5363_911#_c_14792_n 0.015949f $X=30.09 $Y=4.76
+ $X2=25.99 $Y2=0.64
cc_7114 N_Z_c_9077_n N_A_5363_911#_c_14792_n 0.00443806f $X=30.19 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7115 N_Z_c_9077_n N_A_5363_911#_c_14793_n 0.00158445f $X=30.19 $Y=4.225
+ $X2=25.99 $Y2=4.8
cc_7116 N_Z_c_9078_n N_A_6937_66#_c_14867_n 0.00158445f $X=35.13 $Y=1.215 $X2=0
+ $Y2=0
cc_7117 N_Z_M1175_s N_A_6937_66#_c_14868_n 0.00165831f $X=35.095 $Y=0.33 $X2=0
+ $Y2=0
cc_7118 N_Z_c_9028_n N_A_6937_66#_c_14868_n 0.015949f $X=35.23 $Y=0.68 $X2=0
+ $Y2=0
cc_7119 N_Z_c_9030_n N_A_6937_66#_c_14868_n 0.00405549f $X=35.805 $Y=1.215 $X2=0
+ $Y2=0
cc_7120 N_Z_c_9078_n N_A_6937_66#_c_14868_n 0.00443806f $X=35.13 $Y=1.215 $X2=0
+ $Y2=0
cc_7121 N_Z_c_9030_n N_A_6937_66#_c_14889_n 0.00918654f $X=35.805 $Y=1.215 $X2=0
+ $Y2=0
cc_7122 N_Z_M1220_s N_A_6937_66#_c_14870_n 0.00165831f $X=35.935 $Y=0.33 $X2=0
+ $Y2=0
cc_7123 N_Z_c_9030_n N_A_6937_66#_c_14870_n 0.00133192f $X=35.805 $Y=1.215 $X2=0
+ $Y2=0
cc_7124 N_Z_c_9080_n N_A_6937_66#_c_14870_n 0.00293855f $X=35.97 $Y=1.215 $X2=0
+ $Y2=0
cc_7125 N_Z_c_9082_n N_A_6937_66#_c_14870_n 0.0157607f $X=36.07 $Y=0.68 $X2=0
+ $Y2=0
cc_7126 N_Z_c_9082_n N_A_6937_66#_c_14873_n 0.00799417f $X=36.07 $Y=0.68 $X2=0
+ $Y2=0
cc_7127 N_Z_c_9079_n N_A_6937_918#_c_14951_n 0.00158445f $X=35.13 $Y=4.225 $X2=0
+ $Y2=0
cc_7128 N_Z_M1149_s N_A_6937_918#_c_14952_n 0.00165831f $X=35.095 $Y=4.59 $X2=0
+ $Y2=0
cc_7129 N_Z_c_9029_n N_A_6937_918#_c_14952_n 0.015949f $X=35.23 $Y=4.76 $X2=0
+ $Y2=0
cc_7130 N_Z_c_9031_n N_A_6937_918#_c_14952_n 0.00405549f $X=35.805 $Y=4.225
+ $X2=0 $Y2=0
cc_7131 N_Z_c_9079_n N_A_6937_918#_c_14952_n 0.00443806f $X=35.13 $Y=4.225 $X2=0
+ $Y2=0
cc_7132 N_Z_c_9031_n N_A_6937_918#_c_14973_n 0.00918654f $X=35.805 $Y=4.225
+ $X2=0 $Y2=0
cc_7133 N_Z_M1242_s N_A_6937_918#_c_14954_n 0.00165831f $X=35.935 $Y=4.59 $X2=0
+ $Y2=0
cc_7134 N_Z_c_9031_n N_A_6937_918#_c_14954_n 0.00133192f $X=35.805 $Y=4.225
+ $X2=0 $Y2=0
cc_7135 N_Z_c_9081_n N_A_6937_918#_c_14954_n 0.00293855f $X=35.97 $Y=4.225 $X2=0
+ $Y2=0
cc_7136 N_Z_c_9083_n N_A_6937_918#_c_14954_n 0.0157607f $X=36.07 $Y=4.76 $X2=0
+ $Y2=0
cc_7137 N_Z_c_9083_n N_A_6937_918#_c_14957_n 0.00799417f $X=36.07 $Y=4.76 $X2=0
+ $Y2=0
cc_7138 N_Z_c_9085_n N_A_7939_47#_c_15034_n 0.00799417f $X=42.13 $Y=0.68 $X2=0
+ $Y2=0
cc_7139 N_Z_M1202_s N_A_7939_47#_c_15036_n 0.00165831f $X=41.995 $Y=0.33 $X2=0
+ $Y2=0
cc_7140 N_Z_c_9034_n N_A_7939_47#_c_15036_n 0.00133192f $X=42.805 $Y=1.215 $X2=0
+ $Y2=0
cc_7141 N_Z_c_9085_n N_A_7939_47#_c_15036_n 0.0157607f $X=42.13 $Y=0.68 $X2=0
+ $Y2=0
cc_7142 N_Z_c_9088_n N_A_7939_47#_c_15036_n 0.00293855f $X=42.23 $Y=1.215 $X2=0
+ $Y2=0
cc_7143 N_Z_c_9034_n N_A_7939_47#_c_15061_n 0.00918654f $X=42.805 $Y=1.215 $X2=0
+ $Y2=0
cc_7144 N_Z_M1244_s N_A_7939_47#_c_15038_n 0.00165831f $X=42.835 $Y=0.33
+ $X2=25.99 $Y2=4.8
cc_7145 N_Z_c_9034_n N_A_7939_47#_c_15038_n 0.00405549f $X=42.805 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7146 N_Z_c_9036_n N_A_7939_47#_c_15038_n 0.015949f $X=42.97 $Y=0.68 $X2=25.99
+ $Y2=4.8
cc_7147 N_Z_c_9090_n N_A_7939_47#_c_15038_n 0.00443806f $X=43.07 $Y=1.215
+ $X2=25.99 $Y2=4.8
cc_7148 N_Z_c_9090_n N_A_7939_47#_c_15039_n 0.00158445f $X=43.07 $Y=1.215
+ $X2=25.99 $Y2=4.93
cc_7149 N_Z_c_9086_n N_A_7939_911#_c_15116_n 0.00799417f $X=42.13 $Y=4.76 $X2=0
+ $Y2=0
cc_7150 N_Z_M1005_s N_A_7939_911#_c_15118_n 0.00165831f $X=41.995 $Y=4.59 $X2=0
+ $Y2=0
cc_7151 N_Z_c_9035_n N_A_7939_911#_c_15118_n 0.00133192f $X=42.805 $Y=4.225
+ $X2=0 $Y2=0
cc_7152 N_Z_c_9086_n N_A_7939_911#_c_15118_n 0.0157607f $X=42.13 $Y=4.76 $X2=0
+ $Y2=0
cc_7153 N_Z_c_9089_n N_A_7939_911#_c_15118_n 0.00293855f $X=42.23 $Y=4.225 $X2=0
+ $Y2=0
cc_7154 N_Z_c_9035_n N_A_7939_911#_c_15140_n 0.00918654f $X=42.805 $Y=4.225
+ $X2=0 $Y2=0
cc_7155 N_Z_M1162_s N_A_7939_911#_c_15120_n 0.00165831f $X=42.835 $Y=4.59
+ $X2=25.99 $Y2=0.64
cc_7156 N_Z_c_9035_n N_A_7939_911#_c_15120_n 0.00405549f $X=42.805 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7157 N_Z_c_9037_n N_A_7939_911#_c_15120_n 0.015949f $X=42.97 $Y=4.76
+ $X2=25.99 $Y2=0.64
cc_7158 N_Z_c_9091_n N_A_7939_911#_c_15120_n 0.00443806f $X=43.07 $Y=4.225
+ $X2=25.99 $Y2=0.64
cc_7159 N_Z_c_9091_n N_A_7939_911#_c_15121_n 0.00158445f $X=43.07 $Y=4.225
+ $X2=25.99 $Y2=4.8
cc_7160 N_Z_c_9092_n N_A_9513_66#_c_15195_n 0.00158445f $X=48.01 $Y=1.215 $X2=0
+ $Y2=0
cc_7161 N_Z_M1003_s N_A_9513_66#_c_15196_n 0.00165831f $X=47.975 $Y=0.33 $X2=0
+ $Y2=0
cc_7162 N_Z_c_9038_n N_A_9513_66#_c_15196_n 0.015949f $X=48.11 $Y=0.68 $X2=0
+ $Y2=0
cc_7163 N_Z_c_9040_n N_A_9513_66#_c_15196_n 0.00405549f $X=48.685 $Y=1.215 $X2=0
+ $Y2=0
cc_7164 N_Z_c_9092_n N_A_9513_66#_c_15196_n 0.00443806f $X=48.01 $Y=1.215 $X2=0
+ $Y2=0
cc_7165 N_Z_c_9040_n N_A_9513_66#_c_15217_n 0.00918654f $X=48.685 $Y=1.215 $X2=0
+ $Y2=0
cc_7166 N_Z_M1253_s N_A_9513_66#_c_15198_n 0.00165831f $X=48.815 $Y=0.33 $X2=0
+ $Y2=0
cc_7167 N_Z_c_9040_n N_A_9513_66#_c_15198_n 0.00133192f $X=48.685 $Y=1.215 $X2=0
+ $Y2=0
cc_7168 N_Z_c_9094_n N_A_9513_66#_c_15198_n 0.00293855f $X=48.85 $Y=1.215 $X2=0
+ $Y2=0
cc_7169 N_Z_c_9096_n N_A_9513_66#_c_15198_n 0.0157607f $X=48.95 $Y=0.68 $X2=0
+ $Y2=0
cc_7170 N_Z_c_9096_n N_A_9513_66#_c_15201_n 0.00799417f $X=48.95 $Y=0.68 $X2=0
+ $Y2=0
cc_7171 N_Z_c_9093_n N_A_9513_918#_c_15279_n 0.00158445f $X=48.01 $Y=4.225 $X2=0
+ $Y2=0
cc_7172 N_Z_M1104_d N_A_9513_918#_c_15280_n 0.00165831f $X=47.975 $Y=4.59 $X2=0
+ $Y2=0
cc_7173 N_Z_c_9039_n N_A_9513_918#_c_15280_n 0.015949f $X=48.11 $Y=4.76 $X2=0
+ $Y2=0
cc_7174 N_Z_c_9041_n N_A_9513_918#_c_15280_n 0.00405549f $X=48.685 $Y=4.225
+ $X2=0 $Y2=0
cc_7175 N_Z_c_9093_n N_A_9513_918#_c_15280_n 0.00443806f $X=48.01 $Y=4.225 $X2=0
+ $Y2=0
cc_7176 N_Z_c_9041_n N_A_9513_918#_c_15301_n 0.00918654f $X=48.685 $Y=4.225
+ $X2=0 $Y2=0
cc_7177 N_Z_M1197_d N_A_9513_918#_c_15282_n 0.00165831f $X=48.815 $Y=4.59 $X2=0
+ $Y2=0
cc_7178 N_Z_c_9041_n N_A_9513_918#_c_15282_n 0.00133192f $X=48.685 $Y=4.225
+ $X2=0 $Y2=0
cc_7179 N_Z_c_9095_n N_A_9513_918#_c_15282_n 0.00293855f $X=48.85 $Y=4.225 $X2=0
+ $Y2=0
cc_7180 N_Z_c_9097_n N_A_9513_918#_c_15282_n 0.0157607f $X=48.95 $Y=4.76 $X2=0
+ $Y2=0
cc_7181 N_Z_c_9097_n N_A_9513_918#_c_15285_n 0.00799417f $X=48.95 $Y=4.76 $X2=0
+ $Y2=0
cc_7182 N_A_1643_311#_c_10901_n N_A_1643_613#_c_11032_n 0.00460759f $X=9.28
+ $Y=1.7 $X2=0 $Y2=0
cc_7183 N_A_1643_311#_c_10897_n N_A_1693_66#_c_14216_n 0.0147893f $X=11.045
+ $Y=1.58 $X2=0 $Y2=0
cc_7184 N_A_1643_311#_c_10897_n N_A_1693_66#_c_14217_n 0.00239279f $X=11.045
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7185 N_A_1643_311#_c_10898_n N_A_1693_66#_c_14217_n 0.00761509f $X=10.385
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7186 N_A_1643_311#_c_10923_n N_A_1693_66#_c_14219_n 6.95815e-19 $X=11.21
+ $Y=1.66 $X2=0 $Y2=0
cc_7187 N_A_1643_613#_c_11028_n N_A_1693_918#_c_14300_n 0.0147893f $X=11.045
+ $Y=3.86 $X2=0 $Y2=0
cc_7188 N_A_1643_613#_c_11028_n N_A_1693_918#_c_14301_n 0.00239279f $X=11.045
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7189 N_A_1643_613#_c_11029_n N_A_1693_918#_c_14301_n 0.00761509f $X=10.385
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7190 N_A_1643_613#_c_11054_n N_A_1693_918#_c_14302_n 6.95815e-19 $X=11.21
+ $Y=3.78 $X2=0 $Y2=0
cc_7191 N_A_2693_297#_c_11162_n N_A_2693_591#_c_11290_n 0.00460759f $X=16.48
+ $Y=1.7 $X2=0 $Y2=0
cc_7192 N_A_2693_297#_c_11159_n N_A_2695_47#_c_14378_n 0.0247972f $X=15.375
+ $Y=1.58 $X2=25.99 $Y2=1.73
cc_7193 N_A_2693_297#_c_11173_n N_A_2695_47#_c_14384_n 6.95815e-19 $X=14.55
+ $Y=1.66 $X2=0 $Y2=0
cc_7194 N_A_2693_591#_c_11287_n N_A_2695_911#_c_14460_n 0.0247972f $X=15.375
+ $Y=3.86 $X2=0 $Y2=0
cc_7195 N_A_2693_591#_c_11301_n N_A_2695_911#_c_14467_n 6.95815e-19 $X=14.55
+ $Y=3.78 $X2=0 $Y2=0
cc_7196 N_A_4219_311#_c_11419_n N_A_4219_613#_c_11550_n 0.00460759f $X=22.16
+ $Y=1.7 $X2=0 $Y2=0
cc_7197 N_A_4219_311#_c_11415_n N_A_4269_66#_c_14544_n 0.0147893f $X=23.925
+ $Y=1.58 $X2=0 $Y2=0
cc_7198 N_A_4219_311#_c_11415_n N_A_4269_66#_c_14545_n 0.00239279f $X=23.925
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7199 N_A_4219_311#_c_11416_n N_A_4269_66#_c_14545_n 0.00761509f $X=23.265
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7200 N_A_4219_311#_c_11441_n N_A_4269_66#_c_14547_n 6.95815e-19 $X=24.09
+ $Y=1.66 $X2=0 $Y2=0
cc_7201 N_A_4219_613#_c_11546_n N_A_4269_918#_c_14628_n 0.0147893f $X=23.925
+ $Y=3.86 $X2=0 $Y2=0
cc_7202 N_A_4219_613#_c_11546_n N_A_4269_918#_c_14629_n 0.00239279f $X=23.925
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7203 N_A_4219_613#_c_11547_n N_A_4269_918#_c_14629_n 0.00761509f $X=23.265
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7204 N_A_4219_613#_c_11572_n N_A_4269_918#_c_14630_n 6.95815e-19 $X=24.09
+ $Y=3.78 $X2=0 $Y2=0
cc_7205 N_A_5361_297#_c_11680_n N_A_5361_591#_c_11808_n 0.00460759f $X=29.82
+ $Y=1.7 $X2=0 $Y2=0
cc_7206 N_A_5361_297#_c_11677_n N_A_5363_47#_c_14706_n 0.0247972f $X=28.715
+ $Y=1.58 $X2=25.99 $Y2=1.73
cc_7207 N_A_5361_297#_c_11691_n N_A_5363_47#_c_14712_n 6.95815e-19 $X=27.89
+ $Y=1.66 $X2=0 $Y2=0
cc_7208 N_A_5361_591#_c_11805_n N_A_5363_911#_c_14788_n 0.0247972f $X=28.715
+ $Y=3.86 $X2=0 $Y2=0
cc_7209 N_A_5361_591#_c_11819_n N_A_5363_911#_c_14795_n 6.95815e-19 $X=27.89
+ $Y=3.78 $X2=0 $Y2=0
cc_7210 N_A_6887_311#_c_11937_n N_A_6887_613#_c_12068_n 0.00460759f $X=35.5
+ $Y=1.7 $X2=0 $Y2=0
cc_7211 N_A_6887_311#_c_11933_n N_A_6937_66#_c_14872_n 0.0147893f $X=37.265
+ $Y=1.58 $X2=0 $Y2=0
cc_7212 N_A_6887_311#_c_11933_n N_A_6937_66#_c_14873_n 0.00239279f $X=37.265
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7213 N_A_6887_311#_c_11934_n N_A_6937_66#_c_14873_n 0.00761509f $X=36.605
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7214 N_A_6887_311#_c_11959_n N_A_6937_66#_c_14875_n 6.95815e-19 $X=37.43
+ $Y=1.66 $X2=0 $Y2=0
cc_7215 N_A_6887_613#_c_12064_n N_A_6937_918#_c_14956_n 0.0147893f $X=37.265
+ $Y=3.86 $X2=0 $Y2=0
cc_7216 N_A_6887_613#_c_12064_n N_A_6937_918#_c_14957_n 0.00239279f $X=37.265
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7217 N_A_6887_613#_c_12065_n N_A_6937_918#_c_14957_n 0.00761509f $X=36.605
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7218 N_A_6887_613#_c_12090_n N_A_6937_918#_c_14958_n 6.95815e-19 $X=37.43
+ $Y=3.78 $X2=0 $Y2=0
cc_7219 N_A_7937_297#_c_12198_n N_A_7937_591#_c_12326_n 0.00460759f $X=42.7
+ $Y=1.7 $X2=0 $Y2=0
cc_7220 N_A_7937_297#_c_12195_n N_A_7939_47#_c_15034_n 0.0247972f $X=41.595
+ $Y=1.58 $X2=25.99 $Y2=1.73
cc_7221 N_A_7937_297#_c_12209_n N_A_7939_47#_c_15040_n 6.95815e-19 $X=40.77
+ $Y=1.66 $X2=0 $Y2=0
cc_7222 N_A_7937_591#_c_12323_n N_A_7939_911#_c_15116_n 0.0247972f $X=41.595
+ $Y=3.86 $X2=0 $Y2=0
cc_7223 N_A_7937_591#_c_12337_n N_A_7939_911#_c_15123_n 6.95815e-19 $X=40.77
+ $Y=3.78 $X2=0 $Y2=0
cc_7224 N_A_9463_311#_c_12455_n N_A_9463_613#_c_12574_n 0.00460759f $X=48.38
+ $Y=1.7 $X2=0 $Y2=0
cc_7225 N_A_9463_311#_c_12451_n N_A_9513_66#_c_15200_n 0.0147893f $X=50.145
+ $Y=1.58 $X2=0 $Y2=0
cc_7226 N_A_9463_311#_c_12451_n N_A_9513_66#_c_15201_n 0.00239279f $X=50.145
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7227 N_A_9463_311#_c_12452_n N_A_9513_66#_c_15201_n 0.00761509f $X=49.485
+ $Y=1.58 $X2=25.99 $Y2=3.23
cc_7228 N_A_9463_311#_c_12477_n N_A_9513_66#_c_15203_n 6.95815e-19 $X=50.31
+ $Y=1.66 $X2=0 $Y2=0
cc_7229 N_A_9463_613#_c_12570_n N_A_9513_918#_c_15284_n 0.0147893f $X=50.145
+ $Y=3.86 $X2=0 $Y2=0
cc_7230 N_A_9463_613#_c_12570_n N_A_9513_918#_c_15285_n 0.00239279f $X=50.145
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7231 N_A_9463_613#_c_12571_n N_A_9513_918#_c_15285_n 0.00761509f $X=49.485
+ $Y=3.86 $X2=25.99 $Y2=3.23
cc_7232 N_A_9463_613#_c_12596_n N_A_9513_918#_c_15286_n 6.95815e-19 $X=50.31
+ $Y=3.78 $X2=0 $Y2=0
cc_7233 VGND N_A_119_47#_M1084_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7234 VGND N_A_119_47#_M1300_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7235 VGND N_A_119_47#_c_14057_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7236 N_VGND_c_12870_n N_A_119_47#_c_14057_n 0.0188215f $X=1.065 $Y=0 $X2=0
+ $Y2=0
cc_7237 N_VGND_M1219_d N_A_119_47#_c_14060_n 0.00501873f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_7238 N_VGND_c_12693_n N_A_119_47#_c_14060_n 0.0199861f $X=1.2 $Y=0.38 $X2=0
+ $Y2=0
cc_7239 N_VGND_c_12695_n N_A_119_47#_c_14060_n 0.0020257f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_7240 VGND N_A_119_47#_c_14060_n 0.00880092f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7241 N_VGND_c_12870_n N_A_119_47#_c_14060_n 0.0020257f $X=1.065 $Y=0 $X2=0
+ $Y2=0
cc_7242 N_VGND_c_12695_n N_A_119_47#_c_14068_n 0.0188215f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_7243 VGND N_A_119_47#_c_14068_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7244 N_VGND_M1317_d N_A_119_47#_c_14050_n 0.00692362f $X=1.955 $Y=0.235 $X2=0
+ $Y2=0
cc_7245 N_VGND_c_12695_n N_A_119_47#_c_14050_n 0.0020257f $X=2.005 $Y=0 $X2=0
+ $Y2=0
cc_7246 N_VGND_c_12697_n N_A_119_47#_c_14050_n 0.0190091f $X=2.09 $Y=0.38 $X2=0
+ $Y2=0
cc_7247 N_VGND_c_12787_n N_A_119_47#_c_14050_n 0.00262594f $X=4.96 $Y=0 $X2=0
+ $Y2=0
cc_7248 VGND N_A_119_47#_c_14050_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7249 N_VGND_c_12697_n N_A_119_47#_c_14051_n 0.00959666f $X=2.09 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7250 N_VGND_c_12787_n N_A_119_47#_c_14052_n 0.0422314f $X=4.96 $Y=0 $X2=0
+ $Y2=0
cc_7251 VGND N_A_119_47#_c_14052_n 0.0222193f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7252 N_VGND_c_12697_n N_A_119_47#_c_14053_n 0.0147456f $X=2.09 $Y=0.38 $X2=0
+ $Y2=0
cc_7253 N_VGND_c_12787_n N_A_119_47#_c_14053_n 0.0192461f $X=4.96 $Y=0 $X2=0
+ $Y2=0
cc_7254 VGND N_A_119_47#_c_14053_n 0.0103774f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7255 N_VGND_c_12699_n N_A_119_47#_c_14054_n 0.00694621f $X=5.165 $Y=0.445
+ $X2=25.99 $Y2=4.8
cc_7256 N_VGND_c_12787_n N_A_119_47#_c_14054_n 0.0589406f $X=4.96 $Y=0 $X2=25.99
+ $Y2=4.8
cc_7257 VGND N_A_119_47#_c_14054_n 0.030408f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7258 N_VGND_c_12699_n N_A_119_47#_c_14055_n 0.00696245f $X=5.165 $Y=0.445
+ $X2=25.99 $Y2=4.93
cc_7259 N_VGND_c_12787_n N_A_119_47#_c_14090_n 0.0113631f $X=4.96 $Y=0 $X2=0
+ $Y2=0
cc_7260 VGND N_A_119_47#_c_14090_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7261 VGND N_A_119_911#_M1085_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7262 VGND N_A_119_911#_M1235_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7263 N_VGND_M1090_d N_A_119_911#_c_14140_n 0.00501873f $X=1.015 $Y=4.555
+ $X2=0 $Y2=0
cc_7264 N_VGND_c_12694_n N_A_119_911#_c_14140_n 0.0199861f $X=1.2 $Y=5.06 $X2=0
+ $Y2=0
cc_7265 N_VGND_c_12696_n N_A_119_911#_c_14140_n 0.0020257f $X=2.005 $Y=5.44
+ $X2=0 $Y2=0
cc_7266 VGND N_A_119_911#_c_14140_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7267 N_VGND_c_12871_n N_A_119_911#_c_14140_n 0.0020257f $X=1.065 $Y=5.44
+ $X2=0 $Y2=0
cc_7268 N_VGND_M1240_d N_A_119_911#_c_14132_n 0.00692362f $X=1.955 $Y=4.555
+ $X2=0 $Y2=0
cc_7269 N_VGND_c_12696_n N_A_119_911#_c_14132_n 0.0020257f $X=2.005 $Y=5.44
+ $X2=0 $Y2=0
cc_7270 N_VGND_c_12698_n N_A_119_911#_c_14132_n 0.0190091f $X=2.09 $Y=5.06 $X2=0
+ $Y2=0
cc_7271 N_VGND_c_12789_n N_A_119_911#_c_14132_n 0.00262594f $X=4.96 $Y=5.44
+ $X2=0 $Y2=0
cc_7272 VGND N_A_119_911#_c_14132_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7273 N_VGND_c_12698_n N_A_119_911#_c_14133_n 0.00959666f $X=2.09 $Y=5.06
+ $X2=0 $Y2=0
cc_7274 N_VGND_c_12789_n N_A_119_911#_c_14134_n 0.0422314f $X=4.96 $Y=5.44 $X2=0
+ $Y2=0
cc_7275 VGND N_A_119_911#_c_14134_n 0.0222193f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7276 N_VGND_c_12698_n N_A_119_911#_c_14135_n 0.0147456f $X=2.09 $Y=5.06 $X2=0
+ $Y2=0
cc_7277 N_VGND_c_12789_n N_A_119_911#_c_14135_n 0.0192461f $X=4.96 $Y=5.44 $X2=0
+ $Y2=0
cc_7278 VGND N_A_119_911#_c_14135_n 0.0103774f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7279 N_VGND_c_12700_n N_A_119_911#_c_14136_n 0.00694621f $X=5.165 $Y=4.995
+ $X2=25.99 $Y2=0.64
cc_7280 N_VGND_c_12789_n N_A_119_911#_c_14136_n 0.0589406f $X=4.96 $Y=5.44
+ $X2=25.99 $Y2=0.64
cc_7281 VGND N_A_119_911#_c_14136_n 0.030408f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=0.64
cc_7282 N_VGND_c_12700_n N_A_119_911#_c_14137_n 0.00696245f $X=5.165 $Y=4.995
+ $X2=25.99 $Y2=4.8
cc_7283 VGND N_A_119_911#_c_14138_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7284 N_VGND_c_12871_n N_A_119_911#_c_14138_n 0.0188215f $X=1.065 $Y=5.44
+ $X2=0 $Y2=0
cc_7285 N_VGND_c_12696_n N_A_119_911#_c_14139_n 0.0188215f $X=2.005 $Y=5.44
+ $X2=0 $Y2=0
cc_7286 VGND N_A_119_911#_c_14139_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7287 N_VGND_c_12789_n N_A_119_911#_c_14169_n 0.0113631f $X=4.96 $Y=5.44 $X2=0
+ $Y2=0
cc_7288 VGND N_A_119_911#_c_14169_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7289 VGND N_A_1693_66#_M1049_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7290 VGND N_A_1693_66#_M1167_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7291 N_VGND_c_12705_n N_A_1693_66#_c_14211_n 0.00696245f $X=7.715 $Y=0.445
+ $X2=0 $Y2=0
cc_7292 N_VGND_c_12803_n N_A_1693_66#_c_14212_n 0.0422314f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_7293 VGND N_A_1693_66#_c_14212_n 0.0219908f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7294 N_VGND_c_12705_n N_A_1693_66#_c_14213_n 0.00694621f $X=7.715 $Y=0.445
+ $X2=0 $Y2=0
cc_7295 N_VGND_c_12803_n N_A_1693_66#_c_14213_n 0.0167092f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_7296 VGND N_A_1693_66#_c_14213_n 0.00841721f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7297 N_VGND_c_12707_n N_A_1693_66#_c_14214_n 0.0147456f $X=10.79 $Y=0.38
+ $X2=0 $Y2=0
cc_7298 N_VGND_c_12803_n N_A_1693_66#_c_14214_n 0.0614775f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_7299 VGND N_A_1693_66#_c_14214_n 0.0325967f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7300 N_VGND_c_12707_n N_A_1693_66#_c_14215_n 0.00959666f $X=10.79 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7301 N_VGND_M1049_d N_A_1693_66#_c_14216_n 0.00692362f $X=10.665 $Y=0.235
+ $X2=0 $Y2=0
cc_7302 N_VGND_c_12707_n N_A_1693_66#_c_14216_n 0.0190091f $X=10.79 $Y=0.38
+ $X2=0 $Y2=0
cc_7303 N_VGND_c_12803_n N_A_1693_66#_c_14216_n 0.00262594f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_7304 VGND N_A_1693_66#_c_14216_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7305 N_VGND_c_12872_n N_A_1693_66#_c_14216_n 0.0020257f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_7306 VGND N_A_1693_66#_c_14236_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7307 N_VGND_c_12872_n N_A_1693_66#_c_14236_n 0.0188215f $X=11.545 $Y=0 $X2=0
+ $Y2=0
cc_7308 N_VGND_M1098_d N_A_1693_66#_c_14218_n 0.00501873f $X=11.495 $Y=0.235
+ $X2=25.99 $Y2=4.8
cc_7309 N_VGND_c_12709_n N_A_1693_66#_c_14218_n 0.0199861f $X=11.68 $Y=0.38
+ $X2=25.99 $Y2=4.8
cc_7310 VGND N_A_1693_66#_c_14218_n 0.00880092f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7311 N_VGND_c_12872_n N_A_1693_66#_c_14218_n 0.0020257f $X=11.545 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7312 N_VGND_c_12874_n N_A_1693_66#_c_14218_n 0.0020257f $X=12.485 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7313 VGND N_A_1693_66#_c_14245_n 0.0121968f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.93
cc_7314 N_VGND_c_12874_n N_A_1693_66#_c_14245_n 0.0188215f $X=12.485 $Y=0
+ $X2=25.99 $Y2=4.93
cc_7315 N_VGND_c_12803_n N_A_1693_66#_c_14230_n 0.0113631f $X=10.625 $Y=0 $X2=0
+ $Y2=0
cc_7316 VGND N_A_1693_66#_c_14230_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7317 VGND N_A_1693_918#_M1019_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7318 VGND N_A_1693_918#_M1178_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7319 N_VGND_c_12706_n N_A_1693_918#_c_14295_n 0.00696245f $X=7.715 $Y=4.995
+ $X2=0 $Y2=0
cc_7320 N_VGND_c_12805_n N_A_1693_918#_c_14296_n 0.0422314f $X=10.625 $Y=5.44
+ $X2=0 $Y2=0
cc_7321 VGND N_A_1693_918#_c_14296_n 0.0219908f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7322 N_VGND_c_12706_n N_A_1693_918#_c_14297_n 0.00694621f $X=7.715 $Y=4.995
+ $X2=0 $Y2=0
cc_7323 N_VGND_c_12805_n N_A_1693_918#_c_14297_n 0.0167092f $X=10.625 $Y=5.44
+ $X2=0 $Y2=0
cc_7324 VGND N_A_1693_918#_c_14297_n 0.00841721f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7325 N_VGND_c_12708_n N_A_1693_918#_c_14298_n 0.0147456f $X=10.79 $Y=5.06
+ $X2=0 $Y2=0
cc_7326 N_VGND_c_12805_n N_A_1693_918#_c_14298_n 0.0614775f $X=10.625 $Y=5.44
+ $X2=0 $Y2=0
cc_7327 VGND N_A_1693_918#_c_14298_n 0.0325967f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7328 N_VGND_c_12708_n N_A_1693_918#_c_14299_n 0.00959666f $X=10.79 $Y=5.06
+ $X2=25.99 $Y2=0.51
cc_7329 N_VGND_M1019_d N_A_1693_918#_c_14300_n 0.00692362f $X=10.665 $Y=4.555
+ $X2=0 $Y2=0
cc_7330 N_VGND_c_12708_n N_A_1693_918#_c_14300_n 0.0190091f $X=10.79 $Y=5.06
+ $X2=0 $Y2=0
cc_7331 N_VGND_c_12805_n N_A_1693_918#_c_14300_n 0.00262594f $X=10.625 $Y=5.44
+ $X2=0 $Y2=0
cc_7332 VGND N_A_1693_918#_c_14300_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7333 N_VGND_c_12873_n N_A_1693_918#_c_14300_n 0.0020257f $X=11.545 $Y=5.44
+ $X2=0 $Y2=0
cc_7334 N_VGND_M1111_d N_A_1693_918#_c_14320_n 0.00501873f $X=11.495 $Y=4.555
+ $X2=0 $Y2=0
cc_7335 N_VGND_c_12710_n N_A_1693_918#_c_14320_n 0.0199861f $X=11.68 $Y=5.06
+ $X2=0 $Y2=0
cc_7336 VGND N_A_1693_918#_c_14320_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7337 N_VGND_c_12873_n N_A_1693_918#_c_14320_n 0.0020257f $X=11.545 $Y=5.44
+ $X2=0 $Y2=0
cc_7338 N_VGND_c_12875_n N_A_1693_918#_c_14320_n 0.0020257f $X=12.485 $Y=5.44
+ $X2=0 $Y2=0
cc_7339 N_VGND_c_12805_n N_A_1693_918#_c_14314_n 0.0113631f $X=10.625 $Y=5.44
+ $X2=0 $Y2=0
cc_7340 VGND N_A_1693_918#_c_14314_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7341 VGND N_A_1693_918#_c_14302_n 0.0121968f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=4.93
cc_7342 N_VGND_c_12873_n N_A_1693_918#_c_14302_n 0.0188215f $X=11.545 $Y=5.44
+ $X2=25.99 $Y2=4.93
cc_7343 VGND N_A_1693_918#_c_14303_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7344 N_VGND_c_12875_n N_A_1693_918#_c_14303_n 0.0188215f $X=12.485 $Y=5.44
+ $X2=0 $Y2=0
cc_7345 VGND N_A_2695_47#_M1001_d 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7346 VGND N_A_2695_47#_M1110_d 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7347 VGND N_A_2695_47#_c_14385_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7348 N_VGND_c_12876_n N_A_2695_47#_c_14385_n 0.0188215f $X=13.945 $Y=0 $X2=0
+ $Y2=0
cc_7349 N_VGND_M1062_s N_A_2695_47#_c_14388_n 0.00501873f $X=13.895 $Y=0.235
+ $X2=0 $Y2=0
cc_7350 N_VGND_c_12717_n N_A_2695_47#_c_14388_n 0.0199861f $X=14.08 $Y=0.38
+ $X2=0 $Y2=0
cc_7351 N_VGND_c_12719_n N_A_2695_47#_c_14388_n 0.0020257f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_7352 VGND N_A_2695_47#_c_14388_n 0.00880092f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7353 N_VGND_c_12876_n N_A_2695_47#_c_14388_n 0.0020257f $X=13.945 $Y=0 $X2=0
+ $Y2=0
cc_7354 N_VGND_c_12719_n N_A_2695_47#_c_14396_n 0.0188215f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_7355 VGND N_A_2695_47#_c_14396_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7356 N_VGND_M1182_s N_A_2695_47#_c_14378_n 0.00692362f $X=14.835 $Y=0.235
+ $X2=0 $Y2=0
cc_7357 N_VGND_c_12719_n N_A_2695_47#_c_14378_n 0.0020257f $X=14.885 $Y=0 $X2=0
+ $Y2=0
cc_7358 N_VGND_c_12721_n N_A_2695_47#_c_14378_n 0.0190091f $X=14.97 $Y=0.38
+ $X2=0 $Y2=0
cc_7359 N_VGND_c_12807_n N_A_2695_47#_c_14378_n 0.00262594f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_7360 VGND N_A_2695_47#_c_14378_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7361 N_VGND_c_12721_n N_A_2695_47#_c_14379_n 0.00959666f $X=14.97 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7362 N_VGND_c_12807_n N_A_2695_47#_c_14380_n 0.0422314f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_7363 VGND N_A_2695_47#_c_14380_n 0.0222193f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7364 N_VGND_c_12721_n N_A_2695_47#_c_14381_n 0.0147456f $X=14.97 $Y=0.38
+ $X2=0 $Y2=0
cc_7365 N_VGND_c_12807_n N_A_2695_47#_c_14381_n 0.0192461f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_7366 VGND N_A_2695_47#_c_14381_n 0.0103774f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7367 N_VGND_c_12723_n N_A_2695_47#_c_14382_n 0.00694621f $X=18.045 $Y=0.445
+ $X2=25.99 $Y2=4.8
cc_7368 N_VGND_c_12807_n N_A_2695_47#_c_14382_n 0.0589406f $X=17.84 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7369 VGND N_A_2695_47#_c_14382_n 0.030408f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7370 N_VGND_c_12723_n N_A_2695_47#_c_14383_n 0.00696245f $X=18.045 $Y=0.445
+ $X2=25.99 $Y2=4.93
cc_7371 N_VGND_c_12807_n N_A_2695_47#_c_14418_n 0.0113631f $X=17.84 $Y=0 $X2=0
+ $Y2=0
cc_7372 VGND N_A_2695_47#_c_14418_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7373 VGND N_A_2695_911#_M1033_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7374 VGND N_A_2695_911#_M1195_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7375 N_VGND_M1143_d N_A_2695_911#_c_14468_n 0.00501873f $X=13.895 $Y=4.555
+ $X2=0 $Y2=0
cc_7376 N_VGND_c_12718_n N_A_2695_911#_c_14468_n 0.0199861f $X=14.08 $Y=5.06
+ $X2=0 $Y2=0
cc_7377 N_VGND_c_12720_n N_A_2695_911#_c_14468_n 0.0020257f $X=14.885 $Y=5.44
+ $X2=0 $Y2=0
cc_7378 VGND N_A_2695_911#_c_14468_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7379 N_VGND_c_12877_n N_A_2695_911#_c_14468_n 0.0020257f $X=13.945 $Y=5.44
+ $X2=0 $Y2=0
cc_7380 N_VGND_M1307_d N_A_2695_911#_c_14460_n 0.00692362f $X=14.835 $Y=4.555
+ $X2=0 $Y2=0
cc_7381 N_VGND_c_12720_n N_A_2695_911#_c_14460_n 0.0020257f $X=14.885 $Y=5.44
+ $X2=0 $Y2=0
cc_7382 N_VGND_c_12722_n N_A_2695_911#_c_14460_n 0.0190091f $X=14.97 $Y=5.06
+ $X2=0 $Y2=0
cc_7383 N_VGND_c_12809_n N_A_2695_911#_c_14460_n 0.00262594f $X=17.84 $Y=5.44
+ $X2=0 $Y2=0
cc_7384 VGND N_A_2695_911#_c_14460_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7385 N_VGND_c_12722_n N_A_2695_911#_c_14461_n 0.00959666f $X=14.97 $Y=5.06
+ $X2=0 $Y2=0
cc_7386 N_VGND_c_12809_n N_A_2695_911#_c_14462_n 0.0422314f $X=17.84 $Y=5.44
+ $X2=0 $Y2=0
cc_7387 VGND N_A_2695_911#_c_14462_n 0.0222193f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7388 N_VGND_c_12722_n N_A_2695_911#_c_14463_n 0.0147456f $X=14.97 $Y=5.06
+ $X2=0 $Y2=0
cc_7389 N_VGND_c_12809_n N_A_2695_911#_c_14463_n 0.0192461f $X=17.84 $Y=5.44
+ $X2=0 $Y2=0
cc_7390 VGND N_A_2695_911#_c_14463_n 0.0103774f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7391 N_VGND_c_12724_n N_A_2695_911#_c_14464_n 0.00694621f $X=18.045 $Y=4.995
+ $X2=25.99 $Y2=0.64
cc_7392 N_VGND_c_12809_n N_A_2695_911#_c_14464_n 0.0589406f $X=17.84 $Y=5.44
+ $X2=25.99 $Y2=0.64
cc_7393 VGND N_A_2695_911#_c_14464_n 0.030408f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=0.64
cc_7394 N_VGND_c_12724_n N_A_2695_911#_c_14465_n 0.00696245f $X=18.045 $Y=4.995
+ $X2=25.99 $Y2=4.8
cc_7395 VGND N_A_2695_911#_c_14466_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7396 N_VGND_c_12877_n N_A_2695_911#_c_14466_n 0.0188215f $X=13.945 $Y=5.44
+ $X2=0 $Y2=0
cc_7397 N_VGND_c_12720_n N_A_2695_911#_c_14467_n 0.0188215f $X=14.885 $Y=5.44
+ $X2=0 $Y2=0
cc_7398 VGND N_A_2695_911#_c_14467_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7399 N_VGND_c_12809_n N_A_2695_911#_c_14497_n 0.0113631f $X=17.84 $Y=5.44
+ $X2=0 $Y2=0
cc_7400 VGND N_A_2695_911#_c_14497_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7401 VGND N_A_4269_66#_M1041_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7402 VGND N_A_4269_66#_M1135_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7403 N_VGND_c_12729_n N_A_4269_66#_c_14539_n 0.00696245f $X=20.595 $Y=0.445
+ $X2=0 $Y2=0
cc_7404 N_VGND_c_12823_n N_A_4269_66#_c_14540_n 0.0422314f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_7405 VGND N_A_4269_66#_c_14540_n 0.0219908f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7406 N_VGND_c_12729_n N_A_4269_66#_c_14541_n 0.00694621f $X=20.595 $Y=0.445
+ $X2=0 $Y2=0
cc_7407 N_VGND_c_12823_n N_A_4269_66#_c_14541_n 0.0167092f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_7408 VGND N_A_4269_66#_c_14541_n 0.00841721f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7409 N_VGND_c_12731_n N_A_4269_66#_c_14542_n 0.0147456f $X=23.67 $Y=0.38
+ $X2=0 $Y2=0
cc_7410 N_VGND_c_12823_n N_A_4269_66#_c_14542_n 0.0614775f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_7411 VGND N_A_4269_66#_c_14542_n 0.0325967f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7412 N_VGND_c_12731_n N_A_4269_66#_c_14543_n 0.00959666f $X=23.67 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7413 N_VGND_M1041_d N_A_4269_66#_c_14544_n 0.00692362f $X=23.545 $Y=0.235
+ $X2=0 $Y2=0
cc_7414 N_VGND_c_12731_n N_A_4269_66#_c_14544_n 0.0190091f $X=23.67 $Y=0.38
+ $X2=0 $Y2=0
cc_7415 N_VGND_c_12823_n N_A_4269_66#_c_14544_n 0.00262594f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_7416 VGND N_A_4269_66#_c_14544_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7417 N_VGND_c_12878_n N_A_4269_66#_c_14544_n 0.0020257f $X=24.425 $Y=0 $X2=0
+ $Y2=0
cc_7418 VGND N_A_4269_66#_c_14564_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7419 N_VGND_c_12878_n N_A_4269_66#_c_14564_n 0.0188215f $X=24.425 $Y=0 $X2=0
+ $Y2=0
cc_7420 N_VGND_M1100_d N_A_4269_66#_c_14546_n 0.00501873f $X=24.375 $Y=0.235
+ $X2=25.99 $Y2=4.8
cc_7421 N_VGND_c_12733_n N_A_4269_66#_c_14546_n 0.0199861f $X=24.56 $Y=0.38
+ $X2=25.99 $Y2=4.8
cc_7422 VGND N_A_4269_66#_c_14546_n 0.00880092f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7423 N_VGND_c_12878_n N_A_4269_66#_c_14546_n 0.0020257f $X=24.425 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7424 N_VGND_c_12880_n N_A_4269_66#_c_14546_n 0.0020257f $X=25.365 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7425 VGND N_A_4269_66#_c_14573_n 0.0121968f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.93
cc_7426 N_VGND_c_12880_n N_A_4269_66#_c_14573_n 0.0188215f $X=25.365 $Y=0
+ $X2=25.99 $Y2=4.93
cc_7427 N_VGND_c_12823_n N_A_4269_66#_c_14558_n 0.0113631f $X=23.505 $Y=0 $X2=0
+ $Y2=0
cc_7428 VGND N_A_4269_66#_c_14558_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7429 VGND N_A_4269_918#_M1245_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7430 VGND N_A_4269_918#_M1310_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7431 N_VGND_c_12730_n N_A_4269_918#_c_14623_n 0.00696245f $X=20.595 $Y=4.995
+ $X2=0 $Y2=0
cc_7432 N_VGND_c_12825_n N_A_4269_918#_c_14624_n 0.0422314f $X=23.505 $Y=5.44
+ $X2=0 $Y2=0
cc_7433 VGND N_A_4269_918#_c_14624_n 0.0219908f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7434 N_VGND_c_12730_n N_A_4269_918#_c_14625_n 0.00694621f $X=20.595 $Y=4.995
+ $X2=0 $Y2=0
cc_7435 N_VGND_c_12825_n N_A_4269_918#_c_14625_n 0.0167092f $X=23.505 $Y=5.44
+ $X2=0 $Y2=0
cc_7436 VGND N_A_4269_918#_c_14625_n 0.00841721f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7437 N_VGND_c_12732_n N_A_4269_918#_c_14626_n 0.0147456f $X=23.67 $Y=5.06
+ $X2=0 $Y2=0
cc_7438 N_VGND_c_12825_n N_A_4269_918#_c_14626_n 0.0614775f $X=23.505 $Y=5.44
+ $X2=0 $Y2=0
cc_7439 VGND N_A_4269_918#_c_14626_n 0.0325967f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7440 N_VGND_c_12732_n N_A_4269_918#_c_14627_n 0.00959666f $X=23.67 $Y=5.06
+ $X2=25.99 $Y2=0.51
cc_7441 N_VGND_M1245_s N_A_4269_918#_c_14628_n 0.00692362f $X=23.545 $Y=4.555
+ $X2=0 $Y2=0
cc_7442 N_VGND_c_12732_n N_A_4269_918#_c_14628_n 0.0190091f $X=23.67 $Y=5.06
+ $X2=0 $Y2=0
cc_7443 N_VGND_c_12825_n N_A_4269_918#_c_14628_n 0.00262594f $X=23.505 $Y=5.44
+ $X2=0 $Y2=0
cc_7444 VGND N_A_4269_918#_c_14628_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7445 N_VGND_c_12879_n N_A_4269_918#_c_14628_n 0.0020257f $X=24.425 $Y=5.44
+ $X2=0 $Y2=0
cc_7446 N_VGND_M1296_s N_A_4269_918#_c_14648_n 0.00501873f $X=24.375 $Y=4.555
+ $X2=0 $Y2=0
cc_7447 N_VGND_c_12734_n N_A_4269_918#_c_14648_n 0.0199861f $X=24.56 $Y=5.06
+ $X2=0 $Y2=0
cc_7448 VGND N_A_4269_918#_c_14648_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7449 N_VGND_c_12879_n N_A_4269_918#_c_14648_n 0.0020257f $X=24.425 $Y=5.44
+ $X2=0 $Y2=0
cc_7450 N_VGND_c_12881_n N_A_4269_918#_c_14648_n 0.0020257f $X=25.365 $Y=5.44
+ $X2=0 $Y2=0
cc_7451 N_VGND_c_12825_n N_A_4269_918#_c_14642_n 0.0113631f $X=23.505 $Y=5.44
+ $X2=0 $Y2=0
cc_7452 VGND N_A_4269_918#_c_14642_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7453 VGND N_A_4269_918#_c_14630_n 0.0121968f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=4.93
cc_7454 N_VGND_c_12879_n N_A_4269_918#_c_14630_n 0.0188215f $X=24.425 $Y=5.44
+ $X2=25.99 $Y2=4.93
cc_7455 VGND N_A_4269_918#_c_14631_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7456 N_VGND_c_12881_n N_A_4269_918#_c_14631_n 0.0188215f $X=25.365 $Y=5.44
+ $X2=0 $Y2=0
cc_7457 VGND N_A_5363_47#_M1021_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7458 VGND N_A_5363_47#_M1232_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7459 VGND N_A_5363_47#_c_14713_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7460 N_VGND_c_12885_n N_A_5363_47#_c_14713_n 0.0188215f $X=27.285 $Y=0 $X2=0
+ $Y2=0
cc_7461 N_VGND_M1177_d N_A_5363_47#_c_14716_n 0.00501873f $X=27.235 $Y=0.235
+ $X2=0 $Y2=0
cc_7462 N_VGND_c_12741_n N_A_5363_47#_c_14716_n 0.0199861f $X=27.42 $Y=0.38
+ $X2=0 $Y2=0
cc_7463 N_VGND_c_12743_n N_A_5363_47#_c_14716_n 0.0020257f $X=28.225 $Y=0 $X2=0
+ $Y2=0
cc_7464 VGND N_A_5363_47#_c_14716_n 0.00880092f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7465 N_VGND_c_12885_n N_A_5363_47#_c_14716_n 0.0020257f $X=27.285 $Y=0 $X2=0
+ $Y2=0
cc_7466 N_VGND_c_12743_n N_A_5363_47#_c_14724_n 0.0188215f $X=28.225 $Y=0 $X2=0
+ $Y2=0
cc_7467 VGND N_A_5363_47#_c_14724_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7468 N_VGND_M1275_d N_A_5363_47#_c_14706_n 0.00692362f $X=28.175 $Y=0.235
+ $X2=0 $Y2=0
cc_7469 N_VGND_c_12743_n N_A_5363_47#_c_14706_n 0.0020257f $X=28.225 $Y=0 $X2=0
+ $Y2=0
cc_7470 N_VGND_c_12745_n N_A_5363_47#_c_14706_n 0.0190091f $X=28.31 $Y=0.38
+ $X2=0 $Y2=0
cc_7471 N_VGND_c_12827_n N_A_5363_47#_c_14706_n 0.00262594f $X=31.18 $Y=0 $X2=0
+ $Y2=0
cc_7472 VGND N_A_5363_47#_c_14706_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7473 N_VGND_c_12745_n N_A_5363_47#_c_14707_n 0.00959666f $X=28.31 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7474 N_VGND_c_12827_n N_A_5363_47#_c_14708_n 0.0422314f $X=31.18 $Y=0 $X2=0
+ $Y2=0
cc_7475 VGND N_A_5363_47#_c_14708_n 0.0222193f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7476 N_VGND_c_12745_n N_A_5363_47#_c_14709_n 0.0147456f $X=28.31 $Y=0.38
+ $X2=0 $Y2=0
cc_7477 N_VGND_c_12827_n N_A_5363_47#_c_14709_n 0.0192461f $X=31.18 $Y=0 $X2=0
+ $Y2=0
cc_7478 VGND N_A_5363_47#_c_14709_n 0.0103774f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7479 N_VGND_c_12747_n N_A_5363_47#_c_14710_n 0.00694621f $X=31.385 $Y=0.445
+ $X2=25.99 $Y2=4.8
cc_7480 N_VGND_c_12827_n N_A_5363_47#_c_14710_n 0.0589406f $X=31.18 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7481 VGND N_A_5363_47#_c_14710_n 0.030408f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7482 N_VGND_c_12747_n N_A_5363_47#_c_14711_n 0.00696245f $X=31.385 $Y=0.445
+ $X2=25.99 $Y2=4.93
cc_7483 N_VGND_c_12827_n N_A_5363_47#_c_14746_n 0.0113631f $X=31.18 $Y=0 $X2=0
+ $Y2=0
cc_7484 VGND N_A_5363_47#_c_14746_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7485 VGND N_A_5363_911#_M1012_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7486 VGND N_A_5363_911#_M1187_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7487 N_VGND_M1128_d N_A_5363_911#_c_14796_n 0.00501873f $X=27.235 $Y=4.555
+ $X2=0 $Y2=0
cc_7488 N_VGND_c_12742_n N_A_5363_911#_c_14796_n 0.0199861f $X=27.42 $Y=5.06
+ $X2=0 $Y2=0
cc_7489 N_VGND_c_12744_n N_A_5363_911#_c_14796_n 0.0020257f $X=28.225 $Y=5.44
+ $X2=0 $Y2=0
cc_7490 VGND N_A_5363_911#_c_14796_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7491 N_VGND_c_12886_n N_A_5363_911#_c_14796_n 0.0020257f $X=27.285 $Y=5.44
+ $X2=0 $Y2=0
cc_7492 N_VGND_M1267_d N_A_5363_911#_c_14788_n 0.00692362f $X=28.175 $Y=4.555
+ $X2=0 $Y2=0
cc_7493 N_VGND_c_12744_n N_A_5363_911#_c_14788_n 0.0020257f $X=28.225 $Y=5.44
+ $X2=0 $Y2=0
cc_7494 N_VGND_c_12746_n N_A_5363_911#_c_14788_n 0.0190091f $X=28.31 $Y=5.06
+ $X2=0 $Y2=0
cc_7495 N_VGND_c_12829_n N_A_5363_911#_c_14788_n 0.00262594f $X=31.18 $Y=5.44
+ $X2=0 $Y2=0
cc_7496 VGND N_A_5363_911#_c_14788_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7497 N_VGND_c_12746_n N_A_5363_911#_c_14789_n 0.00959666f $X=28.31 $Y=5.06
+ $X2=0 $Y2=0
cc_7498 N_VGND_c_12829_n N_A_5363_911#_c_14790_n 0.0422314f $X=31.18 $Y=5.44
+ $X2=0 $Y2=0
cc_7499 VGND N_A_5363_911#_c_14790_n 0.0222193f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7500 N_VGND_c_12746_n N_A_5363_911#_c_14791_n 0.0147456f $X=28.31 $Y=5.06
+ $X2=0 $Y2=0
cc_7501 N_VGND_c_12829_n N_A_5363_911#_c_14791_n 0.0192461f $X=31.18 $Y=5.44
+ $X2=0 $Y2=0
cc_7502 VGND N_A_5363_911#_c_14791_n 0.0103774f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7503 N_VGND_c_12748_n N_A_5363_911#_c_14792_n 0.00694621f $X=31.385 $Y=4.995
+ $X2=25.99 $Y2=0.64
cc_7504 N_VGND_c_12829_n N_A_5363_911#_c_14792_n 0.0589406f $X=31.18 $Y=5.44
+ $X2=25.99 $Y2=0.64
cc_7505 VGND N_A_5363_911#_c_14792_n 0.030408f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=0.64
cc_7506 N_VGND_c_12748_n N_A_5363_911#_c_14793_n 0.00696245f $X=31.385 $Y=4.995
+ $X2=25.99 $Y2=4.8
cc_7507 VGND N_A_5363_911#_c_14794_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7508 N_VGND_c_12886_n N_A_5363_911#_c_14794_n 0.0188215f $X=27.285 $Y=5.44
+ $X2=0 $Y2=0
cc_7509 N_VGND_c_12744_n N_A_5363_911#_c_14795_n 0.0188215f $X=28.225 $Y=5.44
+ $X2=0 $Y2=0
cc_7510 VGND N_A_5363_911#_c_14795_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7511 N_VGND_c_12829_n N_A_5363_911#_c_14825_n 0.0113631f $X=31.18 $Y=5.44
+ $X2=0 $Y2=0
cc_7512 VGND N_A_5363_911#_c_14825_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7513 VGND N_A_6937_66#_M1029_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7514 VGND N_A_6937_66#_M1247_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7515 N_VGND_c_12753_n N_A_6937_66#_c_14867_n 0.00696245f $X=33.935 $Y=0.445
+ $X2=0 $Y2=0
cc_7516 N_VGND_c_12843_n N_A_6937_66#_c_14868_n 0.0422314f $X=36.845 $Y=0 $X2=0
+ $Y2=0
cc_7517 VGND N_A_6937_66#_c_14868_n 0.0219908f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7518 N_VGND_c_12753_n N_A_6937_66#_c_14869_n 0.00694621f $X=33.935 $Y=0.445
+ $X2=0 $Y2=0
cc_7519 N_VGND_c_12843_n N_A_6937_66#_c_14869_n 0.0167092f $X=36.845 $Y=0 $X2=0
+ $Y2=0
cc_7520 VGND N_A_6937_66#_c_14869_n 0.00841721f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7521 N_VGND_c_12755_n N_A_6937_66#_c_14870_n 0.0147456f $X=37.01 $Y=0.38
+ $X2=0 $Y2=0
cc_7522 N_VGND_c_12843_n N_A_6937_66#_c_14870_n 0.0614775f $X=36.845 $Y=0 $X2=0
+ $Y2=0
cc_7523 VGND N_A_6937_66#_c_14870_n 0.0325967f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7524 N_VGND_c_12755_n N_A_6937_66#_c_14871_n 0.00959666f $X=37.01 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7525 N_VGND_M1029_d N_A_6937_66#_c_14872_n 0.00692362f $X=36.885 $Y=0.235
+ $X2=0 $Y2=0
cc_7526 N_VGND_c_12755_n N_A_6937_66#_c_14872_n 0.0190091f $X=37.01 $Y=0.38
+ $X2=0 $Y2=0
cc_7527 N_VGND_c_12843_n N_A_6937_66#_c_14872_n 0.00262594f $X=36.845 $Y=0 $X2=0
+ $Y2=0
cc_7528 VGND N_A_6937_66#_c_14872_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7529 N_VGND_c_12887_n N_A_6937_66#_c_14872_n 0.0020257f $X=37.765 $Y=0 $X2=0
+ $Y2=0
cc_7530 VGND N_A_6937_66#_c_14892_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7531 N_VGND_c_12887_n N_A_6937_66#_c_14892_n 0.0188215f $X=37.765 $Y=0 $X2=0
+ $Y2=0
cc_7532 N_VGND_M1057_d N_A_6937_66#_c_14874_n 0.00501873f $X=37.715 $Y=0.235
+ $X2=25.99 $Y2=4.8
cc_7533 N_VGND_c_12757_n N_A_6937_66#_c_14874_n 0.0199861f $X=37.9 $Y=0.38
+ $X2=25.99 $Y2=4.8
cc_7534 VGND N_A_6937_66#_c_14874_n 0.00880092f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7535 N_VGND_c_12887_n N_A_6937_66#_c_14874_n 0.0020257f $X=37.765 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7536 N_VGND_c_12889_n N_A_6937_66#_c_14874_n 0.0020257f $X=38.705 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7537 VGND N_A_6937_66#_c_14901_n 0.0121968f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.93
cc_7538 N_VGND_c_12889_n N_A_6937_66#_c_14901_n 0.0188215f $X=38.705 $Y=0
+ $X2=25.99 $Y2=4.93
cc_7539 N_VGND_c_12843_n N_A_6937_66#_c_14886_n 0.0113631f $X=36.845 $Y=0 $X2=0
+ $Y2=0
cc_7540 VGND N_A_6937_66#_c_14886_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7541 VGND N_A_6937_918#_M1132_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7542 VGND N_A_6937_918#_M1274_s 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7543 N_VGND_c_12754_n N_A_6937_918#_c_14951_n 0.00696245f $X=33.935 $Y=4.995
+ $X2=0 $Y2=0
cc_7544 N_VGND_c_12845_n N_A_6937_918#_c_14952_n 0.0422314f $X=36.845 $Y=5.44
+ $X2=0 $Y2=0
cc_7545 VGND N_A_6937_918#_c_14952_n 0.0219908f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7546 N_VGND_c_12754_n N_A_6937_918#_c_14953_n 0.00694621f $X=33.935 $Y=4.995
+ $X2=0 $Y2=0
cc_7547 N_VGND_c_12845_n N_A_6937_918#_c_14953_n 0.0167092f $X=36.845 $Y=5.44
+ $X2=0 $Y2=0
cc_7548 VGND N_A_6937_918#_c_14953_n 0.00841721f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7549 N_VGND_c_12756_n N_A_6937_918#_c_14954_n 0.0147456f $X=37.01 $Y=5.06
+ $X2=0 $Y2=0
cc_7550 N_VGND_c_12845_n N_A_6937_918#_c_14954_n 0.0614775f $X=36.845 $Y=5.44
+ $X2=0 $Y2=0
cc_7551 VGND N_A_6937_918#_c_14954_n 0.0325967f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7552 N_VGND_c_12756_n N_A_6937_918#_c_14955_n 0.00959666f $X=37.01 $Y=5.06
+ $X2=25.99 $Y2=0.51
cc_7553 N_VGND_M1132_d N_A_6937_918#_c_14956_n 0.00692362f $X=36.885 $Y=4.555
+ $X2=0 $Y2=0
cc_7554 N_VGND_c_12756_n N_A_6937_918#_c_14956_n 0.0190091f $X=37.01 $Y=5.06
+ $X2=0 $Y2=0
cc_7555 N_VGND_c_12845_n N_A_6937_918#_c_14956_n 0.00262594f $X=36.845 $Y=5.44
+ $X2=0 $Y2=0
cc_7556 VGND N_A_6937_918#_c_14956_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7557 N_VGND_c_12888_n N_A_6937_918#_c_14956_n 0.0020257f $X=37.765 $Y=5.44
+ $X2=0 $Y2=0
cc_7558 N_VGND_M1136_d N_A_6937_918#_c_14976_n 0.00501873f $X=37.715 $Y=4.555
+ $X2=0 $Y2=0
cc_7559 N_VGND_c_12758_n N_A_6937_918#_c_14976_n 0.0199861f $X=37.9 $Y=5.06
+ $X2=0 $Y2=0
cc_7560 VGND N_A_6937_918#_c_14976_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7561 N_VGND_c_12888_n N_A_6937_918#_c_14976_n 0.0020257f $X=37.765 $Y=5.44
+ $X2=0 $Y2=0
cc_7562 N_VGND_c_12890_n N_A_6937_918#_c_14976_n 0.0020257f $X=38.705 $Y=5.44
+ $X2=0 $Y2=0
cc_7563 N_VGND_c_12845_n N_A_6937_918#_c_14970_n 0.0113631f $X=36.845 $Y=5.44
+ $X2=0 $Y2=0
cc_7564 VGND N_A_6937_918#_c_14970_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7565 VGND N_A_6937_918#_c_14958_n 0.0121968f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=4.93
cc_7566 N_VGND_c_12888_n N_A_6937_918#_c_14958_n 0.0188215f $X=37.765 $Y=5.44
+ $X2=25.99 $Y2=4.93
cc_7567 VGND N_A_6937_918#_c_14959_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7568 N_VGND_c_12890_n N_A_6937_918#_c_14959_n 0.0188215f $X=38.705 $Y=5.44
+ $X2=0 $Y2=0
cc_7569 VGND N_A_7939_47#_M1069_d 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7570 VGND N_A_7939_47#_M1147_d 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7571 VGND N_A_7939_47#_c_15041_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7572 N_VGND_c_12891_n N_A_7939_47#_c_15041_n 0.0188215f $X=40.165 $Y=0 $X2=0
+ $Y2=0
cc_7573 N_VGND_M1122_s N_A_7939_47#_c_15044_n 0.00501873f $X=40.115 $Y=0.235
+ $X2=0 $Y2=0
cc_7574 N_VGND_c_12765_n N_A_7939_47#_c_15044_n 0.0199861f $X=40.3 $Y=0.38 $X2=0
+ $Y2=0
cc_7575 N_VGND_c_12767_n N_A_7939_47#_c_15044_n 0.0020257f $X=41.105 $Y=0 $X2=0
+ $Y2=0
cc_7576 VGND N_A_7939_47#_c_15044_n 0.00880092f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7577 N_VGND_c_12891_n N_A_7939_47#_c_15044_n 0.0020257f $X=40.165 $Y=0 $X2=0
+ $Y2=0
cc_7578 N_VGND_c_12767_n N_A_7939_47#_c_15052_n 0.0188215f $X=41.105 $Y=0 $X2=0
+ $Y2=0
cc_7579 VGND N_A_7939_47#_c_15052_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7580 N_VGND_M1258_s N_A_7939_47#_c_15034_n 0.00692362f $X=41.055 $Y=0.235
+ $X2=0 $Y2=0
cc_7581 N_VGND_c_12767_n N_A_7939_47#_c_15034_n 0.0020257f $X=41.105 $Y=0 $X2=0
+ $Y2=0
cc_7582 N_VGND_c_12769_n N_A_7939_47#_c_15034_n 0.0190091f $X=41.19 $Y=0.38
+ $X2=0 $Y2=0
cc_7583 N_VGND_c_12847_n N_A_7939_47#_c_15034_n 0.00262594f $X=44.06 $Y=0 $X2=0
+ $Y2=0
cc_7584 VGND N_A_7939_47#_c_15034_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7585 N_VGND_c_12769_n N_A_7939_47#_c_15035_n 0.00959666f $X=41.19 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7586 N_VGND_c_12847_n N_A_7939_47#_c_15036_n 0.0422314f $X=44.06 $Y=0 $X2=0
+ $Y2=0
cc_7587 VGND N_A_7939_47#_c_15036_n 0.0222193f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7588 N_VGND_c_12769_n N_A_7939_47#_c_15037_n 0.0147456f $X=41.19 $Y=0.38
+ $X2=0 $Y2=0
cc_7589 N_VGND_c_12847_n N_A_7939_47#_c_15037_n 0.0192461f $X=44.06 $Y=0 $X2=0
+ $Y2=0
cc_7590 VGND N_A_7939_47#_c_15037_n 0.0103774f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7591 N_VGND_c_12771_n N_A_7939_47#_c_15038_n 0.00694621f $X=44.265 $Y=0.445
+ $X2=25.99 $Y2=4.8
cc_7592 N_VGND_c_12847_n N_A_7939_47#_c_15038_n 0.0589406f $X=44.06 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7593 VGND N_A_7939_47#_c_15038_n 0.030408f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7594 N_VGND_c_12771_n N_A_7939_47#_c_15039_n 0.00696245f $X=44.265 $Y=0.445
+ $X2=25.99 $Y2=4.93
cc_7595 N_VGND_c_12847_n N_A_7939_47#_c_15074_n 0.0113631f $X=44.06 $Y=0 $X2=0
+ $Y2=0
cc_7596 VGND N_A_7939_47#_c_15074_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7597 VGND N_A_7939_911#_M1004_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7598 VGND N_A_7939_911#_M1189_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7599 N_VGND_M1179_s N_A_7939_911#_c_15124_n 0.00501873f $X=40.115 $Y=4.555
+ $X2=0 $Y2=0
cc_7600 N_VGND_c_12766_n N_A_7939_911#_c_15124_n 0.0199861f $X=40.3 $Y=5.06
+ $X2=0 $Y2=0
cc_7601 N_VGND_c_12768_n N_A_7939_911#_c_15124_n 0.0020257f $X=41.105 $Y=5.44
+ $X2=0 $Y2=0
cc_7602 VGND N_A_7939_911#_c_15124_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7603 N_VGND_c_12892_n N_A_7939_911#_c_15124_n 0.0020257f $X=40.165 $Y=5.44
+ $X2=0 $Y2=0
cc_7604 N_VGND_M1305_s N_A_7939_911#_c_15116_n 0.00692362f $X=41.055 $Y=4.555
+ $X2=0 $Y2=0
cc_7605 N_VGND_c_12768_n N_A_7939_911#_c_15116_n 0.0020257f $X=41.105 $Y=5.44
+ $X2=0 $Y2=0
cc_7606 N_VGND_c_12770_n N_A_7939_911#_c_15116_n 0.0190091f $X=41.19 $Y=5.06
+ $X2=0 $Y2=0
cc_7607 N_VGND_c_12849_n N_A_7939_911#_c_15116_n 0.00262594f $X=44.06 $Y=5.44
+ $X2=0 $Y2=0
cc_7608 VGND N_A_7939_911#_c_15116_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7609 N_VGND_c_12770_n N_A_7939_911#_c_15117_n 0.00959666f $X=41.19 $Y=5.06
+ $X2=0 $Y2=0
cc_7610 N_VGND_c_12849_n N_A_7939_911#_c_15118_n 0.0422314f $X=44.06 $Y=5.44
+ $X2=0 $Y2=0
cc_7611 VGND N_A_7939_911#_c_15118_n 0.0222193f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7612 N_VGND_c_12770_n N_A_7939_911#_c_15119_n 0.0147456f $X=41.19 $Y=5.06
+ $X2=0 $Y2=0
cc_7613 N_VGND_c_12849_n N_A_7939_911#_c_15119_n 0.0192461f $X=44.06 $Y=5.44
+ $X2=0 $Y2=0
cc_7614 VGND N_A_7939_911#_c_15119_n 0.0103774f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7615 N_VGND_c_12772_n N_A_7939_911#_c_15120_n 0.00694621f $X=44.265 $Y=4.995
+ $X2=25.99 $Y2=0.64
cc_7616 N_VGND_c_12849_n N_A_7939_911#_c_15120_n 0.0589406f $X=44.06 $Y=5.44
+ $X2=25.99 $Y2=0.64
cc_7617 VGND N_A_7939_911#_c_15120_n 0.030408f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=0.64
cc_7618 N_VGND_c_12772_n N_A_7939_911#_c_15121_n 0.00696245f $X=44.265 $Y=4.995
+ $X2=25.99 $Y2=4.8
cc_7619 VGND N_A_7939_911#_c_15122_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7620 N_VGND_c_12892_n N_A_7939_911#_c_15122_n 0.0188215f $X=40.165 $Y=5.44
+ $X2=0 $Y2=0
cc_7621 N_VGND_c_12768_n N_A_7939_911#_c_15123_n 0.0188215f $X=41.105 $Y=5.44
+ $X2=0 $Y2=0
cc_7622 VGND N_A_7939_911#_c_15123_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7623 N_VGND_c_12849_n N_A_7939_911#_c_15153_n 0.0113631f $X=44.06 $Y=5.44
+ $X2=0 $Y2=0
cc_7624 VGND N_A_7939_911#_c_15153_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7625 VGND N_A_9513_66#_M1068_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7626 VGND N_A_9513_66#_M1216_s 0.00215201f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7627 N_VGND_c_12777_n N_A_9513_66#_c_15195_n 0.00696245f $X=46.815 $Y=0.445
+ $X2=0 $Y2=0
cc_7628 N_VGND_c_12863_n N_A_9513_66#_c_15196_n 0.0422314f $X=49.725 $Y=0 $X2=0
+ $Y2=0
cc_7629 VGND N_A_9513_66#_c_15196_n 0.0219908f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7630 N_VGND_c_12777_n N_A_9513_66#_c_15197_n 0.00694621f $X=46.815 $Y=0.445
+ $X2=0 $Y2=0
cc_7631 N_VGND_c_12863_n N_A_9513_66#_c_15197_n 0.0167092f $X=49.725 $Y=0 $X2=0
+ $Y2=0
cc_7632 VGND N_A_9513_66#_c_15197_n 0.00841721f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7633 N_VGND_c_12779_n N_A_9513_66#_c_15198_n 0.0147456f $X=49.89 $Y=0.38
+ $X2=0 $Y2=0
cc_7634 N_VGND_c_12863_n N_A_9513_66#_c_15198_n 0.0614775f $X=49.725 $Y=0 $X2=0
+ $Y2=0
cc_7635 VGND N_A_9513_66#_c_15198_n 0.0325967f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7636 N_VGND_c_12779_n N_A_9513_66#_c_15199_n 0.00959666f $X=49.89 $Y=0.38
+ $X2=25.99 $Y2=0.51
cc_7637 N_VGND_M1068_d N_A_9513_66#_c_15200_n 0.00692362f $X=49.765 $Y=0.235
+ $X2=0 $Y2=0
cc_7638 N_VGND_c_12779_n N_A_9513_66#_c_15200_n 0.0190091f $X=49.89 $Y=0.38
+ $X2=0 $Y2=0
cc_7639 N_VGND_c_12863_n N_A_9513_66#_c_15200_n 0.00262594f $X=49.725 $Y=0 $X2=0
+ $Y2=0
cc_7640 VGND N_A_9513_66#_c_15200_n 0.00940109f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7641 N_VGND_c_12893_n N_A_9513_66#_c_15200_n 0.0020257f $X=50.645 $Y=0 $X2=0
+ $Y2=0
cc_7642 VGND N_A_9513_66#_c_15220_n 0.0121968f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7643 N_VGND_c_12893_n N_A_9513_66#_c_15220_n 0.0188215f $X=50.645 $Y=0 $X2=0
+ $Y2=0
cc_7644 N_VGND_M1115_d N_A_9513_66#_c_15202_n 0.00501873f $X=50.595 $Y=0.235
+ $X2=25.99 $Y2=4.8
cc_7645 N_VGND_c_12781_n N_A_9513_66#_c_15202_n 0.0199861f $X=50.78 $Y=0.38
+ $X2=25.99 $Y2=4.8
cc_7646 VGND N_A_9513_66#_c_15202_n 0.00880092f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.8
cc_7647 N_VGND_c_12893_n N_A_9513_66#_c_15202_n 0.0020257f $X=50.645 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7648 N_VGND_c_12895_n N_A_9513_66#_c_15202_n 0.0020257f $X=51.585 $Y=0
+ $X2=25.99 $Y2=4.8
cc_7649 VGND N_A_9513_66#_c_15229_n 0.0121968f $X=51.665 $Y=-0.085 $X2=25.99
+ $Y2=4.93
cc_7650 N_VGND_c_12895_n N_A_9513_66#_c_15229_n 0.0188215f $X=51.585 $Y=0
+ $X2=25.99 $Y2=4.93
cc_7651 N_VGND_c_12863_n N_A_9513_66#_c_15214_n 0.0113631f $X=49.725 $Y=0 $X2=0
+ $Y2=0
cc_7652 VGND N_A_9513_66#_c_15214_n 0.00572388f $X=51.665 $Y=-0.085 $X2=0 $Y2=0
cc_7653 VGND N_A_9513_918#_M1073_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7654 VGND N_A_9513_918#_M1190_d 0.00215201f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7655 N_VGND_c_12778_n N_A_9513_918#_c_15279_n 0.00696245f $X=46.815 $Y=4.995
+ $X2=0 $Y2=0
cc_7656 N_VGND_c_12865_n N_A_9513_918#_c_15280_n 0.0422314f $X=49.725 $Y=5.44
+ $X2=0 $Y2=0
cc_7657 VGND N_A_9513_918#_c_15280_n 0.0219908f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7658 N_VGND_c_12778_n N_A_9513_918#_c_15281_n 0.00694621f $X=46.815 $Y=4.995
+ $X2=0 $Y2=0
cc_7659 N_VGND_c_12865_n N_A_9513_918#_c_15281_n 0.0167092f $X=49.725 $Y=5.44
+ $X2=0 $Y2=0
cc_7660 VGND N_A_9513_918#_c_15281_n 0.00841721f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7661 N_VGND_c_12780_n N_A_9513_918#_c_15282_n 0.0147456f $X=49.89 $Y=5.06
+ $X2=0 $Y2=0
cc_7662 N_VGND_c_12865_n N_A_9513_918#_c_15282_n 0.0614775f $X=49.725 $Y=5.44
+ $X2=0 $Y2=0
cc_7663 VGND N_A_9513_918#_c_15282_n 0.0325967f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7664 N_VGND_c_12780_n N_A_9513_918#_c_15283_n 0.00959666f $X=49.89 $Y=5.06
+ $X2=25.99 $Y2=0.51
cc_7665 N_VGND_M1073_s N_A_9513_918#_c_15284_n 0.00692362f $X=49.765 $Y=4.555
+ $X2=0 $Y2=0
cc_7666 N_VGND_c_12780_n N_A_9513_918#_c_15284_n 0.0190091f $X=49.89 $Y=5.06
+ $X2=0 $Y2=0
cc_7667 N_VGND_c_12865_n N_A_9513_918#_c_15284_n 0.00262594f $X=49.725 $Y=5.44
+ $X2=0 $Y2=0
cc_7668 VGND N_A_9513_918#_c_15284_n 0.00940109f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7669 N_VGND_c_12894_n N_A_9513_918#_c_15284_n 0.0020257f $X=50.645 $Y=5.44
+ $X2=0 $Y2=0
cc_7670 N_VGND_M1144_s N_A_9513_918#_c_15304_n 0.00501873f $X=50.595 $Y=4.555
+ $X2=0 $Y2=0
cc_7671 N_VGND_c_12782_n N_A_9513_918#_c_15304_n 0.0199861f $X=50.78 $Y=5.06
+ $X2=0 $Y2=0
cc_7672 VGND N_A_9513_918#_c_15304_n 0.00880092f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7673 N_VGND_c_12894_n N_A_9513_918#_c_15304_n 0.0020257f $X=50.645 $Y=5.44
+ $X2=0 $Y2=0
cc_7674 N_VGND_c_12896_n N_A_9513_918#_c_15304_n 0.0020257f $X=51.585 $Y=5.44
+ $X2=0 $Y2=0
cc_7675 N_VGND_c_12865_n N_A_9513_918#_c_15298_n 0.0113631f $X=49.725 $Y=5.44
+ $X2=0 $Y2=0
cc_7676 VGND N_A_9513_918#_c_15298_n 0.00572388f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7677 VGND N_A_9513_918#_c_15286_n 0.0121968f $X=51.665 $Y=5.355 $X2=25.99
+ $Y2=4.93
cc_7678 N_VGND_c_12894_n N_A_9513_918#_c_15286_n 0.0188215f $X=50.645 $Y=5.44
+ $X2=25.99 $Y2=4.93
cc_7679 VGND N_A_9513_918#_c_15287_n 0.0121968f $X=51.665 $Y=5.355 $X2=0 $Y2=0
cc_7680 N_VGND_c_12896_n N_A_9513_918#_c_15287_n 0.0188215f $X=51.585 $Y=5.44
+ $X2=0 $Y2=0
