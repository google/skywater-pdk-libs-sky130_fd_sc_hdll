* File: sky130_fd_sc_hdll__nor2b_1.pxi.spice
* Created: Thu Aug 27 19:15:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%B_N N_B_N_M1005_g N_B_N_c_38_n N_B_N_M1001_g B_N
+ B_N B_N PM_SKY130_FD_SC_HDLL__NOR2B_1%B_N
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%A N_A_c_63_n N_A_M1003_g N_A_c_64_n N_A_M1000_g
+ A PM_SKY130_FD_SC_HDLL__NOR2B_1%A
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_95_n N_A_27_47#_M1002_g N_A_27_47#_c_96_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_97_n N_A_27_47#_c_100_n N_A_27_47#_c_101_n N_A_27_47#_c_128_p
+ N_A_27_47#_c_102_n N_A_27_47#_c_129_p N_A_27_47#_c_103_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%VPWR N_VPWR_M1001_d N_VPWR_c_151_n
+ N_VPWR_c_152_n N_VPWR_c_153_n VPWR N_VPWR_c_154_n N_VPWR_c_150_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%Y N_Y_M1003_d N_Y_M1004_d N_Y_c_185_n
+ N_Y_c_180_n N_Y_c_181_n Y N_Y_c_183_n N_Y_c_182_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR2B_1%VGND N_VGND_M1005_d N_VGND_M1002_d
+ N_VGND_c_220_n N_VGND_c_221_n N_VGND_c_222_n VGND N_VGND_c_223_n
+ N_VGND_c_224_n N_VGND_c_225_n PM_SKY130_FD_SC_HDLL__NOR2B_1%VGND
cc_1 VNB N_B_N_M1005_g 0.0348101f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.445
cc_2 VNB N_B_N_c_38_n 0.029001f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB B_N 0.00911129f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.105
cc_4 VNB N_A_c_63_n 0.0182422f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.975
cc_5 VNB N_A_c_64_n 0.0229012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB A 0.00404492f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_7 VNB N_A_27_47#_c_95_n 0.0198334f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_8 VNB N_A_27_47#_c_96_n 0.0307354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_97_n 0.0481569f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_10 VNB N_VPWR_c_150_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_180_n 0.0187035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_181_n 0.00447608f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_13 VNB N_Y_c_182_n 0.0200443f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.62
cc_14 VNB N_VGND_c_220_n 0.00537507f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_221_n 0.0149656f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_16 VNB N_VGND_c_222_n 0.0216692f $X=-0.19 $Y=-0.24 $X2=0.65 $Y2=1.16
cc_17 VNB N_VGND_c_223_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.62
cc_18 VNB N_VGND_c_224_n 0.0269944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_225_n 0.14317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VPB N_B_N_c_38_n 0.0301157f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_21 VPB B_N 0.00192025f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.105
cc_22 VPB N_A_c_64_n 0.0278377f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_23 VPB A 0.0022879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_24 VPB N_A_27_47#_c_96_n 0.031382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_27_47#_c_97_n 0.0253182f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.16
cc_26 VPB N_A_27_47#_c_100_n 0.0105896f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.62
cc_27 VPB N_A_27_47#_c_101_n 0.0110324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_102_n 7.36918e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_103_n 0.00267601f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_151_n 0.0120199f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_31 VPB N_VPWR_c_152_n 0.0237696f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.495
cc_32 VPB N_VPWR_c_153_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_154_n 0.0320631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_150_n 0.0528939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_Y_c_183_n 0.0361418f $X=-0.19 $Y=1.305 $X2=0.65 $Y2=1.62
cc_36 VPB N_Y_c_182_n 0.0273389f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.62
cc_37 N_B_N_M1005_g N_A_c_63_n 0.0148191f $X=0.47 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_38 N_B_N_c_38_n N_A_c_63_n 6.53552e-19 $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_39 B_N N_A_c_63_n 4.02551e-19 $X=0.56 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_40 N_B_N_c_38_n N_A_c_64_n 0.0326374f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_41 B_N N_A_c_64_n 0.0083951f $X=0.56 $Y=1.105 $X2=0 $Y2=0
cc_42 N_B_N_c_38_n A 7.87155e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_43 B_N A 0.0213193f $X=0.56 $Y=1.105 $X2=0 $Y2=0
cc_44 N_B_N_M1005_g N_A_27_47#_c_97_n 0.0244057f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_45 N_B_N_c_38_n N_A_27_47#_c_97_n 0.00727842f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_46 B_N N_A_27_47#_c_97_n 0.0583295f $X=0.56 $Y=1.105 $X2=0 $Y2=0
cc_47 N_B_N_c_38_n N_A_27_47#_c_100_n 0.0158386f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_48 B_N N_A_27_47#_c_100_n 0.019153f $X=0.56 $Y=1.105 $X2=0 $Y2=0
cc_49 B_N N_VPWR_M1001_d 0.00551439f $X=0.56 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_50 N_B_N_c_38_n N_VPWR_c_152_n 6.43543e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_B_N_M1005_g N_Y_c_185_n 5.34268e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_52 N_B_N_M1005_g N_Y_c_181_n 7.95218e-19 $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_53 N_B_N_M1005_g N_VGND_c_220_n 0.00779852f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_54 N_B_N_c_38_n N_VGND_c_220_n 4.24353e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 B_N N_VGND_c_220_n 0.00564805f $X=0.56 $Y=1.105 $X2=0 $Y2=0
cc_56 N_B_N_M1005_g N_VGND_c_224_n 0.00585385f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_57 N_B_N_M1005_g N_VGND_c_225_n 0.0123468f $X=0.47 $Y=0.445 $X2=0 $Y2=0
cc_58 N_A_c_63_n N_A_27_47#_c_95_n 0.0124776f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A_c_64_n N_A_27_47#_c_96_n 0.0914717f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_60 A N_A_27_47#_c_96_n 0.00167429f $X=1.03 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A_c_64_n N_A_27_47#_c_100_n 0.0165236f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_62 A N_A_27_47#_c_100_n 0.00762929f $X=1.03 $Y=1.105 $X2=0 $Y2=0
cc_63 N_A_c_64_n N_A_27_47#_c_102_n 0.00202023f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_64_n N_A_27_47#_c_103_n 3.09497e-19 $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_65 A N_A_27_47#_c_103_n 0.0176977f $X=1.03 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A_c_64_n N_VPWR_c_151_n 0.0101724f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_c_64_n N_VPWR_c_154_n 0.00452725f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_c_64_n N_VPWR_c_150_n 0.00505132f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_c_63_n N_Y_c_185_n 0.00847537f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_c_63_n N_Y_c_181_n 0.00593404f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_c_64_n N_Y_c_181_n 0.00173954f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_72 A N_Y_c_181_n 0.0120409f $X=1.03 $Y=1.105 $X2=0 $Y2=0
cc_73 N_A_c_64_n N_Y_c_183_n 0.00151471f $X=1.175 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_63_n N_VGND_c_220_n 0.00456426f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_75 A N_VGND_c_220_n 3.46307e-19 $X=1.03 $Y=1.105 $X2=0 $Y2=0
cc_76 N_A_c_63_n N_VGND_c_223_n 0.00465454f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_c_63_n N_VGND_c_225_n 0.00832637f $X=1.14 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_100_n N_VPWR_M1001_d 0.00969636f $X=1.315 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_27_47#_c_96_n N_VPWR_c_151_n 0.00169453f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_100_n N_VPWR_c_151_n 0.0206557f $X=1.315 $Y=2 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_100_n N_VPWR_c_152_n 0.00784038f $X=1.315 $Y=2 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_101_n N_VPWR_c_152_n 0.0050551f $X=0.345 $Y=2 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_96_n N_VPWR_c_154_n 0.00673617f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_100_n N_VPWR_c_154_n 0.00579285f $X=1.315 $Y=2 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_96_n N_VPWR_c_150_n 0.0129495f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_100_n N_VPWR_c_150_n 0.023851f $X=1.315 $Y=2 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_101_n N_VPWR_c_150_n 0.00750746f $X=0.345 $Y=2 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_100_n A_253_297# 0.00208567f $X=1.315 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_27_47#_c_128_p A_253_297# 3.43001e-19 $X=1.4 $Y=1.915 $X2=-0.19
+ $Y2=-0.24
cc_90 N_A_27_47#_c_129_p A_253_297# 0.00265027f $X=1.57 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_27_47#_c_95_n N_Y_c_185_n 0.0114377f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_95_n N_Y_c_180_n 0.010459f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_96_n N_Y_c_180_n 0.00582747f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_103_n N_Y_c_180_n 0.0246339f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_95_n N_Y_c_181_n 9.82755e-19 $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_129_p N_Y_c_181_n 0.00491873f $X=1.57 $Y=1.58 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_103_n N_Y_c_181_n 0.00225036f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_96_n N_Y_c_183_n 0.0109734f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_103_n N_Y_c_183_n 0.00580676f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_95_n N_Y_c_182_n 0.00267478f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_96_n N_Y_c_182_n 0.0177208f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_102_n N_Y_c_182_n 0.00668124f $X=1.57 $Y=1.495 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_129_p N_Y_c_182_n 0.00698945f $X=1.57 $Y=1.58 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_103_n N_Y_c_182_n 0.019076f $X=1.65 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_95_n N_VGND_c_222_n 0.00578121f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_95_n N_VGND_c_223_n 0.00423334f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_27_47#_c_97_n N_VGND_c_224_n 0.0141133f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1005_s N_VGND_c_225_n 0.00388646f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_c_95_n N_VGND_c_225_n 0.00699781f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_97_n N_VGND_c_225_n 0.00938686f $X=0.26 $Y=0.455 $X2=0 $Y2=0
cc_111 N_VPWR_c_150_n A_253_297# 0.00299419f $X=2.07 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_112 N_VPWR_c_150_n N_Y_M1004_d 0.00217517f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_113 N_VPWR_c_151_n N_Y_c_183_n 0.0062597f $X=0.94 $Y=2.34 $X2=0 $Y2=0
cc_114 N_VPWR_c_154_n N_Y_c_183_n 0.0373819f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_c_150_n N_Y_c_183_n 0.0212921f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_116 N_Y_c_180_n N_VGND_M1002_d 0.00413739f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_117 N_Y_c_185_n N_VGND_c_220_n 0.0287408f $X=1.35 $Y=0.39 $X2=0 $Y2=0
cc_118 N_Y_c_180_n N_VGND_c_221_n 0.00162138f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_119 N_Y_c_185_n N_VGND_c_222_n 0.0195332f $X=1.35 $Y=0.39 $X2=0 $Y2=0
cc_120 N_Y_c_180_n N_VGND_c_222_n 0.0311856f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_121 N_Y_c_185_n N_VGND_c_223_n 0.0222324f $X=1.35 $Y=0.39 $X2=0 $Y2=0
cc_122 N_Y_c_180_n N_VGND_c_223_n 0.00265794f $X=2.035 $Y=0.81 $X2=0 $Y2=0
cc_123 N_Y_M1003_d N_VGND_c_225_n 0.00215201f $X=1.215 $Y=0.235 $X2=0 $Y2=0
cc_124 N_Y_c_185_n N_VGND_c_225_n 0.0138958f $X=1.35 $Y=0.39 $X2=0 $Y2=0
cc_125 N_Y_c_180_n N_VGND_c_225_n 0.0094271f $X=2.035 $Y=0.81 $X2=0 $Y2=0
