* File: sky130_fd_sc_hdll__mux2i_1.pex.spice
* Created: Wed Sep  2 08:34:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A0 1 3 4 6 7 12
c27 12 0 6.12641e-20 $X=0.515 $Y=1.202
r28 12 13 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r29 10 12 34.5234 $w=3.63e-07 $l=2.6e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.515 $Y2=1.202
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r31 4 13 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r32 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r33 1 12 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r34 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A1 1 3 4 6 9 13 14
c35 13 0 6.12641e-20 $X=1.15 $Y=1.53
c36 9 0 1.72057e-19 $X=1.09 $Y=1.16
c37 4 0 1.20436e-19 $X=0.985 $Y=1.41
r38 13 14 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=1.165 $Y=1.53
+ $X2=1.165 $Y2=1.87
r39 12 13 11.3682 $w=1.98e-07 $l=2.05e-07 $layer=LI1_cond $X=1.165 $Y=1.325
+ $X2=1.165 $Y2=1.53
r40 9 12 7.95677 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=1.16
+ $X2=1.135 $Y2=1.325
r41 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.09
+ $Y=1.16 $X2=1.09 $Y2=1.16
r42 4 10 46.6797 $w=3.23e-07 $l=2.8592e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=1.062 $Y2=1.16
r43 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r44 1 10 38.5615 $w=3.23e-07 $l=2.09893e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=1.062 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A_303_205# 1 2 7 9 12 14 17 21 25 27
r67 23 27 4.98924 $w=2.45e-07 $l=1.27609e-07 $layer=LI1_cond $X=3.082 $Y=1.31
+ $X2=3.062 $Y2=1.192
r68 23 25 33.2928 $w=2.23e-07 $l=6.5e-07 $layer=LI1_cond $X=3.082 $Y=1.31
+ $X2=3.082 $Y2=1.96
r69 19 27 4.98924 $w=2.45e-07 $l=1.17e-07 $layer=LI1_cond $X=3.062 $Y=1.075
+ $X2=3.062 $Y2=1.192
r70 19 21 28.4849 $w=2.63e-07 $l=6.55e-07 $layer=LI1_cond $X=3.062 $Y=1.075
+ $X2=3.062 $Y2=0.42
r71 17 30 33.1375 $w=3.2e-07 $l=2.2e-07 $layer=POLY_cond $X=1.68 $Y=1.217
+ $X2=1.9 $Y2=1.217
r72 17 28 9.79062 $w=3.2e-07 $l=6.5e-08 $layer=POLY_cond $X=1.68 $Y=1.217
+ $X2=1.615 $Y2=1.217
r73 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.68
+ $Y=1.16 $X2=1.68 $Y2=1.16
r74 14 27 1.49305 $w=2.35e-07 $l=1.32e-07 $layer=LI1_cond $X=2.93 $Y=1.192
+ $X2=3.062 $Y2=1.192
r75 14 16 61.3002 $w=2.33e-07 $l=1.25e-06 $layer=LI1_cond $X=2.93 $Y=1.192
+ $X2=1.68 $Y2=1.192
r76 10 30 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.9 $Y=1.025
+ $X2=1.9 $Y2=1.217
r77 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.9 $Y=1.025
+ $X2=1.9 $Y2=0.56
r78 7 28 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.615 $Y=1.41
+ $X2=1.615 $Y2=1.217
r79 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.615 $Y=1.41
+ $X2=1.615 $Y2=1.985
r80 2 25 300 $w=1.7e-07 $l=5.38284e-07 $layer=licon1_PDIFF $count=2 $X=2.975
+ $Y=1.485 $X2=3.11 $Y2=1.96
r81 1 21 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.965
+ $Y=0.235 $X2=3.11 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%S 3 5 7 8 10 12 13 15 16 17 18 19
r57 24 26 11.9882 $w=3.9e-07 $l=9.7e-08 $layer=POLY_cond $X=3.497 $Y=1.16
+ $X2=3.497 $Y2=1.257
r58 18 19 11.0754 $w=3.83e-07 $l=3.7e-07 $layer=LI1_cond $X=3.557 $Y=1.16
+ $X2=3.557 $Y2=1.53
r59 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.59
+ $Y=1.16 $X2=3.59 $Y2=1.16
r60 17 18 9.27941 $w=3.83e-07 $l=3.1e-07 $layer=LI1_cond $X=3.557 $Y=0.85
+ $X2=3.557 $Y2=1.16
r61 13 24 40.0132 $w=3.9e-07 $l=2.17002e-07 $layer=POLY_cond $X=3.39 $Y=0.99
+ $X2=3.497 $Y2=1.16
r62 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.39 $Y=0.99
+ $X2=3.39 $Y2=0.56
r63 10 26 33.0095 $w=3.9e-07 $l=2.08818e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.497 $Y2=1.257
r64 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r65 9 16 3.69004 $w=1.85e-07 $l=1.14018e-07 $layer=POLY_cond $X=2.445 $Y=1.257
+ $X2=2.345 $Y2=1.287
r66 8 26 20.2722 $w=1.85e-07 $l=2.32e-07 $layer=POLY_cond $X=3.265 $Y=1.257
+ $X2=3.497 $Y2=1.257
r67 8 9 302.927 $w=1.85e-07 $l=8.2e-07 $layer=POLY_cond $X=3.265 $Y=1.257
+ $X2=2.445 $Y2=1.257
r68 5 16 22.4247 $w=1.65e-07 $l=1.23e-07 $layer=POLY_cond $X=2.345 $Y=1.41
+ $X2=2.345 $Y2=1.287
r69 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.345 $Y=1.41
+ $X2=2.345 $Y2=1.985
r70 1 16 22.4247 $w=1.65e-07 $l=1.33918e-07 $layer=POLY_cond $X=2.32 $Y=1.165
+ $X2=2.345 $Y2=1.287
r71 1 3 310.223 $w=1.5e-07 $l=6.05e-07 $layer=POLY_cond $X=2.32 $Y=1.165
+ $X2=2.32 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_297# 1 2 7 9 11 14 15 16 17 19
c45 16 0 1.20436e-19 $X=1.725 $Y=1.565
r46 17 24 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=1.65
+ $X2=2.555 $Y2=1.565
r47 17 19 20.3194 $w=3.78e-07 $l=6.7e-07 $layer=LI1_cond $X=2.555 $Y=1.65
+ $X2=2.555 $Y2=2.32
r48 15 24 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.365 $Y=1.565
+ $X2=2.555 $Y2=1.565
r49 15 16 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.365 $Y=1.565
+ $X2=1.725 $Y2=1.565
r50 13 16 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.615 $Y=1.65
+ $X2=1.725 $Y2=1.565
r51 13 14 33.7875 $w=2.18e-07 $l=6.45e-07 $layer=LI1_cond $X=1.615 $Y=1.65
+ $X2=1.615 $Y2=2.295
r52 12 22 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.42 $Y=2.38 $X2=0.27
+ $Y2=2.38
r53 11 14 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.505 $Y=2.38
+ $X2=1.615 $Y2=2.295
r54 11 12 70.7861 $w=1.68e-07 $l=1.085e-06 $layer=LI1_cond $X=1.505 $Y=2.38
+ $X2=0.42 $Y2=2.38
r55 7 22 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.27 $Y=2.295 $X2=0.27
+ $Y2=2.38
r56 7 9 25.93 $w=2.98e-07 $l=6.75e-07 $layer=LI1_cond $X=0.27 $Y=2.295 $X2=0.27
+ $Y2=1.62
r57 2 24 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.485 $X2=2.58 $Y2=1.64
r58 2 19 400 $w=1.7e-07 $l=9.04599e-07 $layer=licon1_PDIFF $count=1 $X=2.435
+ $Y=1.485 $X2=2.58 $Y2=2.32
r59 1 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r60 1 9 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%Y 1 2 7 8 15
r21 7 18 2.871 $w=2.83e-07 $l=7.1e-08 $layer=LI1_cond $X=0.747 $Y=1.526
+ $X2=0.747 $Y2=1.597
r22 7 25 3.33382 $w=2.83e-07 $l=7.1e-08 $layer=LI1_cond $X=0.747 $Y=1.526
+ $X2=0.747 $Y2=1.455
r23 7 8 10.6753 $w=2.83e-07 $l=2.64e-07 $layer=LI1_cond $X=0.747 $Y=1.606
+ $X2=0.747 $Y2=1.87
r24 7 18 0.363929 $w=2.83e-07 $l=9e-09 $layer=LI1_cond $X=0.747 $Y=1.606
+ $X2=0.747 $Y2=1.597
r25 7 25 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=0.72 $Y=1.45 $X2=0.72
+ $Y2=1.455
r26 7 15 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=0.72 $Y=1.45 $X2=0.72
+ $Y2=0.76
r27 2 7 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.62
r28 1 15 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%VPWR 1 2 9 13 16 17 18 20 36 37 40
r40 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r42 34 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r43 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r45 31 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 30 33 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 28 40 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.175 $Y=2.72
+ $X2=2.035 $Y2=2.72
r49 28 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=2.175 $Y=2.72
+ $X2=2.53 $Y2=2.72
r50 27 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 22 26 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r53 20 40 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.035 $Y2=2.72
r54 20 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r55 18 27 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r56 18 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 16 33 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 16 17 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=3.475 $Y=2.72
+ $X2=3.622 $Y2=2.72
r59 15 36 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=3.77 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 15 17 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.77 $Y=2.72
+ $X2=3.622 $Y2=2.72
r61 11 17 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.622 $Y=2.635
+ $X2=3.622 $Y2=2.72
r62 11 13 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=3.622 $Y=2.635
+ $X2=3.622 $Y2=2
r63 7 40 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=2.635
+ $X2=2.035 $Y2=2.72
r64 7 9 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.035 $Y=2.635
+ $X2=2.035 $Y2=2
r65 2 13 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2
r66 1 9 300 $w=1.7e-07 $l=6.37848e-07 $layer=licon1_PDIFF $count=2 $X=1.705
+ $Y=1.485 $X2=1.98 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A_27_47# 1 2 9 13 15 20 21
r27 20 21 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=0.44 $Y=0.34
+ $X2=1.065 $Y2=0.34
r28 13 21 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=1.275 $Y=0.36
+ $X2=1.065 $Y2=0.36
r29 13 15 21.9177 $w=2.08e-07 $l=4.15e-07 $layer=LI1_cond $X=1.275 $Y=0.36
+ $X2=1.69 $Y2=0.36
r30 7 20 12.318 $w=2.08e-07 $l=2.25e-07 $layer=LI1_cond $X=0.215 $Y=0.36
+ $X2=0.44 $Y2=0.36
r31 7 9 11.3028 $w=2.58e-07 $l=2.55e-07 $layer=LI1_cond $X=0.215 $Y=0.465
+ $X2=0.215 $Y2=0.72
r32 2 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.69 $Y2=0.38
r33 1 7 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r34 1 9 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%A_207_47# 1 2 11 15 17 18
r36 17 18 8.76859 $w=2.28e-07 $l=1.75e-07 $layer=LI1_cond $X=1.575 $Y=0.77
+ $X2=1.75 $Y2=0.77
r37 13 15 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=2.582 $Y=0.715
+ $X2=2.582 $Y2=0.55
r38 11 13 7.04737 $w=1.7e-07 $l=1.53734e-07 $layer=LI1_cond $X=2.465 $Y=0.8
+ $X2=2.582 $Y2=0.715
r39 11 18 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.465 $Y=0.8
+ $X2=1.75 $Y2=0.8
r40 9 17 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=1.17 $Y=0.74
+ $X2=1.575 $Y2=0.74
r41 2 15 182 $w=1.7e-07 $l=3.88844e-07 $layer=licon1_NDIFF $count=1 $X=2.395
+ $Y=0.235 $X2=2.56 $Y2=0.55
r42 1 9 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.17 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_1%VGND 1 2 9 13 16 17 18 20 33 34 37
r44 37 38 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r46 31 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r47 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r48 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r49 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r50 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r51 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 25 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.11
+ $Y2=0
r53 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.53
+ $Y2=0
r54 20 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.11
+ $Y2=0
r55 20 22 117.107 $w=1.68e-07 $l=1.795e-06 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=0.23 $Y2=0
r56 18 38 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.07
+ $Y2=0
r57 18 22 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 16 30 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.45
+ $Y2=0
r59 16 17 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.625
+ $Y2=0
r60 15 33 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.91
+ $Y2=0
r61 15 17 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=3.735 $Y=0 $X2=3.625
+ $Y2=0
r62 11 17 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0
r63 11 13 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.625 $Y=0.085
+ $X2=3.625 $Y2=0.38
r64 7 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=0.085 $X2=2.11
+ $Y2=0
r65 7 9 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.11 $Y=0.085
+ $X2=2.11 $Y2=0.36
r66 2 13 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.235 $X2=3.6 $Y2=0.38
r67 1 9 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=1.975
+ $Y=0.235 $X2=2.11 $Y2=0.36
.ends

