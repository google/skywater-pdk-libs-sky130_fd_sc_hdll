# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a22oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a22oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 1.075000 3.535000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.770000 1.075000 4.620000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 1.075000 1.745000 1.275000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.150000 1.075000 0.830000 1.275000 ;
    END
  END B2
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 5.250000 2.910000 ;
    END
  END VPB
  PIN Y
    ANTENNADIFFAREA  1.278500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.485000 2.360000 1.655000 ;
        RECT 0.095000 1.655000 0.345000 2.465000 ;
        RECT 0.985000 1.655000 1.365000 2.125000 ;
        RECT 1.455000 0.675000 3.295000 0.845000 ;
        RECT 1.925000 1.655000 2.360000 2.125000 ;
        RECT 1.930000 0.845000 2.360000 1.485000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.060000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.510000 ;
        RECT 3.980000  0.085000 4.360000 0.510000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.060000 2.805000 ;
        RECT 3.045000 1.825000 3.215000 2.635000 ;
        RECT 4.085000 1.825000 4.255000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.095000 0.255000 0.345000 0.680000 ;
      RECT 0.095000 0.680000 1.285000 0.850000 ;
      RECT 0.515000 1.825000 0.815000 2.295000 ;
      RECT 0.515000 2.295000 2.825000 2.465000 ;
      RECT 1.115000 0.255000 2.305000 0.505000 ;
      RECT 1.115000 0.505000 1.285000 0.680000 ;
      RECT 1.585000 1.825000 1.755000 2.295000 ;
      RECT 2.495000 0.255000 3.785000 0.505000 ;
      RECT 2.575000 1.485000 4.805000 1.655000 ;
      RECT 2.575000 1.655000 2.825000 2.295000 ;
      RECT 3.385000 1.655000 3.865000 2.465000 ;
      RECT 3.615000 0.505000 3.785000 0.680000 ;
      RECT 3.615000 0.680000 4.875000 0.850000 ;
      RECT 4.425000 1.655000 4.805000 2.465000 ;
      RECT 4.555000 0.255000 4.875000 0.680000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a22oi_2
END LIBRARY
