* File: sky130_fd_sc_hdll__dlygate4sd1_1.spice
* Created: Wed Sep  2 08:30:15 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__dlygate4sd1_1.pex.spice"
.subckt sky130_fd_sc_hdll__dlygate4sd1_1  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1000 N_A_213_47#_M1000_d N_A_27_47#_M1000_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0672 PD=1.36 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_A_213_47#_M1006_g N_A_319_93#_M1006_s VNB NSHORT L=0.15
+ W=0.42 AD=0.145037 AS=0.1344 PD=0.977383 PS=1.48 NRD=82.944 NRS=15.708 M=1
+ R=2.8 SA=75000.2 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_319_93#_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.224463 PD=1.82 PS=1.51262 NRD=0 NRS=31.38 M=1 R=4.33333
+ SA=75000.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1176 PD=0.71 PS=1.4 NRD=0 NRS=7.0329 M=1 R=2.33333 SA=90000.2
+ SB=90000.6 A=0.0756 P=1.2 MULT=1
MM1004 N_A_213_47#_M1004_d N_A_27_47#_M1004_g N_VPWR_M1007_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1092 AS=0.0609 PD=1.36 PS=0.71 NRD=0 NRS=7.0329 M=1 R=2.33333
+ SA=90000.7 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1002 N_VPWR_M1002_d N_A_213_47#_M1002_g N_A_319_93#_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.148331 AS=0.1176 PD=0.913944 PS=1.4 NRD=58.6272 NRS=7.0329 M=1
+ R=2.33333 SA=90000.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1003 N_X_M1003_d N_A_319_93#_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.28 AS=0.353169 PD=2.56 PS=2.17606 NRD=2.9353 NRS=27.5603 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hdll__dlygate4sd1_1.pxi.spice"
*
.ends
*
*
