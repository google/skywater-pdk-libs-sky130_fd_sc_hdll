* File: sky130_fd_sc_hdll__a21bo_1.spice
* Created: Thu Aug 27 18:52:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21bo_1.pex.spice"
.subckt sky130_fd_sc_hdll__a21bo_1  VNB VPB B1_N A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_B1_N_M1004_g N_A_27_413#_M1004_s VNB NSHORT L=0.15
+ W=0.42 AD=0.127688 AS=0.1323 PD=0.942056 PS=1.47 NRD=36.42 NRS=14.28 M=1 R=2.8
+ SA=75000.2 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1003 N_A_235_297#_M1003_d N_A_27_413#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.197612 PD=0.92 PS=1.45794 NRD=0 NRS=26.76 M=1 R=4.33333
+ SA=75000.7 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1001 A_412_47# N_A1_M1001_g N_A_235_297#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.08775 PD=0.98 PS=0.92 NRD=20.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A2_M1006_g A_412_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.290875 AS=0.10725 PD=1.545 PS=0.98 NRD=23.988 NRS=20.304 M=1 R=4.33333
+ SA=75001.6 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1005_d N_A_235_297#_M1005_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.24375 AS=0.290875 PD=2.05 PS=1.545 NRD=20.304 NRS=24.912 M=1 R=4.33333
+ SA=75002.7 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_B1_N_M1002_g N_A_27_413#_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1008 N_A_326_297#_M1008_d N_A_27_413#_M1008_g N_A_235_297#_M1008_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.275 PD=1.29 PS=2.55 NRD=0.9653 NRS=1.9503 M=1
+ R=5.55556 SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A1_M1007_g N_A_326_297#_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.145 PD=1.3 PS=1.29 NRD=1.9503 NRS=0.9653 M=1 R=5.55556 SA=90000.7
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_326_297#_M1000_d N_A2_M1000_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1009 N_X_M1009_d N_A_235_297#_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.385 AS=0.27 PD=2.77 PS=2.54 NRD=23.6203 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__a21bo_1.pxi.spice"
*
.ends
*
*
