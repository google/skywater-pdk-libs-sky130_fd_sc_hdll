# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dlxtn_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  6.440000 BY  2.720000 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.465000 0.955000 1.890000 1.325000 ;
    END
  END D
  PIN GATE_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.985000 0.330000 1.625000 ;
    END
  END GATE_N
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.625000 0.415000 5.910000 0.825000 ;
        RECT 5.625000 1.495000 5.910000 2.455000 ;
        RECT 5.740000 0.825000 5.910000 0.995000 ;
        RECT 5.740000 0.995000 6.345000 1.325000 ;
        RECT 5.740000 1.325000 5.910000 1.495000 ;
    END
  END Q
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.175000  0.345000 0.345000 0.635000 ;
      RECT 0.175000  0.635000 0.830000 0.805000 ;
      RECT 0.175000  1.795000 0.830000 1.965000 ;
      RECT 0.175000  1.965000 0.345000 2.465000 ;
      RECT 0.515000  0.085000 0.895000 0.465000 ;
      RECT 0.515000  2.135000 0.895000 2.635000 ;
      RECT 0.660000  0.805000 0.830000 1.070000 ;
      RECT 0.660000  1.070000 0.890000 1.400000 ;
      RECT 0.660000  1.400000 0.830000 1.795000 ;
      RECT 1.115000  0.345000 1.285000 1.685000 ;
      RECT 1.115000  1.685000 1.340000 2.465000 ;
      RECT 1.555000  1.495000 2.290000 1.665000 ;
      RECT 1.555000  1.665000 1.885000 2.415000 ;
      RECT 1.635000  0.345000 1.805000 0.615000 ;
      RECT 1.635000  0.615000 2.290000 0.765000 ;
      RECT 1.635000  0.765000 2.540000 0.785000 ;
      RECT 1.975000  0.085000 2.355000 0.445000 ;
      RECT 2.105000  1.835000 2.420000 2.635000 ;
      RECT 2.120000  0.785000 2.540000 1.095000 ;
      RECT 2.120000  1.095000 2.290000 1.495000 ;
      RECT 2.670000  1.355000 2.955000 2.005000 ;
      RECT 2.915000  0.705000 3.340000 1.035000 ;
      RECT 3.085000  0.365000 3.795000 0.535000 ;
      RECT 3.145000  2.255000 3.945000 2.425000 ;
      RECT 3.170000  1.035000 3.340000 1.415000 ;
      RECT 3.170000  1.415000 3.510000 1.995000 ;
      RECT 3.625000  0.535000 3.795000 0.995000 ;
      RECT 3.625000  0.995000 4.545000 1.165000 ;
      RECT 3.775000  1.165000 4.545000 1.325000 ;
      RECT 3.775000  1.325000 3.945000 2.255000 ;
      RECT 4.035000  0.085000 4.415000 0.825000 ;
      RECT 4.165000  2.135000 4.465000 2.635000 ;
      RECT 4.185000  1.535000 4.905000 1.865000 ;
      RECT 4.685000  0.415000 4.905000 0.825000 ;
      RECT 4.685000  1.865000 4.905000 2.435000 ;
      RECT 4.735000  0.825000 4.905000 0.995000 ;
      RECT 4.735000  0.995000 5.535000 1.325000 ;
      RECT 4.735000  1.325000 4.905000 1.535000 ;
      RECT 5.135000  0.085000 5.405000 0.825000 ;
      RECT 5.135000  1.495000 5.405000 2.635000 ;
      RECT 6.095000  0.085000 6.355000 0.550000 ;
      RECT 6.095000  1.755000 6.345000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 0.660000  1.445000 0.830000 1.615000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.170000  1.785000 1.340000 1.955000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.670000  1.785000 2.840000 1.955000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.175000  1.445000 3.345000 1.615000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 0.600000 1.415000 0.890000 1.460000 ;
      RECT 0.600000 1.460000 3.405000 1.600000 ;
      RECT 0.600000 1.600000 0.890000 1.645000 ;
      RECT 1.110000 1.755000 1.400000 1.800000 ;
      RECT 1.110000 1.800000 2.900000 1.940000 ;
      RECT 1.110000 1.940000 1.400000 1.985000 ;
      RECT 2.610000 1.755000 2.900000 1.800000 ;
      RECT 2.610000 1.940000 2.900000 1.985000 ;
      RECT 3.115000 1.415000 3.405000 1.460000 ;
      RECT 3.115000 1.600000 3.405000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlxtn_2
