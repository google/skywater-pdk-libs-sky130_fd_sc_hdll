* File: sky130_fd_sc_hdll__o22ai_1.pxi.spice
* Created: Thu Aug 27 19:21:21 2020
* 
x_PM_SKY130_FD_SC_HDLL__O22AI_1%B1 N_B1_c_43_n N_B1_M1004_g N_B1_c_40_n
+ N_B1_M1005_g B1 N_B1_c_42_n PM_SKY130_FD_SC_HDLL__O22AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O22AI_1%B2 N_B2_c_72_n N_B2_M1003_g N_B2_c_73_n
+ N_B2_M1007_g B2 N_B2_c_74_n PM_SKY130_FD_SC_HDLL__O22AI_1%B2
x_PM_SKY130_FD_SC_HDLL__O22AI_1%A2 N_A2_c_108_n N_A2_M1000_g N_A2_c_109_n
+ N_A2_M1002_g N_A2_c_110_n N_A2_c_111_n N_A2_c_114_n A2
+ PM_SKY130_FD_SC_HDLL__O22AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O22AI_1%A1 N_A1_c_153_n N_A1_M1006_g N_A1_c_154_n
+ N_A1_M1001_g A1 A1 PM_SKY130_FD_SC_HDLL__O22AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O22AI_1%VPWR N_VPWR_M1004_s N_VPWR_M1001_d
+ N_VPWR_c_179_n N_VPWR_c_180_n N_VPWR_c_181_n N_VPWR_c_182_n VPWR
+ N_VPWR_c_183_n N_VPWR_c_178_n PM_SKY130_FD_SC_HDLL__O22AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O22AI_1%Y N_Y_M1005_d N_Y_M1007_d N_Y_c_216_n
+ N_Y_c_230_n N_Y_c_221_n N_Y_c_223_n Y N_Y_c_225_n
+ PM_SKY130_FD_SC_HDLL__O22AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O22AI_1%A_27_47# N_A_27_47#_M1005_s N_A_27_47#_M1003_d
+ N_A_27_47#_M1006_d N_A_27_47#_c_255_n N_A_27_47#_c_268_n N_A_27_47#_c_265_n
+ N_A_27_47#_c_256_n N_A_27_47#_c_257_n PM_SKY130_FD_SC_HDLL__O22AI_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O22AI_1%VGND N_VGND_M1000_d N_VGND_c_302_n
+ N_VGND_c_303_n N_VGND_c_304_n VGND N_VGND_c_305_n N_VGND_c_306_n
+ PM_SKY130_FD_SC_HDLL__O22AI_1%VGND
cc_1 VNB N_B1_c_40_n 0.0198746f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB B1 0.0242951f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_B1_c_42_n 0.0404923f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B2_c_72_n 0.0195857f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B2_c_73_n 0.0277171f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B2_c_74_n 0.00539232f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_7 VNB N_A2_c_108_n 0.0189333f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A2_c_109_n 0.0234643f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB N_A2_c_110_n 0.00394442f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_10 VNB N_A2_c_111_n 6.20736e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_153_n 0.0225937f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_A1_c_154_n 0.0375572f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_13 VNB A1 0.00951235f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_14 VNB N_VPWR_c_178_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Y_c_216_n 0.00356348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_255_n 0.00836668f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_17 VNB N_A_27_47#_c_256_n 0.00773281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_257_n 0.0168702f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_302_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_20 VNB N_VGND_c_303_n 0.047888f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.202
cc_21 VNB N_VGND_c_304_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_22 VNB N_VGND_c_305_n 0.0201058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_306_n 0.162397f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VPB N_B1_c_43_n 0.0197502f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_25 VPB B1 0.0270924f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_26 VPB N_B1_c_42_n 0.0178061f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_27 VPB N_B2_c_73_n 0.0300782f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_28 VPB N_B2_c_74_n 0.00164462f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_29 VPB N_A2_c_109_n 0.0292735f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_30 VPB N_A2_c_111_n 0.00155329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A2_c_114_n 0.00274595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A1_c_154_n 0.0355007f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_33 VPB N_VPWR_c_179_n 0.0103382f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_34 VPB N_VPWR_c_180_n 0.00496839f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.202
cc_35 VPB N_VPWR_c_181_n 0.0115201f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_36 VPB N_VPWR_c_182_n 0.0482466f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_37 VPB N_VPWR_c_183_n 0.0534128f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_178_n 0.0437094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_216_n 0.00136858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_B1_c_40_n N_B2_c_72_n 0.0160471f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_41 N_B1_c_43_n N_B2_c_73_n 0.03229f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_42 N_B1_c_42_n N_B2_c_73_n 0.0160471f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_43 N_B1_c_43_n N_B2_c_74_n 2.31286e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_B1_c_42_n N_B2_c_74_n 3.72959e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_45 B1 N_VPWR_M1004_s 0.0111021f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_46 B1 N_VPWR_c_179_n 8.28574e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_47 N_B1_c_43_n N_VPWR_c_180_n 0.0107271f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_48 B1 N_VPWR_c_180_n 0.0151133f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_49 N_B1_c_43_n N_VPWR_c_183_n 0.00609683f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_50 N_B1_c_43_n N_VPWR_c_178_n 0.0108989f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 B1 N_VPWR_c_178_n 0.00223595f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_52 N_B1_c_43_n N_Y_c_216_n 0.0115629f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_B1_c_40_n N_Y_c_216_n 0.00380314f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 N_B1_c_42_n N_Y_c_216_n 0.0138893f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_55 N_B1_c_43_n N_Y_c_221_n 0.0107468f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 B1 N_Y_c_221_n 0.0124152f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_B1_c_40_n N_Y_c_223_n 0.0049099f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 B1 N_Y_c_223_n 0.0875823f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_59 N_B1_c_43_n N_Y_c_225_n 0.00203769f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 B1 N_A_27_47#_M1005_s 0.00545782f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_61 N_B1_c_40_n N_A_27_47#_c_255_n 0.0103292f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_62 B1 N_A_27_47#_c_255_n 0.0168836f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_63 N_B1_c_42_n N_A_27_47#_c_255_n 0.00335784f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_64 N_B1_c_40_n N_VGND_c_303_n 0.00366111f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_65 N_B1_c_40_n N_VGND_c_306_n 0.00655441f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_66 N_B2_c_72_n N_A2_c_108_n 0.0162293f $X=1.065 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_67 N_B2_c_73_n N_A2_c_109_n 0.0364542f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_68 N_B2_c_74_n N_A2_c_109_n 0.00568876f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_69 N_B2_c_73_n N_A2_c_110_n 6.14849e-19 $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B2_c_74_n N_A2_c_110_n 0.0120307f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_71 N_B2_c_74_n N_A2_c_111_n 0.00808297f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_72 N_B2_c_74_n N_A2_c_114_n 0.00690015f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_73 N_B2_c_73_n N_VPWR_c_183_n 0.00494183f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_74 N_B2_c_73_n N_VPWR_c_178_n 0.00757232f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_75 N_B2_c_74_n N_Y_M1007_d 0.00375042f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_76 N_B2_c_72_n N_Y_c_216_n 0.00700731f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_77 N_B2_c_73_n N_Y_c_216_n 0.00597983f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B2_c_74_n N_Y_c_216_n 0.0377172f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_79 N_B2_c_73_n N_Y_c_230_n 0.0129831f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B2_c_74_n N_Y_c_230_n 0.00609922f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_81 N_B2_c_72_n N_Y_c_223_n 0.0021173f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_82 N_B2_c_73_n N_Y_c_225_n 0.0244362f $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B2_c_74_n N_Y_c_225_n 0.0141494f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B2_c_72_n N_A_27_47#_c_255_n 0.0148335f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B2_c_73_n N_A_27_47#_c_255_n 6.23237e-19 $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B2_c_74_n N_A_27_47#_c_255_n 0.00670874f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B2_c_72_n N_A_27_47#_c_265_n 0.00724849f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B2_c_73_n N_A_27_47#_c_265_n 2.69856e-19 $X=1.09 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B2_c_74_n N_A_27_47#_c_265_n 0.00516312f $X=1.14 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B2_c_72_n N_VGND_c_303_n 0.00366111f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B2_c_72_n N_VGND_c_306_n 0.0061708f $X=1.065 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A2_c_108_n N_A1_c_153_n 0.0236799f $X=1.755 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_A2_c_109_n N_A1_c_154_n 0.0926683f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A2_c_110_n N_A1_c_154_n 0.00101971f $X=1.865 $Y=1.245 $X2=0 $Y2=0
cc_95 N_A2_c_111_n N_A1_c_154_n 0.00387989f $X=1.865 $Y=1.445 $X2=0 $Y2=0
cc_96 N_A2_c_114_n N_A1_c_154_n 0.00452382f $X=2.045 $Y=1.615 $X2=0 $Y2=0
cc_97 A2 N_A1_c_154_n 0.0153131f $X=1.92 $Y=1.785 $X2=0 $Y2=0
cc_98 N_A2_c_109_n A1 2.17669e-19 $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A2_c_110_n A1 0.0141102f $X=1.865 $Y=1.245 $X2=0 $Y2=0
cc_100 N_A2_c_111_n A1 0.0023167f $X=1.865 $Y=1.445 $X2=0 $Y2=0
cc_101 N_A2_c_114_n A1 0.00137277f $X=2.045 $Y=1.615 $X2=0 $Y2=0
cc_102 N_A2_c_114_n N_VPWR_c_182_n 0.00743016f $X=2.045 $Y=1.615 $X2=0 $Y2=0
cc_103 N_A2_c_109_n N_VPWR_c_183_n 0.00702461f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_104 A2 N_VPWR_c_183_n 0.00977827f $X=1.92 $Y=1.785 $X2=0 $Y2=0
cc_105 N_A2_c_109_n N_VPWR_c_178_n 0.0131878f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_106 A2 N_VPWR_c_178_n 0.00917077f $X=1.92 $Y=1.785 $X2=0 $Y2=0
cc_107 N_A2_c_109_n N_Y_c_225_n 0.00966705f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A2_c_110_n N_Y_c_225_n 0.00354355f $X=1.865 $Y=1.245 $X2=0 $Y2=0
cc_109 N_A2_c_114_n A_384_297# 3.43001e-19 $X=2.045 $Y=1.615 $X2=-0.19 $Y2=-0.24
cc_110 A2 A_384_297# 0.00162195f $X=1.92 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_111 N_A2_c_108_n N_A_27_47#_c_268_n 0.00234488f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A2_c_108_n N_A_27_47#_c_265_n 0.00350665f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_109_n N_A_27_47#_c_265_n 2.49489e-19 $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A2_c_110_n N_A_27_47#_c_265_n 0.00380802f $X=1.865 $Y=1.245 $X2=0 $Y2=0
cc_115 N_A2_c_108_n N_A_27_47#_c_256_n 0.0131095f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A2_c_109_n N_A_27_47#_c_256_n 0.00261799f $X=1.83 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A2_c_110_n N_A_27_47#_c_256_n 0.0176769f $X=1.865 $Y=1.245 $X2=0 $Y2=0
cc_118 N_A2_c_114_n N_A_27_47#_c_256_n 0.00434787f $X=2.045 $Y=1.615 $X2=0 $Y2=0
cc_119 N_A2_c_108_n N_A_27_47#_c_257_n 5.31342e-19 $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A2_c_108_n N_VGND_c_302_n 0.00477457f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_121 N_A2_c_108_n N_VGND_c_303_n 0.00433717f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A2_c_108_n N_VGND_c_306_n 0.00658113f $X=1.755 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A1_c_154_n N_VPWR_c_182_n 0.0113255f $X=2.24 $Y=1.41 $X2=0 $Y2=0
cc_124 A1 N_VPWR_c_182_n 0.0251868f $X=2.43 $Y=1.105 $X2=0 $Y2=0
cc_125 N_A1_c_154_n N_VPWR_c_183_n 0.00675169f $X=2.24 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A1_c_154_n N_VPWR_c_178_n 0.0125655f $X=2.24 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A1_c_153_n N_A_27_47#_c_256_n 0.0100006f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A1_c_154_n N_A_27_47#_c_256_n 0.00695008f $X=2.24 $Y=1.41 $X2=0 $Y2=0
cc_129 A1 N_A_27_47#_c_256_n 0.0312585f $X=2.43 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A1_c_153_n N_A_27_47#_c_257_n 0.00603703f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A1_c_153_n N_VGND_c_302_n 0.00418719f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A1_c_153_n N_VGND_c_305_n 0.00425752f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A1_c_153_n N_VGND_c_306_n 0.00692541f $X=2.215 $Y=0.995 $X2=0 $Y2=0
cc_134 N_VPWR_c_178_n A_117_297# 0.00509442f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_135 N_VPWR_c_178_n N_Y_M1007_d 0.00664802f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_136 N_VPWR_c_183_n N_Y_c_230_n 0.0049551f $X=2.34 $Y=2.72 $X2=0 $Y2=0
cc_137 N_VPWR_c_178_n N_Y_c_230_n 0.00876066f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_138 N_VPWR_c_183_n N_Y_c_221_n 0.00459378f $X=2.34 $Y=2.72 $X2=0 $Y2=0
cc_139 N_VPWR_c_178_n N_Y_c_221_n 0.00814258f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_140 N_VPWR_c_183_n N_Y_c_225_n 0.036253f $X=2.34 $Y=2.72 $X2=0 $Y2=0
cc_141 N_VPWR_c_178_n N_Y_c_225_n 0.0208382f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_142 N_VPWR_c_178_n A_384_297# 0.00187687f $X=2.53 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_143 A_117_297# N_Y_c_216_n 0.00440527f $X=0.585 $Y=1.485 $X2=0.24 $Y2=2.34
cc_144 A_117_297# N_Y_c_230_n 0.00907655f $X=0.585 $Y=1.485 $X2=0.26 $Y2=2.34
cc_145 A_117_297# N_Y_c_221_n 0.00310243f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_146 N_Y_M1005_d N_A_27_47#_c_255_n 0.00730016f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_147 N_Y_c_223_n N_A_27_47#_c_255_n 0.0250764f $X=0.73 $Y=0.73 $X2=0 $Y2=0
cc_148 N_Y_c_216_n N_A_27_47#_c_265_n 0.0011777f $X=0.642 $Y=1.835 $X2=0 $Y2=0
cc_149 N_Y_c_223_n N_A_27_47#_c_265_n 0.00817314f $X=0.73 $Y=0.73 $X2=0 $Y2=0
cc_150 N_Y_M1005_d N_VGND_c_306_n 0.00320739f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_256_n N_VGND_M1000_d 0.00509943f $X=2.27 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_152 N_A_27_47#_c_268_n N_VGND_c_302_n 0.0103958f $X=1.455 $Y=0.475 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_265_n N_VGND_c_302_n 0.00268853f $X=1.455 $Y=0.695 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_256_n N_VGND_c_302_n 0.0130459f $X=2.27 $Y=0.78 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_257_n N_VGND_c_302_n 0.0155727f $X=2.485 $Y=0.39 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_255_n N_VGND_c_303_n 0.0556024f $X=1.29 $Y=0.385 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_268_n N_VGND_c_303_n 0.018167f $X=1.455 $Y=0.475 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_256_n N_VGND_c_303_n 0.00316092f $X=2.27 $Y=0.78 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_256_n N_VGND_c_305_n 0.00267473f $X=2.27 $Y=0.78 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_257_n N_VGND_c_305_n 0.0215962f $X=2.485 $Y=0.39 $X2=0 $Y2=0
cc_161 N_A_27_47#_M1005_s N_VGND_c_306_n 0.00253093f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_M1003_d N_VGND_c_306_n 0.00468006f $X=1.14 $Y=0.235 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_M1006_d N_VGND_c_306_n 0.0025987f $X=2.29 $Y=0.235 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_255_n N_VGND_c_306_n 0.0423816f $X=1.29 $Y=0.385 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_268_n N_VGND_c_306_n 0.0123794f $X=1.455 $Y=0.475 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_256_n N_VGND_c_306_n 0.0122354f $X=2.27 $Y=0.78 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_257_n N_VGND_c_306_n 0.0145395f $X=2.485 $Y=0.39 $X2=0 $Y2=0
