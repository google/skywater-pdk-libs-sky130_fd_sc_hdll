* NGSPICE file created from sky130_fd_sc_hdll__a2bb2o_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
M1000 a_525_413# a_243_47# a_79_21# VPB phighvt w=420000u l=180000u
+  ad=2.352e+11p pd=2.8e+06u as=1.134e+11p ps=1.38e+06u
M1001 a_611_47# B2 a_79_21# VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=1.134e+11p ps=1.38e+06u
M1002 a_79_21# a_243_47# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=7.746e+11p ps=6.34e+06u
M1003 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=4.674e+11p pd=4.32e+06u as=2.7e+11p ps=2.54e+06u
M1004 a_241_297# A1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.029e+11p pd=1.33e+06u as=0p ps=0u
M1005 a_525_413# B1 VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND A2_N a_243_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1007 VGND B1 a_611_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_243_47# A1_N VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_243_47# A2_N a_241_297# VPB phighvt w=420000u l=180000u
+  ad=1.155e+11p pd=1.39e+06u as=0p ps=0u
M1010 VPWR B2 a_525_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
.ends

