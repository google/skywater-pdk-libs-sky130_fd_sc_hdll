* File: sky130_fd_sc_hdll__sdfstp_1.pxi.spice
* Created: Wed Sep  2 08:51:42 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCD N_SCD_c_263_n N_SCD_c_267_n N_SCD_c_268_n
+ N_SCD_M1008_g N_SCD_c_264_n N_SCD_M1022_g SCD SCD
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCD
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCE N_SCE_M1030_g N_SCE_c_303_n N_SCE_c_304_n
+ N_SCE_M1033_g N_SCE_c_305_n N_SCE_c_306_n N_SCE_M1012_g N_SCE_M1005_g
+ N_SCE_c_298_n N_SCE_c_318_n N_SCE_c_343_p SCE N_SCE_c_299_n N_SCE_c_300_n
+ N_SCE_c_301_n N_SCE_c_302_n SCE PM_SKY130_FD_SC_HDLL__SDFSTP_1%SCE
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%D N_D_c_406_n N_D_c_411_n N_D_M1036_g
+ N_D_M1029_g D D N_D_c_408_n N_D_c_409_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%D
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_349_21# N_A_349_21#_M1005_s
+ N_A_349_21#_M1012_s N_A_349_21#_M1001_g N_A_349_21#_c_461_n
+ N_A_349_21#_c_462_n N_A_349_21#_M1021_g N_A_349_21#_c_456_n
+ N_A_349_21#_c_457_n N_A_349_21#_c_458_n N_A_349_21#_c_459_n
+ N_A_349_21#_c_460_n N_A_349_21#_c_466_n N_A_349_21#_c_467_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_349_21#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%CLK N_CLK_M1039_g N_CLK_c_534_n N_CLK_M1017_g
+ N_CLK_c_535_n N_CLK_c_539_n N_CLK_c_540_n CLK N_CLK_c_536_n N_CLK_c_537_n
+ N_CLK_c_538_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%CLK
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_693_369# N_A_693_369#_M1017_s
+ N_A_693_369#_M1039_s N_A_693_369#_c_609_n N_A_693_369#_c_610_n
+ N_A_693_369#_M1025_g N_A_693_369#_c_592_n N_A_693_369#_M1015_g
+ N_A_693_369#_c_593_n N_A_693_369#_c_594_n N_A_693_369#_M1026_g
+ N_A_693_369#_c_611_n N_A_693_369#_M1037_g N_A_693_369#_c_612_n
+ N_A_693_369#_c_613_n N_A_693_369#_M1013_g N_A_693_369#_M1003_g
+ N_A_693_369#_c_596_n N_A_693_369#_c_625_n N_A_693_369#_c_597_n
+ N_A_693_369#_c_614_n N_A_693_369#_c_615_n N_A_693_369#_c_598_n
+ N_A_693_369#_c_599_n N_A_693_369#_c_690_p N_A_693_369#_c_600_n
+ N_A_693_369#_c_601_n N_A_693_369#_c_602_n N_A_693_369#_c_603_n
+ N_A_693_369#_c_604_n N_A_693_369#_c_605_n N_A_693_369#_c_606_n
+ N_A_693_369#_c_607_n N_A_693_369#_c_681_p N_A_693_369#_c_620_n
+ N_A_693_369#_c_621_n N_A_693_369#_c_622_n N_A_693_369#_c_623_n
+ N_A_693_369#_c_714_p N_A_693_369#_c_608_n N_A_693_369#_c_624_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_693_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_877_369# N_A_877_369#_M1015_d
+ N_A_877_369#_M1025_d N_A_877_369#_c_892_n N_A_877_369#_c_881_n
+ N_A_877_369#_c_893_n N_A_877_369#_c_894_n N_A_877_369#_c_895_n
+ N_A_877_369#_M1006_g N_A_877_369#_M1023_g N_A_877_369#_M1007_g
+ N_A_877_369#_c_897_n N_A_877_369#_M1010_g N_A_877_369#_c_884_n
+ N_A_877_369#_c_898_n N_A_877_369#_c_899_n N_A_877_369#_c_885_n
+ N_A_877_369#_c_886_n N_A_877_369#_c_887_n N_A_877_369#_c_888_n
+ N_A_877_369#_c_889_n N_A_877_369#_c_890_n N_A_877_369#_c_891_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_877_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1229_21# N_A_1229_21#_M1020_s
+ N_A_1229_21#_M1009_d N_A_1229_21#_M1016_g N_A_1229_21#_c_1066_n
+ N_A_1229_21#_c_1072_n N_A_1229_21#_M1038_g N_A_1229_21#_c_1073_n
+ N_A_1229_21#_c_1067_n N_A_1229_21#_c_1074_n N_A_1229_21#_c_1075_n
+ N_A_1229_21#_c_1068_n N_A_1229_21#_c_1128_p N_A_1229_21#_c_1069_n
+ N_A_1229_21#_c_1070_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1229_21#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1075_413# N_A_1075_413#_M1026_d
+ N_A_1075_413#_M1006_d N_A_1075_413#_c_1160_n N_A_1075_413#_c_1172_n
+ N_A_1075_413#_c_1173_n N_A_1075_413#_M1009_g N_A_1075_413#_c_1161_n
+ N_A_1075_413#_M1020_g N_A_1075_413#_c_1174_n N_A_1075_413#_c_1175_n
+ N_A_1075_413#_M1028_g N_A_1075_413#_M1018_g N_A_1075_413#_c_1162_n
+ N_A_1075_413#_c_1190_n N_A_1075_413#_c_1163_n N_A_1075_413#_c_1176_n
+ N_A_1075_413#_c_1164_n N_A_1075_413#_c_1165_n N_A_1075_413#_c_1166_n
+ N_A_1075_413#_c_1167_n N_A_1075_413#_c_1168_n N_A_1075_413#_c_1169_n
+ N_A_1075_413#_c_1170_n N_A_1075_413#_c_1171_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1075_413#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%SET_B N_SET_B_c_1317_n N_SET_B_M1000_g
+ N_SET_B_M1024_g N_SET_B_c_1319_n N_SET_B_M1011_g N_SET_B_M1031_g
+ N_SET_B_c_1321_n N_SET_B_c_1322_n N_SET_B_c_1323_n N_SET_B_c_1324_n
+ N_SET_B_c_1325_n N_SET_B_c_1326_n N_SET_B_c_1327_n SET_B N_SET_B_c_1328_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%SET_B
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1921_295# N_A_1921_295#_M1034_d
+ N_A_1921_295#_M1014_d N_A_1921_295#_c_1456_n N_A_1921_295#_c_1457_n
+ N_A_1921_295#_M1019_g N_A_1921_295#_c_1458_n N_A_1921_295#_c_1459_n
+ N_A_1921_295#_M1027_g N_A_1921_295#_c_1449_n N_A_1921_295#_c_1450_n
+ N_A_1921_295#_c_1451_n N_A_1921_295#_c_1452_n N_A_1921_295#_c_1462_n
+ N_A_1921_295#_c_1463_n N_A_1921_295#_c_1453_n N_A_1921_295#_c_1454_n
+ N_A_1921_295#_c_1455_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1921_295#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1725_329# N_A_1725_329#_M1007_d
+ N_A_1725_329#_M1013_d N_A_1725_329#_M1011_d N_A_1725_329#_M1034_g
+ N_A_1725_329#_c_1552_n N_A_1725_329#_M1014_g N_A_1725_329#_c_1553_n
+ N_A_1725_329#_M1032_g N_A_1725_329#_c_1564_n N_A_1725_329#_M1004_g
+ N_A_1725_329#_c_1555_n N_A_1725_329#_c_1556_n N_A_1725_329#_c_1557_n
+ N_A_1725_329#_c_1566_n N_A_1725_329#_c_1574_n N_A_1725_329#_c_1575_n
+ N_A_1725_329#_c_1567_n N_A_1725_329#_c_1665_p N_A_1725_329#_c_1558_n
+ N_A_1725_329#_c_1568_n N_A_1725_329#_c_1559_n N_A_1725_329#_c_1560_n
+ N_A_1725_329#_c_1561_n N_A_1725_329#_c_1569_n N_A_1725_329#_c_1608_n
+ N_A_1725_329#_c_1570_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_1725_329#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_2381_47# N_A_2381_47#_M1032_s
+ N_A_2381_47#_M1004_s N_A_2381_47#_c_1707_n N_A_2381_47#_M1035_g
+ N_A_2381_47#_c_1708_n N_A_2381_47#_M1002_g N_A_2381_47#_c_1709_n
+ N_A_2381_47#_c_1713_n N_A_2381_47#_c_1710_n N_A_2381_47#_c_1711_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_2381_47#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_27_369# N_A_27_369#_M1008_s
+ N_A_27_369#_M1021_d N_A_27_369#_c_1757_n N_A_27_369#_c_1758_n
+ N_A_27_369#_c_1759_n N_A_27_369#_c_1774_n N_A_27_369#_c_1771_n
+ N_A_27_369#_c_1760_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_27_369#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%VPWR N_VPWR_M1008_d N_VPWR_M1012_d
+ N_VPWR_M1039_d N_VPWR_M1038_d N_VPWR_M1000_d N_VPWR_M1019_d N_VPWR_M1014_s
+ N_VPWR_M1004_d N_VPWR_c_1804_n N_VPWR_c_1805_n N_VPWR_c_1806_n N_VPWR_c_1807_n
+ N_VPWR_c_1808_n N_VPWR_c_1809_n N_VPWR_c_1810_n N_VPWR_c_1811_n
+ N_VPWR_c_1812_n N_VPWR_c_1813_n VPWR N_VPWR_c_1814_n N_VPWR_c_1815_n
+ N_VPWR_c_1816_n N_VPWR_c_1817_n N_VPWR_c_1818_n N_VPWR_c_1803_n
+ N_VPWR_c_1820_n N_VPWR_c_1821_n N_VPWR_c_1822_n N_VPWR_c_1823_n
+ N_VPWR_c_1824_n N_VPWR_c_1825_n N_VPWR_c_1826_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_201_47# N_A_201_47#_M1030_d
+ N_A_201_47#_M1026_s N_A_201_47#_M1036_d N_A_201_47#_M1006_s
+ N_A_201_47#_c_2006_n N_A_201_47#_c_1995_n N_A_201_47#_c_1999_n
+ N_A_201_47#_c_2000_n N_A_201_47#_c_2009_n N_A_201_47#_c_1996_n
+ N_A_201_47#_c_2001_n N_A_201_47#_c_2002_n N_A_201_47#_c_1997_n
+ N_A_201_47#_c_2004_n N_A_201_47#_c_1998_n
+ PM_SKY130_FD_SC_HDLL__SDFSTP_1%A_201_47#
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%Q N_Q_M1002_d N_Q_M1035_d Q Q Q Q Q Q
+ N_Q_c_2130_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%Q
x_PM_SKY130_FD_SC_HDLL__SDFSTP_1%VGND N_VGND_M1022_s N_VGND_M1001_d
+ N_VGND_M1005_d N_VGND_M1017_d N_VGND_M1016_d N_VGND_M1024_d N_VGND_M1031_d
+ N_VGND_M1032_d N_VGND_c_2141_n N_VGND_c_2142_n N_VGND_c_2143_n N_VGND_c_2144_n
+ N_VGND_c_2145_n N_VGND_c_2146_n N_VGND_c_2147_n N_VGND_c_2148_n
+ N_VGND_c_2149_n N_VGND_c_2150_n N_VGND_c_2151_n N_VGND_c_2152_n
+ N_VGND_c_2153_n N_VGND_c_2154_n VGND N_VGND_c_2155_n N_VGND_c_2156_n
+ N_VGND_c_2157_n N_VGND_c_2158_n N_VGND_c_2159_n N_VGND_c_2160_n
+ N_VGND_c_2161_n PM_SKY130_FD_SC_HDLL__SDFSTP_1%VGND
cc_1 VNB N_SCD_c_263_n 0.0614876f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.325
cc_2 VNB N_SCD_c_264_n 0.017667f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_3 VNB SCD 0.0208496f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_SCE_M1030_g 0.0333651f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.77
cc_5 VNB N_SCE_M1005_g 0.0386452f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_6 VNB N_SCE_c_298_n 0.00641659f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_7 VNB N_SCE_c_299_n 0.0221836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_300_n 0.0327362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_301_n 0.00121258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_302_n 0.0063767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_c_406_n 0.00973242f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.62
cc_12 VNB D 0.00603948f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_13 VNB N_D_c_408_n 0.0284342f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_14 VNB N_D_c_409_n 0.0169241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_349_21#_M1001_g 0.030387f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_16 VNB N_A_349_21#_c_456_n 0.013066f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_17 VNB N_A_349_21#_c_457_n 0.00449025f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_349_21#_c_458_n 0.0322814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_349_21#_c_459_n 0.0144986f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_20 VNB N_A_349_21#_c_460_n 0.00694339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_CLK_c_534_n 0.0175885f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_22 VNB N_CLK_c_535_n 0.0179572f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_23 VNB N_CLK_c_536_n 0.0169771f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_24 VNB N_CLK_c_537_n 0.016278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_CLK_c_538_n 0.0139632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_693_369#_c_592_n 0.0177594f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_27 VNB N_A_693_369#_c_593_n 0.0561083f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_28 VNB N_A_693_369#_c_594_n 0.0178231f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_29 VNB N_A_693_369#_M1003_g 0.0241359f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_693_369#_c_596_n 0.0083546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_693_369#_c_597_n 0.00135304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_693_369#_c_598_n 0.00796372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_693_369#_c_599_n 0.0036336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_693_369#_c_600_n 0.00345628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_693_369#_c_601_n 0.0175281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_693_369#_c_602_n 0.00364477f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_693_369#_c_603_n 0.0267582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_693_369#_c_604_n 0.0103737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_693_369#_c_605_n 3.65794e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_693_369#_c_606_n 0.00452671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_693_369#_c_607_n 0.0280277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_693_369#_c_608_n 0.012173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_877_369#_c_881_n 0.0497739f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_44 VNB N_A_877_369#_M1023_g 0.0325688f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_45 VNB N_A_877_369#_M1007_g 0.0372799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_877_369#_c_884_n 0.00471247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_877_369#_c_885_n 0.020596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_877_369#_c_886_n 0.00121103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_877_369#_c_887_n 0.00458377f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_877_369#_c_888_n 0.00286083f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_877_369#_c_889_n 0.00332697f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_877_369#_c_890_n 0.00274772f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_877_369#_c_891_n 0.017185f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1229_21#_M1016_g 0.0191216f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.695
cc_55 VNB N_A_1229_21#_c_1066_n 0.0139193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1229_21#_c_1067_n 0.0078726f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1229_21#_c_1068_n 0.00452229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1229_21#_c_1069_n 0.0031057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1229_21#_c_1070_n 0.028204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_A_1075_413#_c_1160_n 0.0136329f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_61 VNB N_A_1075_413#_c_1161_n 0.0159786f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=1.445
cc_62 VNB N_A_1075_413#_c_1162_n 0.026685f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1075_413#_c_1163_n 0.0097997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1075_413#_c_1164_n 0.00369281f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1075_413#_c_1165_n 0.00204312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1075_413#_c_1166_n 0.00232092f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1075_413#_c_1167_n 0.0043999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1075_413#_c_1168_n 0.0193407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1075_413#_c_1169_n 0.0126327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_A_1075_413#_c_1170_n 0.0207684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_A_1075_413#_c_1171_n 0.0196198f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_SET_B_M1024_g 0.0424006f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_73 VNB N_SET_B_M1031_g 0.0428059f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_74 VNB N_A_1921_295#_M1027_g 0.0217251f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_1921_295#_c_1449_n 0.0070995f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_76 VNB N_A_1921_295#_c_1450_n 0.00169818f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_1921_295#_c_1451_n 0.0298569f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_78 VNB N_A_1921_295#_c_1452_n 0.00925103f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1921_295#_c_1453_n 0.0121382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1921_295#_c_1454_n 0.00332436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_A_1921_295#_c_1455_n 5.01057e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_1725_329#_c_1552_n 0.00678593f $X=-0.19 $Y=-0.24 $X2=0.145
+ $Y2=0.765
cc_83 VNB N_A_1725_329#_c_1553_n 0.0314804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1725_329#_M1032_g 0.0460153f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_85 VNB N_A_1725_329#_c_1555_n 0.0168625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1725_329#_c_1556_n 0.0209563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1725_329#_c_1557_n 0.00260706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1725_329#_c_1558_n 0.00137968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1725_329#_c_1559_n 0.00218903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1725_329#_c_1560_n 0.00924423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1725_329#_c_1561_n 0.0213379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2381_47#_c_1707_n 0.0298935f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_93 VNB N_A_2381_47#_c_1708_n 0.0206947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_2381_47#_c_1709_n 0.0122539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2381_47#_c_1710_n 0.00291179f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=1.16
cc_96 VNB N_A_2381_47#_c_1711_n 0.00378233f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VPWR_c_1803_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_201_47#_c_1995_n 0.00432851f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_99 VNB N_A_201_47#_c_1996_n 0.00130739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_201_47#_c_1997_n 0.00392628f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_201_47#_c_1998_n 0.00439899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_Q_c_2130_n 0.0487456f $X=-0.19 $Y=-0.24 $X2=0.212 $Y2=0.85
cc_103 VNB N_VGND_c_2141_n 0.0312931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_2142_n 0.0352326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_2143_n 0.00803967f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_2144_n 0.0164899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2145_n 0.00820979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2146_n 0.0027219f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2147_n 0.00518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2148_n 0.00322211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2149_n 0.0146232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2150_n 0.00507625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2151_n 0.0629005f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2152_n 0.00478085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2153_n 0.031469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2154_n 0.0065186f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2155_n 0.0619169f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2156_n 0.0199054f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2157_n 0.624496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2158_n 0.00506925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2159_n 0.00664466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2160_n 0.0167152f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2161_n 0.0187556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VPB N_SCD_c_263_n 0.00540609f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.325
cc_125 VPB N_SCD_c_267_n 0.0175267f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_126 VPB N_SCD_c_268_n 0.0494007f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_127 VPB SCD 0.0148037f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_128 VPB N_SCE_c_303_n 0.0133941f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_129 VPB N_SCE_c_304_n 0.0221672f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_130 VPB N_SCE_c_305_n 0.026286f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_131 VPB N_SCE_c_306_n 0.0343446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_SCE_c_299_n 0.0134821f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_SCE_c_300_n 0.00642596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_SCE_c_301_n 0.00419291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_SCE_c_302_n 0.00484581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_D_c_406_n 0.0161429f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.62
cc_137 VPB N_D_c_411_n 0.0222417f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_138 VPB D 0.0044569f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.695
cc_139 VPB N_A_349_21#_c_461_n 0.0220272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_349_21#_c_462_n 0.0251734f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_141 VPB N_A_349_21#_c_456_n 6.82321e-19 $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_142 VPB N_A_349_21#_c_457_n 0.0101942f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_349_21#_c_458_n 0.0147247f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_349_21#_c_466_n 0.00409949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_349_21#_c_467_n 0.0122482f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_CLK_c_539_n 0.0121836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_CLK_c_540_n 0.040301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_CLK_c_536_n 0.0107275f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_149 VPB N_CLK_c_537_n 0.0204466f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_693_369#_c_609_n 0.0149449f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_151 VPB N_A_693_369#_c_610_n 0.0251151f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.695
cc_152 VPB N_A_693_369#_c_611_n 0.0571336f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_693_369#_c_612_n 0.00776925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_693_369#_c_613_n 0.0206139f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_693_369#_c_614_n 0.0015983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_693_369#_c_615_n 0.00133399f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_693_369#_c_600_n 0.00372107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_693_369#_c_601_n 0.0107422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_693_369#_c_602_n 0.00172895f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_693_369#_c_603_n 0.00317743f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_693_369#_c_620_n 0.00671353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_693_369#_c_621_n 3.87498e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_693_369#_c_622_n 0.00682522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_693_369#_c_623_n 0.0022021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_693_369#_c_624_n 0.00224736f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_877_369#_c_892_n 0.0246271f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_167 VPB N_A_877_369#_c_893_n 0.0201586f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_168 VPB N_A_877_369#_c_894_n 0.0107019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_877_369#_c_895_n 0.0193133f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_170 VPB N_A_877_369#_M1007_g 0.0154403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_877_369#_c_897_n 0.0562401f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.53
cc_172 VPB N_A_877_369#_c_898_n 0.004892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_877_369#_c_899_n 0.00997068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_877_369#_c_887_n 2.44563e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_877_369#_c_888_n 0.00747903f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_877_369#_c_889_n 0.00122725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_A_877_369#_c_891_n 0.0170356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_A_1229_21#_c_1066_n 0.0183639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_1229_21#_c_1072_n 0.064302f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_180 VPB N_A_1229_21#_c_1073_n 0.00179081f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_181 VPB N_A_1229_21#_c_1074_n 0.00606886f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.16
cc_182 VPB N_A_1229_21#_c_1075_n 7.95296e-19 $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_183 VPB N_A_1075_413#_c_1172_n 0.0313223f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_1075_413#_c_1173_n 0.0242898f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_185 VPB N_A_1075_413#_c_1174_n 0.00830856f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_186 VPB N_A_1075_413#_c_1175_n 0.0205109f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_187 VPB N_A_1075_413#_c_1176_n 0.0165451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1075_413#_c_1164_n 0.00646138f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1075_413#_c_1165_n 0.0035338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_A_1075_413#_c_1166_n 0.00131078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_A_1075_413#_c_1167_n 0.00164703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_A_1075_413#_c_1168_n 0.00291439f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_A_1075_413#_c_1170_n 0.00993351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_SET_B_c_1317_n 0.061939f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.325
cc_195 VPB N_SET_B_M1024_g 0.0116708f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_196 VPB N_SET_B_c_1319_n 0.0496045f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_197 VPB N_SET_B_M1031_g 0.00817628f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_198 VPB N_SET_B_c_1321_n 0.0108242f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_199 VPB N_SET_B_c_1322_n 0.00791097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_SET_B_c_1323_n 0.0154598f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_201 VPB N_SET_B_c_1324_n 0.0129672f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_SET_B_c_1325_n 0.00253952f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_SET_B_c_1326_n 0.00590741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_SET_B_c_1327_n 0.00437155f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_SET_B_c_1328_n 0.00959939f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_A_1921_295#_c_1456_n 0.0164597f $X=-0.19 $Y=1.305 $X2=0.52
+ $Y2=0.445
cc_207 VPB N_A_1921_295#_c_1457_n 0.0232178f $X=-0.19 $Y=1.305 $X2=0.315
+ $Y2=1.695
cc_208 VPB N_A_1921_295#_c_1458_n 0.0251076f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_A_1921_295#_c_1459_n 0.00834964f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_210 VPB N_A_1921_295#_c_1449_n 0.0118186f $X=-0.19 $Y=1.305 $X2=0.255
+ $Y2=1.16
cc_211 VPB N_A_1921_295#_c_1452_n 0.00658197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_A_1921_295#_c_1462_n 6.86822e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_A_1921_295#_c_1463_n 0.0187809f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_1725_329#_c_1552_n 0.0887952f $X=-0.19 $Y=1.305 $X2=0.145
+ $Y2=0.765
cc_215 VPB N_A_1725_329#_c_1553_n 0.0248059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_A_1725_329#_c_1564_n 0.0390343f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.53
cc_217 VPB N_A_1725_329#_c_1557_n 0.00169698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_A_1725_329#_c_1566_n 0.0119844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_A_1725_329#_c_1567_n 0.00614394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1725_329#_c_1568_n 0.00705837f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_A_1725_329#_c_1569_n 0.00256005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_A_1725_329#_c_1570_n 0.00172568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_2381_47#_c_1707_n 0.0330052f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_224 VPB N_A_2381_47#_c_1713_n 0.0109395f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_225 VPB N_A_2381_47#_c_1710_n 0.00451528f $X=-0.19 $Y=1.305 $X2=0.212
+ $Y2=1.16
cc_226 VPB N_A_27_369#_c_1757_n 0.0170416f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_227 VPB N_A_27_369#_c_1758_n 0.00100316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_27_369#_c_1759_n 0.00945761f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_229 VPB N_A_27_369#_c_1760_n 0.00263317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1804_n 0.00252882f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1805_n 0.00907525f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1806_n 0.0164751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1807_n 0.00282938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1808_n 0.0058842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1809_n 0.00520779f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_VPWR_c_1810_n 0.0167909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1811_n 0.005797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1812_n 0.0307067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1813_n 0.00487897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1814_n 0.0143786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1815_n 0.0512333f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1816_n 0.0566134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1817_n 0.0290079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_VPWR_c_1818_n 0.0198767f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_VPWR_c_1803_n 0.0731487f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_VPWR_c_1820_n 0.00464622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_VPWR_c_1821_n 0.00564769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_VPWR_c_1822_n 0.00547148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_VPWR_c_1823_n 0.0133607f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1824_n 0.0240535f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1825_n 0.0176704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1826_n 0.0051304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_A_201_47#_c_1999_n 8.90825e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_A_201_47#_c_2000_n 0.00245242f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=1.16
cc_255 VPB N_A_201_47#_c_2001_n 0.025058f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_A_201_47#_c_2002_n 0.0031429f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_A_201_47#_c_1997_n 0.00330318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_A_201_47#_c_2004_n 0.00776824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_A_201_47#_c_1998_n 0.00386251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_Q_c_2130_n 0.0502012f $X=-0.19 $Y=1.305 $X2=0.212 $Y2=0.85
cc_261 N_SCD_c_263_n N_SCE_M1030_g 0.00227875f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_262 N_SCD_c_264_n N_SCE_M1030_g 0.0377993f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_263 SCD N_SCE_M1030_g 3.82641e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_264 N_SCD_c_267_n N_SCE_c_303_n 0.00212959f $X=0.315 $Y=1.62 $X2=0 $Y2=0
cc_265 N_SCD_c_268_n N_SCE_c_303_n 0.00802922f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_266 SCD N_SCE_c_303_n 3.4065e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_267 N_SCD_c_268_n N_SCE_c_304_n 0.0232945f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_268 SCD N_SCE_c_318_n 0.00144346f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_269 N_SCD_c_263_n N_SCE_c_299_n 0.0152623f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_270 SCD N_SCE_c_299_n 3.22701e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_271 N_SCD_c_263_n N_SCE_c_302_n 0.0100034f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_272 N_SCD_c_268_n N_SCE_c_302_n 0.00381492f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_273 SCD N_SCE_c_302_n 0.0602867f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_274 N_SCD_c_268_n N_A_27_369#_c_1757_n 0.00843386f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_275 N_SCD_c_268_n N_A_27_369#_c_1758_n 0.0153318f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_276 N_SCD_c_263_n N_A_27_369#_c_1759_n 5.05332e-19 $X=0.315 $Y=1.325 $X2=0
+ $Y2=0
cc_277 N_SCD_c_268_n N_A_27_369#_c_1759_n 0.00332576f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_278 SCD N_A_27_369#_c_1759_n 0.0227399f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_279 N_SCD_c_268_n N_VPWR_c_1804_n 0.011563f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_280 N_SCD_c_268_n N_VPWR_c_1814_n 0.00317293f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_281 N_SCD_c_268_n N_VPWR_c_1803_n 0.0048112f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_282 N_SCD_c_264_n N_A_201_47#_c_2006_n 2.9719e-19 $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_283 N_SCD_c_263_n N_VGND_c_2142_n 0.00690102f $X=0.315 $Y=1.325 $X2=0 $Y2=0
cc_284 N_SCD_c_264_n N_VGND_c_2142_n 0.0210021f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_285 SCD N_VGND_c_2142_n 0.0221805f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_286 SCD N_VGND_c_2157_n 9.88088e-19 $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_287 N_SCE_c_299_n N_D_c_406_n 0.0247422f $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_288 N_SCE_c_302_n N_D_c_406_n 4.55957e-19 $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_289 N_SCE_c_303_n N_D_c_411_n 0.016356f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_290 N_SCE_c_304_n N_D_c_411_n 0.0461727f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_291 N_SCE_M1030_g D 0.00355142f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_292 N_SCE_c_303_n D 0.00637589f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_293 N_SCE_c_304_n D 3.91386e-19 $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_294 N_SCE_c_298_n D 0.0313118f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_295 N_SCE_c_318_n D 0.00223888f $X=0.87 $Y=1.19 $X2=0 $Y2=0
cc_296 N_SCE_c_299_n D 0.00430657f $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_297 N_SCE_c_302_n D 0.0690236f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_298 N_SCE_M1030_g N_D_c_408_n 0.0192751f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_299 N_SCE_c_298_n N_D_c_408_n 0.00134139f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_300 N_SCE_c_302_n N_D_c_408_n 2.52791e-19 $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_301 N_SCE_M1030_g N_D_c_409_n 0.0134262f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_302 N_SCE_c_298_n N_A_349_21#_c_456_n 0.00480032f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_303 N_SCE_c_305_n N_A_349_21#_c_457_n 0.00674156f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_304 N_SCE_M1005_g N_A_349_21#_c_457_n 0.0025686f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_305 N_SCE_c_298_n N_A_349_21#_c_457_n 0.0173777f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_306 N_SCE_c_343_p N_A_349_21#_c_457_n 6.89964e-19 $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_307 N_SCE_c_300_n N_A_349_21#_c_457_n 0.00247942f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_308 N_SCE_c_301_n N_A_349_21#_c_457_n 0.0400811f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_309 N_SCE_c_298_n N_A_349_21#_c_458_n 0.0040858f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_310 N_SCE_c_300_n N_A_349_21#_c_458_n 0.0213661f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_311 N_SCE_c_301_n N_A_349_21#_c_458_n 7.19229e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_312 N_SCE_M1005_g N_A_349_21#_c_459_n 0.00827962f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_313 N_SCE_c_298_n N_A_349_21#_c_459_n 0.00905152f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_314 N_SCE_c_343_p N_A_349_21#_c_459_n 0.00104259f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_315 N_SCE_c_300_n N_A_349_21#_c_459_n 0.002964f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_316 N_SCE_c_301_n N_A_349_21#_c_459_n 0.00979853f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_317 N_SCE_M1005_g N_A_349_21#_c_460_n 0.00585491f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_318 N_SCE_c_306_n N_A_349_21#_c_467_n 0.00355437f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_319 N_SCE_c_300_n N_A_349_21#_c_467_n 4.82439e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_320 N_SCE_c_301_n N_A_349_21#_c_467_n 0.0105043f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_321 N_SCE_M1005_g N_CLK_c_535_n 0.00287881f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_322 N_SCE_c_305_n N_CLK_c_536_n 0.00124305f $X=2.835 $Y=1.67 $X2=0 $Y2=0
cc_323 N_SCE_c_300_n N_CLK_c_536_n 0.00331448f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_324 N_SCE_c_301_n N_CLK_c_536_n 3.6692e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_325 N_SCE_c_305_n N_CLK_c_537_n 0.00357902f $X=2.835 $Y=1.67 $X2=0 $Y2=0
cc_326 N_SCE_c_343_p N_CLK_c_537_n 0.00158915f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_327 N_SCE_c_300_n N_CLK_c_537_n 0.0033024f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_328 N_SCE_c_301_n N_CLK_c_537_n 0.0356601f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_329 N_SCE_c_300_n N_CLK_c_538_n 0.00287881f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_330 N_SCE_c_306_n N_A_693_369#_c_625_n 0.00347988f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_331 N_SCE_M1005_g N_A_693_369#_c_597_n 0.00346504f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_332 N_SCE_c_306_n N_A_693_369#_c_615_n 0.00464142f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_333 N_SCE_M1005_g N_A_693_369#_c_599_n 0.00350126f $X=2.89 $Y=0.445 $X2=0
+ $Y2=0
cc_334 N_SCE_c_304_n N_A_27_369#_c_1758_n 0.0148547f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_335 N_SCE_c_298_n N_A_27_369#_c_1758_n 0.00494807f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_336 N_SCE_c_318_n N_A_27_369#_c_1758_n 0.00104089f $X=0.87 $Y=1.19 $X2=0
+ $Y2=0
cc_337 N_SCE_c_299_n N_A_27_369#_c_1758_n 7.84018e-19 $X=0.93 $Y=1.25 $X2=0
+ $Y2=0
cc_338 N_SCE_c_302_n N_A_27_369#_c_1758_n 0.0226263f $X=0.725 $Y=1.19 $X2=0
+ $Y2=0
cc_339 N_SCE_c_304_n N_A_27_369#_c_1771_n 0.00202367f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_340 N_SCE_c_304_n N_VPWR_c_1804_n 0.00296668f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_341 N_SCE_c_306_n N_VPWR_c_1805_n 0.0049892f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_342 N_SCE_c_304_n N_VPWR_c_1815_n 0.0052046f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_343 N_SCE_c_306_n N_VPWR_c_1815_n 0.00702461f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_344 N_SCE_c_304_n N_VPWR_c_1803_n 0.00671789f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_345 N_SCE_c_306_n N_VPWR_c_1803_n 0.0150885f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_346 N_SCE_M1030_g N_A_201_47#_c_2006_n 0.00782662f $X=0.93 $Y=0.445 $X2=0
+ $Y2=0
cc_347 N_SCE_c_298_n N_A_201_47#_c_2006_n 0.0112441f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_348 N_SCE_c_298_n N_A_201_47#_c_2009_n 0.00450485f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_349 N_SCE_c_305_n N_A_201_47#_c_2001_n 0.00811567f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_350 N_SCE_c_298_n N_A_201_47#_c_2001_n 0.0490896f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_351 N_SCE_c_343_p N_A_201_47#_c_2001_n 0.0249445f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_352 N_SCE_c_300_n N_A_201_47#_c_2001_n 4.55029e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_353 N_SCE_c_301_n N_A_201_47#_c_2001_n 0.0213105f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_SCE_c_298_n N_A_201_47#_c_2002_n 0.030535f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_355 N_SCE_c_298_n N_A_201_47#_c_1997_n 0.0185596f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_356 N_SCE_M1030_g N_VGND_c_2141_n 0.00456464f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_357 N_SCE_M1030_g N_VGND_c_2142_n 0.00569751f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_358 N_SCE_c_318_n N_VGND_c_2142_n 7.54179e-19 $X=0.87 $Y=1.19 $X2=0 $Y2=0
cc_359 N_SCE_c_299_n N_VGND_c_2142_n 3.94412e-19 $X=0.93 $Y=1.25 $X2=0 $Y2=0
cc_360 N_SCE_c_302_n N_VGND_c_2142_n 0.0152769f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_361 N_SCE_M1005_g N_VGND_c_2143_n 0.00178988f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_362 N_SCE_c_298_n N_VGND_c_2143_n 0.00127321f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_363 N_SCE_M1005_g N_VGND_c_2144_n 0.00486043f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_364 N_SCE_M1005_g N_VGND_c_2145_n 0.0100904f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_365 N_SCE_c_301_n N_VGND_c_2145_n 2.63385e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_366 N_SCE_M1030_g N_VGND_c_2157_n 0.00734604f $X=0.93 $Y=0.445 $X2=0 $Y2=0
cc_367 N_SCE_M1005_g N_VGND_c_2157_n 0.00965187f $X=2.89 $Y=0.445 $X2=0 $Y2=0
cc_368 N_SCE_c_302_n N_VGND_c_2157_n 0.00570024f $X=0.725 $Y=1.19 $X2=0 $Y2=0
cc_369 D N_A_349_21#_M1001_g 3.18064e-19 $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_370 N_D_c_408_n N_A_349_21#_M1001_g 0.0203756f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_371 N_D_c_409_n N_A_349_21#_M1001_g 0.0310629f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_372 N_D_c_411_n N_A_349_21#_c_461_n 0.0157634f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_373 N_D_c_411_n N_A_349_21#_c_462_n 0.0234679f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_374 N_D_c_406_n N_A_349_21#_c_456_n 0.0157634f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_375 D N_A_349_21#_c_456_n 0.00160886f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_376 N_D_c_411_n N_A_27_369#_c_1758_n 0.00136438f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_377 D N_A_27_369#_c_1758_n 0.0137059f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_378 N_D_c_411_n N_A_27_369#_c_1774_n 0.00431987f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_379 N_D_c_411_n N_A_27_369#_c_1760_n 0.0135654f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_380 D N_A_27_369#_c_1760_n 0.00422562f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_381 N_D_c_411_n N_VPWR_c_1815_n 0.00429453f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_382 N_D_c_411_n N_VPWR_c_1803_n 0.0060009f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_383 D N_A_201_47#_c_2006_n 0.0313325f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_384 N_D_c_408_n N_A_201_47#_c_2006_n 0.00175893f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_385 N_D_c_409_n N_A_201_47#_c_2006_n 0.012197f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_386 N_D_c_411_n N_A_201_47#_c_2009_n 0.00519966f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_387 D N_A_201_47#_c_2009_n 0.00614145f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_388 D N_A_201_47#_c_2002_n 0.00778368f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_389 N_D_c_406_n N_A_201_47#_c_1997_n 0.00161643f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_390 N_D_c_411_n N_A_201_47#_c_1997_n 0.00355157f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_391 D N_A_201_47#_c_1997_n 0.0689424f $X=1.065 $Y=0.765 $X2=0 $Y2=0
cc_392 N_D_c_408_n N_A_201_47#_c_1997_n 0.00193715f $X=1.35 $Y=0.93 $X2=0 $Y2=0
cc_393 N_D_c_409_n N_A_201_47#_c_1997_n 0.00351003f $X=1.375 $Y=0.765 $X2=0
+ $Y2=0
cc_394 N_D_c_409_n N_VGND_c_2141_n 0.00357877f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_395 N_D_c_409_n N_VGND_c_2157_n 0.00539883f $X=1.375 $Y=0.765 $X2=0 $Y2=0
cc_396 N_A_349_21#_c_467_n N_A_27_369#_M1021_d 0.00555261f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_397 N_A_349_21#_c_462_n N_A_27_369#_c_1760_n 0.011002f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_398 N_A_349_21#_c_466_n N_A_27_369#_c_1760_n 0.0148152f $X=2.595 $Y=1.927
+ $X2=0 $Y2=0
cc_399 N_A_349_21#_c_467_n N_A_27_369#_c_1760_n 0.0132953f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_400 N_A_349_21#_c_462_n N_VPWR_c_1815_n 0.00429453f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_401 N_A_349_21#_c_466_n N_VPWR_c_1815_n 0.0157393f $X=2.595 $Y=1.927 $X2=0
+ $Y2=0
cc_402 N_A_349_21#_c_467_n N_VPWR_c_1815_n 0.00432835f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_403 N_A_349_21#_M1012_s N_VPWR_c_1803_n 0.00304306f $X=2.475 $Y=1.845 $X2=0
+ $Y2=0
cc_404 N_A_349_21#_c_462_n N_VPWR_c_1803_n 0.00737353f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_405 N_A_349_21#_c_466_n N_VPWR_c_1803_n 0.00941222f $X=2.595 $Y=1.927 $X2=0
+ $Y2=0
cc_406 N_A_349_21#_c_467_n N_VPWR_c_1803_n 0.00699224f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_407 N_A_349_21#_M1001_g N_A_201_47#_c_2006_n 0.0106694f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_408 N_A_349_21#_c_460_n N_A_201_47#_c_2006_n 0.00154368f $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_409 N_A_349_21#_c_462_n N_A_201_47#_c_2009_n 0.00556528f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_410 N_A_349_21#_c_467_n N_A_201_47#_c_2009_n 0.0164794f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_411 N_A_349_21#_c_457_n N_A_201_47#_c_2001_n 0.0172766f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_412 N_A_349_21#_c_458_n N_A_201_47#_c_2001_n 0.00172463f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_413 N_A_349_21#_c_467_n N_A_201_47#_c_2001_n 0.0111897f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_414 N_A_349_21#_c_461_n N_A_201_47#_c_2002_n 0.00546081f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_415 N_A_349_21#_c_457_n N_A_201_47#_c_2002_n 0.00296292f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_416 N_A_349_21#_M1001_g N_A_201_47#_c_1997_n 0.00973696f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_417 N_A_349_21#_c_461_n N_A_201_47#_c_1997_n 0.0072174f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_418 N_A_349_21#_c_462_n N_A_201_47#_c_1997_n 0.00456775f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_419 N_A_349_21#_c_456_n N_A_201_47#_c_1997_n 0.00911472f $X=1.845 $Y=1.16
+ $X2=0 $Y2=0
cc_420 N_A_349_21#_c_457_n N_A_201_47#_c_1997_n 0.0488018f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_421 N_A_349_21#_c_459_n N_A_201_47#_c_1997_n 0.0125621f $X=2.59 $Y=0.715
+ $X2=0 $Y2=0
cc_422 N_A_349_21#_c_460_n N_A_201_47#_c_1997_n 0.00338006f $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_423 N_A_349_21#_c_467_n N_A_201_47#_c_1997_n 0.00494415f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_424 N_A_349_21#_M1001_g N_VGND_c_2141_n 0.00433573f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_425 N_A_349_21#_M1001_g N_VGND_c_2143_n 0.0105214f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_426 N_A_349_21#_c_458_n N_VGND_c_2143_n 0.00128608f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_427 N_A_349_21#_c_459_n N_VGND_c_2143_n 0.0174596f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_428 N_A_349_21#_c_460_n N_VGND_c_2143_n 0.0233257f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_429 N_A_349_21#_c_459_n N_VGND_c_2144_n 0.00268684f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_430 N_A_349_21#_c_460_n N_VGND_c_2144_n 0.0176923f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_431 N_A_349_21#_c_460_n N_VGND_c_2145_n 0.0190636f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_432 N_A_349_21#_M1005_s N_VGND_c_2157_n 0.00580108f $X=2.505 $Y=0.235 $X2=0
+ $Y2=0
cc_433 N_A_349_21#_M1001_g N_VGND_c_2157_n 0.00851845f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_434 N_A_349_21#_c_459_n N_VGND_c_2157_n 0.00551711f $X=2.59 $Y=0.715 $X2=0
+ $Y2=0
cc_435 N_A_349_21#_c_460_n N_VGND_c_2157_n 0.00983733f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_436 N_CLK_c_539_n N_A_693_369#_c_609_n 0.0059319f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_437 N_CLK_c_540_n N_A_693_369#_c_609_n 0.00655864f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_438 N_CLK_c_537_n N_A_693_369#_c_609_n 3.04599e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_439 N_CLK_c_540_n N_A_693_369#_c_610_n 0.0222028f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_440 N_CLK_c_534_n N_A_693_369#_c_592_n 0.0116086f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_441 N_CLK_c_535_n N_A_693_369#_c_596_n 0.00767961f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_442 N_CLK_c_534_n N_A_693_369#_c_597_n 0.0056285f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_443 N_CLK_c_540_n N_A_693_369#_c_614_n 0.0161161f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_444 N_CLK_c_537_n N_A_693_369#_c_614_n 0.00934927f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_445 N_CLK_c_540_n N_A_693_369#_c_615_n 3.10042e-19 $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_446 N_CLK_c_536_n N_A_693_369#_c_615_n 5.4866e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_447 N_CLK_c_537_n N_A_693_369#_c_615_n 0.0133612f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_448 N_CLK_c_534_n N_A_693_369#_c_598_n 0.00401517f $X=3.88 $Y=0.73 $X2=0
+ $Y2=0
cc_449 N_CLK_c_535_n N_A_693_369#_c_598_n 0.00847863f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_450 N_CLK_c_537_n N_A_693_369#_c_598_n 0.00801255f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_451 N_CLK_c_538_n N_A_693_369#_c_598_n 0.00151794f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_452 N_CLK_c_535_n N_A_693_369#_c_599_n 0.00352145f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_453 N_CLK_c_536_n N_A_693_369#_c_599_n 8.54762e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_454 N_CLK_c_537_n N_A_693_369#_c_599_n 0.016187f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_455 N_CLK_c_538_n N_A_693_369#_c_599_n 5.61645e-19 $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_456 N_CLK_c_540_n N_A_693_369#_c_600_n 0.00461373f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_457 N_CLK_c_537_n N_A_693_369#_c_600_n 0.0379355f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_458 N_CLK_c_538_n N_A_693_369#_c_600_n 0.00572652f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_459 N_CLK_c_536_n N_A_693_369#_c_601_n 0.0164171f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_460 N_CLK_c_537_n N_A_693_369#_c_601_n 3.92042e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_461 N_CLK_c_538_n N_A_693_369#_c_608_n 0.0053784f $X=3.68 $Y=1.09 $X2=0 $Y2=0
cc_462 N_CLK_c_540_n N_VPWR_c_1805_n 0.00397623f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_463 N_CLK_c_537_n N_VPWR_c_1805_n 0.00278244f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_464 N_CLK_c_540_n N_VPWR_c_1806_n 0.00320592f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_465 N_CLK_c_540_n N_VPWR_c_1803_n 0.00524235f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_466 N_CLK_c_540_n N_VPWR_c_1822_n 0.0111353f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_467 N_CLK_c_539_n N_A_201_47#_c_2001_n 0.0011232f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_468 N_CLK_c_540_n N_A_201_47#_c_2001_n 0.00327618f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_469 N_CLK_c_537_n N_A_201_47#_c_2001_n 0.0533918f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_470 N_CLK_c_534_n N_VGND_c_2145_n 0.00207759f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_471 N_CLK_c_537_n N_VGND_c_2145_n 0.00829842f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_472 N_CLK_c_534_n N_VGND_c_2146_n 0.00817351f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_473 N_CLK_c_534_n N_VGND_c_2149_n 0.00348405f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_474 N_CLK_c_535_n N_VGND_c_2149_n 4.55781e-19 $X=3.88 $Y=0.805 $X2=0 $Y2=0
cc_475 N_CLK_c_534_n N_VGND_c_2157_n 0.00552264f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_476 N_A_693_369#_c_620_n N_A_877_369#_M1025_d 7.76593e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_477 N_A_693_369#_c_621_n N_A_877_369#_M1025_d 6.28941e-19 $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_478 N_A_693_369#_c_609_n N_A_877_369#_c_892_n 0.00683981f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_479 N_A_693_369#_c_610_n N_A_877_369#_c_892_n 0.0051976f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_480 N_A_693_369#_c_611_n N_A_877_369#_c_892_n 0.00286715f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_481 N_A_693_369#_c_620_n N_A_877_369#_c_892_n 0.00113464f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_482 N_A_693_369#_c_611_n N_A_877_369#_c_881_n 0.010354f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_483 N_A_693_369#_c_620_n N_A_877_369#_c_881_n 8.44234e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_484 N_A_693_369#_c_624_n N_A_877_369#_c_881_n 2.5741e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_485 N_A_693_369#_c_611_n N_A_877_369#_c_893_n 0.00899979f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_486 N_A_693_369#_c_620_n N_A_877_369#_c_893_n 0.00501369f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_487 N_A_693_369#_c_623_n N_A_877_369#_c_893_n 7.59275e-19 $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_488 N_A_693_369#_c_624_n N_A_877_369#_c_893_n 6.19475e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_489 N_A_693_369#_c_620_n N_A_877_369#_c_894_n 0.00175018f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_490 N_A_693_369#_c_611_n N_A_877_369#_c_895_n 0.0111876f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_491 N_A_693_369#_c_594_n N_A_877_369#_M1023_g 0.0150319f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_492 N_A_693_369#_c_612_n N_A_877_369#_M1007_g 0.00729154f $X=8.535 $Y=1.47
+ $X2=0 $Y2=0
cc_493 N_A_693_369#_c_613_n N_A_877_369#_M1007_g 0.0122389f $X=8.535 $Y=1.57
+ $X2=0 $Y2=0
cc_494 N_A_693_369#_M1003_g N_A_877_369#_M1007_g 0.0173162f $X=9.7 $Y=0.445
+ $X2=0 $Y2=0
cc_495 N_A_693_369#_c_602_n N_A_877_369#_M1007_g 0.00652006f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_496 N_A_693_369#_c_603_n N_A_877_369#_M1007_g 0.0127789f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_497 N_A_693_369#_c_604_n N_A_877_369#_M1007_g 0.0139816f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_498 N_A_693_369#_c_606_n N_A_877_369#_M1007_g 0.00145044f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_499 N_A_693_369#_c_607_n N_A_877_369#_M1007_g 0.0116495f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_500 N_A_693_369#_c_613_n N_A_877_369#_c_897_n 0.013501f $X=8.535 $Y=1.57
+ $X2=0 $Y2=0
cc_501 N_A_693_369#_c_604_n N_A_877_369#_c_897_n 0.00117792f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_502 N_A_693_369#_c_681_p N_A_877_369#_c_897_n 0.00222399f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_503 N_A_693_369#_c_592_n N_A_877_369#_c_884_n 0.00346646f $X=4.35 $Y=0.73
+ $X2=0 $Y2=0
cc_504 N_A_693_369#_c_593_n N_A_877_369#_c_884_n 0.015478f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_505 N_A_693_369#_c_598_n N_A_877_369#_c_884_n 0.0125458f $X=4.035 $Y=0.8
+ $X2=0 $Y2=0
cc_506 N_A_693_369#_c_600_n N_A_877_369#_c_884_n 0.0662039f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_507 N_A_693_369#_c_608_n N_A_877_369#_c_884_n 0.00343131f $X=4.235 $Y=1.09
+ $X2=0 $Y2=0
cc_508 N_A_693_369#_c_620_n N_A_877_369#_c_898_n 9.60456e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_509 N_A_693_369#_c_609_n N_A_877_369#_c_899_n 0.00343131f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_510 N_A_693_369#_c_610_n N_A_877_369#_c_899_n 0.00697298f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_511 N_A_693_369#_c_690_p N_A_877_369#_c_899_n 0.0109474f $X=4.165 $Y=1.83
+ $X2=0 $Y2=0
cc_512 N_A_693_369#_c_620_n N_A_877_369#_c_899_n 0.0215922f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_513 N_A_693_369#_c_621_n N_A_877_369#_c_899_n 0.00302262f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_514 N_A_693_369#_c_593_n N_A_877_369#_c_885_n 0.00209217f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_515 N_A_693_369#_c_602_n N_A_877_369#_c_885_n 0.0263552f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_516 N_A_693_369#_c_603_n N_A_877_369#_c_885_n 0.00288312f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_517 N_A_693_369#_c_604_n N_A_877_369#_c_885_n 0.0067427f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_518 N_A_693_369#_c_620_n N_A_877_369#_c_885_n 0.014567f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_519 N_A_693_369#_c_622_n N_A_877_369#_c_885_n 0.0617634f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_520 N_A_693_369#_c_623_n N_A_877_369#_c_885_n 0.0147711f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_521 N_A_693_369#_c_624_n N_A_877_369#_c_885_n 8.34727e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_522 N_A_693_369#_c_602_n N_A_877_369#_c_886_n 0.00279016f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_523 N_A_693_369#_c_604_n N_A_877_369#_c_886_n 0.00325976f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_524 N_A_693_369#_c_604_n N_A_877_369#_c_887_n 0.00197051f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_525 N_A_693_369#_c_606_n N_A_877_369#_c_887_n 0.00585937f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_526 N_A_693_369#_c_607_n N_A_877_369#_c_887_n 0.00352288f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_527 N_A_693_369#_c_612_n N_A_877_369#_c_888_n 5.81998e-19 $X=8.535 $Y=1.47
+ $X2=0 $Y2=0
cc_528 N_A_693_369#_c_613_n N_A_877_369#_c_888_n 8.63357e-19 $X=8.535 $Y=1.57
+ $X2=0 $Y2=0
cc_529 N_A_693_369#_c_602_n N_A_877_369#_c_888_n 0.0449022f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_530 N_A_693_369#_c_603_n N_A_877_369#_c_888_n 5.88608e-19 $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_531 N_A_693_369#_c_604_n N_A_877_369#_c_888_n 0.021647f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_532 N_A_693_369#_c_606_n N_A_877_369#_c_888_n 0.00862888f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_533 N_A_693_369#_c_607_n N_A_877_369#_c_888_n 0.00114446f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_534 N_A_693_369#_c_681_p N_A_877_369#_c_888_n 0.0198966f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_535 N_A_693_369#_c_714_p N_A_877_369#_c_888_n 6.2334e-19 $X=8.295 $Y=1.87
+ $X2=0 $Y2=0
cc_536 N_A_693_369#_c_593_n N_A_877_369#_c_889_n 0.00266973f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_537 N_A_693_369#_c_601_n N_A_877_369#_c_889_n 0.00343131f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_538 N_A_693_369#_c_593_n N_A_877_369#_c_890_n 0.00247177f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_539 N_A_693_369#_c_600_n N_A_877_369#_c_890_n 0.00125608f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_540 N_A_693_369#_c_593_n N_A_877_369#_c_891_n 0.0528355f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_541 N_A_693_369#_c_600_n N_A_877_369#_c_891_n 2.72753e-19 $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_542 N_A_693_369#_c_601_n N_A_877_369#_c_891_n 0.0186987f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_543 N_A_693_369#_c_611_n N_A_1229_21#_c_1072_n 0.0334006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_544 N_A_693_369#_c_622_n N_A_1229_21#_c_1072_n 0.00848583f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_545 N_A_693_369#_c_622_n N_A_1229_21#_c_1073_n 0.0111901f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_546 N_A_693_369#_c_681_p N_A_1229_21#_c_1074_n 7.41551e-19 $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_547 N_A_693_369#_c_622_n N_A_1229_21#_c_1074_n 0.0287031f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_548 N_A_693_369#_c_622_n N_A_1229_21#_c_1075_n 0.0032337f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_549 N_A_693_369#_c_622_n N_A_1075_413#_c_1172_n 0.0037979f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_550 N_A_693_369#_c_622_n N_A_1075_413#_c_1173_n 7.54942e-19 $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_551 N_A_693_369#_c_612_n N_A_1075_413#_c_1174_n 0.0123892f $X=8.535 $Y=1.47
+ $X2=0 $Y2=0
cc_552 N_A_693_369#_c_613_n N_A_1075_413#_c_1175_n 0.0734532f $X=8.535 $Y=1.57
+ $X2=0 $Y2=0
cc_553 N_A_693_369#_c_602_n N_A_1075_413#_c_1175_n 7.14688e-19 $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_554 N_A_693_369#_c_681_p N_A_1075_413#_c_1175_n 0.0155414f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_555 N_A_693_369#_c_714_p N_A_1075_413#_c_1175_n 0.00128013f $X=8.295 $Y=1.87
+ $X2=0 $Y2=0
cc_556 N_A_693_369#_c_611_n N_A_1075_413#_c_1190_n 0.0154392f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_557 N_A_693_369#_c_620_n N_A_1075_413#_c_1190_n 0.00362812f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_558 N_A_693_369#_c_622_n N_A_1075_413#_c_1190_n 0.00492445f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_559 N_A_693_369#_c_623_n N_A_1075_413#_c_1190_n 0.00557824f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_560 N_A_693_369#_c_624_n N_A_1075_413#_c_1190_n 0.013294f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_561 N_A_693_369#_c_594_n N_A_1075_413#_c_1163_n 0.0028029f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_562 N_A_693_369#_c_611_n N_A_1075_413#_c_1176_n 0.00612006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_563 N_A_693_369#_c_622_n N_A_1075_413#_c_1176_n 0.0144347f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_564 N_A_693_369#_c_623_n N_A_1075_413#_c_1176_n 0.00314702f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_565 N_A_693_369#_c_624_n N_A_1075_413#_c_1176_n 0.0267088f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_566 N_A_693_369#_c_611_n N_A_1075_413#_c_1164_n 0.00266776f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_567 N_A_693_369#_c_620_n N_A_1075_413#_c_1164_n 0.00188086f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_568 N_A_693_369#_c_622_n N_A_1075_413#_c_1164_n 0.00794771f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_569 N_A_693_369#_c_623_n N_A_1075_413#_c_1164_n 0.00277252f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_570 N_A_693_369#_c_624_n N_A_1075_413#_c_1164_n 0.0162857f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_571 N_A_693_369#_c_622_n N_A_1075_413#_c_1165_n 0.00447966f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_572 N_A_693_369#_c_602_n N_A_1075_413#_c_1167_n 0.0271196f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_573 N_A_693_369#_c_603_n N_A_1075_413#_c_1167_n 0.00191634f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_574 N_A_693_369#_c_681_p N_A_1075_413#_c_1167_n 0.00856289f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_575 N_A_693_369#_c_602_n N_A_1075_413#_c_1168_n 0.00228701f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_576 N_A_693_369#_c_603_n N_A_1075_413#_c_1168_n 0.0123892f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_577 N_A_693_369#_c_681_p N_A_1075_413#_c_1168_n 0.00125282f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_578 N_A_693_369#_c_681_p N_A_1075_413#_c_1169_n 4.30034e-19 $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_579 N_A_693_369#_c_622_n N_A_1075_413#_c_1169_n 0.00254971f $X=8.15 $Y=1.87
+ $X2=0 $Y2=0
cc_580 N_A_693_369#_c_602_n N_A_1075_413#_c_1171_n 0.00245369f $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_581 N_A_693_369#_c_605_n N_A_1075_413#_c_1171_n 0.00430471f $X=8.785 $Y=0.812
+ $X2=0 $Y2=0
cc_582 N_A_693_369#_c_681_p N_SET_B_c_1317_n 0.00412673f $X=8.485 $Y=1.812
+ $X2=-0.19 $Y2=-0.24
cc_583 N_A_693_369#_c_622_n N_SET_B_c_1317_n 0.0103971f $X=8.15 $Y=1.87
+ $X2=-0.19 $Y2=-0.24
cc_584 N_A_693_369#_c_612_n N_SET_B_c_1324_n 5.55856e-19 $X=8.535 $Y=1.47 $X2=0
+ $Y2=0
cc_585 N_A_693_369#_c_613_n N_SET_B_c_1324_n 9.40989e-19 $X=8.535 $Y=1.57 $X2=0
+ $Y2=0
cc_586 N_A_693_369#_c_602_n N_SET_B_c_1324_n 0.0244877f $X=8.57 $Y=1.16 $X2=0
+ $Y2=0
cc_587 N_A_693_369#_c_604_n N_SET_B_c_1324_n 0.00607822f $X=9.52 $Y=0.812 $X2=0
+ $Y2=0
cc_588 N_A_693_369#_c_606_n N_SET_B_c_1324_n 0.00133335f $X=9.64 $Y=1.09 $X2=0
+ $Y2=0
cc_589 N_A_693_369#_c_607_n N_SET_B_c_1324_n 3.78285e-19 $X=9.64 $Y=1.09 $X2=0
+ $Y2=0
cc_590 N_A_693_369#_c_681_p N_SET_B_c_1324_n 0.00962309f $X=8.485 $Y=1.812 $X2=0
+ $Y2=0
cc_591 N_A_693_369#_c_622_n N_SET_B_c_1324_n 0.0347133f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_592 N_A_693_369#_c_714_p N_SET_B_c_1324_n 0.0306434f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_593 N_A_693_369#_c_622_n N_SET_B_c_1325_n 0.0304949f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_594 N_A_693_369#_c_606_n N_SET_B_c_1326_n 0.00810822f $X=9.64 $Y=1.09 $X2=0
+ $Y2=0
cc_595 N_A_693_369#_c_606_n N_SET_B_c_1327_n 0.0188656f $X=9.64 $Y=1.09 $X2=0
+ $Y2=0
cc_596 N_A_693_369#_c_607_n N_SET_B_c_1327_n 6.03712e-19 $X=9.64 $Y=1.09 $X2=0
+ $Y2=0
cc_597 N_A_693_369#_c_681_p N_SET_B_c_1328_n 0.00839448f $X=8.485 $Y=1.812 $X2=0
+ $Y2=0
cc_598 N_A_693_369#_c_622_n N_SET_B_c_1328_n 0.0114229f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_599 N_A_693_369#_c_606_n N_A_1921_295#_c_1459_n 6.86421e-19 $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_600 N_A_693_369#_c_607_n N_A_1921_295#_c_1459_n 0.0104898f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_601 N_A_693_369#_M1003_g N_A_1921_295#_M1027_g 0.0363566f $X=9.7 $Y=0.445
+ $X2=0 $Y2=0
cc_602 N_A_693_369#_c_604_n N_A_1921_295#_M1027_g 0.00202447f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_603 N_A_693_369#_M1003_g N_A_1921_295#_c_1450_n 3.42575e-19 $X=9.7 $Y=0.445
+ $X2=0 $Y2=0
cc_604 N_A_693_369#_c_604_n N_A_1921_295#_c_1450_n 0.00387786f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_605 N_A_693_369#_c_606_n N_A_1921_295#_c_1450_n 0.0209776f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_606 N_A_693_369#_c_606_n N_A_1921_295#_c_1451_n 0.00215477f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_607 N_A_693_369#_c_607_n N_A_1921_295#_c_1451_n 0.0363566f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_608 N_A_693_369#_c_606_n N_A_1921_295#_c_1462_n 0.00472209f $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_609 N_A_693_369#_c_604_n N_A_1725_329#_M1007_d 0.00212707f $X=9.52 $Y=0.812
+ $X2=-0.19 $Y2=-0.24
cc_610 N_A_693_369#_c_602_n N_A_1725_329#_M1013_d 2.08924e-19 $X=8.57 $Y=1.16
+ $X2=0 $Y2=0
cc_611 N_A_693_369#_c_681_p N_A_1725_329#_M1013_d 0.00508388f $X=8.485 $Y=1.812
+ $X2=0 $Y2=0
cc_612 N_A_693_369#_c_613_n N_A_1725_329#_c_1574_n 0.00145523f $X=8.535 $Y=1.57
+ $X2=0 $Y2=0
cc_613 N_A_693_369#_M1003_g N_A_1725_329#_c_1575_n 0.0142183f $X=9.7 $Y=0.445
+ $X2=0 $Y2=0
cc_614 N_A_693_369#_c_604_n N_A_1725_329#_c_1575_n 0.0505779f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_615 N_A_693_369#_c_607_n N_A_1725_329#_c_1575_n 4.18621e-19 $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_616 N_A_693_369#_c_604_n N_A_1725_329#_c_1558_n 0.0022632f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_617 N_A_693_369#_c_604_n N_A_1725_329#_c_1559_n 0.0026858f $X=9.52 $Y=0.812
+ $X2=0 $Y2=0
cc_618 N_A_693_369#_c_606_n N_A_1725_329#_c_1569_n 7.3466e-19 $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_619 N_A_693_369#_c_607_n N_A_1725_329#_c_1569_n 3.84956e-19 $X=9.64 $Y=1.09
+ $X2=0 $Y2=0
cc_620 N_A_693_369#_c_614_n N_VPWR_M1039_d 7.92879e-19 $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_621 N_A_693_369#_c_690_p N_VPWR_M1039_d 0.00150754f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_622 N_A_693_369#_c_681_p N_VPWR_M1000_d 0.00600677f $X=8.485 $Y=1.812 $X2=0
+ $Y2=0
cc_623 N_A_693_369#_c_622_n N_VPWR_M1000_d 0.00149961f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_624 N_A_693_369#_c_625_n N_VPWR_c_1805_n 0.0102695f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_625 N_A_693_369#_c_625_n N_VPWR_c_1806_n 0.00603303f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_626 N_A_693_369#_c_614_n N_VPWR_c_1806_n 0.00195426f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_627 N_A_693_369#_c_610_n N_VPWR_c_1816_n 0.0055518f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_628 N_A_693_369#_c_611_n N_VPWR_c_1816_n 0.00429453f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_629 N_A_693_369#_c_690_p N_VPWR_c_1816_n 0.00103674f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_630 N_A_693_369#_M1039_s N_VPWR_c_1803_n 0.00400999f $X=3.465 $Y=1.845 $X2=0
+ $Y2=0
cc_631 N_A_693_369#_c_610_n N_VPWR_c_1803_n 0.00657032f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_632 N_A_693_369#_c_611_n N_VPWR_c_1803_n 0.00620168f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_633 N_A_693_369#_c_613_n N_VPWR_c_1803_n 0.00112675f $X=8.535 $Y=1.57 $X2=0
+ $Y2=0
cc_634 N_A_693_369#_c_625_n N_VPWR_c_1803_n 0.00591039f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_635 N_A_693_369#_c_614_n N_VPWR_c_1803_n 0.004831f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_636 N_A_693_369#_c_690_p N_VPWR_c_1803_n 0.00153627f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_637 N_A_693_369#_c_681_p N_VPWR_c_1803_n 0.00802397f $X=8.485 $Y=1.812 $X2=0
+ $Y2=0
cc_638 N_A_693_369#_c_620_n N_VPWR_c_1803_n 0.0552922f $X=5.545 $Y=1.87 $X2=0
+ $Y2=0
cc_639 N_A_693_369#_c_621_n N_VPWR_c_1803_n 0.0167052f $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_640 N_A_693_369#_c_622_n N_VPWR_c_1803_n 0.103241f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_641 N_A_693_369#_c_623_n N_VPWR_c_1803_n 0.018311f $X=5.885 $Y=1.87 $X2=0
+ $Y2=0
cc_642 N_A_693_369#_c_714_p N_VPWR_c_1803_n 0.0168958f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_643 N_A_693_369#_c_610_n N_VPWR_c_1822_n 0.00815097f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_644 N_A_693_369#_c_625_n N_VPWR_c_1822_n 0.00373276f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_645 N_A_693_369#_c_614_n N_VPWR_c_1822_n 0.00632657f $X=4.035 $Y=1.915 $X2=0
+ $Y2=0
cc_646 N_A_693_369#_c_690_p N_VPWR_c_1822_n 0.00632896f $X=4.165 $Y=1.83 $X2=0
+ $Y2=0
cc_647 N_A_693_369#_c_621_n N_VPWR_c_1822_n 8.52709e-19 $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_648 N_A_693_369#_c_622_n N_VPWR_c_1823_n 0.00139085f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_649 N_A_693_369#_c_613_n N_VPWR_c_1825_n 0.0203001f $X=8.535 $Y=1.57 $X2=0
+ $Y2=0
cc_650 N_A_693_369#_c_681_p N_VPWR_c_1825_n 0.0428021f $X=8.485 $Y=1.812 $X2=0
+ $Y2=0
cc_651 N_A_693_369#_c_622_n N_VPWR_c_1825_n 0.00788962f $X=8.15 $Y=1.87 $X2=0
+ $Y2=0
cc_652 N_A_693_369#_c_714_p N_VPWR_c_1825_n 0.00402866f $X=8.295 $Y=1.87 $X2=0
+ $Y2=0
cc_653 N_A_693_369#_c_594_n N_A_201_47#_c_1995_n 0.00439649f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_654 N_A_693_369#_c_611_n N_A_201_47#_c_2000_n 3.6876e-19 $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_655 N_A_693_369#_c_620_n N_A_201_47#_c_2000_n 0.0162746f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_656 N_A_693_369#_c_623_n N_A_201_47#_c_2000_n 0.00274259f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_657 N_A_693_369#_c_593_n N_A_201_47#_c_1996_n 0.0110036f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_658 N_A_693_369#_c_609_n N_A_201_47#_c_2001_n 0.00641873f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_659 N_A_693_369#_c_596_n N_A_201_47#_c_2001_n 0.00176142f $X=4.317 $Y=0.805
+ $X2=0 $Y2=0
cc_660 N_A_693_369#_c_614_n N_A_201_47#_c_2001_n 0.0099266f $X=4.035 $Y=1.915
+ $X2=0 $Y2=0
cc_661 N_A_693_369#_c_615_n N_A_201_47#_c_2001_n 0.00126159f $X=3.675 $Y=1.915
+ $X2=0 $Y2=0
cc_662 N_A_693_369#_c_598_n N_A_201_47#_c_2001_n 0.00714535f $X=4.035 $Y=0.8
+ $X2=0 $Y2=0
cc_663 N_A_693_369#_c_599_n N_A_201_47#_c_2001_n 7.07979e-19 $X=3.705 $Y=0.8
+ $X2=0 $Y2=0
cc_664 N_A_693_369#_c_600_n N_A_201_47#_c_2001_n 0.0221679f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_665 N_A_693_369#_c_620_n N_A_201_47#_c_2001_n 0.0423006f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_666 N_A_693_369#_c_621_n N_A_201_47#_c_2001_n 0.030156f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_667 N_A_693_369#_c_611_n N_A_201_47#_c_2004_n 0.00118188f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_668 N_A_693_369#_c_620_n N_A_201_47#_c_2004_n 0.0257219f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_669 N_A_693_369#_c_624_n N_A_201_47#_c_2004_n 0.00187515f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_670 N_A_693_369#_c_593_n N_A_201_47#_c_1998_n 0.0062731f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_671 N_A_693_369#_c_611_n N_A_201_47#_c_1998_n 0.00244962f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_672 N_A_693_369#_c_624_n N_A_201_47#_c_1998_n 0.0103278f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_673 N_A_693_369#_c_681_p A_1643_329# 0.00203855f $X=8.485 $Y=1.812 $X2=-0.19
+ $Y2=-0.24
cc_674 N_A_693_369#_c_714_p A_1643_329# 0.001538f $X=8.295 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_675 N_A_693_369#_c_597_n N_VGND_c_2145_n 0.0239409f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_676 N_A_693_369#_c_592_n N_VGND_c_2146_n 0.00312892f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_677 N_A_693_369#_c_596_n N_VGND_c_2146_n 2.23286e-19 $X=4.317 $Y=0.805 $X2=0
+ $Y2=0
cc_678 N_A_693_369#_c_597_n N_VGND_c_2146_n 0.0176685f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_679 N_A_693_369#_c_598_n N_VGND_c_2146_n 0.0235008f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_680 N_A_693_369#_c_601_n N_VGND_c_2146_n 4.8449e-19 $X=4.21 $Y=1.255 $X2=0
+ $Y2=0
cc_681 N_A_693_369#_c_597_n N_VGND_c_2149_n 0.0127969f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_682 N_A_693_369#_c_598_n N_VGND_c_2149_n 0.00317989f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_683 N_A_693_369#_M1003_g N_VGND_c_2151_n 0.00362032f $X=9.7 $Y=0.445 $X2=0
+ $Y2=0
cc_684 N_A_693_369#_c_604_n N_VGND_c_2151_n 0.00312232f $X=9.52 $Y=0.812 $X2=0
+ $Y2=0
cc_685 N_A_693_369#_c_605_n N_VGND_c_2151_n 0.00486578f $X=8.785 $Y=0.812 $X2=0
+ $Y2=0
cc_686 N_A_693_369#_c_592_n N_VGND_c_2155_n 0.00565513f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_687 N_A_693_369#_c_593_n N_VGND_c_2155_n 0.00394222f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_688 N_A_693_369#_c_594_n N_VGND_c_2155_n 0.00585385f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_689 N_A_693_369#_c_598_n N_VGND_c_2155_n 6.403e-19 $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_690 N_A_693_369#_M1017_s N_VGND_c_2157_n 0.00388795f $X=3.495 $Y=0.235 $X2=0
+ $Y2=0
cc_691 N_A_693_369#_c_592_n N_VGND_c_2157_n 0.0113329f $X=4.35 $Y=0.73 $X2=0
+ $Y2=0
cc_692 N_A_693_369#_c_593_n N_VGND_c_2157_n 0.00371212f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_693 N_A_693_369#_c_594_n N_VGND_c_2157_n 0.0121314f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_694 N_A_693_369#_M1003_g N_VGND_c_2157_n 0.00557586f $X=9.7 $Y=0.445 $X2=0
+ $Y2=0
cc_695 N_A_693_369#_c_597_n N_VGND_c_2157_n 0.00703355f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_696 N_A_693_369#_c_598_n N_VGND_c_2157_n 0.00765233f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_697 N_A_693_369#_c_604_n N_VGND_c_2157_n 0.00715642f $X=9.52 $Y=0.812 $X2=0
+ $Y2=0
cc_698 N_A_693_369#_c_605_n N_VGND_c_2157_n 0.00847772f $X=8.785 $Y=0.812 $X2=0
+ $Y2=0
cc_699 N_A_693_369#_c_605_n N_VGND_c_2161_n 0.00757352f $X=8.785 $Y=0.812 $X2=0
+ $Y2=0
cc_700 N_A_693_369#_c_604_n A_1645_47# 0.00355082f $X=9.52 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_701 N_A_693_369#_c_605_n A_1645_47# 0.00939028f $X=8.785 $Y=0.812 $X2=-0.19
+ $Y2=-0.24
cc_702 N_A_877_369#_M1023_g N_A_1229_21#_M1016_g 0.0469974f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_703 N_A_877_369#_M1023_g N_A_1229_21#_c_1066_n 0.00658605f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_704 N_A_877_369#_c_885_n N_A_1229_21#_c_1066_n 0.0031108f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_705 N_A_877_369#_c_885_n N_A_1229_21#_c_1073_n 5.84337e-19 $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_706 N_A_877_369#_c_885_n N_A_1229_21#_c_1067_n 0.00911256f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_707 N_A_877_369#_M1023_g N_A_1229_21#_c_1069_n 0.00133724f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_708 N_A_877_369#_c_885_n N_A_1229_21#_c_1069_n 0.00983807f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_709 N_A_877_369#_c_885_n N_A_1229_21#_c_1070_n 0.00306049f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_710 N_A_877_369#_c_881_n N_A_1075_413#_c_1163_n 0.0141556f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_711 N_A_877_369#_M1023_g N_A_1075_413#_c_1163_n 0.0220882f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_712 N_A_877_369#_c_885_n N_A_1075_413#_c_1163_n 0.0327905f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_713 N_A_877_369#_c_885_n N_A_1075_413#_c_1176_n 3.47492e-19 $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_714 N_A_877_369#_c_881_n N_A_1075_413#_c_1164_n 0.00570521f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_715 N_A_877_369#_c_885_n N_A_1075_413#_c_1164_n 0.0218948f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_716 N_A_877_369#_c_891_n N_A_1075_413#_c_1164_n 3.61543e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_717 N_A_877_369#_c_885_n N_A_1075_413#_c_1165_n 0.0189259f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_718 N_A_877_369#_c_885_n N_A_1075_413#_c_1166_n 0.0111401f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_719 N_A_877_369#_c_885_n N_A_1075_413#_c_1167_n 0.0165793f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_720 N_A_877_369#_c_885_n N_A_1075_413#_c_1169_n 0.0392923f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_721 N_A_877_369#_c_885_n N_A_1075_413#_c_1170_n 0.00146646f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_722 N_A_877_369#_c_897_n N_SET_B_c_1324_n 0.00128196f $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_723 N_A_877_369#_c_885_n N_SET_B_c_1324_n 0.0959458f $X=8.94 $Y=1.19 $X2=0
+ $Y2=0
cc_724 N_A_877_369#_c_886_n N_SET_B_c_1324_n 0.0341086f $X=9.055 $Y=1.19 $X2=0
+ $Y2=0
cc_725 N_A_877_369#_c_888_n N_SET_B_c_1324_n 0.0191646f $X=9.135 $Y=1.19 $X2=0
+ $Y2=0
cc_726 N_A_877_369#_c_885_n N_SET_B_c_1325_n 0.0308357f $X=8.94 $Y=1.19 $X2=0
+ $Y2=0
cc_727 N_A_877_369#_c_897_n N_SET_B_c_1326_n 7.0679e-19 $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_728 N_A_877_369#_c_888_n N_SET_B_c_1326_n 0.00271248f $X=9.135 $Y=1.19 $X2=0
+ $Y2=0
cc_729 N_A_877_369#_M1007_g N_SET_B_c_1327_n 4.40484e-19 $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_730 N_A_877_369#_c_897_n N_SET_B_c_1327_n 9.25038e-19 $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_731 N_A_877_369#_c_888_n N_SET_B_c_1327_n 0.0131909f $X=9.135 $Y=1.19 $X2=0
+ $Y2=0
cc_732 N_A_877_369#_c_885_n N_SET_B_c_1328_n 0.00141286f $X=8.94 $Y=1.19 $X2=0
+ $Y2=0
cc_733 N_A_877_369#_c_888_n N_A_1921_295#_c_1456_n 9.93036e-19 $X=9.135 $Y=1.19
+ $X2=0 $Y2=0
cc_734 N_A_877_369#_c_897_n N_A_1921_295#_c_1457_n 0.0196293f $X=9.115 $Y=1.99
+ $X2=0 $Y2=0
cc_735 N_A_877_369#_M1007_g N_A_1921_295#_c_1459_n 0.00238957f $X=9.09 $Y=0.555
+ $X2=0 $Y2=0
cc_736 N_A_877_369#_c_897_n N_A_1921_295#_c_1459_n 0.0163679f $X=9.115 $Y=1.99
+ $X2=0 $Y2=0
cc_737 N_A_877_369#_c_888_n N_A_1921_295#_c_1459_n 4.84072e-19 $X=9.135 $Y=1.19
+ $X2=0 $Y2=0
cc_738 N_A_877_369#_c_888_n N_A_1921_295#_c_1449_n 0.00357125f $X=9.135 $Y=1.19
+ $X2=0 $Y2=0
cc_739 N_A_877_369#_c_897_n N_A_1725_329#_c_1574_n 0.0168408f $X=9.115 $Y=1.99
+ $X2=0 $Y2=0
cc_740 N_A_877_369#_c_888_n N_A_1725_329#_c_1574_n 0.0164674f $X=9.135 $Y=1.19
+ $X2=0 $Y2=0
cc_741 N_A_877_369#_M1007_g N_A_1725_329#_c_1575_n 0.0183431f $X=9.09 $Y=0.555
+ $X2=0 $Y2=0
cc_742 N_A_877_369#_c_897_n N_A_1725_329#_c_1569_n 0.00445422f $X=9.115 $Y=1.99
+ $X2=0 $Y2=0
cc_743 N_A_877_369#_c_888_n N_A_1725_329#_c_1569_n 5.99952e-19 $X=9.135 $Y=1.19
+ $X2=0 $Y2=0
cc_744 N_A_877_369#_c_893_n N_VPWR_c_1816_n 4.12218e-19 $X=5.195 $Y=1.915 $X2=0
+ $Y2=0
cc_745 N_A_877_369#_c_894_n N_VPWR_c_1816_n 0.00206689f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_746 N_A_877_369#_c_895_n N_VPWR_c_1816_n 0.00702461f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_747 N_A_877_369#_c_898_n N_VPWR_c_1816_n 0.0242014f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_748 N_A_877_369#_c_897_n N_VPWR_c_1817_n 0.00430708f $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_749 N_A_877_369#_M1025_d N_VPWR_c_1803_n 0.00224652f $X=4.385 $Y=1.845 $X2=0
+ $Y2=0
cc_750 N_A_877_369#_c_894_n N_VPWR_c_1803_n 0.00154765f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_751 N_A_877_369#_c_895_n N_VPWR_c_1803_n 0.00872443f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_752 N_A_877_369#_c_897_n N_VPWR_c_1803_n 0.00662364f $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_753 N_A_877_369#_c_898_n N_VPWR_c_1803_n 0.00627246f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_754 N_A_877_369#_c_898_n N_VPWR_c_1822_n 0.0122663f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_755 N_A_877_369#_c_897_n N_VPWR_c_1825_n 0.00124505f $X=9.115 $Y=1.99 $X2=0
+ $Y2=0
cc_756 N_A_877_369#_c_884_n N_A_201_47#_c_1995_n 0.041221f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_757 N_A_877_369#_c_892_n N_A_201_47#_c_1999_n 0.00358193f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_758 N_A_877_369#_c_899_n N_A_201_47#_c_1999_n 0.0324615f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_759 N_A_877_369#_c_885_n N_A_201_47#_c_1999_n 6.11234e-19 $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_760 N_A_877_369#_c_892_n N_A_201_47#_c_2000_n 0.00244422f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_761 N_A_877_369#_c_893_n N_A_201_47#_c_2000_n 0.00940185f $X=5.195 $Y=1.915
+ $X2=0 $Y2=0
cc_762 N_A_877_369#_c_894_n N_A_201_47#_c_2000_n 0.00335679f $X=5.04 $Y=1.915
+ $X2=0 $Y2=0
cc_763 N_A_877_369#_c_895_n N_A_201_47#_c_2000_n 0.00398401f $X=5.285 $Y=1.99
+ $X2=0 $Y2=0
cc_764 N_A_877_369#_c_898_n N_A_201_47#_c_2000_n 0.0324615f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_765 N_A_877_369#_c_885_n N_A_201_47#_c_1996_n 0.00517494f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_766 N_A_877_369#_c_890_n N_A_201_47#_c_1996_n 3.91268e-19 $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_767 N_A_877_369#_c_891_n N_A_201_47#_c_1996_n 9.17329e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_768 N_A_877_369#_c_892_n N_A_201_47#_c_2001_n 0.00251435f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_769 N_A_877_369#_c_899_n N_A_201_47#_c_2001_n 0.0189338f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_770 N_A_877_369#_c_885_n N_A_201_47#_c_2001_n 0.00685911f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_771 N_A_877_369#_c_889_n N_A_201_47#_c_2001_n 0.0014563f $X=4.72 $Y=1.185
+ $X2=0 $Y2=0
cc_772 N_A_877_369#_c_890_n N_A_201_47#_c_2001_n 0.0250391f $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_773 N_A_877_369#_c_891_n N_A_201_47#_c_2001_n 8.40015e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_774 N_A_877_369#_c_892_n N_A_201_47#_c_2004_n 8.26579e-19 $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_775 N_A_877_369#_c_899_n N_A_201_47#_c_2004_n 0.00217539f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_776 N_A_877_369#_c_885_n N_A_201_47#_c_2004_n 0.0260799f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_777 N_A_877_369#_c_891_n N_A_201_47#_c_2004_n 5.52268e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_778 N_A_877_369#_c_892_n N_A_201_47#_c_1998_n 0.00416664f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_779 N_A_877_369#_c_881_n N_A_201_47#_c_1998_n 0.00791292f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_780 N_A_877_369#_M1023_g N_A_201_47#_c_1998_n 8.1098e-19 $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_781 N_A_877_369#_c_884_n N_A_201_47#_c_1998_n 0.0138333f $X=4.56 $Y=0.42
+ $X2=0 $Y2=0
cc_782 N_A_877_369#_c_899_n N_A_201_47#_c_1998_n 0.00871828f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_783 N_A_877_369#_c_885_n N_A_201_47#_c_1998_n 0.0126669f $X=8.94 $Y=1.19
+ $X2=0 $Y2=0
cc_784 N_A_877_369#_c_889_n N_A_201_47#_c_1998_n 0.0222258f $X=4.72 $Y=1.185
+ $X2=0 $Y2=0
cc_785 N_A_877_369#_c_890_n N_A_201_47#_c_1998_n 0.0023779f $X=4.865 $Y=1.185
+ $X2=0 $Y2=0
cc_786 N_A_877_369#_c_891_n N_A_201_47#_c_1998_n 0.00621958f $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_787 N_A_877_369#_M1007_g N_VGND_c_2151_n 0.00367042f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_788 N_A_877_369#_M1023_g N_VGND_c_2155_n 0.00717785f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_789 N_A_877_369#_c_884_n N_VGND_c_2155_n 0.0144177f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_790 N_A_877_369#_M1015_d N_VGND_c_2157_n 0.00382094f $X=4.425 $Y=0.235 $X2=0
+ $Y2=0
cc_791 N_A_877_369#_M1023_g N_VGND_c_2157_n 0.00537275f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_792 N_A_877_369#_M1007_g N_VGND_c_2157_n 0.00708667f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_793 N_A_877_369#_c_884_n N_VGND_c_2157_n 0.00801045f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_794 N_A_877_369#_M1007_g N_VGND_c_2161_n 0.0132789f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_795 N_A_877_369#_c_885_n N_VGND_c_2161_n 0.00635838f $X=8.94 $Y=1.19 $X2=0
+ $Y2=0
cc_796 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1160_n 5.62208e-19 $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_797 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1172_n 0.00632289f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_798 N_A_1229_21#_c_1072_n N_A_1075_413#_c_1172_n 0.0171889f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_799 N_A_1229_21#_c_1073_n N_A_1075_413#_c_1172_n 0.00183365f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_800 N_A_1229_21#_c_1072_n N_A_1075_413#_c_1173_n 0.0150522f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_801 N_A_1229_21#_c_1073_n N_A_1075_413#_c_1173_n 4.03149e-19 $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_802 N_A_1229_21#_c_1074_n N_A_1075_413#_c_1173_n 0.0160003f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_803 N_A_1229_21#_c_1067_n N_A_1075_413#_c_1161_n 0.00198418f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_804 N_A_1229_21#_c_1068_n N_A_1075_413#_c_1161_n 0.0077537f $X=6.95 $Y=0.51
+ $X2=0 $Y2=0
cc_805 N_A_1229_21#_M1016_g N_A_1075_413#_c_1162_n 8.49245e-19 $X=6.22 $Y=0.445
+ $X2=0 $Y2=0
cc_806 N_A_1229_21#_c_1067_n N_A_1075_413#_c_1162_n 0.00806227f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_807 N_A_1229_21#_c_1069_n N_A_1075_413#_c_1162_n 0.00110084f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_808 N_A_1229_21#_c_1070_n N_A_1075_413#_c_1162_n 0.00784562f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_809 N_A_1229_21#_M1016_g N_A_1075_413#_c_1163_n 0.00122809f $X=6.22 $Y=0.445
+ $X2=0 $Y2=0
cc_810 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1163_n 0.00261079f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_811 N_A_1229_21#_c_1069_n N_A_1075_413#_c_1163_n 0.0269973f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_812 N_A_1229_21#_c_1070_n N_A_1075_413#_c_1163_n 0.00113583f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_813 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1176_n 0.011517f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_814 N_A_1229_21#_c_1072_n N_A_1075_413#_c_1176_n 0.00116159f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_815 N_A_1229_21#_c_1073_n N_A_1075_413#_c_1176_n 0.0201747f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_816 N_A_1229_21#_c_1075_n N_A_1075_413#_c_1176_n 0.00880623f $X=6.595 $Y=2.02
+ $X2=0 $Y2=0
cc_817 N_A_1229_21#_c_1069_n N_A_1075_413#_c_1164_n 0.0192437f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_818 N_A_1229_21#_c_1070_n N_A_1075_413#_c_1164_n 0.0018579f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_819 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1165_n 0.0152311f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_820 N_A_1229_21#_c_1072_n N_A_1075_413#_c_1165_n 0.00260846f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_821 N_A_1229_21#_c_1073_n N_A_1075_413#_c_1165_n 0.0109804f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_822 N_A_1229_21#_c_1067_n N_A_1075_413#_c_1165_n 0.00808722f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_823 N_A_1229_21#_c_1074_n N_A_1075_413#_c_1165_n 0.00696445f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_824 N_A_1229_21#_c_1070_n N_A_1075_413#_c_1165_n 5.30627e-19 $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_825 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1166_n 0.0017292f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_826 N_A_1229_21#_c_1067_n N_A_1075_413#_c_1166_n 0.0178097f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_827 N_A_1229_21#_c_1069_n N_A_1075_413#_c_1166_n 0.0020275f $X=6.285 $Y=0.72
+ $X2=0 $Y2=0
cc_828 N_A_1229_21#_c_1070_n N_A_1075_413#_c_1166_n 0.00156611f $X=6.31 $Y=0.93
+ $X2=0 $Y2=0
cc_829 N_A_1229_21#_c_1074_n N_A_1075_413#_c_1169_n 0.00267752f $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_830 N_A_1229_21#_c_1066_n N_A_1075_413#_c_1170_n 0.0115036f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_831 N_A_1229_21#_c_1067_n N_A_1075_413#_c_1170_n 0.00227132f $X=6.785 $Y=0.72
+ $X2=0 $Y2=0
cc_832 N_A_1229_21#_c_1074_n N_A_1075_413#_c_1170_n 6.97279e-19 $X=7.155 $Y=2.02
+ $X2=0 $Y2=0
cc_833 N_A_1229_21#_c_1074_n N_SET_B_c_1317_n 0.00719198f $X=7.155 $Y=2.02
+ $X2=-0.19 $Y2=-0.24
cc_834 N_A_1229_21#_c_1128_p N_SET_B_c_1317_n 0.00390541f $X=7.265 $Y=2.285
+ $X2=-0.19 $Y2=-0.24
cc_835 N_A_1229_21#_c_1073_n N_SET_B_c_1328_n 0.005781f $X=6.51 $Y=1.74 $X2=0
+ $Y2=0
cc_836 N_A_1229_21#_c_1074_n N_SET_B_c_1328_n 0.0155982f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_837 N_A_1229_21#_c_1074_n N_VPWR_M1038_d 0.00298622f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_838 N_A_1229_21#_c_1075_n N_VPWR_M1038_d 0.00153636f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_839 N_A_1229_21#_c_1072_n N_VPWR_c_1816_n 0.00743866f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_840 N_A_1229_21#_M1009_d N_VPWR_c_1803_n 0.00331536f $X=7.095 $Y=2.065 $X2=0
+ $Y2=0
cc_841 N_A_1229_21#_c_1072_n N_VPWR_c_1803_n 0.00849347f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_842 N_A_1229_21#_c_1074_n N_VPWR_c_1803_n 0.0042909f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_843 N_A_1229_21#_c_1075_n N_VPWR_c_1803_n 7.82982e-19 $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_844 N_A_1229_21#_c_1128_p N_VPWR_c_1803_n 0.00471488f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_845 N_A_1229_21#_c_1072_n N_VPWR_c_1823_n 0.0056962f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_846 N_A_1229_21#_c_1074_n N_VPWR_c_1823_n 0.0164669f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_847 N_A_1229_21#_c_1075_n N_VPWR_c_1823_n 0.0102436f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_848 N_A_1229_21#_c_1128_p N_VPWR_c_1823_n 0.00867119f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_849 N_A_1229_21#_c_1074_n N_VPWR_c_1824_n 0.00479971f $X=7.155 $Y=2.02 $X2=0
+ $Y2=0
cc_850 N_A_1229_21#_c_1128_p N_VPWR_c_1824_n 0.0165337f $X=7.265 $Y=2.285 $X2=0
+ $Y2=0
cc_851 N_A_1229_21#_c_1067_n N_VGND_M1016_d 8.64202e-19 $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_852 N_A_1229_21#_c_1069_n N_VGND_M1016_d 0.00133208f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_853 N_A_1229_21#_M1016_g N_VGND_c_2155_n 0.014377f $X=6.22 $Y=0.445 $X2=0
+ $Y2=0
cc_854 N_A_1229_21#_c_1067_n N_VGND_c_2155_n 0.00919218f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_855 N_A_1229_21#_c_1068_n N_VGND_c_2155_n 0.0164501f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_856 N_A_1229_21#_c_1069_n N_VGND_c_2155_n 0.0212099f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_857 N_A_1229_21#_c_1070_n N_VGND_c_2155_n 8.18098e-19 $X=6.31 $Y=0.93 $X2=0
+ $Y2=0
cc_858 N_A_1229_21#_M1020_s N_VGND_c_2157_n 0.00468266f $X=6.825 $Y=0.235 $X2=0
+ $Y2=0
cc_859 N_A_1229_21#_c_1067_n N_VGND_c_2157_n 0.00594673f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_860 N_A_1229_21#_c_1068_n N_VGND_c_2157_n 0.00949852f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_861 N_A_1229_21#_c_1069_n N_VGND_c_2157_n 0.00174322f $X=6.285 $Y=0.72 $X2=0
+ $Y2=0
cc_862 N_A_1229_21#_c_1067_n N_VGND_c_2160_n 0.00346394f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_863 N_A_1229_21#_c_1068_n N_VGND_c_2160_n 0.0172232f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_864 N_A_1229_21#_c_1067_n N_VGND_c_2161_n 0.0118068f $X=6.785 $Y=0.72 $X2=0
+ $Y2=0
cc_865 N_A_1229_21#_c_1068_n N_VGND_c_2161_n 0.0251021f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_866 N_A_1075_413#_c_1172_n N_SET_B_c_1317_n 0.0252095f $X=7.005 $Y=1.89
+ $X2=-0.19 $Y2=-0.24
cc_867 N_A_1075_413#_c_1173_n N_SET_B_c_1317_n 0.0108477f $X=7.005 $Y=1.99
+ $X2=-0.19 $Y2=-0.24
cc_868 N_A_1075_413#_c_1175_n N_SET_B_c_1317_n 0.0311852f $X=8.125 $Y=1.57
+ $X2=-0.19 $Y2=-0.24
cc_869 N_A_1075_413#_c_1162_n N_SET_B_c_1317_n 2.44193e-19 $X=7.26 $Y=0.805
+ $X2=-0.19 $Y2=-0.24
cc_870 N_A_1075_413#_c_1169_n N_SET_B_c_1317_n 0.00135225f $X=7.905 $Y=1.15
+ $X2=-0.19 $Y2=-0.24
cc_871 N_A_1075_413#_c_1160_n N_SET_B_M1024_g 0.0171583f $X=7.005 $Y=1.095 $X2=0
+ $Y2=0
cc_872 N_A_1075_413#_c_1161_n N_SET_B_M1024_g 0.0504282f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_873 N_A_1075_413#_c_1174_n N_SET_B_M1024_g 0.00502284f $X=8.125 $Y=1.47 $X2=0
+ $Y2=0
cc_874 N_A_1075_413#_c_1166_n N_SET_B_M1024_g 5.27107e-19 $X=6.975 $Y=1.185
+ $X2=0 $Y2=0
cc_875 N_A_1075_413#_c_1167_n N_SET_B_M1024_g 0.00114053f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_876 N_A_1075_413#_c_1168_n N_SET_B_M1024_g 0.0161502f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_877 N_A_1075_413#_c_1169_n N_SET_B_M1024_g 0.0165077f $X=7.905 $Y=1.15 $X2=0
+ $Y2=0
cc_878 N_A_1075_413#_c_1171_n N_SET_B_M1024_g 0.0184897f $X=8.09 $Y=0.995 $X2=0
+ $Y2=0
cc_879 N_A_1075_413#_c_1174_n N_SET_B_c_1324_n 0.00137145f $X=8.125 $Y=1.47
+ $X2=0 $Y2=0
cc_880 N_A_1075_413#_c_1175_n N_SET_B_c_1324_n 0.00387957f $X=8.125 $Y=1.57
+ $X2=0 $Y2=0
cc_881 N_A_1075_413#_c_1167_n N_SET_B_c_1324_n 0.00383469f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_882 N_A_1075_413#_c_1168_n N_SET_B_c_1324_n 0.00108862f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_883 N_A_1075_413#_c_1169_n N_SET_B_c_1324_n 0.00505042f $X=7.905 $Y=1.15
+ $X2=0 $Y2=0
cc_884 N_A_1075_413#_c_1172_n N_SET_B_c_1325_n 4.79368e-19 $X=7.005 $Y=1.89
+ $X2=0 $Y2=0
cc_885 N_A_1075_413#_c_1174_n N_SET_B_c_1325_n 6.70195e-19 $X=8.125 $Y=1.47
+ $X2=0 $Y2=0
cc_886 N_A_1075_413#_c_1175_n N_SET_B_c_1325_n 6.64941e-19 $X=8.125 $Y=1.57
+ $X2=0 $Y2=0
cc_887 N_A_1075_413#_c_1169_n N_SET_B_c_1325_n 0.00206701f $X=7.905 $Y=1.15
+ $X2=0 $Y2=0
cc_888 N_A_1075_413#_c_1172_n N_SET_B_c_1328_n 0.00633121f $X=7.005 $Y=1.89
+ $X2=0 $Y2=0
cc_889 N_A_1075_413#_c_1174_n N_SET_B_c_1328_n 0.00182229f $X=8.125 $Y=1.47
+ $X2=0 $Y2=0
cc_890 N_A_1075_413#_c_1175_n N_SET_B_c_1328_n 0.00195011f $X=8.125 $Y=1.57
+ $X2=0 $Y2=0
cc_891 N_A_1075_413#_c_1169_n N_SET_B_c_1328_n 0.0358497f $X=7.905 $Y=1.15 $X2=0
+ $Y2=0
cc_892 N_A_1075_413#_c_1190_n N_VPWR_c_1816_n 0.0464661f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_893 N_A_1075_413#_M1006_d N_VPWR_c_1803_n 0.00231251f $X=5.375 $Y=2.065 $X2=0
+ $Y2=0
cc_894 N_A_1075_413#_c_1173_n N_VPWR_c_1803_n 0.00720657f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_895 N_A_1075_413#_c_1190_n N_VPWR_c_1803_n 0.012998f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_896 N_A_1075_413#_c_1173_n N_VPWR_c_1823_n 0.00620668f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_897 N_A_1075_413#_c_1173_n N_VPWR_c_1824_n 0.00512994f $X=7.005 $Y=1.99 $X2=0
+ $Y2=0
cc_898 N_A_1075_413#_c_1175_n N_VPWR_c_1825_n 0.0209123f $X=8.125 $Y=1.57 $X2=0
+ $Y2=0
cc_899 N_A_1075_413#_c_1163_n N_A_201_47#_c_1995_n 0.040178f $X=5.55 $Y=0.42
+ $X2=0 $Y2=0
cc_900 N_A_1075_413#_c_1164_n N_A_201_47#_c_1998_n 0.00906057f $X=6.205 $Y=1.31
+ $X2=0 $Y2=0
cc_901 N_A_1075_413#_c_1190_n A_1169_413# 0.00692155f $X=6.035 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_902 N_A_1075_413#_c_1176_n A_1169_413# 0.00130666f $X=6.12 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_903 N_A_1075_413#_c_1161_n N_VGND_c_2155_n 0.00172114f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_904 N_A_1075_413#_c_1163_n N_VGND_c_2155_n 0.0270576f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_905 N_A_1075_413#_M1026_d N_VGND_c_2157_n 0.00428929f $X=5.415 $Y=0.235 $X2=0
+ $Y2=0
cc_906 N_A_1075_413#_c_1161_n N_VGND_c_2157_n 0.00630011f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_907 N_A_1075_413#_c_1162_n N_VGND_c_2157_n 0.00363714f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_908 N_A_1075_413#_c_1163_n N_VGND_c_2157_n 0.0155321f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_909 N_A_1075_413#_c_1161_n N_VGND_c_2160_n 0.00271402f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_910 N_A_1075_413#_c_1162_n N_VGND_c_2160_n 0.00305109f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_911 N_A_1075_413#_c_1161_n N_VGND_c_2161_n 0.017478f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_912 N_A_1075_413#_c_1162_n N_VGND_c_2161_n 0.00301799f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_913 N_A_1075_413#_c_1168_n N_VGND_c_2161_n 7.27879e-19 $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_914 N_A_1075_413#_c_1169_n N_VGND_c_2161_n 0.0788733f $X=7.905 $Y=1.15 $X2=0
+ $Y2=0
cc_915 N_A_1075_413#_c_1171_n N_VGND_c_2161_n 0.0314809f $X=8.09 $Y=0.995 $X2=0
+ $Y2=0
cc_916 N_SET_B_c_1319_n N_A_1921_295#_c_1456_n 0.00590071f $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_917 N_SET_B_c_1322_n N_A_1921_295#_c_1456_n 3.59733e-19 $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_918 N_SET_B_c_1323_n N_A_1921_295#_c_1456_n 0.00440707f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_919 N_SET_B_c_1327_n N_A_1921_295#_c_1456_n 0.00596796f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_920 N_SET_B_c_1319_n N_A_1921_295#_c_1457_n 0.0136437f $X=10.26 $Y=1.99 $X2=0
+ $Y2=0
cc_921 N_SET_B_c_1319_n N_A_1921_295#_c_1458_n 0.00158074f $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_922 N_SET_B_c_1322_n N_A_1921_295#_c_1458_n 0.0162082f $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_923 N_SET_B_c_1323_n N_A_1921_295#_c_1458_n 0.00547816f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_924 N_SET_B_c_1326_n N_A_1921_295#_c_1458_n 0.00178525f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_925 N_SET_B_c_1327_n N_A_1921_295#_c_1458_n 0.00395328f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_926 N_SET_B_c_1327_n N_A_1921_295#_c_1459_n 0.00465625f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_927 N_SET_B_M1031_g N_A_1921_295#_M1027_g 0.0227341f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_928 N_SET_B_M1031_g N_A_1921_295#_c_1449_n 0.0108005f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_929 N_SET_B_c_1321_n N_A_1921_295#_c_1449_n 0.00547816f $X=10.53 $Y=1.6 $X2=0
+ $Y2=0
cc_930 N_SET_B_c_1326_n N_A_1921_295#_c_1449_n 0.00165716f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_931 N_SET_B_c_1327_n N_A_1921_295#_c_1449_n 0.00171402f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_932 N_SET_B_M1031_g N_A_1921_295#_c_1450_n 0.0014323f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_933 N_SET_B_c_1319_n N_A_1921_295#_c_1451_n 0.00138929f $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_934 N_SET_B_M1031_g N_A_1921_295#_c_1451_n 0.0208264f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_935 N_SET_B_c_1322_n N_A_1921_295#_c_1451_n 2.9881e-19 $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_936 N_SET_B_M1031_g N_A_1921_295#_c_1452_n 0.0107344f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_937 N_SET_B_c_1321_n N_A_1921_295#_c_1452_n 0.00322511f $X=10.53 $Y=1.6 $X2=0
+ $Y2=0
cc_938 N_SET_B_c_1322_n N_A_1921_295#_c_1452_n 0.028507f $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_939 N_SET_B_c_1322_n N_A_1921_295#_c_1462_n 0.0182139f $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_940 N_SET_B_c_1321_n N_A_1725_329#_c_1552_n 0.0178474f $X=10.53 $Y=1.6 $X2=0
+ $Y2=0
cc_941 N_SET_B_c_1322_n N_A_1725_329#_c_1552_n 0.00236806f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_942 N_SET_B_c_1323_n N_A_1725_329#_c_1552_n 0.00294313f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_943 N_SET_B_M1031_g N_A_1725_329#_c_1555_n 0.0201382f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_944 N_SET_B_M1031_g N_A_1725_329#_c_1556_n 0.0126062f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_945 N_SET_B_c_1324_n N_A_1725_329#_c_1574_n 0.0148412f $X=9.565 $Y=1.53 $X2=0
+ $Y2=0
cc_946 N_SET_B_M1031_g N_A_1725_329#_c_1575_n 0.0101264f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_947 N_SET_B_c_1319_n N_A_1725_329#_c_1567_n 0.0138916f $X=10.26 $Y=1.99 $X2=0
+ $Y2=0
cc_948 N_SET_B_c_1322_n N_A_1725_329#_c_1567_n 0.03927f $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_949 N_SET_B_c_1326_n N_A_1725_329#_c_1567_n 0.00127121f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_950 N_SET_B_c_1327_n N_A_1725_329#_c_1567_n 0.0115337f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_951 N_SET_B_M1031_g N_A_1725_329#_c_1558_n 0.00829661f $X=10.59 $Y=0.445
+ $X2=0 $Y2=0
cc_952 N_SET_B_c_1319_n N_A_1725_329#_c_1568_n 0.00376998f $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_953 N_SET_B_c_1322_n N_A_1725_329#_c_1568_n 0.00700059f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_954 N_SET_B_M1031_g N_A_1725_329#_c_1559_n 0.00596999f $X=10.59 $Y=0.445
+ $X2=0 $Y2=0
cc_955 N_SET_B_M1031_g N_A_1725_329#_c_1560_n 0.0034132f $X=10.59 $Y=0.445 $X2=0
+ $Y2=0
cc_956 N_SET_B_c_1321_n N_A_1725_329#_c_1561_n 0.0201382f $X=10.53 $Y=1.6 $X2=0
+ $Y2=0
cc_957 N_SET_B_c_1319_n N_A_1725_329#_c_1569_n 7.06352e-19 $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_958 N_SET_B_c_1324_n N_A_1725_329#_c_1569_n 0.0012603f $X=9.565 $Y=1.53 $X2=0
+ $Y2=0
cc_959 N_SET_B_c_1326_n N_A_1725_329#_c_1569_n 0.00122335f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1327_n N_A_1725_329#_c_1569_n 0.00798024f $X=9.71 $Y=1.53 $X2=0
+ $Y2=0
cc_961 N_SET_B_c_1319_n N_A_1725_329#_c_1608_n 0.00893486f $X=10.26 $Y=1.99
+ $X2=0 $Y2=0
cc_962 N_SET_B_c_1322_n N_A_1725_329#_c_1608_n 0.0150414f $X=10.53 $Y=1.63 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1322_n N_A_1725_329#_c_1570_n 0.00970636f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_964 N_SET_B_c_1323_n N_A_1725_329#_c_1570_n 0.00273595f $X=10.53 $Y=1.63
+ $X2=0 $Y2=0
cc_965 N_SET_B_c_1319_n N_VPWR_c_1807_n 0.00888095f $X=10.26 $Y=1.99 $X2=0 $Y2=0
cc_966 N_SET_B_c_1319_n N_VPWR_c_1808_n 0.00298416f $X=10.26 $Y=1.99 $X2=0 $Y2=0
cc_967 N_SET_B_c_1319_n N_VPWR_c_1810_n 0.0054346f $X=10.26 $Y=1.99 $X2=0 $Y2=0
cc_968 N_SET_B_c_1317_n N_VPWR_c_1803_n 0.00847755f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_969 N_SET_B_c_1319_n N_VPWR_c_1803_n 0.00655278f $X=10.26 $Y=1.99 $X2=0 $Y2=0
cc_970 N_SET_B_c_1317_n N_VPWR_c_1824_n 0.00742527f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_971 N_SET_B_c_1317_n N_VPWR_c_1825_n 0.00364248f $X=7.595 $Y=1.99 $X2=0 $Y2=0
cc_972 N_SET_B_c_1324_n N_VPWR_c_1825_n 5.22073e-19 $X=9.565 $Y=1.53 $X2=0 $Y2=0
cc_973 N_SET_B_M1031_g N_VGND_c_2147_n 0.00533087f $X=10.59 $Y=0.445 $X2=0 $Y2=0
cc_974 N_SET_B_M1031_g N_VGND_c_2151_n 0.00384182f $X=10.59 $Y=0.445 $X2=0 $Y2=0
cc_975 N_SET_B_M1031_g N_VGND_c_2157_n 0.00605525f $X=10.59 $Y=0.445 $X2=0 $Y2=0
cc_976 N_SET_B_M1024_g N_VGND_c_2161_n 0.0265529f $X=7.62 $Y=0.445 $X2=0 $Y2=0
cc_977 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1552_n 0.020908f $X=11.425 $Y=1.28
+ $X2=0 $Y2=0
cc_978 N_A_1921_295#_c_1463_n N_A_1725_329#_c_1552_n 0.0278731f $X=11.51
+ $Y=2.285 $X2=0 $Y2=0
cc_979 N_A_1921_295#_c_1454_n N_A_1725_329#_c_1552_n 6.04442e-19 $X=11.51
+ $Y=0.42 $X2=0 $Y2=0
cc_980 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1553_n 0.00134819f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_981 N_A_1921_295#_c_1455_n N_A_1725_329#_c_1553_n 0.0170978f $X=11.555
+ $Y=1.28 $X2=0 $Y2=0
cc_982 N_A_1921_295#_c_1453_n N_A_1725_329#_M1032_g 7.43555e-19 $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_983 N_A_1921_295#_c_1463_n N_A_1725_329#_c_1564_n 0.00110434f $X=11.51
+ $Y=2.285 $X2=0 $Y2=0
cc_984 N_A_1921_295#_c_1453_n N_A_1725_329#_c_1555_n 0.00150633f $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_985 N_A_1921_295#_c_1453_n N_A_1725_329#_c_1556_n 0.00693654f $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_986 N_A_1921_295#_c_1454_n N_A_1725_329#_c_1556_n 0.0082592f $X=11.51 $Y=0.42
+ $X2=0 $Y2=0
cc_987 N_A_1921_295#_c_1463_n N_A_1725_329#_c_1566_n 0.00151882f $X=11.51
+ $Y=2.285 $X2=0 $Y2=0
cc_988 N_A_1921_295#_c_1457_n N_A_1725_329#_c_1574_n 6.76132e-19 $X=9.705
+ $Y=1.99 $X2=0 $Y2=0
cc_989 N_A_1921_295#_M1027_g N_A_1725_329#_c_1575_n 0.0158652f $X=10.06 $Y=0.445
+ $X2=0 $Y2=0
cc_990 N_A_1921_295#_c_1450_n N_A_1725_329#_c_1575_n 0.00935668f $X=10.12
+ $Y=1.02 $X2=0 $Y2=0
cc_991 N_A_1921_295#_c_1451_n N_A_1725_329#_c_1575_n 0.00137429f $X=10.12
+ $Y=1.02 $X2=0 $Y2=0
cc_992 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1575_n 0.00488861f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_993 N_A_1921_295#_c_1457_n N_A_1725_329#_c_1567_n 0.00876434f $X=9.705
+ $Y=1.99 $X2=0 $Y2=0
cc_994 N_A_1921_295#_c_1458_n N_A_1725_329#_c_1567_n 0.00194629f $X=9.985
+ $Y=1.55 $X2=0 $Y2=0
cc_995 N_A_1921_295#_M1027_g N_A_1725_329#_c_1558_n 0.00381803f $X=10.06
+ $Y=0.445 $X2=0 $Y2=0
cc_996 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1568_n 0.00616622f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_997 N_A_1921_295#_M1027_g N_A_1725_329#_c_1559_n 7.21921e-19 $X=10.06
+ $Y=0.445 $X2=0 $Y2=0
cc_998 N_A_1921_295#_c_1450_n N_A_1725_329#_c_1559_n 0.0132237f $X=10.12 $Y=1.02
+ $X2=0 $Y2=0
cc_999 N_A_1921_295#_c_1451_n N_A_1725_329#_c_1559_n 0.00102789f $X=10.12
+ $Y=1.02 $X2=0 $Y2=0
cc_1000 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1559_n 0.015092f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_1001 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1560_n 0.0443791f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_1002 N_A_1921_295#_c_1453_n N_A_1725_329#_c_1560_n 0.0196589f $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_1003 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1561_n 0.00501833f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_1004 N_A_1921_295#_c_1453_n N_A_1725_329#_c_1561_n 0.0067596f $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_1005 N_A_1921_295#_c_1457_n N_A_1725_329#_c_1569_n 0.0156991f $X=9.705
+ $Y=1.99 $X2=0 $Y2=0
cc_1006 N_A_1921_295#_c_1452_n N_A_1725_329#_c_1570_n 0.0213588f $X=11.425
+ $Y=1.28 $X2=0 $Y2=0
cc_1007 N_A_1921_295#_c_1463_n N_A_1725_329#_c_1570_n 0.0360588f $X=11.51
+ $Y=2.285 $X2=0 $Y2=0
cc_1008 N_A_1921_295#_c_1454_n N_A_2381_47#_c_1709_n 0.0596011f $X=11.51 $Y=0.42
+ $X2=0 $Y2=0
cc_1009 N_A_1921_295#_c_1463_n N_A_2381_47#_c_1713_n 0.0901388f $X=11.51
+ $Y=2.285 $X2=0 $Y2=0
cc_1010 N_A_1921_295#_c_1455_n N_A_2381_47#_c_1713_n 0.00324854f $X=11.555
+ $Y=1.28 $X2=0 $Y2=0
cc_1011 N_A_1921_295#_c_1453_n N_A_2381_47#_c_1711_n 0.0172076f $X=11.57
+ $Y=1.195 $X2=0 $Y2=0
cc_1012 N_A_1921_295#_c_1455_n N_A_2381_47#_c_1711_n 0.0110951f $X=11.555
+ $Y=1.28 $X2=0 $Y2=0
cc_1013 N_A_1921_295#_c_1457_n N_VPWR_c_1807_n 0.0055538f $X=9.705 $Y=1.99 $X2=0
+ $Y2=0
cc_1014 N_A_1921_295#_c_1463_n N_VPWR_c_1808_n 0.0177194f $X=11.51 $Y=2.285
+ $X2=0 $Y2=0
cc_1015 N_A_1921_295#_c_1463_n N_VPWR_c_1812_n 0.0182101f $X=11.51 $Y=2.285
+ $X2=0 $Y2=0
cc_1016 N_A_1921_295#_c_1457_n N_VPWR_c_1817_n 0.00486131f $X=9.705 $Y=1.99
+ $X2=0 $Y2=0
cc_1017 N_A_1921_295#_M1014_d N_VPWR_c_1803_n 0.00404917f $X=11.365 $Y=2.065
+ $X2=0 $Y2=0
cc_1018 N_A_1921_295#_c_1457_n N_VPWR_c_1803_n 0.00699047f $X=9.705 $Y=1.99
+ $X2=0 $Y2=0
cc_1019 N_A_1921_295#_c_1463_n N_VPWR_c_1803_n 0.00993603f $X=11.51 $Y=2.285
+ $X2=0 $Y2=0
cc_1020 N_A_1921_295#_M1027_g N_VGND_c_2151_n 0.00362032f $X=10.06 $Y=0.445
+ $X2=0 $Y2=0
cc_1021 N_A_1921_295#_c_1454_n N_VGND_c_2153_n 0.0234496f $X=11.51 $Y=0.42 $X2=0
+ $Y2=0
cc_1022 N_A_1921_295#_M1034_d N_VGND_c_2157_n 0.00537869f $X=11.255 $Y=0.235
+ $X2=0 $Y2=0
cc_1023 N_A_1921_295#_M1027_g N_VGND_c_2157_n 0.00541928f $X=10.06 $Y=0.445
+ $X2=0 $Y2=0
cc_1024 N_A_1921_295#_c_1454_n N_VGND_c_2157_n 0.0129422f $X=11.51 $Y=0.42 $X2=0
+ $Y2=0
cc_1025 N_A_1725_329#_M1032_g N_A_2381_47#_c_1707_n 0.0213829f $X=12.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1026 N_A_1725_329#_c_1564_n N_A_2381_47#_c_1707_n 0.0156176f $X=12.265
+ $Y=1.77 $X2=0 $Y2=0
cc_1027 N_A_1725_329#_c_1557_n N_A_2381_47#_c_1707_n 0.00265456f $X=12.24
+ $Y=1.28 $X2=0 $Y2=0
cc_1028 N_A_1725_329#_c_1566_n N_A_2381_47#_c_1707_n 0.00356778f $X=12.265
+ $Y=1.535 $X2=0 $Y2=0
cc_1029 N_A_1725_329#_M1032_g N_A_2381_47#_c_1708_n 0.0219521f $X=12.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1030 N_A_1725_329#_M1032_g N_A_2381_47#_c_1709_n 0.0145903f $X=12.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1031 N_A_1725_329#_c_1552_n N_A_2381_47#_c_1713_n 9.56144e-19 $X=11.275
+ $Y=1.99 $X2=0 $Y2=0
cc_1032 N_A_1725_329#_c_1553_n N_A_2381_47#_c_1713_n 0.00652469f $X=12.165
+ $Y=1.28 $X2=0 $Y2=0
cc_1033 N_A_1725_329#_c_1564_n N_A_2381_47#_c_1713_n 0.0205437f $X=12.265
+ $Y=1.77 $X2=0 $Y2=0
cc_1034 N_A_1725_329#_c_1557_n N_A_2381_47#_c_1713_n 5.85784e-19 $X=12.24
+ $Y=1.28 $X2=0 $Y2=0
cc_1035 N_A_1725_329#_c_1566_n N_A_2381_47#_c_1713_n 0.00722127f $X=12.265
+ $Y=1.535 $X2=0 $Y2=0
cc_1036 N_A_1725_329#_M1032_g N_A_2381_47#_c_1710_n 0.00918507f $X=12.24
+ $Y=0.445 $X2=0 $Y2=0
cc_1037 N_A_1725_329#_c_1564_n N_A_2381_47#_c_1710_n 0.00207256f $X=12.265
+ $Y=1.77 $X2=0 $Y2=0
cc_1038 N_A_1725_329#_c_1557_n N_A_2381_47#_c_1710_n 0.00810845f $X=12.24
+ $Y=1.28 $X2=0 $Y2=0
cc_1039 N_A_1725_329#_c_1553_n N_A_2381_47#_c_1711_n 0.0105257f $X=12.165
+ $Y=1.28 $X2=0 $Y2=0
cc_1040 N_A_1725_329#_M1032_g N_A_2381_47#_c_1711_n 0.00638627f $X=12.24
+ $Y=0.445 $X2=0 $Y2=0
cc_1041 N_A_1725_329#_c_1557_n N_A_2381_47#_c_1711_n 3.38992e-19 $X=12.24
+ $Y=1.28 $X2=0 $Y2=0
cc_1042 N_A_1725_329#_c_1561_n N_A_2381_47#_c_1711_n 2.95577e-19 $X=11.07
+ $Y=0.93 $X2=0 $Y2=0
cc_1043 N_A_1725_329#_c_1570_n N_VPWR_M1014_s 0.0028505f $X=11.04 $Y=1.69 $X2=0
+ $Y2=0
cc_1044 N_A_1725_329#_c_1567_n N_VPWR_c_1807_n 0.0228296f $X=10.395 $Y=1.98
+ $X2=0 $Y2=0
cc_1045 N_A_1725_329#_c_1569_n N_VPWR_c_1807_n 0.0166483f $X=9.605 $Y=1.98 $X2=0
+ $Y2=0
cc_1046 N_A_1725_329#_c_1552_n N_VPWR_c_1808_n 0.0135992f $X=11.275 $Y=1.99
+ $X2=0 $Y2=0
cc_1047 N_A_1725_329#_c_1665_p N_VPWR_c_1808_n 0.0120083f $X=10.495 $Y=2.285
+ $X2=0 $Y2=0
cc_1048 N_A_1725_329#_c_1570_n N_VPWR_c_1808_n 0.0284102f $X=11.04 $Y=1.69 $X2=0
+ $Y2=0
cc_1049 N_A_1725_329#_c_1564_n N_VPWR_c_1809_n 0.00557621f $X=12.265 $Y=1.77
+ $X2=0 $Y2=0
cc_1050 N_A_1725_329#_c_1567_n N_VPWR_c_1810_n 0.00327146f $X=10.395 $Y=1.98
+ $X2=0 $Y2=0
cc_1051 N_A_1725_329#_c_1665_p N_VPWR_c_1810_n 0.0121777f $X=10.495 $Y=2.285
+ $X2=0 $Y2=0
cc_1052 N_A_1725_329#_c_1568_n N_VPWR_c_1810_n 0.00488937f $X=10.875 $Y=1.98
+ $X2=0 $Y2=0
cc_1053 N_A_1725_329#_c_1552_n N_VPWR_c_1812_n 0.00448207f $X=11.275 $Y=1.99
+ $X2=0 $Y2=0
cc_1054 N_A_1725_329#_c_1564_n N_VPWR_c_1812_n 0.00673617f $X=12.265 $Y=1.77
+ $X2=0 $Y2=0
cc_1055 N_A_1725_329#_c_1574_n N_VPWR_c_1817_n 0.0428408f $X=9.52 $Y=2.292 $X2=0
+ $Y2=0
cc_1056 N_A_1725_329#_c_1567_n N_VPWR_c_1817_n 0.00277068f $X=10.395 $Y=1.98
+ $X2=0 $Y2=0
cc_1057 N_A_1725_329#_c_1569_n N_VPWR_c_1817_n 0.00927152f $X=9.605 $Y=1.98
+ $X2=0 $Y2=0
cc_1058 N_A_1725_329#_M1013_d N_VPWR_c_1803_n 0.00444786f $X=8.625 $Y=1.645
+ $X2=0 $Y2=0
cc_1059 N_A_1725_329#_M1011_d N_VPWR_c_1803_n 0.002435f $X=10.35 $Y=2.065 $X2=0
+ $Y2=0
cc_1060 N_A_1725_329#_c_1552_n N_VPWR_c_1803_n 0.00895167f $X=11.275 $Y=1.99
+ $X2=0 $Y2=0
cc_1061 N_A_1725_329#_c_1564_n N_VPWR_c_1803_n 0.0133267f $X=12.265 $Y=1.77
+ $X2=0 $Y2=0
cc_1062 N_A_1725_329#_c_1574_n N_VPWR_c_1803_n 0.0264464f $X=9.52 $Y=2.292 $X2=0
+ $Y2=0
cc_1063 N_A_1725_329#_c_1567_n N_VPWR_c_1803_n 0.0105634f $X=10.395 $Y=1.98
+ $X2=0 $Y2=0
cc_1064 N_A_1725_329#_c_1665_p N_VPWR_c_1803_n 0.00752885f $X=10.495 $Y=2.285
+ $X2=0 $Y2=0
cc_1065 N_A_1725_329#_c_1568_n N_VPWR_c_1803_n 0.0078048f $X=10.875 $Y=1.98
+ $X2=0 $Y2=0
cc_1066 N_A_1725_329#_c_1569_n N_VPWR_c_1803_n 0.00608385f $X=9.605 $Y=1.98
+ $X2=0 $Y2=0
cc_1067 N_A_1725_329#_c_1570_n N_VPWR_c_1803_n 0.0017435f $X=11.04 $Y=1.69 $X2=0
+ $Y2=0
cc_1068 N_A_1725_329#_c_1574_n N_VPWR_c_1825_n 0.0291057f $X=9.52 $Y=2.292 $X2=0
+ $Y2=0
cc_1069 N_A_1725_329#_c_1574_n A_1841_413# 0.00846189f $X=9.52 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1070 N_A_1725_329#_c_1569_n A_1841_413# 0.00200501f $X=9.605 $Y=1.98
+ $X2=-0.19 $Y2=-0.24
cc_1071 N_A_1725_329#_c_1555_n N_VGND_c_2147_n 0.00383167f $X=11.095 $Y=0.925
+ $X2=0 $Y2=0
cc_1072 N_A_1725_329#_c_1556_n N_VGND_c_2147_n 0.00322049f $X=11.095 $Y=0.765
+ $X2=0 $Y2=0
cc_1073 N_A_1725_329#_c_1575_n N_VGND_c_2147_n 0.0204189f $X=10.45 $Y=0.41 $X2=0
+ $Y2=0
cc_1074 N_A_1725_329#_c_1560_n N_VGND_c_2147_n 0.0134367f $X=11.07 $Y=0.93 $X2=0
+ $Y2=0
cc_1075 N_A_1725_329#_M1032_g N_VGND_c_2148_n 0.0145605f $X=12.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1076 N_A_1725_329#_c_1575_n N_VGND_c_2151_n 0.084725f $X=10.45 $Y=0.41 $X2=0
+ $Y2=0
cc_1077 N_A_1725_329#_M1032_g N_VGND_c_2153_n 0.0046653f $X=12.24 $Y=0.445 $X2=0
+ $Y2=0
cc_1078 N_A_1725_329#_c_1555_n N_VGND_c_2153_n 3.91476e-19 $X=11.095 $Y=0.925
+ $X2=0 $Y2=0
cc_1079 N_A_1725_329#_c_1556_n N_VGND_c_2153_n 0.00585385f $X=11.095 $Y=0.765
+ $X2=0 $Y2=0
cc_1080 N_A_1725_329#_M1007_d N_VGND_c_2157_n 0.00371781f $X=9.165 $Y=0.235
+ $X2=0 $Y2=0
cc_1081 N_A_1725_329#_M1032_g N_VGND_c_2157_n 0.00921786f $X=12.24 $Y=0.445
+ $X2=0 $Y2=0
cc_1082 N_A_1725_329#_c_1555_n N_VGND_c_2157_n 5.20533e-19 $X=11.095 $Y=0.925
+ $X2=0 $Y2=0
cc_1083 N_A_1725_329#_c_1556_n N_VGND_c_2157_n 0.00777067f $X=11.095 $Y=0.765
+ $X2=0 $Y2=0
cc_1084 N_A_1725_329#_c_1575_n N_VGND_c_2157_n 0.0579097f $X=10.45 $Y=0.41 $X2=0
+ $Y2=0
cc_1085 N_A_1725_329#_c_1560_n N_VGND_c_2157_n 0.013916f $X=11.07 $Y=0.93 $X2=0
+ $Y2=0
cc_1086 N_A_1725_329#_c_1575_n A_1955_47# 0.00429931f $X=10.45 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1087 N_A_1725_329#_c_1575_n A_2027_47# 0.00737326f $X=10.45 $Y=0.41 $X2=-0.19
+ $Y2=-0.24
cc_1088 N_A_1725_329#_c_1558_n A_2027_47# 0.00144878f $X=10.55 $Y=0.785
+ $X2=-0.19 $Y2=-0.24
cc_1089 N_A_2381_47#_c_1707_n N_VPWR_c_1809_n 0.00598634f $X=12.79 $Y=1.41 $X2=0
+ $Y2=0
cc_1090 N_A_2381_47#_c_1713_n N_VPWR_c_1809_n 0.0362894f $X=12.03 $Y=1.99 $X2=0
+ $Y2=0
cc_1091 N_A_2381_47#_c_1710_n N_VPWR_c_1809_n 0.00822336f $X=12.66 $Y=1.16 $X2=0
+ $Y2=0
cc_1092 N_A_2381_47#_c_1713_n N_VPWR_c_1812_n 0.0217765f $X=12.03 $Y=1.99 $X2=0
+ $Y2=0
cc_1093 N_A_2381_47#_c_1707_n N_VPWR_c_1818_n 0.00702461f $X=12.79 $Y=1.41 $X2=0
+ $Y2=0
cc_1094 N_A_2381_47#_M1004_s N_VPWR_c_1803_n 0.00217517f $X=11.905 $Y=1.845
+ $X2=0 $Y2=0
cc_1095 N_A_2381_47#_c_1707_n N_VPWR_c_1803_n 0.0135619f $X=12.79 $Y=1.41 $X2=0
+ $Y2=0
cc_1096 N_A_2381_47#_c_1713_n N_VPWR_c_1803_n 0.0128576f $X=12.03 $Y=1.99 $X2=0
+ $Y2=0
cc_1097 N_A_2381_47#_c_1707_n N_Q_c_2130_n 0.015587f $X=12.79 $Y=1.41 $X2=0
+ $Y2=0
cc_1098 N_A_2381_47#_c_1708_n N_Q_c_2130_n 0.0226531f $X=12.815 $Y=0.995 $X2=0
+ $Y2=0
cc_1099 N_A_2381_47#_c_1710_n N_Q_c_2130_n 0.0274885f $X=12.66 $Y=1.16 $X2=0
+ $Y2=0
cc_1100 N_A_2381_47#_c_1707_n N_VGND_c_2148_n 0.00315676f $X=12.79 $Y=1.41 $X2=0
+ $Y2=0
cc_1101 N_A_2381_47#_c_1708_n N_VGND_c_2148_n 0.00506737f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1102 N_A_2381_47#_c_1710_n N_VGND_c_2148_n 0.0151608f $X=12.66 $Y=1.16 $X2=0
+ $Y2=0
cc_1103 N_A_2381_47#_c_1709_n N_VGND_c_2153_n 0.018001f $X=12.03 $Y=0.425 $X2=0
+ $Y2=0
cc_1104 N_A_2381_47#_c_1708_n N_VGND_c_2156_n 0.00585385f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1105 N_A_2381_47#_M1032_s N_VGND_c_2157_n 0.00382897f $X=11.905 $Y=0.235
+ $X2=0 $Y2=0
cc_1106 N_A_2381_47#_c_1708_n N_VGND_c_2157_n 0.0121054f $X=12.815 $Y=0.995
+ $X2=0 $Y2=0
cc_1107 N_A_2381_47#_c_1709_n N_VGND_c_2157_n 0.00993603f $X=12.03 $Y=0.425
+ $X2=0 $Y2=0
cc_1108 N_A_27_369#_c_1758_n N_VPWR_M1008_d 0.00342966f $X=1.055 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_1109 N_A_27_369#_c_1757_n N_VPWR_c_1804_n 0.0205323f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1110 N_A_27_369#_c_1758_n N_VPWR_c_1804_n 0.0187115f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1111 N_A_27_369#_c_1757_n N_VPWR_c_1814_n 0.0180865f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1112 N_A_27_369#_c_1758_n N_VPWR_c_1814_n 0.00206566f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1113 N_A_27_369#_c_1758_n N_VPWR_c_1815_n 0.00290212f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1114 N_A_27_369#_c_1771_n N_VPWR_c_1815_n 0.00991509f $X=1.225 $Y=2.36 $X2=0
+ $Y2=0
cc_1115 N_A_27_369#_c_1760_n N_VPWR_c_1815_n 0.0582047f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1116 N_A_27_369#_M1008_s N_VPWR_c_1803_n 0.00244672f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1117 N_A_27_369#_M1021_d N_VPWR_c_1803_n 0.00217543f $X=1.935 $Y=1.845 $X2=0
+ $Y2=0
cc_1118 N_A_27_369#_c_1757_n N_VPWR_c_1803_n 0.00991202f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1119 N_A_27_369#_c_1758_n N_VPWR_c_1803_n 0.0103345f $X=1.055 $Y=1.935 $X2=0
+ $Y2=0
cc_1120 N_A_27_369#_c_1771_n N_VPWR_c_1803_n 0.00653118f $X=1.225 $Y=2.36 $X2=0
+ $Y2=0
cc_1121 N_A_27_369#_c_1760_n N_VPWR_c_1803_n 0.0364411f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1122 N_A_27_369#_c_1758_n A_211_369# 0.00274315f $X=1.055 $Y=1.935 $X2=-0.19
+ $Y2=1.305
cc_1123 N_A_27_369#_c_1774_n A_211_369# 0.00234118f $X=1.14 $Y=2.255 $X2=-0.19
+ $Y2=1.305
cc_1124 N_A_27_369#_c_1771_n A_211_369# 0.00110197f $X=1.225 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1125 N_A_27_369#_c_1760_n N_A_201_47#_M1036_d 0.0035404f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1126 N_A_27_369#_c_1758_n N_A_201_47#_c_2009_n 0.0151838f $X=1.055 $Y=1.935
+ $X2=0 $Y2=0
cc_1127 N_A_27_369#_c_1774_n N_A_201_47#_c_2009_n 0.00444947f $X=1.14 $Y=2.255
+ $X2=0 $Y2=0
cc_1128 N_A_27_369#_c_1760_n N_A_201_47#_c_2009_n 0.0229871f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1129 N_A_27_369#_c_1760_n N_A_201_47#_c_2002_n 0.00286705f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1130 N_VPWR_c_1803_n A_211_369# 0.00184693f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1131 N_VPWR_c_1803_n N_A_201_47#_M1036_d 0.00232895f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1132 N_VPWR_c_1803_n N_A_201_47#_M1006_s 0.0020949f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1133 N_VPWR_c_1816_n N_A_201_47#_c_2000_n 0.0135499f $X=6.445 $Y=2.72 $X2=0
+ $Y2=0
cc_1134 N_VPWR_c_1803_n N_A_201_47#_c_2000_n 0.00390749f $X=13.11 $Y=2.72 $X2=0
+ $Y2=0
cc_1135 N_VPWR_c_1805_n N_A_201_47#_c_2001_n 0.00826221f $X=3.07 $Y=2.34 $X2=0
+ $Y2=0
cc_1136 N_VPWR_c_1803_n A_1169_413# 0.00263276f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1137 N_VPWR_c_1825_n A_1643_329# 0.00116125f $X=8.625 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1138 N_VPWR_c_1803_n A_1841_413# 0.00329526f $X=13.11 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1139 N_VPWR_c_1803_n N_Q_M1035_d 0.00339514f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1140 N_VPWR_c_1818_n N_Q_c_2130_n 0.0201751f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1141 N_VPWR_c_1803_n N_Q_c_2130_n 0.0123504f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_1142 N_A_201_47#_c_2006_n N_VGND_c_2141_n 0.0541179f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1143 N_A_201_47#_c_2006_n N_VGND_c_2142_n 0.0294921f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1144 N_A_201_47#_c_2006_n N_VGND_c_2143_n 0.0224969f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1145 N_A_201_47#_c_1995_n N_VGND_c_2155_n 0.0226408f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1146 N_A_201_47#_M1030_d N_VGND_c_2157_n 0.00255381f $X=1.005 $Y=0.235 $X2=0
+ $Y2=0
cc_1147 N_A_201_47#_M1026_s N_VGND_c_2157_n 0.0054218f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_1148 N_A_201_47#_c_2006_n N_VGND_c_2157_n 0.0334433f $X=1.655 $Y=0.425 $X2=0
+ $Y2=0
cc_1149 N_A_201_47#_c_1995_n N_VGND_c_2157_n 0.0123998f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1150 N_A_201_47#_c_2006_n A_295_47# 0.00393714f $X=1.655 $Y=0.425 $X2=-0.19
+ $Y2=-0.24
cc_1151 N_A_201_47#_c_1997_n A_295_47# 6.98288e-19 $X=1.76 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1152 N_Q_c_2130_n N_VGND_c_2156_n 0.0192978f $X=13.025 $Y=0.44 $X2=0 $Y2=0
cc_1153 N_Q_M1002_d N_VGND_c_2157_n 0.00301111f $X=12.89 $Y=0.235 $X2=0 $Y2=0
cc_1154 N_Q_c_2130_n N_VGND_c_2157_n 0.0123198f $X=13.025 $Y=0.44 $X2=0 $Y2=0
cc_1155 N_VGND_c_2142_n A_119_47# 0.00411471f $X=0.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1156 N_VGND_c_2157_n A_119_47# 0.00142631f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1157 N_VGND_c_2157_n A_295_47# 0.00216824f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1158 N_VGND_c_2155_n A_1177_47# 0.00329703f $X=6.06 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1159 N_VGND_c_2157_n A_1177_47# 0.00735224f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1160 N_VGND_c_2157_n A_1645_47# 0.0141841f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1161 N_VGND_c_2161_n A_1645_47# 0.0115658f $X=8.315 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1162 N_VGND_c_2157_n A_1955_47# 0.00169327f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1163 N_VGND_c_2157_n A_2027_47# 0.00306387f $X=13.11 $Y=0 $X2=-0.19 $Y2=-0.24
