* NGSPICE file created from sky130_fd_sc_hdll__or4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or4_2 A B C D VGND VNB VPB VPWR X
M1000 a_27_297# D VGND VNB nshort w=420000u l=150000u
+  ad=2.94e+11p pd=3.08e+06u as=6.666e+11p ps=6.83e+06u
M1001 VGND A a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=3.4775e+11p pd=2.37e+06u as=0p ps=0u
M1003 a_117_297# D a_27_297# VPB phighvt w=420000u l=180000u
+  ad=1.47e+11p pd=1.54e+06u as=1.134e+11p ps=1.38e+06u
M1004 VPWR A a_305_297# VPB phighvt w=420000u l=180000u
+  ad=6.257e+11p pd=5.35e+06u as=1.47e+11p ps=1.54e+06u
M1005 a_27_297# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND C a_27_297# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_27_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=4.55e+11p ps=2.91e+06u
M1008 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_223_297# C a_117_297# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1011 a_305_297# B a_223_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

