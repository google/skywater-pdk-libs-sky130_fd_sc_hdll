* File: sky130_fd_sc_hdll__o211a_4.spice
* Created: Wed Sep  2 08:42:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o211a_4.pex.spice"
.subckt sky130_fd_sc_hdll__o211a_4  VNB VPB B1 C1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* C1	C1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1009 N_X_M1009_d N_A_80_21#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.17225 PD=0.97 PS=1.83 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1009_d N_A_80_21#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1021 N_X_M1021_d N_A_80_21#_M1021_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=7.38 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1022 N_X_M1021_d N_A_80_21#_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.221 PD=0.97 PS=1.98 NRD=0 NRS=7.38 M=1 R=4.33333 SA=75001.6
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1008 A_818_47# N_B1_M1008_g N_A_524_47#_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.17225 PD=0.86 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1023 N_A_80_21#_M1023_d N_C1_M1023_g A_818_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.177125 AS=0.06825 PD=1.195 PS=0.86 NRD=12.912 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75003.3 A=0.0975 P=1.6 MULT=1
MM1019 N_A_80_21#_M1023_d N_C1_M1019_g A_607_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.177125 AS=0.076375 PD=1.195 PS=0.885 NRD=36 NRS=11.532 M=1 R=4.33333
+ SA=75001.2 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1015 A_607_47# N_B1_M1015_g N_A_524_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.076375 AS=0.105625 PD=0.885 PS=0.975 NRD=11.532 NRS=4.608 M=1 R=4.33333
+ SA=75001.6 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_524_47#_M1015_s N_A1_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.105625 AS=0.12675 PD=0.975 PS=1.04 NRD=3.684 NRS=7.38 M=1 R=4.33333
+ SA=75002.1 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1000 N_A_524_47#_M1000_d N_A2_M1000_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.12675 PD=0.98 PS=1.04 NRD=9.228 NRS=12.912 M=1 R=4.33333
+ SA=75002.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1003 N_A_524_47#_M1000_d N_A2_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75003.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1016 N_A_524_47#_M1016_d N_A1_M1016_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.10725 PD=1.93 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 N_VPWR_M1005_d N_A_80_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.33 AS=0.15 PD=2.66 PS=1.3 NRD=2.9353 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90005.6 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_80_21#_M1010_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90000.7
+ SB=90005.2 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1010_d N_A_80_21#_M1012_g N_X_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=2.9353 NRS=0.9653 M=1 R=5.55556 SA=90001.2
+ SB=90004.7 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A_80_21#_M1017_g N_X_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1475 AS=0.15 PD=1.295 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556
+ SA=90001.7 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_80_21#_M1001_d N_B1_M1001_g N_VPWR_M1017_d VPB PHIGHVT L=0.18 W=1
+ AD=0.2375 AS=0.1475 PD=1.475 PS=1.295 NRD=21.67 NRS=1.9503 M=1 R=5.55556
+ SA=90002.2 SB=90003.7 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_C1_M1004_g N_A_80_21#_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.2375 PD=1.3 PS=1.475 NRD=1.9503 NRS=16.7253 M=1 R=5.55556
+ SA=90002.8 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1004_d N_C1_M1014_g N_A_80_21#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1575 PD=1.3 PS=1.315 NRD=1.9503 NRS=5.8903 M=1 R=5.55556
+ SA=90003.3 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1002 N_A_80_21#_M1014_s N_B1_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1575 AS=0.1475 PD=1.315 PS=1.295 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90003.8 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1002_s N_A1_M1018_g A_1010_297# VPB PHIGHVT L=0.18 W=1 AD=0.1475
+ AS=0.15 PD=1.295 PS=1.3 NRD=0.9653 NRS=18.6953 M=1 R=5.55556 SA=90004.3
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 A_1010_297# N_A2_M1006_g N_A_80_21#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=18.6953 NRS=1.9503 M=1 R=5.55556 SA=90004.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1020 A_1202_297# N_A2_M1020_g N_A_80_21#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=18.6953 NRS=1.9503 M=1 R=5.55556 SA=90005.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A1_M1011_g A_1202_297# VPB PHIGHVT L=0.18 W=1 AD=0.275
+ AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=18.6953 M=1 R=5.55556 SA=90005.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=11.6844 P=17.77
c_694 A_1010_297# 0 1.15076e-19 $X=5.05 $Y=1.485
*
.include "sky130_fd_sc_hdll__o211a_4.pxi.spice"
*
.ends
*
*
