* File: sky130_fd_sc_hdll__o221ai_2.pex.spice
* Created: Thu Aug 27 19:20:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%C1 1 3 4 6 7 9 10 12 13 20
r43 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.97 $Y=1.202
+ $X2=0.995 $Y2=1.202
r44 19 20 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.525 $Y=1.202
+ $X2=0.97 $Y2=1.202
r45 18 19 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.5 $Y=1.202
+ $X2=0.525 $Y2=1.202
r46 16 18 30.3726 $w=3.65e-07 $l=2.3e-07 $layer=POLY_cond $X=0.27 $Y=1.202
+ $X2=0.5 $Y2=1.202
r47 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r48 10 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=0.56
r50 7 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.97 $Y=1.41
+ $X2=0.97 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.97 $Y=1.41 $X2=0.97
+ $Y2=1.985
r52 4 19 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=1.202
r53 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.56
r54 1 18 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.202
r55 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%B1 1 3 4 6 7 9 10 12 13 15 19 21 26 31
c77 10 0 1.91072e-19 $X=3.395 $Y=0.995
r78 26 31 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=1.6 $Y=1.345 $X2=1.57
+ $Y2=1.345
r79 21 24 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.37 $Y=1.16
+ $X2=3.37 $Y2=1.53
r80 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.345
+ $Y=1.16 $X2=3.345 $Y2=1.16
r81 17 19 11.6507 $w=5.38e-07 $l=2.5e-07 $layer=LI1_cond $X=1.935 $Y=1.345
+ $X2=2.185 $Y2=1.345
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.935
+ $Y=1.16 $X2=1.935 $Y2=1.16
r83 15 26 6.97712 $w=5.38e-07 $l=3.15e-07 $layer=LI1_cond $X=1.915 $Y=1.345
+ $X2=1.6 $Y2=1.345
r84 15 17 0.442992 $w=5.38e-07 $l=2e-08 $layer=LI1_cond $X=1.915 $Y=1.345
+ $X2=1.935 $Y2=1.345
r85 13 24 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.18 $Y=1.53 $X2=3.37
+ $Y2=1.53
r86 13 19 64.9144 $w=1.68e-07 $l=9.95e-07 $layer=LI1_cond $X=3.18 $Y=1.53
+ $X2=2.185 $Y2=1.53
r87 10 22 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.395 $Y=0.995
+ $X2=3.37 $Y2=1.16
r88 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.395 $Y=0.995
+ $X2=3.395 $Y2=0.56
r89 7 22 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.37 $Y=1.41
+ $X2=3.37 $Y2=1.16
r90 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.37 $Y=1.41 $X2=3.37
+ $Y2=1.985
r91 4 18 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.96 $Y2=1.16
r92 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.985 $Y=0.995
+ $X2=1.985 $Y2=0.56
r93 1 18 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.16
r94 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.96 $Y=1.41 $X2=1.96
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%B2 1 3 4 6 7 9 10 12 13 19 20 25
r43 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.9 $Y=1.202
+ $X2=2.925 $Y2=1.202
r44 19 25 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.665 $Y=1.175
+ $X2=2.55 $Y2=1.175
r45 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.665 $Y=1.202
+ $X2=2.9 $Y2=1.202
r46 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.665
+ $Y=1.16 $X2=2.665 $Y2=1.16
r47 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=2.43 $Y=1.202
+ $X2=2.665 $Y2=1.202
r48 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.43 $Y2=1.202
r49 13 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=2.535 $Y=1.175
+ $X2=2.55 $Y2=1.175
r50 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.925 $Y=0.995
+ $X2=2.925 $Y2=1.202
r51 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.925 $Y=0.995
+ $X2=2.925 $Y2=0.56
r52 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.9 $Y=1.41 $X2=2.9
+ $Y2=1.202
r53 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.9 $Y=1.41 $X2=2.9
+ $Y2=1.985
r54 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.202
r55 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.41 $X2=2.43
+ $Y2=1.985
r56 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.405 $Y=0.995
+ $X2=2.405 $Y2=1.202
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.405 $Y=0.995
+ $X2=2.405 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A1 1 3 4 6 7 9 10 12 13 16 18 23 24 31
c73 7 0 3.32201e-19 $X=5.33 $Y=1.41
c74 4 0 2.98731e-20 $X=3.945 $Y=0.995
r75 28 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.305
+ $Y=1.16 $X2=5.305 $Y2=1.16
r76 24 31 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=5.705 $Y=1.175
+ $X2=5.29 $Y2=1.175
r77 23 31 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.265 $Y=1.175
+ $X2=5.29 $Y2=1.175
r78 18 21 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.92 $Y=1.16
+ $X2=3.92 $Y2=1.53
r79 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.895
+ $Y=1.16 $X2=3.895 $Y2=1.16
r80 15 23 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.18 $Y=1.275
+ $X2=5.265 $Y2=1.175
r81 15 16 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.18 $Y=1.275
+ $X2=5.18 $Y2=1.445
r82 14 21 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.11 $Y=1.53 $X2=3.92
+ $Y2=1.53
r83 13 16 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.095 $Y=1.53
+ $X2=5.18 $Y2=1.445
r84 13 14 64.262 $w=1.68e-07 $l=9.85e-07 $layer=LI1_cond $X=5.095 $Y=1.53
+ $X2=4.11 $Y2=1.53
r85 10 28 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.33 $Y2=1.16
r86 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.355 $Y=0.995
+ $X2=5.355 $Y2=0.56
r87 7 28 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.33 $Y=1.41
+ $X2=5.33 $Y2=1.16
r88 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.33 $Y=1.41 $X2=5.33
+ $Y2=1.985
r89 4 19 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.92 $Y2=1.16
r90 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=0.56
r91 1 19 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.92 $Y=1.41
+ $X2=3.92 $Y2=1.16
r92 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.92 $Y=1.41 $X2=3.92
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A2 1 3 4 6 7 9 10 12 13 20 25
c47 13 0 1.89398e-19 $X=4.705 $Y=1.105
r48 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=4.885 $Y2=1.202
r49 19 25 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=4.625 $Y=1.175
+ $X2=4.745 $Y2=1.175
r50 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.625 $Y=1.202
+ $X2=4.86 $Y2=1.202
r51 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.625
+ $Y=1.16 $X2=4.625 $Y2=1.16
r52 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.39 $Y=1.202
+ $X2=4.625 $Y2=1.202
r53 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.365 $Y=1.202
+ $X2=4.39 $Y2=1.202
r54 13 25 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=4.79 $Y=1.175
+ $X2=4.745 $Y2=1.175
r55 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.885 $Y=0.995
+ $X2=4.885 $Y2=1.202
r56 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.885 $Y=0.995
+ $X2=4.885 $Y2=0.56
r57 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.202
r58 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.86 $Y=1.41 $X2=4.86
+ $Y2=1.985
r59 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.39 $Y=1.41
+ $X2=4.39 $Y2=1.202
r60 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.39 $Y=1.41 $X2=4.39
+ $Y2=1.985
r61 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.365 $Y2=1.202
r62 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.365 $Y=0.995
+ $X2=4.365 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%VPWR 1 2 3 4 13 15 23 27 32 33 35 36 37
+ 53 54 62 68
r73 67 68 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=1.725 $Y=2.465
+ $X2=1.85 $Y2=2.465
r74 64 67 2.02278 $w=6.78e-07 $l=1.15e-07 $layer=LI1_cond $X=1.61 $Y=2.465
+ $X2=1.725 $Y2=2.465
r75 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 61 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 60 64 8.09112 $w=6.78e-07 $l=4.6e-07 $layer=LI1_cond $X=1.15 $Y=2.465
+ $X2=1.61 $Y2=2.465
r78 60 62 9.00537 $w=6.78e-07 $l=7e-08 $layer=LI1_cond $X=1.15 $Y=2.465 $X2=1.08
+ $Y2=2.465
r79 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r80 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r81 51 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r82 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r83 48 51 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r84 47 50 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r85 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r86 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r87 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r88 42 45 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r89 42 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r90 41 44 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r91 41 68 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=1.85 $Y2=2.72
r92 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 37 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r94 37 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 35 50 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.29 $Y2=2.72
r96 35 36 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.485 $Y=2.72
+ $X2=5.587 $Y2=2.72
r97 34 53 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=2.72 $X2=5.75
+ $Y2=2.72
r98 34 36 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=5.69 $Y=2.72
+ $X2=5.587 $Y2=2.72
r99 32 44 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.48 $Y=2.72 $X2=3.45
+ $Y2=2.72
r100 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.48 $Y=2.72
+ $X2=3.645 $Y2=2.72
r101 31 47 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.81 $Y=2.72 $X2=3.91
+ $Y2=2.72
r102 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.81 $Y=2.72
+ $X2=3.645 $Y2=2.72
r103 27 30 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=5.587 $Y=1.62
+ $X2=5.587 $Y2=2.3
r104 25 36 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.587 $Y=2.635
+ $X2=5.587 $Y2=2.72
r105 25 30 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=5.587 $Y=2.635
+ $X2=5.587 $Y2=2.3
r106 21 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.645 $Y=2.635
+ $X2=3.645 $Y2=2.72
r107 21 23 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.645 $Y=2.635
+ $X2=3.645 $Y2=2.3
r108 20 57 3.97976 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r109 20 62 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=1.08 $Y2=2.72
r110 15 18 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.265 $Y=1.65
+ $X2=0.265 $Y2=2.33
r111 13 57 3.1634 $w=2.5e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.195 $Y2=2.72
r112 13 18 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.33
r113 4 30 400 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.485 $X2=5.57 $Y2=2.3
r114 4 27 400 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.485 $X2=5.57 $Y2=1.62
r115 3 23 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.46
+ $Y=1.485 $X2=3.605 $Y2=2.3
r116 2 67 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.485 $X2=1.725 $Y2=2.3
r117 1 18 400 $w=1.7e-07 $l=9.05345e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=2.33
r118 1 15 400 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=1 $X=0.14
+ $Y=1.485 $X2=0.265 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%Y 1 2 3 4 13 16 19 23 28 30 32 33 34 39
+ 44 48
r65 44 48 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=1.61 $Y=1.87 $X2=1.63
+ $Y2=1.87
r66 39 42 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.625 $Y=1.87
+ $X2=4.625 $Y2=1.96
r67 34 48 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=2.54 $Y=1.87 $X2=1.63
+ $Y2=1.87
r68 33 37 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=2.665 $Y=1.87
+ $X2=2.665 $Y2=1.96
r69 33 34 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.665 $Y=1.87
+ $X2=2.54 $Y2=1.87
r70 31 44 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.9 $Y=1.87 $X2=1.61
+ $Y2=1.87
r71 31 32 3.05049 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.9 $Y=1.87
+ $X2=0.755 $Y2=1.87
r72 26 28 2.20012 $w=2.18e-07 $l=4.2e-08 $layer=LI1_cond $X=0.735 $Y=0.755
+ $X2=0.777 $Y2=0.755
r73 24 33 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.79 $Y=1.87
+ $X2=2.665 $Y2=1.87
r74 23 39 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.5 $Y=1.87
+ $X2=4.625 $Y2=1.87
r75 23 24 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=4.5 $Y=1.87
+ $X2=2.79 $Y2=1.87
r76 21 28 0.0766963 $w=2.45e-07 $l=1.1e-07 $layer=LI1_cond $X=0.777 $Y=0.865
+ $X2=0.777 $Y2=0.755
r77 21 30 27.2823 $w=2.43e-07 $l=5.8e-07 $layer=LI1_cond $X=0.777 $Y=0.865
+ $X2=0.777 $Y2=1.445
r78 17 32 3.46198 $w=2.7e-07 $l=9.44722e-08 $layer=LI1_cond $X=0.735 $Y=1.955
+ $X2=0.755 $Y2=1.87
r79 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.735 $Y=1.955
+ $X2=0.735 $Y2=1.96
r80 14 32 3.46198 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.755 $Y2=1.87
r81 14 16 6.557 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.755 $Y=1.785
+ $X2=0.755 $Y2=1.62
r82 13 30 6.07313 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=0.755 $Y=1.59
+ $X2=0.755 $Y2=1.445
r83 13 16 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=0.755 $Y=1.59
+ $X2=0.755 $Y2=1.62
r84 4 42 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.485 $X2=4.625 $Y2=1.96
r85 3 37 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.485 $X2=2.665 $Y2=1.96
r86 2 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.735 $Y2=1.96
r87 2 16 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.485 $X2=0.735 $Y2=1.62
r88 1 26 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.735 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A_410_297# 1 2 7 10 15
r22 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.135 $Y=2.3 $X2=3.135
+ $Y2=2.38
r23 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=2.195 $Y=2.3 $X2=2.195
+ $Y2=2.38
r24 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.32 $Y=2.38
+ $X2=2.195 $Y2=2.38
r25 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.01 $Y=2.38
+ $X2=3.135 $Y2=2.38
r26 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.01 $Y=2.38 $X2=2.32
+ $Y2=2.38
r27 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.485 $X2=3.135 $Y2=2.3
r28 1 10 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.485 $X2=2.195 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A_802_297# 1 2 7 11 14
c17 11 0 1.42804e-19 $X=5.095 $Y=1.96
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.155 $Y=2.3 $X2=4.155
+ $Y2=2.38
r19 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.095 $Y=2.295
+ $X2=5.095 $Y2=1.96
r20 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.28 $Y=2.38
+ $X2=4.155 $Y2=2.38
r21 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.97 $Y=2.38
+ $X2=5.095 $Y2=2.295
r22 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.97 $Y=2.38 $X2=4.28
+ $Y2=2.38
r23 2 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.485 $X2=5.095 $Y2=1.96
r24 1 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.485 $X2=4.155 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A_28_47# 1 2 3 4 13 15 17 19 20 25
c49 25 0 1.91072e-19 $X=3.135 $Y=0.73
r50 23 25 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=2.195 $Y=0.775
+ $X2=3.135 $Y2=0.775
r51 21 32 3.34309 $w=2.6e-07 $l=1.25e-07 $layer=LI1_cond $X=1.37 $Y=0.775
+ $X2=1.245 $Y2=0.775
r52 21 23 36.5679 $w=2.58e-07 $l=8.25e-07 $layer=LI1_cond $X=1.37 $Y=0.775
+ $X2=2.195 $Y2=0.775
r53 20 32 3.47681 $w=2.5e-07 $l=1.3e-07 $layer=LI1_cond $X=1.245 $Y=0.645
+ $X2=1.245 $Y2=0.775
r54 19 30 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.245 $Y=0.475
+ $X2=1.245 $Y2=0.365
r55 19 20 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=1.245 $Y=0.475
+ $X2=1.245 $Y2=0.645
r56 18 28 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=0.35 $Y=0.365
+ $X2=0.225 $Y2=0.365
r57 17 30 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.12 $Y=0.365
+ $X2=1.245 $Y2=0.365
r58 17 18 40.3355 $w=2.18e-07 $l=7.7e-07 $layer=LI1_cond $X=1.12 $Y=0.365
+ $X2=0.35 $Y2=0.365
r59 13 28 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=0.225 $Y=0.475
+ $X2=0.225 $Y2=0.365
r60 13 15 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.225 $Y=0.475
+ $X2=0.225 $Y2=0.73
r61 4 25 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3
+ $Y=0.235 $X2=3.135 $Y2=0.73
r62 3 23 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.06
+ $Y=0.235 $X2=2.195 $Y2=0.73
r63 2 32 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.205 $Y2=0.73
r64 2 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.205 $Y2=0.39
r65 1 28 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.39
r66 1 15 182 $w=1.7e-07 $l=5.53986e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%A_320_47# 1 2 3 4 5 16 22 26 27 30 32 36
+ 40
c68 40 0 2.98731e-20 $X=4.6 $Y=0.815
r69 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.54 $Y=0.725
+ $X2=5.54 $Y2=0.39
r70 33 40 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=4.79 $Y=0.815
+ $X2=4.6 $Y2=0.815
r71 32 34 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.35 $Y=0.815
+ $X2=5.54 $Y2=0.725
r72 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.35 $Y=0.815
+ $X2=4.79 $Y2=0.815
r73 28 40 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.6 $Y=0.725 $X2=4.6
+ $Y2=0.815
r74 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.6 $Y=0.725
+ $X2=4.6 $Y2=0.39
r75 26 40 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=4.41 $Y=0.82
+ $X2=4.6 $Y2=0.815
r76 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.41 $Y=0.82
+ $X2=3.85 $Y2=0.82
r77 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.685 $Y=0.735
+ $X2=3.85 $Y2=0.82
r78 23 25 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.685 $Y=0.735
+ $X2=3.685 $Y2=0.73
r79 22 39 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=3.685 $Y=0.475
+ $X2=3.685 $Y2=0.365
r80 22 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3.685 $Y=0.475
+ $X2=3.685 $Y2=0.73
r81 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=1.725 $Y=0.365
+ $X2=2.665 $Y2=0.365
r82 16 39 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=3.685 $Y2=0.365
r83 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=2.665 $Y2=0.365
r84 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.43
+ $Y=0.235 $X2=5.565 $Y2=0.39
r85 4 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.44
+ $Y=0.235 $X2=4.625 $Y2=0.39
r86 3 39 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.235 $X2=3.65 $Y2=0.39
r87 3 25 182 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_NDIFF $count=1 $X=3.47
+ $Y=0.235 $X2=3.65 $Y2=0.73
r88 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.665 $Y2=0.39
r89 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.6
+ $Y=0.235 $X2=1.725 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O221AI_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r70 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r71 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r72 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r73 28 29 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r74 24 28 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r75 21 29 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=3.91
+ $Y2=0
r76 21 24 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r77 19 31 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=5.01 $Y=0 $X2=4.83
+ $Y2=0
r78 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.01 $Y=0 $X2=5.095
+ $Y2=0
r79 18 34 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=5.18 $Y=0 $X2=5.75
+ $Y2=0
r80 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=0 $X2=5.095
+ $Y2=0
r81 16 28 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.07 $Y=0 $X2=3.91
+ $Y2=0
r82 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=0 $X2=4.155
+ $Y2=0
r83 15 31 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.83
+ $Y2=0
r84 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.155
+ $Y2=0
r85 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0
r86 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.095 $Y=0.085
+ $X2=5.095 $Y2=0.39
r87 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=0.085
+ $X2=4.155 $Y2=0
r88 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.155 $Y=0.085
+ $X2=4.155 $Y2=0.39
r89 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.96
+ $Y=0.235 $X2=5.095 $Y2=0.39
r90 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.155 $Y2=0.39
.ends

