* File: sky130_fd_sc_hdll__sdlclkp_1.pxi.spice
* Created: Wed Sep  2 08:52:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%SCE N_SCE_c_142_n N_SCE_c_143_n N_SCE_M1005_g
+ N_SCE_M1015_g SCE SCE N_SCE_c_141_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%SCE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GATE N_GATE_c_171_n N_GATE_c_172_n
+ N_GATE_M1003_g N_GATE_M1021_g GATE GATE N_GATE_c_169_n N_GATE_c_170_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GATE
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_269_21# N_A_269_21#_M1007_d
+ N_A_269_21#_M1002_d N_A_269_21#_M1014_g N_A_269_21#_c_220_n
+ N_A_269_21#_M1009_g N_A_269_21#_M1019_g N_A_269_21#_c_210_n
+ N_A_269_21#_M1020_g N_A_269_21#_c_211_n N_A_269_21#_c_212_n
+ N_A_269_21#_c_213_n N_A_269_21#_c_223_n N_A_269_21#_c_214_n
+ N_A_269_21#_c_215_n N_A_269_21#_c_216_n N_A_269_21#_c_224_n
+ N_A_269_21#_c_217_n N_A_269_21#_c_218_n N_A_269_21#_c_219_n
+ N_A_269_21#_c_226_n N_A_269_21#_c_235_n N_A_269_21#_c_227_n
+ N_A_269_21#_c_228_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_269_21#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_266_243# N_A_266_243#_M1019_s
+ N_A_266_243#_M1020_s N_A_266_243#_c_394_n N_A_266_243#_c_395_n
+ N_A_266_243#_M1017_g N_A_266_243#_c_382_n N_A_266_243#_c_383_n
+ N_A_266_243#_M1006_g N_A_266_243#_c_384_n N_A_266_243#_c_385_n
+ N_A_266_243#_c_386_n N_A_266_243#_c_399_n N_A_266_243#_c_387_n
+ N_A_266_243#_c_388_n N_A_266_243#_c_389_n N_A_266_243#_c_390_n
+ N_A_266_243#_c_391_n N_A_266_243#_c_392_n N_A_266_243#_c_393_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_266_243#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_484_315# N_A_484_315#_M1004_d
+ N_A_484_315#_M1000_d N_A_484_315#_c_503_n N_A_484_315#_M1010_g
+ N_A_484_315#_M1011_g N_A_484_315#_c_505_n N_A_484_315#_c_506_n
+ N_A_484_315#_M1001_g N_A_484_315#_M1008_g N_A_484_315#_c_507_n
+ N_A_484_315#_c_519_n N_A_484_315#_c_500_n N_A_484_315#_c_509_n
+ N_A_484_315#_c_501_n N_A_484_315#_c_530_n N_A_484_315#_c_531_n
+ N_A_484_315#_c_502_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_484_315#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_299_47# N_A_299_47#_M1014_d
+ N_A_299_47#_M1017_d N_A_299_47#_c_628_n N_A_299_47#_M1000_g
+ N_A_299_47#_c_629_n N_A_299_47#_M1004_g N_A_299_47#_c_642_n
+ N_A_299_47#_c_646_n N_A_299_47#_c_636_n N_A_299_47#_c_630_n
+ N_A_299_47#_c_631_n N_A_299_47#_c_632_n N_A_299_47#_c_633_n
+ N_A_299_47#_c_634_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_299_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%CLK N_CLK_M1007_g N_CLK_c_731_n N_CLK_M1002_g
+ N_CLK_c_740_n N_CLK_c_741_n N_CLK_M1016_g N_CLK_M1013_g N_CLK_c_733_n
+ N_CLK_c_761_n N_CLK_c_734_n N_CLK_c_735_n CLK N_CLK_c_736_n N_CLK_c_737_n CLK
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_1%CLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_1089_47# N_A_1089_47#_M1008_s
+ N_A_1089_47#_M1001_d N_A_1089_47#_c_825_n N_A_1089_47#_M1012_g
+ N_A_1089_47#_c_826_n N_A_1089_47#_M1018_g N_A_1089_47#_c_833_n
+ N_A_1089_47#_c_827_n N_A_1089_47#_c_828_n N_A_1089_47#_c_840_n
+ N_A_1089_47#_c_829_n N_A_1089_47#_c_832_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_1089_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VPWR N_VPWR_M1005_s N_VPWR_M1010_d
+ N_VPWR_M1020_d N_VPWR_M1001_s N_VPWR_M1016_d N_VPWR_c_900_n N_VPWR_c_901_n
+ N_VPWR_c_902_n N_VPWR_c_903_n N_VPWR_c_904_n N_VPWR_c_905_n N_VPWR_c_906_n
+ VPWR N_VPWR_c_907_n N_VPWR_c_908_n N_VPWR_c_899_n N_VPWR_c_910_n
+ N_VPWR_c_911_n N_VPWR_c_912_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VPWR
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_27_47# N_A_27_47#_M1015_s N_A_27_47#_M1021_d
+ N_A_27_47#_M1003_d N_A_27_47#_c_996_n N_A_27_47#_c_997_n N_A_27_47#_c_998_n
+ N_A_27_47#_c_999_n N_A_27_47#_c_1009_n N_A_27_47#_c_1018_n N_A_27_47#_c_1022_n
+ PM_SKY130_FD_SC_HDLL__SDLCLKP_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GCLK N_GCLK_M1018_d N_GCLK_M1012_d GCLK GCLK
+ GCLK GCLK PM_SKY130_FD_SC_HDLL__SDLCLKP_1%GCLK
x_PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VGND N_VGND_M1015_d N_VGND_M1011_d
+ N_VGND_M1019_d N_VGND_M1013_d N_VGND_c_1066_n N_VGND_c_1067_n N_VGND_c_1068_n
+ N_VGND_c_1069_n VGND N_VGND_c_1070_n N_VGND_c_1071_n N_VGND_c_1072_n
+ N_VGND_c_1073_n N_VGND_c_1074_n N_VGND_c_1075_n N_VGND_c_1076_n
+ N_VGND_c_1077_n PM_SKY130_FD_SC_HDLL__SDLCLKP_1%VGND
cc_1 VNB N_SCE_M1015_g 0.035163f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB SCE 0.0151026f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_SCE_c_141_n 0.0371984f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_GATE_M1021_g 0.0275553f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_GATE_c_169_n 0.0265721f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_GATE_c_170_n 0.00513867f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_7 VNB N_A_269_21#_M1014_g 0.0199099f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_269_21#_M1019_g 0.0350075f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_9 VNB N_A_269_21#_c_210_n 0.0291982f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_10 VNB N_A_269_21#_c_211_n 0.00753371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_269_21#_c_212_n 0.0299387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_269_21#_c_213_n 0.00330504f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_269_21#_c_214_n 0.00421076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_269_21#_c_215_n 0.011506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_269_21#_c_216_n 0.00165799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_269_21#_c_217_n 0.00409988f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_269_21#_c_218_n 0.00224307f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_269_21#_c_219_n 8.70148e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_266_243#_c_382_n 0.0157472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_266_243#_c_383_n 0.00701797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_266_243#_c_384_n 0.012193f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_22 VNB N_A_266_243#_c_385_n 0.00850373f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_23 VNB N_A_266_243#_c_386_n 0.00765412f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_24 VNB N_A_266_243#_c_387_n 0.0101381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_266_243#_c_388_n 0.00127289f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_266_243#_c_389_n 0.00124593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_266_243#_c_390_n 0.00542601f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_266_243#_c_391_n 0.025854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_266_243#_c_392_n 0.00326317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_266_243#_c_393_n 0.019636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_484_315#_M1011_g 0.045987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_484_315#_M1008_g 0.0389156f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_33 VNB N_A_484_315#_c_500_n 0.0083999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_484_315#_c_501_n 0.0101946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_484_315#_c_502_n 0.0319981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_299_47#_c_628_n 0.0279771f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_37 VNB N_A_299_47#_c_629_n 0.0210956f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_38 VNB N_A_299_47#_c_630_n 0.0023264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_299_47#_c_631_n 0.00229294f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_40 VNB N_A_299_47#_c_632_n 0.00188091f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_299_47#_c_633_n 0.00258328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_299_47#_c_634_n 0.00219952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_CLK_M1007_g 0.0405534f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.77
cc_44 VNB N_CLK_c_731_n 0.0277121f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_45 VNB N_CLK_M1013_g 0.0295754f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_46 VNB N_CLK_c_733_n 0.0165208f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_47 VNB N_CLK_c_734_n 8.13421e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_CLK_c_735_n 0.00535835f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_CLK_c_736_n 0.0182493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_CLK_c_737_n 0.00228925f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_1089_47#_c_825_n 0.0271303f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_52 VNB N_A_1089_47#_c_826_n 0.0196888f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_53 VNB N_A_1089_47#_c_827_n 0.00524678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1089_47#_c_828_n 0.0024418f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_55 VNB N_A_1089_47#_c_829_n 0.00113231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VPWR_c_899_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_27_47#_c_996_n 0.0141581f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_27_47#_c_997_n 0.00395907f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_59 VNB N_A_27_47#_c_998_n 0.0105678f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_60 VNB N_A_27_47#_c_999_n 0.0108603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB GCLK 0.0451979f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_62 VNB N_VGND_c_1066_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_63 VNB N_VGND_c_1067_n 0.00562936f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_64 VNB N_VGND_c_1068_n 0.0083383f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.16
cc_65 VNB N_VGND_c_1069_n 0.0449122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_1070_n 0.0142754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_1071_n 0.048839f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_1072_n 0.0336157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1073_n 0.0207195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_1074_n 0.367396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_VGND_c_1075_n 0.00556536f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_VGND_c_1076_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_VGND_c_1077_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VPB N_SCE_c_142_n 0.0182203f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_75 VPB N_SCE_c_143_n 0.0288642f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_76 VPB SCE 0.0186881f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_77 VPB N_SCE_c_141_n 0.0111298f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_78 VPB N_GATE_c_171_n 0.0179893f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.67
cc_79 VPB N_GATE_c_172_n 0.0218835f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_80 VPB N_GATE_c_169_n 0.00419201f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_81 VPB N_GATE_c_170_n 0.00393713f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_82 VPB N_A_269_21#_c_220_n 0.0517349f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_83 VPB N_A_269_21#_c_210_n 0.013615f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_84 VPB N_A_269_21#_M1020_g 0.0428907f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.16
cc_85 VPB N_A_269_21#_c_223_n 0.0035611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_269_21#_c_224_n 0.0102358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_269_21#_c_218_n 6.69987e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_269_21#_c_226_n 0.017224f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_269_21#_c_227_n 0.00417665f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_269_21#_c_228_n 0.00330281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_266_243#_c_394_n 0.0310551f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_92 VPB N_A_266_243#_c_395_n 0.0241018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_A_266_243#_c_382_n 0.0175257f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_A_266_243#_c_383_n 0.00247433f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_266_243#_c_386_n 0.00481438f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_96 VPB N_A_266_243#_c_399_n 0.00295943f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_484_315#_c_503_n 0.0570583f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_98 VPB N_A_484_315#_M1011_g 0.0168089f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_A_484_315#_c_505_n 0.0236659f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_100 VPB N_A_484_315#_c_506_n 0.0267616f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_101 VPB N_A_484_315#_c_507_n 0.00246621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_484_315#_c_500_n 0.00372381f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_484_315#_c_509_n 0.0181402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_484_315#_c_501_n 0.0085137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_484_315#_c_502_n 0.00814611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_299_47#_c_628_n 0.0320723f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_107 VPB N_A_299_47#_c_636_n 0.0132653f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_A_299_47#_c_630_n 0.00162406f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_A_299_47#_c_631_n 8.46875e-19 $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_110 VPB N_A_299_47#_c_633_n 0.00331303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_A_299_47#_c_634_n 5.36217e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_CLK_c_731_n 0.0138105f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_113 VPB N_CLK_M1002_g 0.0446644f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_114 VPB N_CLK_c_740_n 0.0190768f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_115 VPB N_CLK_c_741_n 0.0217757f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_116 VPB N_CLK_c_734_n 5.58243e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_CLK_c_735_n 0.00183387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_CLK_c_736_n 0.00265165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_A_1089_47#_c_825_n 0.0295703f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_120 VPB N_A_1089_47#_c_829_n 0.001647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_1089_47#_c_832_n 0.00714727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_VPWR_c_900_n 0.0098838f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_123 VPB N_VPWR_c_901_n 0.0319853f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_124 VPB N_VPWR_c_902_n 0.00506198f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_125 VPB N_VPWR_c_903_n 0.0314135f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_VPWR_c_904_n 0.00468864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_VPWR_c_905_n 0.0168195f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_VPWR_c_906_n 0.00631443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_VPWR_c_907_n 0.0111737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_VPWR_c_908_n 0.0198621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_VPWR_c_899_n 0.0488527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_VPWR_c_910_n 0.0540052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_VPWR_c_911_n 0.0135649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_VPWR_c_912_n 0.0201646f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_27_47#_c_997_n 0.00318143f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_136 VPB GCLK 0.0461283f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_137 N_SCE_c_142_n N_GATE_c_171_n 0.0156312f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_138 N_SCE_c_143_n N_GATE_c_172_n 0.0632861f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_139 N_SCE_M1015_g N_GATE_M1021_g 0.025321f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_140 N_SCE_c_141_n N_GATE_c_169_n 0.0156312f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_141 N_SCE_c_141_n N_GATE_c_170_n 7.45308e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_142 N_SCE_c_143_n N_VPWR_c_901_n 0.00695514f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_143 SCE N_VPWR_c_901_n 0.0228425f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_144 N_SCE_c_141_n N_VPWR_c_901_n 0.0013127f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_145 N_SCE_c_143_n N_VPWR_c_899_n 0.0107787f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_146 N_SCE_c_143_n N_VPWR_c_910_n 0.00596194f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_147 N_SCE_c_142_n N_A_27_47#_c_997_n 0.00689877f $X=0.495 $Y=1.67 $X2=0 $Y2=0
cc_148 N_SCE_c_143_n N_A_27_47#_c_997_n 0.0139589f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_149 N_SCE_M1015_g N_A_27_47#_c_997_n 0.00963306f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_150 SCE N_A_27_47#_c_997_n 0.0477147f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_151 N_SCE_c_141_n N_A_27_47#_c_997_n 0.00850344f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_152 N_SCE_M1015_g N_A_27_47#_c_999_n 0.0136308f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_153 SCE N_A_27_47#_c_999_n 0.020595f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_154 N_SCE_c_141_n N_A_27_47#_c_999_n 0.00574324f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_155 N_SCE_c_143_n N_A_27_47#_c_1009_n 0.00888327f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_156 N_SCE_M1015_g N_VGND_c_1070_n 0.00196986f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_157 N_SCE_M1015_g N_VGND_c_1074_n 0.00356708f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_158 N_SCE_M1015_g N_VGND_c_1075_n 0.0109522f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_159 N_GATE_M1021_g N_A_269_21#_M1014_g 0.0193371f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_160 N_GATE_M1021_g N_A_269_21#_c_211_n 9.10923e-19 $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_161 N_GATE_c_169_n N_A_269_21#_c_211_n 0.00114135f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_GATE_c_170_n N_A_269_21#_c_211_n 0.0641903f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_163 N_GATE_c_169_n N_A_269_21#_c_212_n 5.40897e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_164 N_GATE_c_170_n N_A_269_21#_c_212_n 4.46444e-19 $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_GATE_c_170_n N_A_269_21#_c_235_n 0.00143054f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_166 N_GATE_c_172_n N_A_269_21#_c_227_n 3.10662e-19 $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_167 N_GATE_c_172_n N_A_266_243#_c_394_n 0.0147937f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_168 N_GATE_c_172_n N_A_266_243#_c_395_n 0.0162305f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_169 N_GATE_c_171_n N_A_266_243#_c_383_n 0.00747498f $X=0.905 $Y=1.67 $X2=0
+ $Y2=0
cc_170 N_GATE_c_169_n N_A_266_243#_c_383_n 0.0067961f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_GATE_c_170_n N_A_266_243#_c_383_n 0.00653544f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_172 N_GATE_c_172_n N_VPWR_c_899_n 0.00613085f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_173 N_GATE_c_172_n N_VPWR_c_910_n 0.00429453f $X=0.905 $Y=1.77 $X2=0 $Y2=0
cc_174 N_GATE_c_170_n N_A_27_47#_M1003_d 0.00332039f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_175 N_GATE_c_172_n N_A_27_47#_c_997_n 0.00461756f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_176 N_GATE_M1021_g N_A_27_47#_c_997_n 0.00356352f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_177 N_GATE_c_169_n N_A_27_47#_c_997_n 0.00432932f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_178 N_GATE_c_170_n N_A_27_47#_c_997_n 0.0758785f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_179 N_GATE_M1021_g N_A_27_47#_c_998_n 0.0113083f $X=0.945 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_GATE_c_169_n N_A_27_47#_c_998_n 0.00268203f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_181 N_GATE_c_170_n N_A_27_47#_c_998_n 0.0315401f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_182 N_GATE_c_172_n N_A_27_47#_c_1018_n 0.0184335f $X=0.905 $Y=1.77 $X2=0
+ $Y2=0
cc_183 N_GATE_c_170_n N_A_27_47#_c_1018_n 0.0257572f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_184 N_GATE_M1021_g N_VGND_c_1071_n 0.0035176f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_185 N_GATE_M1021_g N_VGND_c_1074_n 0.00420343f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_186 N_GATE_M1021_g N_VGND_c_1075_n 0.00759201f $X=0.945 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_269_21#_c_220_n N_A_266_243#_c_394_n 0.0213218f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_188 N_A_269_21#_c_218_n N_A_266_243#_c_394_n 0.00322667f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_189 N_A_269_21#_c_227_n N_A_266_243#_c_394_n 0.0123339f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_190 N_A_269_21#_c_220_n N_A_266_243#_c_395_n 0.0123925f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_191 N_A_269_21#_c_227_n N_A_266_243#_c_395_n 0.00342606f $X=1.71 $Y=1.53
+ $X2=0 $Y2=0
cc_192 N_A_269_21#_c_220_n N_A_266_243#_c_382_n 0.021863f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_193 N_A_269_21#_c_218_n N_A_266_243#_c_382_n 0.019479f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_194 N_A_269_21#_c_226_n N_A_266_243#_c_382_n 0.00280811f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_195 N_A_269_21#_c_212_n N_A_266_243#_c_383_n 0.0262024f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_196 N_A_269_21#_c_218_n N_A_266_243#_c_383_n 0.0029158f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_197 N_A_269_21#_c_218_n N_A_266_243#_c_384_n 0.00135637f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_198 N_A_269_21#_M1019_g N_A_266_243#_c_385_n 0.00725487f $X=4.19 $Y=0.445
+ $X2=0 $Y2=0
cc_199 N_A_269_21#_c_216_n N_A_266_243#_c_385_n 0.00807489f $X=4.55 $Y=0.7 $X2=0
+ $Y2=0
cc_200 N_A_269_21#_M1019_g N_A_266_243#_c_386_n 0.00393841f $X=4.19 $Y=0.445
+ $X2=0 $Y2=0
cc_201 N_A_269_21#_c_210_n N_A_266_243#_c_386_n 0.0048599f $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_202 N_A_269_21#_M1020_g N_A_266_243#_c_386_n 0.00152654f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_203 N_A_269_21#_c_213_n N_A_266_243#_c_386_n 0.0137757f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_204 N_A_269_21#_c_223_n N_A_266_243#_c_386_n 0.00887327f $X=4.457 $Y=1.495
+ $X2=0 $Y2=0
cc_205 N_A_269_21#_c_214_n N_A_266_243#_c_386_n 0.00537229f $X=4.465 $Y=1.105
+ $X2=0 $Y2=0
cc_206 N_A_269_21#_c_226_n N_A_266_243#_c_386_n 0.0102301f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_207 N_A_269_21#_c_228_n N_A_266_243#_c_386_n 9.52575e-19 $X=4.45 $Y=1.53
+ $X2=0 $Y2=0
cc_208 N_A_269_21#_c_210_n N_A_266_243#_c_399_n 2.6841e-19 $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_209 N_A_269_21#_M1020_g N_A_266_243#_c_399_n 0.00239927f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_210 N_A_269_21#_c_213_n N_A_266_243#_c_399_n 0.00188351f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_211 N_A_269_21#_c_223_n N_A_266_243#_c_399_n 0.0103461f $X=4.457 $Y=1.495
+ $X2=0 $Y2=0
cc_212 N_A_269_21#_c_226_n N_A_266_243#_c_399_n 0.00994167f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_213 N_A_269_21#_c_228_n N_A_266_243#_c_399_n 0.0011663f $X=4.45 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_269_21#_c_226_n N_A_266_243#_c_387_n 0.0623626f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_215 N_A_269_21#_c_211_n N_A_266_243#_c_388_n 0.00137702f $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_216 N_A_269_21#_c_226_n N_A_266_243#_c_388_n 0.0131578f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_217 N_A_269_21#_M1019_g N_A_266_243#_c_389_n 7.51712e-19 $X=4.19 $Y=0.445
+ $X2=0 $Y2=0
cc_218 N_A_269_21#_c_214_n N_A_266_243#_c_389_n 0.00175981f $X=4.465 $Y=1.105
+ $X2=0 $Y2=0
cc_219 N_A_269_21#_c_216_n N_A_266_243#_c_389_n 3.81144e-19 $X=4.55 $Y=0.7 $X2=0
+ $Y2=0
cc_220 N_A_269_21#_c_226_n N_A_266_243#_c_389_n 0.013701f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_221 N_A_269_21#_c_214_n N_A_266_243#_c_390_n 0.00656646f $X=4.465 $Y=1.105
+ $X2=0 $Y2=0
cc_222 N_A_269_21#_c_226_n N_A_266_243#_c_390_n 0.00134723f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_223 N_A_269_21#_c_211_n N_A_266_243#_c_391_n 0.00731088f $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_224 N_A_269_21#_c_212_n N_A_266_243#_c_391_n 0.0165461f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_225 N_A_269_21#_c_220_n N_A_266_243#_c_392_n 2.78293e-19 $X=1.96 $Y=1.99
+ $X2=0 $Y2=0
cc_226 N_A_269_21#_c_211_n N_A_266_243#_c_392_n 0.0247397f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_227 N_A_269_21#_c_212_n N_A_266_243#_c_392_n 2.64542e-19 $X=1.55 $Y=0.87
+ $X2=0 $Y2=0
cc_228 N_A_269_21#_c_226_n N_A_266_243#_c_392_n 0.00523969f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_229 N_A_269_21#_M1014_g N_A_266_243#_c_393_n 0.0132713f $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_230 N_A_269_21#_c_226_n N_A_484_315#_M1000_d 8.06277e-19 $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_231 N_A_269_21#_c_220_n N_A_484_315#_c_503_n 0.0289443f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_232 N_A_269_21#_c_226_n N_A_484_315#_c_503_n 0.00449033f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_233 N_A_269_21#_c_226_n N_A_484_315#_M1011_g 0.00420735f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_234 N_A_269_21#_c_224_n N_A_484_315#_c_505_n 9.98965e-19 $X=5.05 $Y=1.66
+ $X2=0 $Y2=0
cc_235 N_A_269_21#_c_215_n N_A_484_315#_M1008_g 7.46752e-19 $X=4.965 $Y=0.7
+ $X2=0 $Y2=0
cc_236 N_A_269_21#_c_226_n N_A_484_315#_c_507_n 0.0222174f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_237 N_A_269_21#_M1020_g N_A_484_315#_c_519_n 0.00487772f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_238 N_A_269_21#_c_226_n N_A_484_315#_c_500_n 0.022258f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_239 N_A_269_21#_M1002_d N_A_484_315#_c_509_n 0.00518929f $X=4.905 $Y=1.515
+ $X2=0 $Y2=0
cc_240 N_A_269_21#_c_210_n N_A_484_315#_c_509_n 9.1318e-19 $X=4.215 $Y=1.44
+ $X2=0 $Y2=0
cc_241 N_A_269_21#_M1020_g N_A_484_315#_c_509_n 0.0164643f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_242 N_A_269_21#_c_213_n N_A_484_315#_c_509_n 0.00166026f $X=4.365 $Y=1.19
+ $X2=0 $Y2=0
cc_243 N_A_269_21#_c_223_n N_A_484_315#_c_509_n 0.0140488f $X=4.457 $Y=1.495
+ $X2=0 $Y2=0
cc_244 N_A_269_21#_c_224_n N_A_484_315#_c_509_n 0.0397345f $X=5.05 $Y=1.66 $X2=0
+ $Y2=0
cc_245 N_A_269_21#_c_226_n N_A_484_315#_c_509_n 0.013136f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_246 N_A_269_21#_c_228_n N_A_484_315#_c_509_n 0.00314908f $X=4.45 $Y=1.53
+ $X2=0 $Y2=0
cc_247 N_A_269_21#_c_224_n N_A_484_315#_c_501_n 0.0220307f $X=5.05 $Y=1.66 $X2=0
+ $Y2=0
cc_248 N_A_269_21#_c_226_n N_A_484_315#_c_530_n 0.007409f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_249 N_A_269_21#_M1020_g N_A_484_315#_c_531_n 0.00335363f $X=4.215 $Y=1.835
+ $X2=0 $Y2=0
cc_250 N_A_269_21#_c_226_n N_A_484_315#_c_531_n 0.00302634f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_251 N_A_269_21#_c_226_n N_A_299_47#_c_628_n 0.0085668f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_252 N_A_269_21#_M1014_g N_A_299_47#_c_642_n 0.00807723f $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_253 N_A_269_21#_c_211_n N_A_299_47#_c_642_n 0.0249565f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_254 N_A_269_21#_c_212_n N_A_299_47#_c_642_n 0.00135285f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_255 N_A_269_21#_c_218_n N_A_299_47#_c_642_n 0.00401633f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_256 N_A_269_21#_c_220_n N_A_299_47#_c_646_n 0.0152026f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_257 N_A_269_21#_c_226_n N_A_299_47#_c_646_n 0.00562701f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_258 N_A_269_21#_c_235_n N_A_299_47#_c_646_n 0.00102774f $X=1.855 $Y=1.53
+ $X2=0 $Y2=0
cc_259 N_A_269_21#_c_227_n N_A_299_47#_c_646_n 0.0255421f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_260 N_A_269_21#_c_220_n N_A_299_47#_c_636_n 0.0073981f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_261 N_A_269_21#_c_218_n N_A_299_47#_c_636_n 0.0438627f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_262 N_A_269_21#_c_226_n N_A_299_47#_c_636_n 0.0204925f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_263 N_A_269_21#_c_235_n N_A_299_47#_c_636_n 5.16817e-19 $X=1.855 $Y=1.53
+ $X2=0 $Y2=0
cc_264 N_A_269_21#_c_226_n N_A_299_47#_c_630_n 0.005814f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_265 N_A_269_21#_c_218_n N_A_299_47#_c_631_n 0.0147478f $X=1.712 $Y=1.452
+ $X2=0 $Y2=0
cc_266 N_A_269_21#_c_226_n N_A_299_47#_c_633_n 0.00800313f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_267 N_A_269_21#_c_211_n N_A_299_47#_c_634_n 0.00566979f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_268 N_A_269_21#_c_226_n N_A_299_47#_c_634_n 0.00229606f $X=4.305 $Y=1.53
+ $X2=0 $Y2=0
cc_269 N_A_269_21#_M1019_g N_CLK_M1007_g 0.0157264f $X=4.19 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A_269_21#_c_214_n N_CLK_M1007_g 0.00542813f $X=4.465 $Y=1.105 $X2=0
+ $Y2=0
cc_271 N_A_269_21#_c_215_n N_CLK_M1007_g 0.0138617f $X=4.965 $Y=0.7 $X2=0 $Y2=0
cc_272 N_A_269_21#_c_217_n N_CLK_M1007_g 0.0047281f $X=5.05 $Y=0.465 $X2=0 $Y2=0
cc_273 N_A_269_21#_c_210_n N_CLK_c_731_n 0.017606f $X=4.215 $Y=1.44 $X2=0 $Y2=0
cc_274 N_A_269_21#_c_223_n N_CLK_c_731_n 0.00285076f $X=4.457 $Y=1.495 $X2=0
+ $Y2=0
cc_275 N_A_269_21#_c_215_n N_CLK_c_731_n 0.00449177f $X=4.965 $Y=0.7 $X2=0 $Y2=0
cc_276 N_A_269_21#_c_224_n N_CLK_c_731_n 0.00404517f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_277 N_A_269_21#_c_219_n N_CLK_c_731_n 0.00121068f $X=4.457 $Y=1.19 $X2=0
+ $Y2=0
cc_278 N_A_269_21#_c_228_n N_CLK_c_731_n 4.22826e-19 $X=4.45 $Y=1.53 $X2=0 $Y2=0
cc_279 N_A_269_21#_M1020_g N_CLK_M1002_g 0.0345833f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_280 N_A_269_21#_c_223_n N_CLK_M1002_g 0.00100311f $X=4.457 $Y=1.495 $X2=0
+ $Y2=0
cc_281 N_A_269_21#_c_224_n N_CLK_M1002_g 0.0136189f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_282 N_A_269_21#_c_228_n N_CLK_M1002_g 0.00109498f $X=4.45 $Y=1.53 $X2=0 $Y2=0
cc_283 N_A_269_21#_c_215_n N_CLK_c_733_n 0.00691214f $X=4.965 $Y=0.7 $X2=0 $Y2=0
cc_284 N_A_269_21#_c_224_n N_CLK_c_733_n 0.00702604f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_285 N_A_269_21#_c_223_n N_CLK_c_761_n 2.20902e-19 $X=4.457 $Y=1.495 $X2=0
+ $Y2=0
cc_286 N_A_269_21#_c_214_n N_CLK_c_761_n 2.19371e-19 $X=4.465 $Y=1.105 $X2=0
+ $Y2=0
cc_287 N_A_269_21#_c_215_n N_CLK_c_761_n 0.0017699f $X=4.965 $Y=0.7 $X2=0 $Y2=0
cc_288 N_A_269_21#_c_224_n N_CLK_c_761_n 0.00208449f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_289 N_A_269_21#_c_219_n N_CLK_c_761_n 0.00134698f $X=4.457 $Y=1.19 $X2=0
+ $Y2=0
cc_290 N_A_269_21#_c_210_n N_CLK_c_737_n 4.61377e-19 $X=4.215 $Y=1.44 $X2=0
+ $Y2=0
cc_291 N_A_269_21#_c_223_n N_CLK_c_737_n 0.0029265f $X=4.457 $Y=1.495 $X2=0
+ $Y2=0
cc_292 N_A_269_21#_c_214_n N_CLK_c_737_n 0.00697859f $X=4.465 $Y=1.105 $X2=0
+ $Y2=0
cc_293 N_A_269_21#_c_215_n N_CLK_c_737_n 0.0182322f $X=4.965 $Y=0.7 $X2=0 $Y2=0
cc_294 N_A_269_21#_c_224_n N_CLK_c_737_n 0.0216073f $X=5.05 $Y=1.66 $X2=0 $Y2=0
cc_295 N_A_269_21#_c_219_n N_CLK_c_737_n 0.0101522f $X=4.457 $Y=1.19 $X2=0 $Y2=0
cc_296 N_A_269_21#_c_217_n N_A_1089_47#_c_833_n 0.0174382f $X=5.05 $Y=0.465
+ $X2=0 $Y2=0
cc_297 N_A_269_21#_c_215_n N_A_1089_47#_c_828_n 0.0101606f $X=4.965 $Y=0.7 $X2=0
+ $Y2=0
cc_298 N_A_269_21#_c_226_n N_VPWR_M1010_d 0.00203938f $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_299 N_A_269_21#_c_223_n N_VPWR_M1020_d 0.00627377f $X=4.457 $Y=1.495 $X2=0
+ $Y2=0
cc_300 N_A_269_21#_c_224_n N_VPWR_M1020_d 0.00126167f $X=5.05 $Y=1.66 $X2=0
+ $Y2=0
cc_301 N_A_269_21#_c_228_n N_VPWR_M1020_d 5.5836e-19 $X=4.45 $Y=1.53 $X2=0 $Y2=0
cc_302 N_A_269_21#_M1020_g N_VPWR_c_903_n 0.0156985f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_303 N_A_269_21#_M1020_g N_VPWR_c_907_n 0.00974554f $X=4.215 $Y=1.835 $X2=0
+ $Y2=0
cc_304 N_A_269_21#_c_220_n N_VPWR_c_899_n 0.00645844f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_305 N_A_269_21#_c_227_n N_VPWR_c_899_n 0.00621311f $X=1.71 $Y=1.53 $X2=0
+ $Y2=0
cc_306 N_A_269_21#_c_220_n N_VPWR_c_910_n 0.00429453f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_307 N_A_269_21#_c_220_n N_VPWR_c_911_n 0.00138786f $X=1.96 $Y=1.99 $X2=0
+ $Y2=0
cc_308 N_A_269_21#_c_226_n N_VPWR_c_911_n 6.32368e-19 $X=4.305 $Y=1.53 $X2=0
+ $Y2=0
cc_309 N_A_269_21#_M1014_g N_A_27_47#_c_998_n 0.0036696f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_310 N_A_269_21#_c_211_n N_A_27_47#_c_998_n 0.00671481f $X=1.55 $Y=0.87 $X2=0
+ $Y2=0
cc_311 N_A_269_21#_M1014_g N_A_27_47#_c_1022_n 4.57344e-19 $X=1.42 $Y=0.415
+ $X2=0 $Y2=0
cc_312 N_A_269_21#_c_215_n N_VGND_M1019_d 0.00137428f $X=4.965 $Y=0.7 $X2=0
+ $Y2=0
cc_313 N_A_269_21#_c_216_n N_VGND_M1019_d 0.00258762f $X=4.55 $Y=0.7 $X2=0 $Y2=0
cc_314 N_A_269_21#_M1019_g N_VGND_c_1067_n 0.00332046f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_315 N_A_269_21#_c_210_n N_VGND_c_1067_n 0.0018575f $X=4.215 $Y=1.44 $X2=0
+ $Y2=0
cc_316 N_A_269_21#_c_213_n N_VGND_c_1067_n 0.00152098f $X=4.365 $Y=1.19 $X2=0
+ $Y2=0
cc_317 N_A_269_21#_c_215_n N_VGND_c_1067_n 0.00481916f $X=4.965 $Y=0.7 $X2=0
+ $Y2=0
cc_318 N_A_269_21#_c_216_n N_VGND_c_1067_n 0.0142335f $X=4.55 $Y=0.7 $X2=0 $Y2=0
cc_319 N_A_269_21#_c_217_n N_VGND_c_1067_n 0.00877137f $X=5.05 $Y=0.465 $X2=0
+ $Y2=0
cc_320 N_A_269_21#_c_219_n N_VGND_c_1067_n 4.34631e-19 $X=4.457 $Y=1.19 $X2=0
+ $Y2=0
cc_321 N_A_269_21#_c_215_n N_VGND_c_1069_n 0.00529754f $X=4.965 $Y=0.7 $X2=0
+ $Y2=0
cc_322 N_A_269_21#_c_217_n N_VGND_c_1069_n 0.017177f $X=5.05 $Y=0.465 $X2=0
+ $Y2=0
cc_323 N_A_269_21#_M1014_g N_VGND_c_1071_n 0.00539883f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_324 N_A_269_21#_M1019_g N_VGND_c_1072_n 0.00585385f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_325 N_A_269_21#_M1007_d N_VGND_c_1074_n 0.00283928f $X=4.865 $Y=0.235 $X2=0
+ $Y2=0
cc_326 N_A_269_21#_M1014_g N_VGND_c_1074_n 0.0101587f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_327 N_A_269_21#_M1019_g N_VGND_c_1074_n 0.0123217f $X=4.19 $Y=0.445 $X2=0
+ $Y2=0
cc_328 N_A_269_21#_c_215_n N_VGND_c_1074_n 0.0096407f $X=4.965 $Y=0.7 $X2=0
+ $Y2=0
cc_329 N_A_269_21#_c_216_n N_VGND_c_1074_n 8.89004e-19 $X=4.55 $Y=0.7 $X2=0
+ $Y2=0
cc_330 N_A_269_21#_c_217_n N_VGND_c_1074_n 0.00948959f $X=5.05 $Y=0.465 $X2=0
+ $Y2=0
cc_331 N_A_269_21#_M1014_g N_VGND_c_1075_n 0.00108095f $X=1.42 $Y=0.415 $X2=0
+ $Y2=0
cc_332 N_A_266_243#_c_387_n N_A_484_315#_M1004_d 0.00127746f $X=3.74 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_333 N_A_266_243#_c_384_n N_A_484_315#_M1011_g 0.00699103f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_334 N_A_266_243#_c_387_n N_A_484_315#_M1011_g 0.00341307f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_335 N_A_266_243#_c_391_n N_A_484_315#_M1011_g 0.00969942f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_336 N_A_266_243#_c_392_n N_A_484_315#_M1011_g 8.23951e-19 $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_337 N_A_266_243#_c_393_n N_A_484_315#_M1011_g 0.0121621f $X=2.06 $Y=0.705
+ $X2=0 $Y2=0
cc_338 N_A_266_243#_c_385_n N_A_484_315#_c_500_n 0.0907185f $X=3.98 $Y=0.465
+ $X2=0 $Y2=0
cc_339 N_A_266_243#_c_399_n N_A_484_315#_c_500_n 0.00406408f $X=3.98 $Y=1.66
+ $X2=0 $Y2=0
cc_340 N_A_266_243#_c_387_n N_A_484_315#_c_500_n 0.0175797f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_341 N_A_266_243#_c_389_n N_A_484_315#_c_500_n 6.53653e-19 $X=3.885 $Y=0.85
+ $X2=0 $Y2=0
cc_342 N_A_266_243#_M1020_s N_A_484_315#_c_509_n 0.00535544f $X=3.855 $Y=1.515
+ $X2=0 $Y2=0
cc_343 N_A_266_243#_c_399_n N_A_484_315#_c_509_n 0.024093f $X=3.98 $Y=1.66 $X2=0
+ $Y2=0
cc_344 N_A_266_243#_c_399_n N_A_484_315#_c_531_n 0.00889198f $X=3.98 $Y=1.66
+ $X2=0 $Y2=0
cc_345 N_A_266_243#_c_399_n N_A_299_47#_c_628_n 5.9685e-19 $X=3.98 $Y=1.66 $X2=0
+ $Y2=0
cc_346 N_A_266_243#_c_387_n N_A_299_47#_c_628_n 0.00370099f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_347 N_A_266_243#_c_387_n N_A_299_47#_c_629_n 0.00861904f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_348 N_A_266_243#_c_383_n N_A_299_47#_c_642_n 7.38226e-19 $X=1.53 $Y=1.29
+ $X2=0 $Y2=0
cc_349 N_A_266_243#_c_387_n N_A_299_47#_c_642_n 0.00173979f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_350 N_A_266_243#_c_388_n N_A_299_47#_c_642_n 0.00205588f $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_351 N_A_266_243#_c_391_n N_A_299_47#_c_642_n 0.00273817f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_352 N_A_266_243#_c_392_n N_A_299_47#_c_642_n 0.0213864f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_353 N_A_266_243#_c_393_n N_A_299_47#_c_642_n 0.0130546f $X=2.06 $Y=0.705
+ $X2=0 $Y2=0
cc_354 N_A_266_243#_c_394_n N_A_299_47#_c_636_n 6.38369e-19 $X=1.43 $Y=1.89
+ $X2=0 $Y2=0
cc_355 N_A_266_243#_c_387_n N_A_299_47#_c_630_n 0.00153861f $X=3.74 $Y=0.85
+ $X2=0 $Y2=0
cc_356 N_A_266_243#_c_388_n N_A_299_47#_c_630_n 9.40357e-19 $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_357 N_A_266_243#_c_392_n N_A_299_47#_c_630_n 3.1525e-19 $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_358 N_A_266_243#_c_384_n N_A_299_47#_c_631_n 0.00225667f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_359 N_A_266_243#_c_388_n N_A_299_47#_c_631_n 7.66293e-19 $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_360 N_A_266_243#_c_391_n N_A_299_47#_c_631_n 0.00151422f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_361 N_A_266_243#_c_392_n N_A_299_47#_c_631_n 0.0128773f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_362 N_A_266_243#_c_387_n N_A_299_47#_c_632_n 0.0164716f $X=3.74 $Y=0.85 $X2=0
+ $Y2=0
cc_363 N_A_266_243#_c_388_n N_A_299_47#_c_632_n 0.00275249f $X=2.365 $Y=0.85
+ $X2=0 $Y2=0
cc_364 N_A_266_243#_c_391_n N_A_299_47#_c_632_n 6.88042e-19 $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_365 N_A_266_243#_c_392_n N_A_299_47#_c_632_n 0.020669f $X=2.06 $Y=0.87 $X2=0
+ $Y2=0
cc_366 N_A_266_243#_c_393_n N_A_299_47#_c_632_n 0.00291704f $X=2.06 $Y=0.705
+ $X2=0 $Y2=0
cc_367 N_A_266_243#_c_387_n N_A_299_47#_c_633_n 0.016448f $X=3.74 $Y=0.85 $X2=0
+ $Y2=0
cc_368 N_A_266_243#_c_384_n N_A_299_47#_c_634_n 0.00188395f $X=2.022 $Y=1.215
+ $X2=0 $Y2=0
cc_369 N_A_266_243#_c_392_n N_A_299_47#_c_634_n 0.00346908f $X=2.06 $Y=0.87
+ $X2=0 $Y2=0
cc_370 N_A_266_243#_c_395_n N_VPWR_c_899_n 0.0118046f $X=1.43 $Y=1.99 $X2=0
+ $Y2=0
cc_371 N_A_266_243#_c_395_n N_VPWR_c_910_n 0.00743866f $X=1.43 $Y=1.99 $X2=0
+ $Y2=0
cc_372 N_A_266_243#_c_387_n N_VGND_M1011_d 0.00222845f $X=3.74 $Y=0.85 $X2=0
+ $Y2=0
cc_373 N_A_266_243#_c_387_n N_VGND_c_1066_n 0.00775574f $X=3.74 $Y=0.85 $X2=0
+ $Y2=0
cc_374 N_A_266_243#_c_393_n N_VGND_c_1071_n 0.00357877f $X=2.06 $Y=0.705 $X2=0
+ $Y2=0
cc_375 N_A_266_243#_c_385_n N_VGND_c_1072_n 0.0230197f $X=3.98 $Y=0.465 $X2=0
+ $Y2=0
cc_376 N_A_266_243#_M1019_s N_VGND_c_1074_n 0.00358181f $X=3.855 $Y=0.235 $X2=0
+ $Y2=0
cc_377 N_A_266_243#_c_385_n N_VGND_c_1074_n 0.00645346f $X=3.98 $Y=0.465 $X2=0
+ $Y2=0
cc_378 N_A_266_243#_c_387_n N_VGND_c_1074_n 0.0668138f $X=3.74 $Y=0.85 $X2=0
+ $Y2=0
cc_379 N_A_266_243#_c_388_n N_VGND_c_1074_n 0.0148704f $X=2.365 $Y=0.85 $X2=0
+ $Y2=0
cc_380 N_A_266_243#_c_389_n N_VGND_c_1074_n 0.0146243f $X=3.885 $Y=0.85 $X2=0
+ $Y2=0
cc_381 N_A_266_243#_c_393_n N_VGND_c_1074_n 0.00611524f $X=2.06 $Y=0.705 $X2=0
+ $Y2=0
cc_382 N_A_484_315#_c_503_n N_A_299_47#_c_628_n 0.0141627f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_383 N_A_484_315#_M1011_g N_A_299_47#_c_628_n 0.033994f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_384 N_A_484_315#_c_507_n N_A_299_47#_c_628_n 0.0217841f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_385 N_A_484_315#_c_500_n N_A_299_47#_c_628_n 0.0079676f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_386 N_A_484_315#_c_530_n N_A_299_47#_c_628_n 3.54096e-19 $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_387 N_A_484_315#_M1011_g N_A_299_47#_c_629_n 0.0160518f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_388 N_A_484_315#_c_500_n N_A_299_47#_c_629_n 0.0207844f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_389 N_A_484_315#_M1011_g N_A_299_47#_c_642_n 0.00982828f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_390 N_A_484_315#_c_503_n N_A_299_47#_c_646_n 0.00307829f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_391 N_A_484_315#_c_503_n N_A_299_47#_c_636_n 0.00690356f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_392 N_A_484_315#_M1011_g N_A_299_47#_c_636_n 0.00512785f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_393 N_A_484_315#_c_530_n N_A_299_47#_c_636_n 0.0255996f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_394 N_A_484_315#_c_503_n N_A_299_47#_c_630_n 0.00169011f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_395 N_A_484_315#_c_530_n N_A_299_47#_c_630_n 2.34133e-19 $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_396 N_A_484_315#_M1011_g N_A_299_47#_c_632_n 0.0124362f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_397 N_A_484_315#_M1011_g N_A_299_47#_c_633_n 0.00997152f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_398 N_A_484_315#_c_507_n N_A_299_47#_c_633_n 0.0189559f $X=3.325 $Y=1.77
+ $X2=0 $Y2=0
cc_399 N_A_484_315#_c_500_n N_A_299_47#_c_633_n 0.0302043f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_400 N_A_484_315#_c_530_n N_A_299_47#_c_633_n 0.00101123f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_401 N_A_484_315#_c_503_n N_A_299_47#_c_634_n 0.00197841f $X=2.52 $Y=1.99
+ $X2=0 $Y2=0
cc_402 N_A_484_315#_M1011_g N_A_299_47#_c_634_n 0.00804706f $X=2.655 $Y=0.445
+ $X2=0 $Y2=0
cc_403 N_A_484_315#_c_530_n N_A_299_47#_c_634_n 0.00960172f $X=2.665 $Y=1.74
+ $X2=0 $Y2=0
cc_404 N_A_484_315#_c_501_n N_CLK_c_731_n 0.00445883f $X=5.61 $Y=1.16 $X2=0
+ $Y2=0
cc_405 N_A_484_315#_c_502_n N_CLK_c_731_n 0.00872741f $X=5.83 $Y=1.16 $X2=0
+ $Y2=0
cc_406 N_A_484_315#_c_509_n N_CLK_M1002_g 0.0144714f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_407 N_A_484_315#_c_501_n N_CLK_M1002_g 0.00520848f $X=5.61 $Y=1.16 $X2=0
+ $Y2=0
cc_408 N_A_484_315#_c_505_n N_CLK_c_740_n 0.00965828f $X=5.805 $Y=1.67 $X2=0
+ $Y2=0
cc_409 N_A_484_315#_c_501_n N_CLK_c_740_n 9.8199e-19 $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_410 N_A_484_315#_c_506_n N_CLK_c_741_n 0.0271713f $X=5.805 $Y=1.77 $X2=0
+ $Y2=0
cc_411 N_A_484_315#_M1008_g N_CLK_M1013_g 0.0346278f $X=5.83 $Y=0.445 $X2=0
+ $Y2=0
cc_412 N_A_484_315#_c_501_n N_CLK_c_733_n 0.0373194f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_413 N_A_484_315#_c_502_n N_CLK_c_733_n 0.00965113f $X=5.83 $Y=1.16 $X2=0
+ $Y2=0
cc_414 N_A_484_315#_c_501_n N_CLK_c_761_n 6.48982e-19 $X=5.61 $Y=1.16 $X2=0
+ $Y2=0
cc_415 N_A_484_315#_c_501_n N_CLK_c_734_n 0.00253643f $X=5.61 $Y=1.16 $X2=0
+ $Y2=0
cc_416 N_A_484_315#_c_502_n N_CLK_c_734_n 0.00152994f $X=5.83 $Y=1.16 $X2=0
+ $Y2=0
cc_417 N_A_484_315#_c_501_n N_CLK_c_735_n 0.0186286f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_418 N_A_484_315#_c_502_n N_CLK_c_735_n 0.00245494f $X=5.83 $Y=1.16 $X2=0
+ $Y2=0
cc_419 N_A_484_315#_c_501_n N_CLK_c_736_n 3.1611e-19 $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_420 N_A_484_315#_c_502_n N_CLK_c_736_n 0.021501f $X=5.83 $Y=1.16 $X2=0 $Y2=0
cc_421 N_A_484_315#_c_501_n N_CLK_c_737_n 0.0132645f $X=5.61 $Y=1.16 $X2=0 $Y2=0
cc_422 N_A_484_315#_c_502_n N_CLK_c_737_n 4.55837e-19 $X=5.83 $Y=1.16 $X2=0
+ $Y2=0
cc_423 N_A_484_315#_M1008_g N_A_1089_47#_c_827_n 0.0131249f $X=5.83 $Y=0.445
+ $X2=0 $Y2=0
cc_424 N_A_484_315#_c_501_n N_A_1089_47#_c_827_n 0.00177648f $X=5.61 $Y=1.16
+ $X2=0 $Y2=0
cc_425 N_A_484_315#_c_502_n N_A_1089_47#_c_827_n 0.00102546f $X=5.83 $Y=1.16
+ $X2=0 $Y2=0
cc_426 N_A_484_315#_c_501_n N_A_1089_47#_c_828_n 0.0114741f $X=5.61 $Y=1.16
+ $X2=0 $Y2=0
cc_427 N_A_484_315#_c_502_n N_A_1089_47#_c_828_n 0.00127183f $X=5.83 $Y=1.16
+ $X2=0 $Y2=0
cc_428 N_A_484_315#_c_506_n N_A_1089_47#_c_840_n 0.00473478f $X=5.805 $Y=1.77
+ $X2=0 $Y2=0
cc_429 N_A_484_315#_c_505_n N_A_1089_47#_c_832_n 0.00259412f $X=5.805 $Y=1.67
+ $X2=0 $Y2=0
cc_430 N_A_484_315#_c_506_n N_A_1089_47#_c_832_n 0.00224874f $X=5.805 $Y=1.77
+ $X2=0 $Y2=0
cc_431 N_A_484_315#_c_509_n N_A_1089_47#_c_832_n 0.0120899f $X=5.385 $Y=2 $X2=0
+ $Y2=0
cc_432 N_A_484_315#_c_501_n N_A_1089_47#_c_832_n 0.0290204f $X=5.61 $Y=1.16
+ $X2=0 $Y2=0
cc_433 N_A_484_315#_c_507_n N_VPWR_M1010_d 0.00492813f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_434 N_A_484_315#_c_509_n N_VPWR_M1020_d 0.00664869f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_435 N_A_484_315#_c_509_n N_VPWR_M1001_s 0.00310031f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_436 N_A_484_315#_c_501_n N_VPWR_M1001_s 3.05534e-19 $X=5.61 $Y=1.16 $X2=0
+ $Y2=0
cc_437 N_A_484_315#_c_509_n N_VPWR_c_903_n 0.0244473f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_438 N_A_484_315#_c_506_n N_VPWR_c_904_n 0.00854229f $X=5.805 $Y=1.77 $X2=0
+ $Y2=0
cc_439 N_A_484_315#_c_506_n N_VPWR_c_905_n 0.00622633f $X=5.805 $Y=1.77 $X2=0
+ $Y2=0
cc_440 N_A_484_315#_c_519_n N_VPWR_c_907_n 0.0107733f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_441 N_A_484_315#_c_509_n N_VPWR_c_907_n 0.105732f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_442 N_A_484_315#_M1000_d N_VPWR_c_899_n 0.00237624f $X=3.315 $Y=1.485 $X2=0
+ $Y2=0
cc_443 N_A_484_315#_c_503_n N_VPWR_c_899_n 0.00514038f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_444 N_A_484_315#_c_506_n N_VPWR_c_899_n 0.0104813f $X=5.805 $Y=1.77 $X2=0
+ $Y2=0
cc_445 N_A_484_315#_c_507_n N_VPWR_c_899_n 0.00668636f $X=3.325 $Y=1.77 $X2=0
+ $Y2=0
cc_446 N_A_484_315#_c_519_n N_VPWR_c_899_n 0.00839556f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_447 N_A_484_315#_c_509_n N_VPWR_c_899_n 0.0185684f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_448 N_A_484_315#_c_530_n N_VPWR_c_899_n 0.00344844f $X=2.665 $Y=1.74 $X2=0
+ $Y2=0
cc_449 N_A_484_315#_c_503_n N_VPWR_c_910_n 0.00368409f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_450 N_A_484_315#_c_503_n N_VPWR_c_911_n 0.0256563f $X=2.52 $Y=1.99 $X2=0
+ $Y2=0
cc_451 N_A_484_315#_c_530_n N_VPWR_c_911_n 0.0407968f $X=2.665 $Y=1.74 $X2=0
+ $Y2=0
cc_452 N_A_484_315#_c_519_n N_VPWR_c_912_n 0.0137273f $X=3.46 $Y=2.205 $X2=0
+ $Y2=0
cc_453 N_A_484_315#_c_509_n N_VPWR_c_912_n 0.0052614f $X=5.385 $Y=2 $X2=0 $Y2=0
cc_454 N_A_484_315#_M1011_g N_VGND_c_1066_n 0.00720923f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_455 N_A_484_315#_c_500_n N_VGND_c_1066_n 0.0140386f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_456 N_A_484_315#_M1008_g N_VGND_c_1068_n 0.00175127f $X=5.83 $Y=0.445 $X2=0
+ $Y2=0
cc_457 N_A_484_315#_M1008_g N_VGND_c_1069_n 0.00422112f $X=5.83 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_484_315#_M1011_g N_VGND_c_1071_n 0.00486707f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_459 N_A_484_315#_c_500_n N_VGND_c_1072_n 0.0116048f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_460 N_A_484_315#_M1004_d N_VGND_c_1074_n 0.00243215f $X=3.325 $Y=0.235 $X2=0
+ $Y2=0
cc_461 N_A_484_315#_M1011_g N_VGND_c_1074_n 0.0068389f $X=2.655 $Y=0.445 $X2=0
+ $Y2=0
cc_462 N_A_484_315#_M1008_g N_VGND_c_1074_n 0.0073803f $X=5.83 $Y=0.445 $X2=0
+ $Y2=0
cc_463 N_A_484_315#_c_500_n N_VGND_c_1074_n 0.00308197f $X=3.46 $Y=0.42 $X2=0
+ $Y2=0
cc_464 N_A_299_47#_c_628_n N_VPWR_c_907_n 0.00300894f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_465 N_A_299_47#_M1017_d N_VPWR_c_899_n 0.00328896f $X=1.52 $Y=2.065 $X2=0
+ $Y2=0
cc_466 N_A_299_47#_c_628_n N_VPWR_c_899_n 0.00903378f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_A_299_47#_c_646_n N_VPWR_c_899_n 0.0253092f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_468 N_A_299_47#_c_646_n N_VPWR_c_910_n 0.0424693f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_469 N_A_299_47#_c_628_n N_VPWR_c_911_n 0.0067571f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_470 N_A_299_47#_c_646_n N_VPWR_c_911_n 0.0240862f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_471 N_A_299_47#_c_636_n N_VPWR_c_911_n 0.00308511f $X=2.215 $Y=2.125 $X2=0
+ $Y2=0
cc_472 N_A_299_47#_c_628_n N_VPWR_c_912_n 0.0062441f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_473 N_A_299_47#_c_646_n N_A_27_47#_c_1018_n 0.0186379f $X=2.13 $Y=2.295 $X2=0
+ $Y2=0
cc_474 N_A_299_47#_c_646_n A_410_413# 0.00683749f $X=2.13 $Y=2.295 $X2=-0.19
+ $Y2=-0.24
cc_475 N_A_299_47#_c_636_n A_410_413# 0.0014313f $X=2.215 $Y=2.125 $X2=-0.19
+ $Y2=-0.24
cc_476 N_A_299_47#_c_628_n N_VGND_c_1066_n 0.00209689f $X=3.225 $Y=1.41 $X2=0
+ $Y2=0
cc_477 N_A_299_47#_c_629_n N_VGND_c_1066_n 0.0064755f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_478 N_A_299_47#_c_642_n N_VGND_c_1066_n 0.0156107f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_479 N_A_299_47#_c_632_n N_VGND_c_1066_n 0.0138859f $X=2.56 $Y=0.995 $X2=0
+ $Y2=0
cc_480 N_A_299_47#_c_633_n N_VGND_c_1066_n 0.0112879f $X=3.12 $Y=1.16 $X2=0
+ $Y2=0
cc_481 N_A_299_47#_c_642_n N_VGND_c_1071_n 0.0704643f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_482 N_A_299_47#_c_629_n N_VGND_c_1072_n 0.00585385f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_483 N_A_299_47#_M1014_d N_VGND_c_1074_n 0.003457f $X=1.495 $Y=0.235 $X2=0
+ $Y2=0
cc_484 N_A_299_47#_c_629_n N_VGND_c_1074_n 0.00812028f $X=3.25 $Y=0.995 $X2=0
+ $Y2=0
cc_485 N_A_299_47#_c_642_n N_VGND_c_1074_n 0.0318035f $X=2.475 $Y=0.395 $X2=0
+ $Y2=0
cc_486 N_A_299_47#_c_642_n A_415_47# 0.0103317f $X=2.475 $Y=0.395 $X2=-0.19
+ $Y2=-0.24
cc_487 N_A_299_47#_c_632_n A_415_47# 0.00167546f $X=2.56 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_488 N_CLK_c_740_n N_A_1089_47#_c_825_n 0.0155223f $X=6.285 $Y=1.67 $X2=0
+ $Y2=0
cc_489 N_CLK_c_741_n N_A_1089_47#_c_825_n 0.0187655f $X=6.285 $Y=1.77 $X2=0
+ $Y2=0
cc_490 N_CLK_c_735_n N_A_1089_47#_c_825_n 0.00214331f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_491 N_CLK_c_736_n N_A_1089_47#_c_825_n 0.0206471f $X=6.25 $Y=1.16 $X2=0 $Y2=0
cc_492 N_CLK_M1013_g N_A_1089_47#_c_826_n 0.0219147f $X=6.31 $Y=0.445 $X2=0
+ $Y2=0
cc_493 N_CLK_M1013_g N_A_1089_47#_c_827_n 0.012164f $X=6.31 $Y=0.445 $X2=0 $Y2=0
cc_494 N_CLK_c_733_n N_A_1089_47#_c_827_n 0.00694877f $X=5.94 $Y=1.19 $X2=0
+ $Y2=0
cc_495 N_CLK_c_734_n N_A_1089_47#_c_827_n 0.00232634f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_496 N_CLK_c_735_n N_A_1089_47#_c_827_n 0.0265421f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_497 N_CLK_c_736_n N_A_1089_47#_c_827_n 0.00280903f $X=6.25 $Y=1.16 $X2=0
+ $Y2=0
cc_498 N_CLK_M1007_g N_A_1089_47#_c_828_n 6.0552e-19 $X=4.79 $Y=0.445 $X2=0
+ $Y2=0
cc_499 N_CLK_c_733_n N_A_1089_47#_c_828_n 0.00108081f $X=5.94 $Y=1.19 $X2=0
+ $Y2=0
cc_500 N_CLK_c_741_n N_A_1089_47#_c_840_n 0.00477137f $X=6.285 $Y=1.77 $X2=0
+ $Y2=0
cc_501 N_CLK_c_740_n N_A_1089_47#_c_829_n 0.00326424f $X=6.285 $Y=1.67 $X2=0
+ $Y2=0
cc_502 N_CLK_M1013_g N_A_1089_47#_c_829_n 0.00405202f $X=6.31 $Y=0.445 $X2=0
+ $Y2=0
cc_503 N_CLK_c_734_n N_A_1089_47#_c_829_n 0.001051f $X=6.085 $Y=1.19 $X2=0 $Y2=0
cc_504 N_CLK_c_735_n N_A_1089_47#_c_829_n 0.0179762f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_505 N_CLK_c_736_n N_A_1089_47#_c_829_n 3.80665e-19 $X=6.25 $Y=1.16 $X2=0
+ $Y2=0
cc_506 N_CLK_c_740_n N_A_1089_47#_c_832_n 0.0100532f $X=6.285 $Y=1.67 $X2=0
+ $Y2=0
cc_507 N_CLK_c_741_n N_A_1089_47#_c_832_n 0.019834f $X=6.285 $Y=1.77 $X2=0 $Y2=0
cc_508 N_CLK_c_734_n N_A_1089_47#_c_832_n 0.00217896f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_509 N_CLK_c_735_n N_A_1089_47#_c_832_n 0.0340841f $X=6.085 $Y=1.19 $X2=0
+ $Y2=0
cc_510 N_CLK_c_736_n N_A_1089_47#_c_832_n 0.00162024f $X=6.25 $Y=1.16 $X2=0
+ $Y2=0
cc_511 N_CLK_c_741_n N_VPWR_c_902_n 0.00183161f $X=6.285 $Y=1.77 $X2=0 $Y2=0
cc_512 N_CLK_M1002_g N_VPWR_c_903_n 0.0274119f $X=4.815 $Y=1.835 $X2=0 $Y2=0
cc_513 N_CLK_c_741_n N_VPWR_c_904_n 5.67264e-19 $X=6.285 $Y=1.77 $X2=0 $Y2=0
cc_514 N_CLK_c_741_n N_VPWR_c_905_n 0.00510113f $X=6.285 $Y=1.77 $X2=0 $Y2=0
cc_515 N_CLK_c_741_n N_VPWR_c_899_n 0.00677441f $X=6.285 $Y=1.77 $X2=0 $Y2=0
cc_516 N_CLK_M1007_g N_VGND_c_1067_n 0.00548485f $X=4.79 $Y=0.445 $X2=0 $Y2=0
cc_517 N_CLK_M1013_g N_VGND_c_1068_n 0.0111788f $X=6.31 $Y=0.445 $X2=0 $Y2=0
cc_518 N_CLK_M1007_g N_VGND_c_1069_n 0.00422112f $X=4.79 $Y=0.445 $X2=0 $Y2=0
cc_519 N_CLK_M1013_g N_VGND_c_1069_n 0.00253267f $X=6.31 $Y=0.445 $X2=0 $Y2=0
cc_520 N_CLK_M1007_g N_VGND_c_1074_n 0.00762862f $X=4.79 $Y=0.445 $X2=0 $Y2=0
cc_521 N_CLK_M1013_g N_VGND_c_1074_n 0.00329891f $X=6.31 $Y=0.445 $X2=0 $Y2=0
cc_522 N_A_1089_47#_c_832_n N_VPWR_M1016_d 0.00916762f $X=6.73 $Y=1.79 $X2=0
+ $Y2=0
cc_523 N_A_1089_47#_c_825_n N_VPWR_c_902_n 0.00327647f $X=6.81 $Y=1.41 $X2=0
+ $Y2=0
cc_524 N_A_1089_47#_c_832_n N_VPWR_c_902_n 0.0191719f $X=6.73 $Y=1.79 $X2=0
+ $Y2=0
cc_525 N_A_1089_47#_c_840_n N_VPWR_c_904_n 0.013449f $X=6.04 $Y=2.085 $X2=0
+ $Y2=0
cc_526 N_A_1089_47#_c_840_n N_VPWR_c_905_n 0.0113299f $X=6.04 $Y=2.085 $X2=0
+ $Y2=0
cc_527 N_A_1089_47#_c_832_n N_VPWR_c_905_n 0.00411817f $X=6.73 $Y=1.79 $X2=0
+ $Y2=0
cc_528 N_A_1089_47#_c_825_n N_VPWR_c_908_n 0.00600944f $X=6.81 $Y=1.41 $X2=0
+ $Y2=0
cc_529 N_A_1089_47#_c_832_n N_VPWR_c_908_n 0.00171698f $X=6.73 $Y=1.79 $X2=0
+ $Y2=0
cc_530 N_A_1089_47#_M1001_d N_VPWR_c_899_n 0.0047429f $X=5.895 $Y=1.845 $X2=0
+ $Y2=0
cc_531 N_A_1089_47#_c_825_n N_VPWR_c_899_n 0.010503f $X=6.81 $Y=1.41 $X2=0 $Y2=0
cc_532 N_A_1089_47#_c_840_n N_VPWR_c_899_n 0.00637602f $X=6.04 $Y=2.085 $X2=0
+ $Y2=0
cc_533 N_A_1089_47#_c_832_n N_VPWR_c_899_n 0.0109373f $X=6.73 $Y=1.79 $X2=0
+ $Y2=0
cc_534 N_A_1089_47#_c_825_n GCLK 0.0126536f $X=6.81 $Y=1.41 $X2=0 $Y2=0
cc_535 N_A_1089_47#_c_826_n GCLK 0.0223692f $X=6.835 $Y=0.995 $X2=0 $Y2=0
cc_536 N_A_1089_47#_c_827_n GCLK 0.0137304f $X=6.645 $Y=0.7 $X2=0 $Y2=0
cc_537 N_A_1089_47#_c_829_n GCLK 0.0521292f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_538 N_A_1089_47#_c_832_n GCLK 0.0474911f $X=6.73 $Y=1.79 $X2=0 $Y2=0
cc_539 N_A_1089_47#_c_827_n N_VGND_M1013_d 0.00866786f $X=6.645 $Y=0.7 $X2=0
+ $Y2=0
cc_540 N_A_1089_47#_c_829_n N_VGND_M1013_d 0.00122986f $X=6.73 $Y=1.16 $X2=0
+ $Y2=0
cc_541 N_A_1089_47#_c_825_n N_VGND_c_1068_n 2.19196e-19 $X=6.81 $Y=1.41 $X2=0
+ $Y2=0
cc_542 N_A_1089_47#_c_826_n N_VGND_c_1068_n 0.00539507f $X=6.835 $Y=0.995 $X2=0
+ $Y2=0
cc_543 N_A_1089_47#_c_827_n N_VGND_c_1068_n 0.0227671f $X=6.645 $Y=0.7 $X2=0
+ $Y2=0
cc_544 N_A_1089_47#_c_833_n N_VGND_c_1069_n 0.0114f $X=5.62 $Y=0.46 $X2=0 $Y2=0
cc_545 N_A_1089_47#_c_827_n N_VGND_c_1069_n 0.00975466f $X=6.645 $Y=0.7 $X2=0
+ $Y2=0
cc_546 N_A_1089_47#_c_826_n N_VGND_c_1073_n 0.00525463f $X=6.835 $Y=0.995 $X2=0
+ $Y2=0
cc_547 N_A_1089_47#_c_827_n N_VGND_c_1073_n 0.00198779f $X=6.645 $Y=0.7 $X2=0
+ $Y2=0
cc_548 N_A_1089_47#_M1008_s N_VGND_c_1074_n 0.00583031f $X=5.445 $Y=0.235 $X2=0
+ $Y2=0
cc_549 N_A_1089_47#_c_826_n N_VGND_c_1074_n 0.0102389f $X=6.835 $Y=0.995 $X2=0
+ $Y2=0
cc_550 N_A_1089_47#_c_833_n N_VGND_c_1074_n 0.00642843f $X=5.62 $Y=0.46 $X2=0
+ $Y2=0
cc_551 N_A_1089_47#_c_827_n N_VGND_c_1074_n 0.0220442f $X=6.645 $Y=0.7 $X2=0
+ $Y2=0
cc_552 N_A_1089_47#_c_827_n A_1181_47# 0.0036795f $X=6.645 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_553 N_VPWR_c_899_n A_117_369# 0.001847f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_554 N_VPWR_c_899_n N_A_27_47#_M1003_d 0.00460184f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_555 N_VPWR_c_901_n N_A_27_47#_c_997_n 0.0210314f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_556 N_VPWR_c_901_n N_A_27_47#_c_1009_n 0.027538f $X=0.26 $Y=2 $X2=0 $Y2=0
cc_557 N_VPWR_c_899_n N_A_27_47#_c_1009_n 0.00621702f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_558 N_VPWR_c_910_n N_A_27_47#_c_1009_n 0.00975127f $X=2.52 $Y=2.44 $X2=0
+ $Y2=0
cc_559 N_VPWR_c_899_n N_A_27_47#_c_1018_n 0.0216808f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_560 N_VPWR_c_910_n N_A_27_47#_c_1018_n 0.0355985f $X=2.52 $Y=2.44 $X2=0 $Y2=0
cc_561 N_VPWR_c_899_n A_410_413# 0.00736425f $X=7.13 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_562 N_VPWR_c_899_n N_GCLK_M1012_d 0.0053737f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_563 N_VPWR_c_908_n GCLK 0.0174931f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_564 N_VPWR_c_899_n GCLK 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_565 A_117_369# N_A_27_47#_c_997_n 0.00282259f $X=0.585 $Y=1.845 $X2=0 $Y2=0
cc_566 A_117_369# N_A_27_47#_c_1009_n 4.10738e-19 $X=0.585 $Y=1.845 $X2=0.26
+ $Y2=2
cc_567 A_117_369# N_A_27_47#_c_1018_n 0.00367792f $X=0.585 $Y=1.845 $X2=3.885
+ $Y2=2.72
cc_568 N_A_27_47#_c_998_n N_VGND_M1015_d 0.00129376f $X=1.115 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_569 N_A_27_47#_c_999_n N_VGND_M1015_d 3.36173e-19 $X=0.685 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_570 N_A_27_47#_c_996_n N_VGND_c_1070_n 0.0173928f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_571 N_A_27_47#_c_999_n N_VGND_c_1070_n 0.00260613f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_572 N_A_27_47#_c_998_n N_VGND_c_1071_n 0.00341938f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_573 N_A_27_47#_c_1022_n N_VGND_c_1071_n 0.0120906f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_574 N_A_27_47#_M1015_s N_VGND_c_1074_n 0.00286466f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_575 N_A_27_47#_M1021_d N_VGND_c_1074_n 0.00463742f $X=1.02 $Y=0.235 $X2=0
+ $Y2=0
cc_576 N_A_27_47#_c_996_n N_VGND_c_1074_n 0.00977915f $X=0.26 $Y=0.43 $X2=0
+ $Y2=0
cc_577 N_A_27_47#_c_998_n N_VGND_c_1074_n 0.00569248f $X=1.115 $Y=0.7 $X2=0
+ $Y2=0
cc_578 N_A_27_47#_c_999_n N_VGND_c_1074_n 0.00628516f $X=0.685 $Y=0.7 $X2=0
+ $Y2=0
cc_579 N_A_27_47#_c_1022_n N_VGND_c_1074_n 0.00681108f $X=1.2 $Y=0.42 $X2=0
+ $Y2=0
cc_580 N_A_27_47#_c_996_n N_VGND_c_1075_n 0.0146378f $X=0.26 $Y=0.43 $X2=0 $Y2=0
cc_581 N_A_27_47#_c_999_n N_VGND_c_1075_n 0.0193989f $X=0.685 $Y=0.7 $X2=0 $Y2=0
cc_582 N_A_27_47#_c_1022_n N_VGND_c_1075_n 0.0116788f $X=1.2 $Y=0.42 $X2=0 $Y2=0
cc_583 GCLK N_VGND_c_1068_n 0.00989259f $X=7.045 $Y=0.425 $X2=0 $Y2=0
cc_584 GCLK N_VGND_c_1073_n 0.0174931f $X=7.045 $Y=0.425 $X2=0 $Y2=0
cc_585 N_GCLK_M1018_d N_VGND_c_1074_n 0.00494456f $X=6.91 $Y=0.235 $X2=0 $Y2=0
cc_586 GCLK N_VGND_c_1074_n 0.00955092f $X=7.045 $Y=0.425 $X2=0 $Y2=0
cc_587 N_VGND_c_1074_n A_415_47# 0.00329302f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
cc_588 N_VGND_c_1074_n A_1181_47# 0.00378298f $X=7.13 $Y=0 $X2=-0.19 $Y2=-0.24
