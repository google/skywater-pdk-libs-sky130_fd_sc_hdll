* File: sky130_fd_sc_hdll__nor2_4.pex.spice
* Created: Wed Sep  2 08:39:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 26 40 41 47
r79 41 42 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r80 39 41 20.0833 $w=3.72e-07 $l=1.55e-07 $layer=POLY_cond $X=1.77 $Y=1.202
+ $X2=1.925 $Y2=1.202
r81 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.77
+ $Y=1.16 $X2=1.77 $Y2=1.16
r82 37 39 40.8145 $w=3.72e-07 $l=3.15e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.77 $Y2=1.202
r83 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r84 35 36 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r85 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r86 33 47 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.6 $Y=1.175
+ $X2=0.695 $Y2=1.175
r87 32 34 46.6452 $w=3.72e-07 $l=3.6e-07 $layer=POLY_cond $X=0.6 $Y=1.202
+ $X2=0.96 $Y2=1.202
r88 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.6 $Y=1.16
+ $X2=0.6 $Y2=1.16
r89 30 32 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.6 $Y2=1.202
r90 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r91 26 40 56.8409 $w=1.98e-07 $l=1.025e-06 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=1.77 $Y2=1.175
r92 26 47 2.77273 $w=1.98e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.175
+ $X2=0.695 $Y2=1.175
r93 25 33 20.2409 $w=1.98e-07 $l=3.65e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.6 $Y2=1.175
r94 22 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r95 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r96 19 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r97 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r98 16 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r99 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r100 13 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r101 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r102 10 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r103 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r104 7 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r105 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=0.56
r106 4 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r107 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r108 1 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r109 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 38 39 44
c86 10 0 7.78669e-20 $X=2.865 $Y=1.41
r87 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=3.83 $Y2=1.202
r88 37 39 18.1398 $w=3.72e-07 $l=1.4e-07 $layer=POLY_cond $X=3.665 $Y=1.202
+ $X2=3.805 $Y2=1.202
r89 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.665
+ $Y=1.16 $X2=3.665 $Y2=1.16
r90 35 37 42.7581 $w=3.72e-07 $l=3.3e-07 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.665 $Y2=1.202
r91 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.202
+ $X2=3.335 $Y2=1.202
r92 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.865 $Y=1.202
+ $X2=3.31 $Y2=1.202
r93 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r94 31 44 43.8091 $w=1.98e-07 $l=7.9e-07 $layer=LI1_cond $X=2.495 $Y=1.175
+ $X2=3.285 $Y2=1.175
r95 30 32 44.7016 $w=3.72e-07 $l=3.45e-07 $layer=POLY_cond $X=2.495 $Y=1.202
+ $X2=2.84 $Y2=1.202
r96 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.495
+ $Y=1.16 $X2=2.495 $Y2=1.16
r97 28 30 12.957 $w=3.72e-07 $l=1e-07 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.495 $Y2=1.202
r98 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r99 25 38 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=3.295 $Y=1.175
+ $X2=3.665 $Y2=1.175
r100 25 44 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=3.295 $Y=1.175
+ $X2=3.285 $Y2=1.175
r101 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.202
r102 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r103 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r104 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r105 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r106 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r107 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.202
r108 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r109 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r110 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r111 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r112 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r113 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r114 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r115 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r116 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29 30
+ 32 37 43 48
c86 28 0 7.78669e-20 $X=2.135 $Y=1.665
r87 43 45 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.075 $Y2=2.38
r88 33 45 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.265 $Y=2.38
+ $X2=3.075 $Y2=2.38
r89 32 48 9.7744 $w=4.63e-07 $l=3.8e-07 $layer=LI1_cond $X=4.057 $Y=2.38
+ $X2=4.057 $Y2=2
r90 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.825 $Y=2.38
+ $X2=3.265 $Y2=2.38
r91 31 41 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=2.38
+ $X2=2.135 $Y2=2.38
r92 30 45 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=2.38
+ $X2=3.075 $Y2=2.38
r93 30 31 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.885 $Y=2.38
+ $X2=2.325 $Y2=2.38
r94 29 41 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=2.295
+ $X2=2.135 $Y2=2.38
r95 28 39 2.69784 $w=3.8e-07 $l=1.05e-07 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.135 $Y2=1.56
r96 28 29 19.1063 $w=3.78e-07 $l=6.3e-07 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.135 $Y2=2.295
r97 27 37 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=1.56 $X2=1.22
+ $Y2=1.56
r98 26 39 4.88181 $w=2.1e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=1.56
+ $X2=2.135 $Y2=1.56
r99 26 27 33.8009 $w=2.08e-07 $l=6.4e-07 $layer=LI1_cond $X=1.945 $Y=1.56
+ $X2=1.305 $Y2=1.56
r100 22 37 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=1.56
r101 22 24 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.22 $Y=1.665
+ $X2=1.22 $Y2=2.3
r102 21 35 3.96222 $w=2.1e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=1.56
+ $X2=0.227 $Y2=1.56
r103 20 37 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=1.22 $Y2=1.56
r104 20 21 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=1.56
+ $X2=0.365 $Y2=1.56
r105 16 35 3.01473 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=1.56
r106 16 18 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=0.227 $Y=1.665
+ $X2=0.227 $Y2=2.3
r107 5 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=2
r108 4 43 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.02
r109 3 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.34
r110 3 39 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r111 2 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r112 2 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r113 1 35 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r114 1 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%VPWR 1 2 9 13 15 17 22 32 33 36 39
r60 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 32 33 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r63 30 33 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=4.37 $Y2=2.72
r64 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 29 32 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=4.37 $Y2=2.72
r66 29 30 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 27 39 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.625 $Y2=2.72
r68 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 26 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r70 26 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 23 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=0.725 $Y2=2.72
r73 23 25 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=0.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r74 22 39 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.625 $Y2=2.72
r75 22 25 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=1.475 $Y=2.72
+ $X2=1.15 $Y2=2.72
r76 17 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.725 $Y2=2.72
r77 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 15 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r79 15 19 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r80 11 39 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.625 $Y=2.635
+ $X2=1.625 $Y2=2.72
r81 11 13 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=1.625 $Y=2.635
+ $X2=1.625 $Y2=2
r82 7 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2.72
r83 7 9 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.725 $Y=2.635
+ $X2=0.725 $Y2=2
r84 2 13 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2
r85 1 9 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%Y 1 2 3 4 5 6 21 23 24 27 29 33 35 37 39 41
+ 45 49 51 53 55 56 59 61 63
r125 62 63 12.2278 $w=5.63e-07 $l=5.4e-07 $layer=LI1_cond $X=4.292 $Y=0.905
+ $X2=4.292 $Y2=1.445
r126 54 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.735 $Y=0.815
+ $X2=3.545 $Y2=0.815
r127 53 62 8.1363 $w=1.8e-07 $l=2.37779e-07 $layer=LI1_cond $X=4.095 $Y=0.815
+ $X2=4.292 $Y2=0.905
r128 53 54 22.1818 $w=1.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.095 $Y=0.815
+ $X2=3.735 $Y2=0.815
r129 52 61 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=1.595
+ $X2=3.57 $Y2=1.595
r130 51 63 3.96467 $w=3e-07 $l=1.97e-07 $layer=LI1_cond $X=4.095 $Y=1.595
+ $X2=4.292 $Y2=1.595
r131 51 52 16.9025 $w=2.98e-07 $l=4.4e-07 $layer=LI1_cond $X=4.095 $Y=1.595
+ $X2=3.655 $Y2=1.595
r132 47 61 3.44808 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.57 $Y=1.745
+ $X2=3.57 $Y2=1.595
r133 47 49 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.57 $Y=1.745
+ $X2=3.57 $Y2=1.96
r134 43 59 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.815
r135 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.545 $Y=0.725
+ $X2=3.545 $Y2=0.39
r136 42 56 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.795 $Y=0.815
+ $X2=2.605 $Y2=0.815
r137 41 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=3.545 $Y2=0.815
r138 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.355 $Y=0.815
+ $X2=2.795 $Y2=0.815
r139 40 58 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=1.595
+ $X2=2.63 $Y2=1.595
r140 39 61 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=1.595
+ $X2=3.57 $Y2=1.595
r141 39 40 29.5794 $w=2.98e-07 $l=7.7e-07 $layer=LI1_cond $X=3.485 $Y=1.595
+ $X2=2.715 $Y2=1.595
r142 35 58 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.63 $Y=1.745
+ $X2=2.63 $Y2=1.595
r143 35 37 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.63 $Y=1.745
+ $X2=2.63 $Y2=1.96
r144 31 56 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.815
r145 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.605 $Y=0.725
+ $X2=2.605 $Y2=0.39
r146 30 55 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r147 29 56 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=2.605 $Y2=0.815
r148 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.415 $Y=0.815
+ $X2=1.855 $Y2=0.815
r149 25 55 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r150 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r151 23 55 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r152 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r153 19 24 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r154 19 21 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r155 6 61 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
r156 6 49 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.96
r157 5 58 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.62
r158 5 37 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.96
r159 4 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.39
r160 3 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
r161 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r162 1 21 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR2_4%VGND 1 2 3 4 5 16 18 20 24 28 32 36 39 40
+ 42 43 45 46 47 60 61 67
r77 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r78 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r79 58 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r80 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r81 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r82 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r83 52 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r84 52 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r85 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r86 49 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r87 49 51 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r88 47 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r89 47 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r90 45 57 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.955 $Y=0 $X2=3.91
+ $Y2=0
r91 45 46 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.955 $Y=0 $X2=4.097
+ $Y2=0
r92 44 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.37
+ $Y2=0
r93 44 46 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.097
+ $Y2=0
r94 42 54 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=2.99
+ $Y2=0
r95 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.015 $Y=0 $X2=3.1
+ $Y2=0
r96 41 57 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.91
+ $Y2=0
r97 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.185 $Y=0 $X2=3.1
+ $Y2=0
r98 39 51 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.07
+ $Y2=0
r99 39 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.075 $Y=0 $X2=2.16
+ $Y2=0
r100 38 54 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.245 $Y=0
+ $X2=2.99 $Y2=0
r101 38 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.16
+ $Y2=0
r102 34 46 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=4.097 $Y=0.085
+ $X2=4.097 $Y2=0
r103 34 36 12.3332 $w=2.83e-07 $l=3.05e-07 $layer=LI1_cond $X=4.097 $Y=0.085
+ $X2=4.097 $Y2=0.39
r104 30 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=0.085 $X2=3.1
+ $Y2=0
r105 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.1 $Y=0.085
+ $X2=3.1 $Y2=0.39
r106 26 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0
r107 26 28 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.16 $Y=0.085
+ $X2=2.16 $Y2=0.39
r108 22 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r109 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r110 21 64 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0
+ $X2=0.182 $Y2=0
r111 20 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r112 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.365 $Y2=0
r113 16 64 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r114 16 18 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r115 5 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.39
r116 4 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r117 3 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r118 2 24 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r119 1 18 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

