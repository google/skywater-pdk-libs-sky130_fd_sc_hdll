* File: sky130_fd_sc_hdll__xor3_2.pex.spice
* Created: Wed Sep  2 08:54:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_81_21# 1 2 7 9 10 12 13 15 16 18 19 20 21
+ 23 24 26 28 30 31 33 40 41 46
r126 45 46 0.656676 $w=3.67e-07 $l=5e-09 $layer=POLY_cond $X=0.975 $Y=1.202
+ $X2=0.98 $Y2=1.202
r127 44 45 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=0.505 $Y=1.202
+ $X2=0.975 $Y2=1.202
r128 43 44 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.48 $Y=1.202
+ $X2=0.505 $Y2=1.202
r129 40 41 13.5904 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=3.025 $Y=0.355
+ $X2=2.785 $Y2=0.355
r130 38 46 26.267 $w=3.67e-07 $l=2e-07 $layer=POLY_cond $X=1.18 $Y=1.202
+ $X2=0.98 $Y2=1.202
r131 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.18
+ $Y=1.16 $X2=1.18 $Y2=1.16
r132 35 37 25.0595 $w=1.85e-07 $l=3.8e-07 $layer=LI1_cond $X=1.195 $Y=0.78
+ $X2=1.195 $Y2=1.16
r133 31 33 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.865 $Y=2.32
+ $X2=3.025 $Y2=2.32
r134 30 41 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.745 $Y=0.34
+ $X2=2.785 $Y2=0.34
r135 28 31 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.755 $Y=2.235
+ $X2=1.865 $Y2=2.32
r136 27 28 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.755 $Y=2.045
+ $X2=1.755 $Y2=2.235
r137 25 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.635 $Y=0.425
+ $X2=1.745 $Y2=0.34
r138 25 26 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.635 $Y=0.425
+ $X2=1.635 $Y2=0.695
r139 23 27 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.645 $Y=1.96
+ $X2=1.755 $Y2=2.045
r140 23 24 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.645 $Y=1.96
+ $X2=1.295 $Y2=1.96
r141 22 35 1.22693 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=0.78
+ $X2=1.195 $Y2=0.78
r142 21 26 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.525 $Y=0.78
+ $X2=1.635 $Y2=0.695
r143 21 22 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.525 $Y=0.78
+ $X2=1.295 $Y2=0.78
r144 20 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.21 $Y=1.875
+ $X2=1.295 $Y2=1.96
r145 19 37 10.9829 $w=1.85e-07 $l=1.72337e-07 $layer=LI1_cond $X=1.21 $Y=1.325
+ $X2=1.195 $Y2=1.16
r146 19 20 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=1.21 $Y=1.325
+ $X2=1.21 $Y2=1.875
r147 16 46 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.98 $Y=0.995
+ $X2=0.98 $Y2=1.202
r148 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.98 $Y=0.995
+ $X2=0.98 $Y2=0.56
r149 13 45 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.202
r150 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
r151 10 44 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.202
r152 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.985
r153 7 43 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=1.202
r154 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.48 $Y=0.995
+ $X2=0.48 $Y2=0.56
r155 2 33 600 $w=1.7e-07 $l=7.84267e-07 $layer=licon1_PDIFF $count=1 $X=2.835
+ $Y=1.625 $X2=3.025 $Y2=2.32
r156 1 40 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.89
+ $Y=0.245 $X2=3.025 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%C 1 3 7 8 10 12 13 15 16 18 22
r65 18 22 0.52383 $w=6.83e-07 $l=3e-08 $layer=LI1_cond $X=2.597 $Y=1.19
+ $X2=2.597 $Y2=1.16
r66 13 15 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.815 $Y=0.995
+ $X2=2.815 $Y2=0.565
r67 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.745 $Y=1.55
+ $X2=2.745 $Y2=2.045
r68 9 16 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.725 $Y=1.16
+ $X2=1.625 $Y2=1.202
r69 8 10 84.4272 $w=2.29e-07 $l=4.00849e-07 $layer=POLY_cond $X=2.767 $Y=1.16
+ $X2=2.745 $Y2=1.55
r70 8 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.705
+ $Y=1.16 $X2=2.705 $Y2=1.16
r71 8 13 40.4635 $w=2.29e-07 $l=1.8747e-07 $layer=POLY_cond $X=2.767 $Y=1.16
+ $X2=2.815 $Y2=0.995
r72 8 9 160.872 $w=3.3e-07 $l=9.2e-07 $layer=POLY_cond $X=2.645 $Y=1.16
+ $X2=1.725 $Y2=1.16
r73 4 16 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.625 $Y2=1.202
r74 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.625 $Y=1.41
+ $X2=1.625 $Y2=1.805
r75 1 16 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.6 $Y=0.995
+ $X2=1.625 $Y2=1.202
r76 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.6 $Y=0.995 $X2=1.6
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_335_93# 1 2 7 9 10 12 13 18 20 23 24 28
r75 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.3
+ $Y=1.16 $X2=3.3 $Y2=1.16
r76 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=3.195 $Y=1.16
+ $X2=3.3 $Y2=1.16
r77 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.16
r78 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=3.195 $Y=1.325
+ $X2=3.195 $Y2=1.535
r79 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.085 $Y=1.62 $X2=2
+ $Y2=1.62
r80 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.11 $Y=1.62
+ $X2=3.195 $Y2=1.535
r81 20 21 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=3.11 $Y=1.62
+ $X2=2.085 $Y2=1.62
r82 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2 $Y=1.535 $X2=2
+ $Y2=1.62
r83 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=2 $Y=1.535 $X2=2
+ $Y2=0.76
r84 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.915 $Y=1.62 $X2=2
+ $Y2=1.62
r85 13 15 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=1.915 $Y=1.62
+ $X2=1.86 $Y2=1.62
r86 10 29 38.8824 $w=2.71e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.325 $Y2=1.16
r87 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.41 $Y=0.995
+ $X2=3.41 $Y2=0.565
r88 7 29 74.8096 $w=2.71e-07 $l=3.9e-07 $layer=POLY_cond $X=3.325 $Y=1.55
+ $X2=3.325 $Y2=1.16
r89 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.325 $Y=1.55
+ $X2=3.325 $Y2=2.045
r90 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.715
+ $Y=1.485 $X2=1.86 $Y2=1.62
r91 1 18 182 $w=1.7e-07 $l=4.48888e-07 $layer=licon1_NDIFF $count=1 $X=1.675
+ $Y=0.465 $X2=2 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_934_297# 1 2 7 9 12 14 15 16 18 19 21 22
+ 23 27 35 37 38 39 40 47 49 50 58
c180 14 0 8.91061e-20 $X=8.075 $Y=1.28
r181 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.005
+ $Y=1.11 $X2=8.005 $Y2=1.11
r182 50 56 11.5766 $w=2.74e-07 $l=2.6e-07 $layer=LI1_cond $X=7.93 $Y=0.85
+ $X2=7.93 $Y2=1.11
r183 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.875 $Y=0.85
+ $X2=7.875 $Y2=0.85
r184 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.395 $Y=0.85
+ $X2=6.395 $Y2=0.85
r185 42 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.915 $Y=0.85
+ $X2=4.915 $Y2=0.85
r186 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.54 $Y=0.85
+ $X2=6.395 $Y2=0.85
r187 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.73 $Y=0.85
+ $X2=7.875 $Y2=0.85
r188 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=7.73 $Y=0.85
+ $X2=6.54 $Y2=0.85
r189 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.06 $Y=0.85
+ $X2=4.915 $Y2=0.85
r190 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.25 $Y=0.85
+ $X2=6.395 $Y2=0.85
r191 37 38 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=6.25 $Y=0.85
+ $X2=5.06 $Y2=0.85
r192 35 47 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=6.372 $Y=0.995
+ $X2=6.372 $Y2=0.85
r193 31 35 6.36987 $w=2.73e-07 $l=1.52e-07 $layer=LI1_cond $X=6.22 $Y=1.132
+ $X2=6.372 $Y2=1.132
r194 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.22
+ $Y=1.16 $X2=6.22 $Y2=1.16
r195 28 58 28.8111 $w=2.88e-07 $l=7.25e-07 $layer=LI1_cond $X=4.97 $Y=1.445
+ $X2=4.97 $Y2=0.72
r196 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.97 $Y=1.58
+ $X2=4.97 $Y2=1.445
r197 25 27 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.815 $Y=1.58
+ $X2=4.97 $Y2=1.58
r198 22 32 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.485 $Y=1.16
+ $X2=6.22 $Y2=1.16
r199 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=6.485 $Y=1.16
+ $X2=6.585 $Y2=1.202
r200 19 55 38.5326 $w=3.08e-07 $l=2.0106e-07 $layer=POLY_cond $X=8.105 $Y=0.945
+ $X2=8.025 $Y2=1.11
r201 19 21 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=8.105 $Y=0.945
+ $X2=8.105 $Y2=0.535
r202 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.075 $Y=1.57
+ $X2=8.075 $Y2=2.065
r203 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.075 $Y=1.47 $X2=8.075
+ $Y2=1.57
r204 14 55 32.5213 $w=3.08e-07 $l=1.93391e-07 $layer=POLY_cond $X=8.075 $Y=1.28
+ $X2=8.025 $Y2=1.11
r205 14 15 62.9997 $w=2e-07 $l=1.9e-07 $layer=POLY_cond $X=8.075 $Y=1.28
+ $X2=8.075 $Y2=1.47
r206 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=6.61 $Y=0.995
+ $X2=6.585 $Y2=1.202
r207 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.61 $Y=0.995
+ $X2=6.61 $Y2=0.455
r208 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=6.585 $Y=1.41
+ $X2=6.585 $Y2=1.202
r209 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.585 $Y=1.41
+ $X2=6.585 $Y2=1.805
r210 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.67
+ $Y=1.485 $X2=4.815 $Y2=1.63
r211 1 58 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=5.03 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 33
+ 38 39 40 42
c135 42 0 1.94872e-19 $X=7.6 $Y=1.555
r136 38 41 40.3353 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.47 $Y=1.16
+ $X2=7.47 $Y2=1.325
r137 38 40 48.2009 $w=2.8e-07 $l=1.65e-07 $layer=POLY_cond $X=7.47 $Y=1.16
+ $X2=7.47 $Y2=0.995
r138 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.465
+ $Y=1.16 $X2=7.465 $Y2=1.16
r139 33 42 3.40825 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=7.49 $Y=1.555
+ $X2=7.6 $Y2=1.555
r140 33 39 11.5822 $w=3.08e-07 $l=2.85e-07 $layer=LI1_cond $X=7.49 $Y=1.445
+ $X2=7.49 $Y2=1.16
r141 33 42 2.21818 $w=2.2e-07 $l=4e-08 $layer=LI1_cond $X=7.64 $Y=1.555 $X2=7.6
+ $Y2=1.555
r142 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.775 $Y=1.16
+ $X2=5.775 $Y2=1.085
r143 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=7.51 $Y=2.415
+ $X2=7.51 $Y2=1.965
r144 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.51 $Y=1.57
+ $X2=7.51 $Y2=1.965
r145 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.51 $Y=1.47 $X2=7.51
+ $Y2=1.57
r146 24 41 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=7.51 $Y=1.47
+ $X2=7.51 $Y2=1.325
r147 22 40 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.405 $Y=0.565
+ $X2=7.405 $Y2=0.995
r148 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=7.41 $Y=2.54
+ $X2=7.51 $Y2=2.415
r149 18 19 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=7.41 $Y=2.54
+ $X2=5.875 $Y2=2.54
r150 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.8 $Y=0.565
+ $X2=5.8 $Y2=1.085
r151 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=5.775 $Y=2.455
+ $X2=5.875 $Y2=2.54
r152 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=5.775 $Y=2.455
+ $X2=5.775 $Y2=1.905
r153 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=5.775 $Y=1.41
+ $X2=5.775 $Y2=1.16
r154 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.775 $Y=1.41
+ $X2=5.775 $Y2=1.905
r155 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.675 $Y=1.16
+ $X2=5.775 $Y2=1.16
r156 8 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=5.675 $Y=1.16
+ $X2=4.845 $Y2=1.16
r157 4 9 21.9526 $w=2.45e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.77 $Y=1.085
+ $X2=4.845 $Y2=1.16
r158 4 29 37.3796 $w=2.45e-07 $l=2.58612e-07 $layer=POLY_cond $X=4.77 $Y=1.085
+ $X2=4.58 $Y2=1.247
r159 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.77 $Y=1.085
+ $X2=4.77 $Y2=0.56
r160 1 29 10.0521 $w=1.8e-07 $l=1.63e-07 $layer=POLY_cond $X=4.58 $Y=1.41
+ $X2=4.58 $Y2=1.247
r161 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.58 $Y=1.41
+ $X2=4.58 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A 1 3 4 6 7 13
c38 1 0 1.94872e-19 $X=8.63 $Y=1.41
r39 7 13 5.53173 $w=2.48e-07 $l=1.2e-07 $layer=LI1_cond $X=8.515 $Y=1.2
+ $X2=8.395 $Y2=1.2
r40 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.525
+ $Y=1.16 $X2=8.525 $Y2=1.16
r41 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=8.655 $Y=0.995
+ $X2=8.56 $Y2=1.16
r42 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.655 $Y=0.995
+ $X2=8.655 $Y2=0.555
r43 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=8.63 $Y=1.41
+ $X2=8.56 $Y2=1.16
r44 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.63 $Y=1.41 $X2=8.63
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_1050_365# 1 2 3 4 13 15 16 18 21 23 27 28
+ 29 30 36 37 40 43 44
c130 30 0 1.07404e-19 $X=9.015 $Y=1.495
c131 13 0 3.96944e-20 $X=9.1 $Y=1.41
r132 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.385 $Y=0.51
+ $X2=8.385 $Y2=0.51
r133 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.425 $Y=0.51
+ $X2=5.425 $Y2=0.51
r134 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.57 $Y=0.51
+ $X2=5.425 $Y2=0.51
r135 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.24 $Y=0.51
+ $X2=8.385 $Y2=0.51
r136 36 37 3.30445 $w=1.4e-07 $l=2.67e-06 $layer=MET1_cond $X=8.24 $Y=0.51
+ $X2=5.57 $Y2=0.51
r137 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.075
+ $Y=1.16 $X2=9.075 $Y2=1.16
r138 32 34 17.9567 $w=2.31e-07 $l=3.4e-07 $layer=LI1_cond $X=9.07 $Y=0.82
+ $X2=9.07 $Y2=1.16
r139 31 44 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=8.415 $Y=0.735
+ $X2=8.415 $Y2=0.51
r140 29 34 9.58904 $w=2.31e-07 $l=1.90526e-07 $layer=LI1_cond $X=9.015 $Y=1.325
+ $X2=9.07 $Y2=1.16
r141 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.015 $Y=1.325
+ $X2=9.015 $Y2=1.495
r142 28 31 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.56 $Y=0.82
+ $X2=8.415 $Y2=0.735
r143 27 32 2.5345 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.93 $Y=0.82 $X2=9.07
+ $Y2=0.82
r144 27 28 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=8.93 $Y=0.82
+ $X2=8.56 $Y2=0.82
r145 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.93 $Y=1.6
+ $X2=9.015 $Y2=1.495
r146 23 25 28.2554 $w=2.08e-07 $l=5.35e-07 $layer=LI1_cond $X=8.93 $Y=1.6
+ $X2=8.395 $Y2=1.6
r147 19 40 3.61456 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.375 $Y=0.595
+ $X2=5.375 $Y2=0.43
r148 19 21 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.375 $Y=0.595
+ $X2=5.375 $Y2=1.94
r149 16 35 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=9.125 $Y=0.995
+ $X2=9.1 $Y2=1.16
r150 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.125 $Y=0.995
+ $X2=9.125 $Y2=0.555
r151 13 35 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=9.1 $Y=1.41
+ $X2=9.1 $Y2=1.16
r152 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.1 $Y=1.41
+ $X2=9.1 $Y2=1.985
r153 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=8.165
+ $Y=1.645 $X2=8.395 $Y2=1.62
r154 3 21 600 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_PDIFF $count=1 $X=5.25
+ $Y=1.825 $X2=5.375 $Y2=1.94
r155 2 44 182 $w=1.7e-07 $l=4.85747e-07 $layer=licon1_NDIFF $count=1 $X=8.18
+ $Y=0.235 $X2=8.395 $Y2=0.625
r156 1 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.245 $X2=5.54 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%VPWR 1 2 3 4 13 15 17 21 25 28 31 34 36 52
+ 53 59 62
c107 4 0 1.07404e-19 $X=8.72 $Y=1.485
r108 62 63 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r109 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r110 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r111 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r112 49 50 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r113 47 50 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=8.51 $Y2=2.72
r114 47 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 46 49 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=8.51 $Y2=2.72
r116 46 47 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r117 44 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.51 $Y=2.72
+ $X2=4.345 $Y2=2.72
r118 44 46 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=4.51 $Y=2.72
+ $X2=4.83 $Y2=2.72
r119 43 63 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r121 40 43 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r122 40 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r123 39 42 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r125 37 59 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=1.292 $Y2=2.72
r126 37 39 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=1.61 $Y2=2.72
r127 36 62 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.18 $Y=2.72
+ $X2=4.345 $Y2=2.72
r128 36 42 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=4.18 $Y=2.72
+ $X2=3.91 $Y2=2.72
r129 34 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r130 34 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r131 32 52 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=9.035 $Y=2.72
+ $X2=9.43 $Y2=2.72
r132 31 49 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=8.65 $Y=2.72
+ $X2=8.51 $Y2=2.72
r133 31 32 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=8.842 $Y=2.72
+ $X2=9.035 $Y2=2.72
r134 28 31 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=8.842 $Y=2.36
+ $X2=8.842 $Y2=2.72
r135 23 62 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.345 $Y=2.635
+ $X2=4.345 $Y2=2.72
r136 23 25 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.345 $Y=2.635
+ $X2=4.345 $Y2=2.32
r137 19 59 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=1.292 $Y=2.635
+ $X2=1.292 $Y2=2.72
r138 19 21 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.292 $Y=2.635
+ $X2=1.292 $Y2=2.3
r139 18 56 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.217 $Y2=2.72
r140 17 59 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=1.125 $Y=2.72
+ $X2=1.292 $Y2=2.72
r141 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.125 $Y=2.72
+ $X2=0.435 $Y2=2.72
r142 13 56 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.217 $Y2=2.72
r143 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=2.3
r144 4 28 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=8.72
+ $Y=1.485 $X2=8.865 $Y2=2.36
r145 3 25 600 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=4.22
+ $Y=1.485 $X2=4.345 $Y2=2.32
r146 2 21 600 $w=1.7e-07 $l=9.22862e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.485 $X2=1.295 $Y2=2.3
r147 1 15 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%X 1 2 11 13 15 21 24 25
r45 24 25 5.3331 $w=5.73e-07 $l=1.8e-07 $layer=LI1_cond $X=0.617 $Y=1.62
+ $X2=0.617 $Y2=1.44
r46 21 28 7.53038 $w=5.73e-07 $l=1.75e-07 $layer=LI1_cond $X=0.617 $Y=1.87
+ $X2=0.617 $Y2=2.045
r47 21 24 5.20034 $w=5.73e-07 $l=2.5e-07 $layer=LI1_cond $X=0.617 $Y=1.87
+ $X2=0.617 $Y2=1.62
r48 13 15 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=0.805 $Y=0.66
+ $X2=0.805 $Y2=0.56
r49 11 28 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.78 $Y=2.3
+ $X2=0.78 $Y2=2.045
r50 7 13 12.7421 $w=2.63e-07 $l=2.93e-07 $layer=LI1_cond $X=0.512 $Y=0.792
+ $X2=0.805 $Y2=0.792
r51 7 25 16.2605 $w=3.63e-07 $l=5.15e-07 $layer=LI1_cond $X=0.512 $Y=0.925
+ $X2=0.512 $Y2=1.44
r52 2 24 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=1.62
r53 2 11 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=2.3
r54 1 15 182 $w=1.7e-07 $l=4.16983e-07 $layer=licon1_NDIFF $count=1 $X=0.555
+ $Y=0.235 $X2=0.765 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_465_325# 1 2 3 4 13 18 21 23 25 27 30 32
+ 33 35 37 38 39 45 49
c147 35 0 8.91061e-20 $X=7.675 $Y=0.38
r148 48 49 11.956 $w=2.5e-07 $l=2.45e-07 $layer=LI1_cond $X=3.585 $Y=1.535
+ $X2=3.83 $Y2=1.535
r149 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.395 $Y=1.53
+ $X2=6.395 $Y2=1.53
r150 42 49 5.612 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=3.945 $Y=1.535
+ $X2=3.83 $Y2=1.535
r151 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.945 $Y=1.53
+ $X2=3.945 $Y2=1.53
r152 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.09 $Y=1.53
+ $X2=3.945 $Y2=1.53
r153 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.25 $Y=1.53
+ $X2=6.395 $Y2=1.53
r154 38 39 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=6.25 $Y=1.53
+ $X2=4.09 $Y2=1.53
r155 33 37 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.38 $Y2=0.36
r156 33 35 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=7.59 $Y=0.36
+ $X2=7.675 $Y2=0.36
r157 32 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.87 $Y=0.34
+ $X2=7.38 $Y2=0.34
r158 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.785 $Y=0.425
+ $X2=6.87 $Y2=0.34
r159 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.785 $Y=0.425
+ $X2=6.785 $Y2=1.445
r160 28 46 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.455 $Y=1.53
+ $X2=6.247 $Y2=1.53
r161 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.7 $Y=1.53
+ $X2=6.785 $Y2=1.445
r162 27 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.7 $Y=1.53
+ $X2=6.455 $Y2=1.53
r163 23 46 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=6.247 $Y=1.615
+ $X2=6.247 $Y2=1.53
r164 23 25 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=6.247 $Y=1.615
+ $X2=6.247 $Y2=1.62
r165 19 49 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.83 $Y=1.375
+ $X2=3.83 $Y2=1.535
r166 19 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.83 $Y=1.375
+ $X2=3.83 $Y2=0.76
r167 17 48 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.585 $Y=1.695
+ $X2=3.585 $Y2=1.535
r168 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.585 $Y=1.695
+ $X2=3.585 $Y2=1.895
r169 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.5 $Y=1.98
+ $X2=3.585 $Y2=1.895
r170 13 15 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.5 $Y=1.98
+ $X2=2.51 $Y2=1.98
r171 4 25 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.865
+ $Y=1.485 $X2=6.215 $Y2=1.62
r172 3 15 600 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=1 $X=2.325
+ $Y=1.625 $X2=2.51 $Y2=1.98
r173 2 35 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.48
+ $Y=0.245 $X2=7.675 $Y2=0.38
r174 1 21 182 $w=1.7e-07 $l=6.65507e-07 $layer=licon1_NDIFF $count=1 $X=3.485
+ $Y=0.245 $X2=3.83 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_483_49# 1 2 3 4 13 18 19 20 22 23 24 26
+ 28 29 32 33 34 36 39 43 48 52 54 55 57
r187 55 56 17.995 $w=2e-07 $l=2.95e-07 $layer=LI1_cond $X=5.715 $Y=0.772
+ $X2=6.01 $Y2=0.772
r188 50 52 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.17 $Y=1.12
+ $X2=4.285 $Y2=1.12
r189 46 48 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.81 $Y=2.32
+ $X2=3.925 $Y2=2.32
r190 41 56 1.68994 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=6.01 $Y=0.655
+ $X2=6.01 $Y2=0.772
r191 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=6.01 $Y=0.655
+ $X2=6.01 $Y2=0.545
r192 37 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.8 $Y=2.36
+ $X2=5.715 $Y2=2.36
r193 37 39 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=5.8 $Y=2.36
+ $X2=7.83 $Y2=2.36
r194 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=2.275
+ $X2=5.715 $Y2=2.36
r195 35 55 1.68994 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=5.715 $Y=0.89
+ $X2=5.715 $Y2=0.772
r196 35 36 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.715 $Y=0.89
+ $X2=5.715 $Y2=2.275
r197 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=2.36
+ $X2=5.715 $Y2=2.36
r198 33 34 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.63 $Y=2.36
+ $X2=5.115 $Y2=2.36
r199 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.03 $Y=2.275
+ $X2=5.115 $Y2=2.36
r200 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.03 $Y=2.065
+ $X2=5.03 $Y2=2.275
r201 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=1.98
+ $X2=4.285 $Y2=1.98
r202 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.945 $Y=1.98
+ $X2=5.03 $Y2=2.065
r203 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.945 $Y=1.98
+ $X2=4.37 $Y2=1.98
r204 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=1.895
+ $X2=4.285 $Y2=1.98
r205 27 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=1.205
+ $X2=4.285 $Y2=1.12
r206 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.285 $Y=1.205
+ $X2=4.285 $Y2=1.895
r207 26 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=1.035
+ $X2=4.17 $Y2=1.12
r208 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.17 $Y=0.425
+ $X2=4.17 $Y2=1.035
r209 23 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.2 $Y=1.98
+ $X2=4.285 $Y2=1.98
r210 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.2 $Y=1.98
+ $X2=4.01 $Y2=1.98
r211 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.925 $Y=2.235
+ $X2=3.925 $Y2=2.32
r212 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.925 $Y=2.065
+ $X2=4.01 $Y2=1.98
r213 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.925 $Y=2.065
+ $X2=3.925 $Y2=2.235
r214 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=4.17 $Y2=0.425
r215 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.085 $Y=0.34
+ $X2=3.575 $Y2=0.34
r216 17 20 6.93832 $w=1.7e-07 $l=1.44375e-07 $layer=LI1_cond $X=3.467 $Y=0.425
+ $X2=3.575 $Y2=0.34
r217 17 18 12.3285 $w=2.13e-07 $l=2.3e-07 $layer=LI1_cond $X=3.467 $Y=0.425
+ $X2=3.467 $Y2=0.655
r218 13 18 6.93832 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.36 $Y=0.74
+ $X2=3.467 $Y2=0.655
r219 13 15 52.8449 $w=1.68e-07 $l=8.1e-07 $layer=LI1_cond $X=3.36 $Y=0.74
+ $X2=2.55 $Y2=0.74
r220 4 39 600 $w=1.7e-07 $l=8.21995e-07 $layer=licon1_PDIFF $count=1 $X=7.6
+ $Y=1.645 $X2=7.83 $Y2=2.36
r221 3 46 600 $w=1.7e-07 $l=8.70373e-07 $layer=licon1_PDIFF $count=1 $X=3.415
+ $Y=1.625 $X2=3.81 $Y2=2.32
r222 2 43 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.875
+ $Y=0.245 $X2=6.01 $Y2=0.545
r223 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.245 $X2=2.55 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%A_1335_297# 1 2 3 4 15 18 23 26 29 31 36
r66 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.335 $Y=0.42
+ $X2=9.465 $Y2=0.42
r67 28 29 17.0922 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.34 $Y=1.99
+ $X2=9.015 $Y2=1.99
r68 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.465 $Y=1.875
+ $X2=9.465 $Y2=1.99
r69 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.465 $Y=0.585
+ $X2=9.465 $Y2=0.42
r70 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.465 $Y=0.585
+ $X2=9.465 $Y2=1.875
r71 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=9.402 $Y=1.99
+ $X2=9.465 $Y2=1.99
r72 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=9.402 $Y=1.99
+ $X2=9.34 $Y2=1.99
r73 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=9.402 $Y=2.105
+ $X2=9.402 $Y2=2.3
r74 20 29 113.519 $w=1.68e-07 $l=1.74e-06 $layer=LI1_cond $X=7.275 $Y=2.02
+ $X2=9.015 $Y2=2.02
r75 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.21 $Y=2.02
+ $X2=7.275 $Y2=2.02
r76 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.125 $Y=1.935
+ $X2=7.21 $Y2=2.02
r77 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=7.125 $Y=1.935
+ $X2=7.125 $Y2=0.76
r78 4 28 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.485 $X2=9.34 $Y2=1.96
r79 4 23 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=9.19
+ $Y=1.485 $X2=9.34 $Y2=2.3
r80 3 20 600 $w=1.7e-07 $l=8.25227e-07 $layer=licon1_PDIFF $count=1 $X=6.675
+ $Y=1.485 $X2=7.275 $Y2=2.02
r81 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.2
+ $Y=0.235 $X2=9.335 $Y2=0.42
r82 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=6.685
+ $Y=0.245 $X2=7.125 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_2%VGND 1 2 3 4 13 15 17 21 25 29 32 33 35 36
+ 37 53 54 60
c115 29 0 3.96944e-20 $X=8.865 $Y=0.4
r116 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r117 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r118 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=9.43
+ $Y2=0
r119 50 51 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r120 48 51 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.83 $Y=0 $X2=8.51
+ $Y2=0
r121 47 50 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=8.51
+ $Y2=0
r122 47 48 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r123 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r124 44 45 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r125 42 45 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=4.37 $Y2=0
r126 42 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r127 41 44 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.61 $Y=0 $X2=4.37
+ $Y2=0
r128 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r129 39 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.23
+ $Y2=0
r130 39 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.355 $Y=0
+ $X2=1.61 $Y2=0
r131 37 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r132 37 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r133 35 50 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=8.78 $Y=0 $X2=8.51
+ $Y2=0
r134 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.78 $Y=0 $X2=8.865
+ $Y2=0
r135 34 53 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=8.95 $Y=0 $X2=9.43
+ $Y2=0
r136 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.95 $Y=0 $X2=8.865
+ $Y2=0
r137 32 44 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.37
+ $Y2=0
r138 32 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.425 $Y=0 $X2=4.51
+ $Y2=0
r139 31 47 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.595 $Y=0
+ $X2=4.83 $Y2=0
r140 31 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.595 $Y=0 $X2=4.51
+ $Y2=0
r141 27 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.865 $Y=0.085
+ $X2=8.865 $Y2=0
r142 27 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.865 $Y=0.085
+ $X2=8.865 $Y2=0.4
r143 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=0.085
+ $X2=4.51 $Y2=0
r144 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.51 $Y=0.085
+ $X2=4.51 $Y2=0.36
r145 19 60 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r146 19 21 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.36
r147 18 57 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=0
+ $X2=0.217 $Y2=0
r148 17 60 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.23
+ $Y2=0
r149 17 18 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.105 $Y=0
+ $X2=0.435 $Y2=0
r150 13 57 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.217 $Y2=0
r151 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.38
r152 4 29 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=8.73
+ $Y=0.235 $X2=8.865 $Y2=0.4
r153 3 25 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.345
+ $Y=0.235 $X2=4.51 $Y2=0.36
r154 2 21 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=1.055
+ $Y=0.235 $X2=1.27 $Y2=0.36
r155 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

