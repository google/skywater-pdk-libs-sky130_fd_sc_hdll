* File: sky130_fd_sc_hdll__or4_1.pex.spice
* Created: Thu Aug 27 19:24:48 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4_1%D 1 3 6 8 9 15
r29 15 16 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 13 15 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 8 9 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.265 $Y=0.85
+ $X2=0.265 $Y2=1.16
r33 4 16 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r35 1 15 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%C 1 3 6 8 10 22 26
r39 18 26 4.14769 $w=6.18e-07 $l=2.15e-07 $layer=LI1_cond $X=0.94 $Y=1.305
+ $X2=1.155 $Y2=1.305
r40 18 22 2.9902 $w=6.18e-07 $l=1.55e-07 $layer=LI1_cond $X=0.94 $Y=1.305
+ $X2=0.785 $Y2=1.305
r41 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r42 10 26 1.92916 $w=6.18e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=1.305
+ $X2=1.155 $Y2=1.305
r43 8 22 0.771663 $w=6.18e-07 $l=4e-08 $layer=LI1_cond $X=0.745 $Y=1.305
+ $X2=0.785 $Y2=1.305
r44 4 17 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=0.965 $Y2=1.16
r45 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.05 $Y=0.995 $X2=1.05
+ $Y2=0.475
r46 1 17 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=0.965 $Y2=1.16
r47 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=1.025 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%B 1 2 3 4 6 9 10 11 12 13 19 24 27
c42 2 0 8.49032e-20 $X=1.445 $Y=1.31
r43 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.48
+ $Y=2.31 $X2=1.48 $Y2=2.31
r44 13 19 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.255 $Y=2.27
+ $X2=1.48 $Y2=2.27
r45 13 27 3.97394 $w=2.88e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=2.27
+ $X2=1.155 $Y2=2.27
r46 12 27 16.2932 $w=2.88e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=2.27
+ $X2=1.155 $Y2=2.27
r47 12 24 1.98697 $w=2.88e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=2.27
+ $X2=0.695 $Y2=2.27
r48 11 24 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=2.27
+ $X2=0.695 $Y2=2.27
r49 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.47 $Y=0.475 $X2=1.47
+ $Y2=0.76
r50 4 18 56.6054 $w=2.52e-07 $l=2.91976e-07 $layer=POLY_cond $X=1.445 $Y=2.035
+ $X2=1.48 $Y2=2.31
r51 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.445 $Y=2.035
+ $X2=1.445 $Y2=1.695
r52 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.445 $Y=1.41
+ $X2=1.445 $Y2=1.695
r53 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.445 $Y=1.31 $X2=1.445
+ $Y2=1.41
r54 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.445 $Y=0.86 $X2=1.445
+ $Y2=0.76
r55 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=1.445 $Y=0.86 $X2=1.445
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%A 1 3 6 8 12 14
r40 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.93
+ $Y=1.16 $X2=1.93 $Y2=1.16
r41 8 12 5.76222 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.93 $Y2=1.16
r42 8 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.615 $Y2=1.16
r43 4 11 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.93 $Y2=1.16
r44 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.99 $Y=0.995 $X2=1.99
+ $Y2=0.475
r45 1 11 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.93 $Y2=1.16
r46 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%A_27_297# 1 2 3 10 12 13 15 16 20 22 23 26
+ 28 30 35 37 41 42 47 49
c97 47 0 1.16645e-19 $X=2.47 $Y=1.16
c98 35 0 1.07404e-19 $X=2.35 $Y=1.495
r99 47 50 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=1.16
+ $X2=2.41 $Y2=1.325
r100 47 49 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=2.41 $Y=1.16
+ $X2=2.41 $Y2=0.995
r101 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.47
+ $Y=1.16 $X2=2.47 $Y2=1.16
r102 42 44 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.745 $Y=1.58
+ $X2=1.745 $Y2=1.87
r103 37 39 6.66256 $w=3.18e-07 $l=1.85e-07 $layer=LI1_cond $X=0.25 $Y=1.685
+ $X2=0.25 $Y2=1.87
r104 35 50 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.35 $Y=1.495
+ $X2=2.35 $Y2=1.325
r105 32 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.35 $Y=0.825
+ $X2=2.35 $Y2=0.995
r106 31 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=1.58
+ $X2=1.745 $Y2=1.58
r107 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=1.58
+ $X2=2.35 $Y2=1.495
r108 30 31 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.265 $Y=1.58
+ $X2=1.83 $Y2=1.58
r109 29 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=0.74
+ $X2=1.73 $Y2=0.74
r110 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=0.74
+ $X2=2.35 $Y2=0.825
r111 28 29 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.265 $Y=0.74
+ $X2=1.815 $Y2=0.74
r112 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.655
+ $X2=1.73 $Y2=0.74
r113 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.73 $Y=0.655
+ $X2=1.73 $Y2=0.47
r114 22 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.74
+ $X2=1.73 $Y2=0.74
r115 22 23 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.645 $Y=0.74
+ $X2=0.845 $Y2=0.74
r116 18 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.845 $Y2=0.74
r117 18 20 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.76 $Y2=0.47
r118 17 39 4.44149 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.41 $Y=1.87
+ $X2=0.25 $Y2=1.87
r119 16 44 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=1.745 $Y2=1.87
r120 16 17 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=0.41 $Y2=1.87
r121 13 48 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.53 $Y=0.995
+ $X2=2.47 $Y2=1.16
r122 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.53 $Y=0.995
+ $X2=2.53 $Y2=0.56
r123 10 48 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.47 $Y2=1.16
r124 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.985
r125 3 37 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.685
r126 2 26 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.265 $X2=1.73 $Y2=0.47
r127 1 20 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=0.76 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%VPWR 1 6 9 10 11 21 22
c24 1 0 1.07404e-19 $X=2.055 $Y=1.485
r25 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r26 19 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r27 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 14 18 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r29 11 19 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r30 11 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r31 9 18 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 9 10 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.115 $Y=2.72 $X2=2.255
+ $Y2=2.72
r33 8 21 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.99 $Y2=2.72
r34 8 10 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.395 $Y=2.72 $X2=2.255
+ $Y2=2.72
r35 4 10 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2.72
r36 4 6 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2
r37 1 6 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=1.485 $X2=2.265 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%X 1 2 12 14 15 16
r19 14 16 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.94 $Y=1.63
+ $X2=2.94 $Y2=1.845
r20 14 15 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.94 $Y=1.63
+ $X2=2.94 $Y2=1.495
r21 10 12 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=2.89 $Y=0.587 $X2=2.99
+ $Y2=0.587
r22 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.99 $Y=0.76 $X2=2.99
+ $Y2=0.587
r23 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.99 $Y=0.76
+ $X2=2.99 $Y2=1.495
r24 2 16 300 $w=1.7e-07 $l=4.85592e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.485 $X2=2.89 $Y2=1.845
r25 1 10 182 $w=1.7e-07 $l=4.76655e-07 $layer=licon1_NDIFF $count=1 $X=2.605
+ $Y=0.235 $X2=2.89 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_1%VGND 1 2 3 10 12 16 18 20 25 32 33 39 43
r52 43 46 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.2
+ $Y2=0.4
r53 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r54 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r56 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r57 30 43 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.2
+ $Y2=0
r58 30 32 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.99
+ $Y2=0
r59 29 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r60 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r61 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r62 26 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.235
+ $Y2=0
r63 26 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.61
+ $Y2=0
r64 25 43 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.2
+ $Y2=0
r65 25 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.61
+ $Y2=0
r66 24 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r67 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r68 21 36 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r69 21 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r70 20 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.235
+ $Y2=0
r71 20 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.69
+ $Y2=0
r72 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r73 18 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r74 14 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r75 14 16 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.4
r76 10 36 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r77 10 12 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.5
r78 3 46 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.265 $X2=2.25 $Y2=0.4
r79 2 16 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.265 $X2=1.26 $Y2=0.4
r80 1 12 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends

