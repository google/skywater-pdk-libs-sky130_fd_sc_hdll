* File: sky130_fd_sc_hdll__clkinvlp_4.pxi.spice
* Created: Thu Aug 27 19:03:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_4%A N_A_M1000_g N_A_M1003_g N_A_M1001_g
+ N_A_M1002_g N_A_M1005_g N_A_M1006_g N_A_M1004_g N_A_M1007_g A A N_A_c_36_n
+ PM_SKY130_FD_SC_HDLL__CLKINVLP_4%A
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VPWR N_VPWR_M1000_s N_VPWR_M1002_s
+ N_VPWR_M1007_s N_VPWR_c_97_n N_VPWR_c_98_n N_VPWR_c_99_n N_VPWR_c_100_n
+ N_VPWR_c_101_n N_VPWR_c_102_n N_VPWR_c_103_n VPWR N_VPWR_c_104_n N_VPWR_c_96_n
+ PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_4%Y N_Y_M1001_s N_Y_M1000_d N_Y_M1006_d
+ N_Y_c_135_n N_Y_c_136_n Y Y Y Y Y Y Y N_Y_c_152_n
+ PM_SKY130_FD_SC_HDLL__CLKINVLP_4%Y
x_PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VGND N_VGND_M1003_d N_VGND_M1004_d
+ N_VGND_c_171_n N_VGND_c_172_n N_VGND_c_173_n N_VGND_c_174_n N_VGND_c_175_n
+ VGND N_VGND_c_176_n N_VGND_c_177_n PM_SKY130_FD_SC_HDLL__CLKINVLP_4%VGND
cc_1 VNB N_A_M1003_g 0.0242965f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.51
cc_2 VNB N_A_M1001_g 0.018421f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=0.51
cc_3 VNB N_A_M1005_g 0.0202106f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.51
cc_4 VNB N_A_M1004_g 0.0282192f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=0.51
cc_5 VNB A 0.0216425f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_6 VNB N_A_c_36_n 0.126945f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=1.16
cc_7 VNB N_VPWR_c_96_n 0.117919f $X=-0.19 $Y=-0.24 $X2=1.56 $Y2=1.16
cc_8 VNB Y 0.00354801f $X=-0.19 $Y=-0.24 $X2=1.56 $Y2=1.985
cc_9 VNB N_VGND_c_171_n 0.0103065f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.51
cc_10 VNB N_VGND_c_172_n 0.0162274f $X=-0.19 $Y=-0.24 $X2=0.835 $Y2=0.995
cc_11 VNB N_VGND_c_173_n 0.0239037f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.325
cc_12 VNB N_VGND_c_174_n 0.0322153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_175_n 0.00503814f $X=-0.19 $Y=-0.24 $X2=1.265 $Y2=0.995
cc_14 VNB N_VGND_c_176_n 0.026328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_177_n 0.188128f $X=-0.19 $Y=-0.24 $X2=2.08 $Y2=1.325
cc_16 VPB N_A_M1000_g 0.0313004f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.985
cc_17 VPB N_A_M1002_g 0.0242818f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.985
cc_18 VPB N_A_M1006_g 0.0239892f $X=-0.19 $Y=1.305 $X2=1.56 $Y2=1.985
cc_19 VPB N_A_M1007_g 0.0316355f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.985
cc_20 VPB A 0.00394216f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_21 VPB N_A_c_36_n 0.0212686f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.16
cc_22 VPB N_VPWR_c_97_n 0.0102436f $X=-0.19 $Y=1.305 $X2=0.835 $Y2=0.51
cc_23 VPB N_VPWR_c_98_n 0.0412701f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_VPWR_c_99_n 0.00471426f $X=-0.19 $Y=1.305 $X2=1.265 $Y2=0.51
cc_25 VPB N_VPWR_c_100_n 0.0156949f $X=-0.19 $Y=1.305 $X2=1.56 $Y2=1.985
cc_26 VPB N_VPWR_c_101_n 0.055579f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_102_n 0.0198788f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.325
cc_28 VPB N_VPWR_c_103_n 0.0040505f $X=-0.19 $Y=1.305 $X2=2.08 $Y2=1.985
cc_29 VPB N_VPWR_c_104_n 0.0199729f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_30 VPB N_VPWR_c_96_n 0.0495615f $X=-0.19 $Y=1.305 $X2=1.56 $Y2=1.16
cc_31 N_A_M1000_g N_VPWR_c_98_n 0.0224351f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_32 N_A_M1002_g N_VPWR_c_98_n 9.0909e-19 $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_33 A N_VPWR_c_98_n 0.025424f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_34 N_A_c_36_n N_VPWR_c_98_n 0.00196424f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_35 N_A_M1002_g N_VPWR_c_99_n 0.00320986f $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_36 N_A_M1006_g N_VPWR_c_99_n 0.0219833f $X=1.56 $Y=1.985 $X2=0 $Y2=0
cc_37 N_A_M1007_g N_VPWR_c_99_n 0.00116152f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_38 N_A_c_36_n N_VPWR_c_99_n 0.00254056f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_39 N_A_M1007_g N_VPWR_c_101_n 0.00545629f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_40 N_A_M1000_g N_VPWR_c_102_n 0.00817093f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_41 N_A_M1002_g N_VPWR_c_102_n 0.00931616f $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_42 N_A_M1006_g N_VPWR_c_104_n 0.00832274f $X=1.56 $Y=1.985 $X2=0 $Y2=0
cc_43 N_A_M1007_g N_VPWR_c_104_n 0.00931616f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_VPWR_c_96_n 0.0129363f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_45 N_A_M1002_g N_VPWR_c_96_n 0.015569f $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_46 N_A_M1006_g N_VPWR_c_96_n 0.0133061f $X=1.56 $Y=1.985 $X2=0 $Y2=0
cc_47 N_A_M1007_g N_VPWR_c_96_n 0.0166452f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_48 N_A_c_36_n N_Y_c_135_n 0.0920753f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A_M1002_g N_Y_c_136_n 8.62388e-19 $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_50 N_A_M1006_g N_Y_c_136_n 0.0219217f $X=1.56 $Y=1.985 $X2=0 $Y2=0
cc_51 N_A_M1007_g N_Y_c_136_n 0.0234474f $X=2.08 $Y=1.985 $X2=0 $Y2=0
cc_52 N_A_c_36_n N_Y_c_136_n 0.00572328f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_53 N_A_M1000_g Y 0.027701f $X=0.52 $Y=1.985 $X2=0 $Y2=0
cc_54 N_A_M1002_g Y 0.019344f $X=1.04 $Y=1.985 $X2=0 $Y2=0
cc_55 N_A_M1006_g Y 9.23721e-19 $X=1.56 $Y=1.985 $X2=0 $Y2=0
cc_56 A Y 0.00212432f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_c_36_n Y 0.00499639f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_M1003_g Y 0.00174362f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_59 N_A_M1001_g Y 0.00853887f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_60 N_A_M1005_g Y 0.00491562f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_61 A Y 0.0187987f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_c_36_n Y 0.00242316f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_63 A Y 0.0213899f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_c_36_n Y 0.013871f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_65 N_A_M1001_g N_Y_c_152_n 0.0105146f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_66 N_A_c_36_n N_Y_c_152_n 0.00254697f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_67 A N_VGND_M1003_d 0.00242856f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_68 N_A_M1003_g N_VGND_c_172_n 0.00980416f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_69 N_A_M1001_g N_VGND_c_172_n 0.00147043f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_70 A N_VGND_c_172_n 0.0232502f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_71 N_A_c_36_n N_VGND_c_172_n 0.00113123f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_M1005_g N_VGND_c_173_n 0.00288319f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_73 N_A_M1004_g N_VGND_c_173_n 0.018424f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_74 N_A_c_36_n N_VGND_c_173_n 0.00770088f $X=2.08 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1003_g N_VGND_c_174_n 0.00486043f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_76 N_A_M1001_g N_VGND_c_174_n 0.00357877f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_77 N_A_M1005_g N_VGND_c_174_n 0.00585385f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_VGND_c_174_n 0.00486043f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_79 N_A_M1003_g N_VGND_c_177_n 0.00809891f $X=0.475 $Y=0.51 $X2=0 $Y2=0
cc_80 N_A_M1001_g N_VGND_c_177_n 0.00511556f $X=0.835 $Y=0.51 $X2=0 $Y2=0
cc_81 N_A_M1005_g N_VGND_c_177_n 0.0106631f $X=1.265 $Y=0.51 $X2=0 $Y2=0
cc_82 N_A_M1004_g N_VGND_c_177_n 0.00809891f $X=1.625 $Y=0.51 $X2=0 $Y2=0
cc_83 A N_VGND_c_177_n 0.00163141f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_84 N_VPWR_c_96_n N_Y_M1000_d 0.00215201f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_85 N_VPWR_c_96_n N_Y_M1006_d 0.00215201f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_86 N_VPWR_c_99_n N_Y_c_135_n 0.0226618f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_87 N_VPWR_c_99_n N_Y_c_136_n 0.0663107f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_88 N_VPWR_c_101_n N_Y_c_136_n 0.0290915f $X=2.34 $Y=1.63 $X2=0 $Y2=0
cc_89 N_VPWR_c_104_n N_Y_c_136_n 0.0189039f $X=2.225 $Y=2.72 $X2=0 $Y2=0
cc_90 N_VPWR_c_96_n N_Y_c_136_n 0.0122217f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_91 N_VPWR_c_98_n Y 0.0680999f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_92 N_VPWR_c_99_n Y 0.0292203f $X=1.3 $Y=1.63 $X2=0 $Y2=0
cc_93 N_VPWR_c_102_n Y 0.0195857f $X=1.185 $Y=2.72 $X2=0 $Y2=0
cc_94 N_VPWR_c_96_n Y 0.0125611f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_95 N_Y_c_135_n N_VGND_c_173_n 0.0186638f $X=1.655 $Y=1.155 $X2=0 $Y2=0
cc_96 N_Y_c_152_n N_VGND_c_174_n 0.0327013f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_97 N_Y_M1001_s N_VGND_c_177_n 0.00311651f $X=0.91 $Y=0.235 $X2=0 $Y2=0
cc_98 N_Y_c_152_n N_VGND_c_177_n 0.0205935f $X=1.05 $Y=0.445 $X2=0 $Y2=0
cc_99 Y A_110_47# 2.78895e-19 $X=0.66 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_100 N_Y_c_152_n A_110_47# 0.0011988f $X=1.05 $Y=0.445 $X2=-0.19 $Y2=-0.24
cc_101 N_VGND_c_177_n A_110_47# 0.00358776f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_102 N_VGND_c_177_n A_268_47# 0.00897657f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
