* File: sky130_fd_sc_hdll__o2bb2ai_4.pex.spice
* Created: Wed Sep  2 08:46:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A2_N 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 44
c65 22 0 1.98558e-19 $X=1.95 $Y=0.995
r66 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r67 37 39 21.379 $w=3.72e-07 $l=1.65e-07 $layer=POLY_cond $X=1.76 $Y=1.202
+ $X2=1.925 $Y2=1.202
r68 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.76
+ $Y=1.16 $X2=1.76 $Y2=1.16
r69 35 37 39.5188 $w=3.72e-07 $l=3.05e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.76 $Y2=1.202
r70 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r71 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.43 $Y2=1.202
r72 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r73 31 44 29.0476 $w=2.08e-07 $l=5.5e-07 $layer=LI1_cond $X=0.59 $Y=1.18
+ $X2=1.14 $Y2=1.18
r74 30 32 47.9409 $w=3.72e-07 $l=3.7e-07 $layer=POLY_cond $X=0.59 $Y=1.202
+ $X2=0.96 $Y2=1.202
r75 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r76 28 30 9.71774 $w=3.72e-07 $l=7.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.59 $Y2=1.202
r77 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r78 25 38 27.4632 $w=2.08e-07 $l=5.2e-07 $layer=LI1_cond $X=1.24 $Y=1.18
+ $X2=1.76 $Y2=1.18
r79 25 44 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=1.24 $Y=1.18 $X2=1.14
+ $Y2=1.18
r80 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r81 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r82 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r83 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r84 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r85 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r86 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r87 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=0.56
r88 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r89 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r90 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r91 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
r92 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r93 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r94 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r95 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A1_N 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 44
r81 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.805 $Y=1.202
+ $X2=3.83 $Y2=1.202
r82 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=3.63 $Y=1.202
+ $X2=3.805 $Y2=1.202
r83 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r84 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=3.335 $Y=1.202
+ $X2=3.63 $Y2=1.202
r85 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.202
+ $X2=3.335 $Y2=1.202
r86 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.865 $Y=1.202
+ $X2=3.31 $Y2=1.202
r87 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.84 $Y=1.202
+ $X2=2.865 $Y2=1.202
r88 31 44 27.4632 $w=2.08e-07 $l=5.2e-07 $layer=LI1_cond $X=2.46 $Y=1.18
+ $X2=2.98 $Y2=1.18
r89 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=2.46 $Y=1.202
+ $X2=2.84 $Y2=1.202
r90 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r91 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=2.395 $Y=1.202
+ $X2=2.46 $Y2=1.202
r92 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.202
+ $X2=2.395 $Y2=1.202
r93 25 38 18.4848 $w=2.08e-07 $l=3.5e-07 $layer=LI1_cond $X=3.28 $Y=1.18
+ $X2=3.63 $Y2=1.18
r94 25 44 15.8442 $w=2.08e-07 $l=3e-07 $layer=LI1_cond $X=3.28 $Y=1.18 $X2=2.98
+ $Y2=1.18
r95 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=1.202
r96 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.83 $Y=0.995
+ $X2=3.83 $Y2=0.56
r97 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.202
r98 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r99 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.202
r100 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r101 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=1.202
r102 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.31 $Y=0.995
+ $X2=3.31 $Y2=0.56
r103 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.202
r104 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r105 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=1.202
r106 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.84 $Y=0.995
+ $X2=2.84 $Y2=0.56
r107 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.202
r108 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r109 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=1.202
r110 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.37 $Y=0.995
+ $X2=2.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_113_47# 1 2 3 4 5 6 19 21 22 24 25 27
+ 28 30 31 33 34 36 37 39 40 42 44 45 49 51 52 55 57 61 63 67 69 73 75 78 79 84
+ 88 90 92 94 103
r162 103 104 7.14555 $w=3.71e-07 $l=5.5e-08 $layer=POLY_cond $X=6.175 $Y=1.202
+ $X2=6.23 $Y2=1.202
r163 100 101 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=5.705 $Y=1.202
+ $X2=5.71 $Y2=1.202
r164 99 100 60.4124 $w=3.71e-07 $l=4.65e-07 $layer=POLY_cond $X=5.24 $Y=1.202
+ $X2=5.705 $Y2=1.202
r165 98 99 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=5.235 $Y=1.202
+ $X2=5.24 $Y2=1.202
r166 95 96 0.649596 $w=3.71e-07 $l=5e-09 $layer=POLY_cond $X=4.765 $Y=1.202
+ $X2=4.77 $Y2=1.202
r167 85 103 18.8383 $w=3.71e-07 $l=1.45e-07 $layer=POLY_cond $X=6.03 $Y=1.202
+ $X2=6.175 $Y2=1.202
r168 85 101 41.5741 $w=3.71e-07 $l=3.2e-07 $layer=POLY_cond $X=6.03 $Y=1.202
+ $X2=5.71 $Y2=1.202
r169 84 85 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r170 82 98 48.7197 $w=3.71e-07 $l=3.75e-07 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=5.235 $Y2=1.202
r171 82 96 11.6927 $w=3.71e-07 $l=9e-08 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=4.77 $Y2=1.202
r172 81 84 61.7922 $w=2.08e-07 $l=1.17e-06 $layer=LI1_cond $X=4.86 $Y=1.18
+ $X2=6.03 $Y2=1.18
r173 81 82 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.86
+ $Y=1.16 $X2=4.86 $Y2=1.16
r174 79 81 28.7836 $w=2.08e-07 $l=5.45e-07 $layer=LI1_cond $X=4.315 $Y=1.18
+ $X2=4.86 $Y2=1.18
r175 77 79 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=4.23 $Y=1.285
+ $X2=4.315 $Y2=1.18
r176 77 78 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.23 $Y=1.285
+ $X2=4.23 $Y2=1.455
r177 76 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.695 $Y=1.54
+ $X2=3.57 $Y2=1.54
r178 75 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.145 $Y=1.54
+ $X2=4.23 $Y2=1.455
r179 75 76 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.145 $Y=1.54
+ $X2=3.695 $Y2=1.54
r180 71 94 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=1.625
+ $X2=3.57 $Y2=1.54
r181 71 73 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.57 $Y=1.625
+ $X2=3.57 $Y2=2.3
r182 70 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.755 $Y=1.54
+ $X2=2.63 $Y2=1.54
r183 69 94 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=3.57 $Y2=1.54
r184 69 70 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.445 $Y=1.54
+ $X2=2.755 $Y2=1.54
r185 65 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=1.625
+ $X2=2.63 $Y2=1.54
r186 65 67 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.63 $Y=1.625
+ $X2=2.63 $Y2=2.3
r187 64 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=1.54
+ $X2=1.69 $Y2=1.54
r188 63 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.505 $Y=1.54
+ $X2=2.63 $Y2=1.54
r189 63 64 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.505 $Y=1.54
+ $X2=1.815 $Y2=1.54
r190 59 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=1.54
r191 59 61 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.69 $Y=1.625
+ $X2=1.69 $Y2=2.3
r192 58 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=1.54
+ $X2=0.75 $Y2=1.54
r193 57 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.565 $Y=1.54
+ $X2=1.69 $Y2=1.54
r194 57 58 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.565 $Y=1.54
+ $X2=0.875 $Y2=1.54
r195 53 88 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.625
+ $X2=0.75 $Y2=1.54
r196 53 55 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=1.625
+ $X2=0.75 $Y2=2.3
r197 51 88 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.625 $Y=1.54
+ $X2=0.75 $Y2=1.54
r198 51 52 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.625 $Y=1.54
+ $X2=0.255 $Y2=1.54
r199 47 49 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=0.75 $Y=0.775
+ $X2=1.69 $Y2=0.775
r200 45 47 21.9407 $w=2.58e-07 $l=4.95e-07 $layer=LI1_cond $X=0.255 $Y=0.775
+ $X2=0.75 $Y2=0.775
r201 44 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.17 $Y=1.455
+ $X2=0.255 $Y2=1.54
r202 43 45 7.21222 $w=2.6e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.255 $Y2=0.775
r203 43 44 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=0.17 $Y=0.905
+ $X2=0.17 $Y2=1.455
r204 40 104 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.23 $Y2=1.202
r205 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.23 $Y=0.995
+ $X2=6.23 $Y2=0.56
r206 37 103 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.202
r207 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.175 $Y=1.41
+ $X2=6.175 $Y2=1.985
r208 34 101 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=1.202
r209 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.71 $Y=0.995
+ $X2=5.71 $Y2=0.56
r210 31 100 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.705 $Y=1.41
+ $X2=5.705 $Y2=1.202
r211 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.705 $Y=1.41
+ $X2=5.705 $Y2=1.985
r212 28 99 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=1.202
r213 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.24 $Y=0.995
+ $X2=5.24 $Y2=0.56
r214 25 98 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.235 $Y=1.41
+ $X2=5.235 $Y2=1.202
r215 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.235 $Y=1.41
+ $X2=5.235 $Y2=1.985
r216 22 96 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=1.202
r217 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.77 $Y=0.995
+ $X2=4.77 $Y2=0.56
r218 19 95 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.765 $Y=1.41
+ $X2=4.765 $Y2=1.202
r219 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.765 $Y=1.41
+ $X2=4.765 $Y2=1.985
r220 6 94 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.62
r221 6 73 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=2.3
r222 5 92 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.62
r223 5 67 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=2.3
r224 4 90 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r225 4 61 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2.3
r226 3 88 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.62
r227 3 55 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.3
r228 2 49 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.73
r229 1 47 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 45
c85 1 0 2.97897e-20 $X=7.14 $Y=0.995
r86 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.575 $Y=1.202
+ $X2=8.6 $Y2=1.202
r87 38 45 29.3117 $w=2.08e-07 $l=5.55e-07 $layer=LI1_cond $X=8.4 $Y=1.18
+ $X2=7.845 $Y2=1.18
r88 37 39 22.6747 $w=3.72e-07 $l=1.75e-07 $layer=POLY_cond $X=8.4 $Y=1.202
+ $X2=8.575 $Y2=1.202
r89 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.4 $Y=1.16
+ $X2=8.4 $Y2=1.16
r90 35 37 38.2231 $w=3.72e-07 $l=2.95e-07 $layer=POLY_cond $X=8.105 $Y=1.202
+ $X2=8.4 $Y2=1.202
r91 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.08 $Y=1.202
+ $X2=8.105 $Y2=1.202
r92 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=7.635 $Y=1.202
+ $X2=8.08 $Y2=1.202
r93 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.61 $Y=1.202
+ $X2=7.635 $Y2=1.202
r94 30 32 49.2366 $w=3.72e-07 $l=3.8e-07 $layer=POLY_cond $X=7.23 $Y=1.202
+ $X2=7.61 $Y2=1.202
r95 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=7.23
+ $Y=1.16 $X2=7.23 $Y2=1.16
r96 28 30 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=7.165 $Y=1.202
+ $X2=7.23 $Y2=1.202
r97 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.14 $Y=1.202
+ $X2=7.165 $Y2=1.202
r98 25 45 0.792208 $w=2.08e-07 $l=1.5e-08 $layer=LI1_cond $X=7.83 $Y=1.18
+ $X2=7.845 $Y2=1.18
r99 25 31 31.6883 $w=2.08e-07 $l=6e-07 $layer=LI1_cond $X=7.83 $Y=1.18 $X2=7.23
+ $Y2=1.18
r100 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.6 $Y=0.995
+ $X2=8.6 $Y2=1.202
r101 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.6 $Y=0.995
+ $X2=8.6 $Y2=0.56
r102 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.575 $Y=1.41
+ $X2=8.575 $Y2=1.202
r103 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.575 $Y=1.41
+ $X2=8.575 $Y2=1.985
r104 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.105 $Y=1.41
+ $X2=8.105 $Y2=1.202
r105 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.105 $Y=1.41
+ $X2=8.105 $Y2=1.985
r106 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.08 $Y=0.995
+ $X2=8.08 $Y2=1.202
r107 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.08 $Y=0.995
+ $X2=8.08 $Y2=0.56
r108 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.635 $Y=1.41
+ $X2=7.635 $Y2=1.202
r109 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.635 $Y=1.41
+ $X2=7.635 $Y2=1.985
r110 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.61 $Y=0.995
+ $X2=7.61 $Y2=1.202
r111 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.61 $Y=0.995
+ $X2=7.61 $Y2=0.56
r112 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.165 $Y=1.41
+ $X2=7.165 $Y2=1.202
r113 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.165 $Y=1.41
+ $X2=7.165 $Y2=1.985
r114 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.14 $Y=0.995
+ $X2=7.14 $Y2=1.202
r115 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.14 $Y=0.995
+ $X2=7.14 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 38 39 44
r75 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=10.455 $Y=1.202
+ $X2=10.48 $Y2=1.202
r76 37 39 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=10.25 $Y=1.202
+ $X2=10.455 $Y2=1.202
r77 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.25
+ $Y=1.16 $X2=10.25 $Y2=1.16
r78 35 37 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=9.985 $Y=1.202
+ $X2=10.25 $Y2=1.202
r79 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.96 $Y=1.202
+ $X2=9.985 $Y2=1.202
r80 33 34 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=9.515 $Y=1.202
+ $X2=9.96 $Y2=1.202
r81 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.49 $Y=1.202
+ $X2=9.515 $Y2=1.202
r82 31 44 40.4026 $w=2.08e-07 $l=7.65e-07 $layer=LI1_cond $X=9.08 $Y=1.18
+ $X2=9.845 $Y2=1.18
r83 30 32 53.1237 $w=3.72e-07 $l=4.1e-07 $layer=POLY_cond $X=9.08 $Y=1.202
+ $X2=9.49 $Y2=1.202
r84 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.08
+ $Y=1.16 $X2=9.08 $Y2=1.16
r85 28 30 4.53495 $w=3.72e-07 $l=3.5e-08 $layer=POLY_cond $X=9.045 $Y=1.202
+ $X2=9.08 $Y2=1.202
r86 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.02 $Y=1.202
+ $X2=9.045 $Y2=1.202
r87 25 38 19.2771 $w=2.08e-07 $l=3.65e-07 $layer=LI1_cond $X=9.885 $Y=1.18
+ $X2=10.25 $Y2=1.18
r88 25 44 2.11255 $w=2.08e-07 $l=4e-08 $layer=LI1_cond $X=9.885 $Y=1.18
+ $X2=9.845 $Y2=1.18
r89 22 40 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.48 $Y=0.995
+ $X2=10.48 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.48 $Y=0.995
+ $X2=10.48 $Y2=0.56
r91 19 39 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.455 $Y=1.41
+ $X2=10.455 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.455 $Y=1.41
+ $X2=10.455 $Y2=1.985
r93 16 35 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.985 $Y=1.41
+ $X2=9.985 $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.985 $Y=1.41
+ $X2=9.985 $Y2=1.985
r95 13 34 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.96 $Y=0.995
+ $X2=9.96 $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.96 $Y=0.995
+ $X2=9.96 $Y2=0.56
r97 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.515 $Y=1.41
+ $X2=9.515 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.515 $Y=1.41
+ $X2=9.515 $Y2=1.985
r99 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.49 $Y=0.995
+ $X2=9.49 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.49 $Y=0.995
+ $X2=9.49 $Y2=0.56
r101 4 28 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.045 $Y=1.41
+ $X2=9.045 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.045 $Y=1.41
+ $X2=9.045 $Y2=1.985
r103 1 27 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.02 $Y=0.995
+ $X2=9.02 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.02 $Y=0.995
+ $X2=9.02 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VPWR 1 2 3 4 5 6 7 8 9 28 30 32 36 38 42
+ 44 48 52 56 60 64 68 71 72 74 75 77 78 80 81 82 84 106 107 113 116 119 122 127
r150 122 123 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r151 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r152 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r153 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r154 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r155 114 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.23 $Y2=2.72
r156 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r157 110 127 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r158 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r159 104 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r160 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r161 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r162 100 101 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r163 98 101 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.97 $Y2=2.72
r164 97 100 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.97 $Y2=2.72
r165 97 98 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r166 95 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r167 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r168 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r169 92 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r170 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r171 89 122 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=4.285 $Y2=2.72
r172 89 91 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.655 $Y=2.72
+ $X2=5.29 $Y2=2.72
r173 88 123 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r174 88 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r175 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r176 85 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.225 $Y=2.72
+ $X2=3.1 $Y2=2.72
r177 85 87 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.225 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 84 122 14.0645 $w=1.7e-07 $l=3.7e-07 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=4.285 $Y2=2.72
r179 84 87 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.915 $Y=2.72
+ $X2=3.91 $Y2=2.72
r180 82 127 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r181 80 103 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=10.095 $Y=2.72
+ $X2=9.89 $Y2=2.72
r182 80 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.095 $Y=2.72
+ $X2=10.22 $Y2=2.72
r183 79 106 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=10.345 $Y=2.72
+ $X2=10.81 $Y2=2.72
r184 79 81 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=10.345 $Y=2.72
+ $X2=10.22 $Y2=2.72
r185 77 100 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=8.97 $Y2=2.72
r186 77 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.155 $Y=2.72
+ $X2=9.28 $Y2=2.72
r187 76 103 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=9.405 $Y=2.72
+ $X2=9.89 $Y2=2.72
r188 76 78 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.405 $Y=2.72
+ $X2=9.28 $Y2=2.72
r189 74 94 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.21 $Y2=2.72
r190 74 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.41 $Y2=2.72
r191 73 97 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.67 $Y2=2.72
r192 73 75 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.535 $Y=2.72
+ $X2=6.41 $Y2=2.72
r193 71 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r194 71 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.47 $Y2=2.72
r195 70 94 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=6.21 $Y2=2.72
r196 70 72 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.47 $Y2=2.72
r197 66 81 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=2.635
+ $X2=10.22 $Y2=2.72
r198 66 68 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=10.22 $Y=2.635
+ $X2=10.22 $Y2=1.96
r199 62 78 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.28 $Y2=2.72
r200 62 64 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.28 $Y=2.635
+ $X2=9.28 $Y2=1.96
r201 58 75 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=2.635
+ $X2=6.41 $Y2=2.72
r202 58 60 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=6.41 $Y=2.635
+ $X2=6.41 $Y2=1.96
r203 54 72 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.47 $Y=2.635
+ $X2=5.47 $Y2=2.72
r204 54 56 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.47 $Y=2.635
+ $X2=5.47 $Y2=1.96
r205 50 122 2.97738 $w=7.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.285 $Y=2.635
+ $X2=4.285 $Y2=2.72
r206 50 52 10.9102 $w=7.38e-07 $l=6.75e-07 $layer=LI1_cond $X=4.285 $Y=2.635
+ $X2=4.285 $Y2=1.96
r207 46 119 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.1 $Y=2.635
+ $X2=3.1 $Y2=2.72
r208 46 48 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=3.1 $Y=2.635
+ $X2=3.1 $Y2=1.96
r209 45 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.285 $Y=2.72
+ $X2=2.16 $Y2=2.72
r210 44 119 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.975 $Y=2.72
+ $X2=3.1 $Y2=2.72
r211 44 45 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.975 $Y=2.72
+ $X2=2.285 $Y2=2.72
r212 40 116 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=2.635
+ $X2=2.16 $Y2=2.72
r213 40 42 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=2.16 $Y=2.635
+ $X2=2.16 $Y2=1.96
r214 39 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.22 $Y2=2.72
r215 38 116 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=2.16 $Y2=2.72
r216 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=2.72
+ $X2=1.345 $Y2=2.72
r217 34 113 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r218 34 36 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=1.96
r219 33 110 3.96192 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r220 32 113 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=1.22 $Y2=2.72
r221 32 33 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.405 $Y2=2.72
r222 28 110 3.18124 $w=2.5e-07 $l=1.17707e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.202 $Y2=2.72
r223 28 30 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=1.96
r224 9 68 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.075
+ $Y=1.485 $X2=10.22 $Y2=1.96
r225 8 64 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.135
+ $Y=1.485 $X2=9.28 $Y2=1.96
r226 7 60 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.265
+ $Y=1.485 $X2=6.41 $Y2=1.96
r227 6 56 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.325
+ $Y=1.485 $X2=5.47 $Y2=1.96
r228 5 52 150 $w=1.7e-07 $l=8.39553e-07 $layer=licon1_PDIFF $count=4 $X=3.895
+ $Y=1.485 $X2=4.53 $Y2=1.96
r229 4 48 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=1.96
r230 3 42 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.96
r231 2 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.96
r232 1 30 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%Y 1 2 3 4 5 6 19 25 27 29 33 35 37 41 48
+ 51 53 54
r89 54 57 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.64 $Y=1.54 $X2=6.64
+ $Y2=1.455
r90 54 57 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=6.64 $Y=1.45 $X2=6.64
+ $Y2=1.455
r91 49 54 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=6.64 $Y=0.905
+ $X2=6.64 $Y2=1.45
r92 42 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.525 $Y=1.54
+ $X2=7.4 $Y2=1.54
r93 41 53 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.215 $Y=1.54
+ $X2=8.34 $Y2=1.54
r94 41 42 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.215 $Y=1.54
+ $X2=7.525 $Y2=1.54
r95 38 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.805 $Y=1.54
+ $X2=6.64 $Y2=1.54
r96 37 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.275 $Y=1.54
+ $X2=7.4 $Y2=1.54
r97 37 38 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=7.275 $Y=1.54
+ $X2=6.805 $Y2=1.54
r98 36 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.065 $Y=1.54
+ $X2=5.94 $Y2=1.54
r99 35 54 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.475 $Y=1.54
+ $X2=6.64 $Y2=1.54
r100 35 36 26.7487 $w=1.68e-07 $l=4.1e-07 $layer=LI1_cond $X=6.475 $Y=1.54
+ $X2=6.065 $Y2=1.54
r101 31 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.94 $Y=1.625
+ $X2=5.94 $Y2=1.54
r102 31 33 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.94 $Y=1.625
+ $X2=5.94 $Y2=2.3
r103 30 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.125 $Y=1.54 $X2=5
+ $Y2=1.54
r104 29 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.815 $Y=1.54
+ $X2=5.94 $Y2=1.54
r105 29 30 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.815 $Y=1.54
+ $X2=5.125 $Y2=1.54
r106 25 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5 $Y=1.625 $X2=5
+ $Y2=1.54
r107 25 27 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5 $Y=1.625 $X2=5
+ $Y2=2.3
r108 21 24 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=5.03 $Y=0.775
+ $X2=5.97 $Y2=0.775
r109 19 49 6.94204 $w=2.6e-07 $l=2.20624e-07 $layer=LI1_cond $X=6.475 $Y=0.775
+ $X2=6.64 $Y2=0.905
r110 19 24 22.384 $w=2.58e-07 $l=5.05e-07 $layer=LI1_cond $X=6.475 $Y=0.775
+ $X2=5.97 $Y2=0.775
r111 6 53 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.195
+ $Y=1.485 $X2=8.34 $Y2=1.62
r112 5 51 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.255
+ $Y=1.485 $X2=7.4 $Y2=1.62
r113 4 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.795
+ $Y=1.485 $X2=5.94 $Y2=1.62
r114 4 33 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.795
+ $Y=1.485 $X2=5.94 $Y2=2.3
r115 3 46 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.485 $X2=5 $Y2=1.62
r116 3 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.855
+ $Y=1.485 $X2=5 $Y2=2.3
r117 2 24 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=5.785
+ $Y=0.235 $X2=5.97 $Y2=0.73
r118 1 21 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.845
+ $Y=0.235 $X2=5.03 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_1361_297# 1 2 3 4 5 18 20 21 24 26 28
+ 29 30 34 36 38 40 42 48
r64 38 50 2.69138 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=10.72 $Y=1.625
+ $X2=10.72 $Y2=1.54
r65 38 40 25.0935 $w=3.08e-07 $l=6.75e-07 $layer=LI1_cond $X=10.72 $Y=1.625
+ $X2=10.72 $Y2=2.3
r66 37 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.875 $Y=1.54
+ $X2=9.75 $Y2=1.54
r67 36 50 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=10.565 $Y=1.54
+ $X2=10.72 $Y2=1.54
r68 36 37 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=10.565 $Y=1.54
+ $X2=9.875 $Y2=1.54
r69 32 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.75 $Y=1.625
+ $X2=9.75 $Y2=1.54
r70 32 34 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=9.75 $Y=1.625
+ $X2=9.75 $Y2=2.3
r71 31 44 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.935 $Y=1.54
+ $X2=8.81 $Y2=1.54
r72 30 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.625 $Y=1.54
+ $X2=9.75 $Y2=1.54
r73 30 31 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.625 $Y=1.54
+ $X2=8.935 $Y2=1.54
r74 29 46 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=2.295
+ $X2=8.81 $Y2=2.38
r75 28 44 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.81 $Y=1.625
+ $X2=8.81 $Y2=1.54
r76 28 29 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=8.81 $Y=1.625
+ $X2=8.81 $Y2=2.295
r77 27 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.995 $Y=2.38
+ $X2=7.87 $Y2=2.38
r78 26 46 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=8.81 $Y2=2.38
r79 26 27 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=7.995 $Y2=2.38
r80 22 42 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.87 $Y=2.295
+ $X2=7.87 $Y2=2.38
r81 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.87 $Y=2.295
+ $X2=7.87 $Y2=1.96
r82 20 42 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.745 $Y=2.38
+ $X2=7.87 $Y2=2.38
r83 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.745 $Y=2.38
+ $X2=7.055 $Y2=2.38
r84 16 21 7.36005 $w=1.7e-07 $l=1.77482e-07 $layer=LI1_cond $X=6.915 $Y=2.295
+ $X2=7.055 $Y2=2.38
r85 16 18 13.7882 $w=2.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.915 $Y=2.295
+ $X2=6.915 $Y2=1.96
r86 5 50 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=10.545
+ $Y=1.485 $X2=10.69 $Y2=1.62
r87 5 40 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=10.545
+ $Y=1.485 $X2=10.69 $Y2=2.3
r88 4 48 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=9.605
+ $Y=1.485 $X2=9.75 $Y2=1.62
r89 4 34 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=9.605
+ $Y=1.485 $X2=9.75 $Y2=2.3
r90 3 46 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=8.665
+ $Y=1.485 $X2=8.81 $Y2=2.3
r91 3 44 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=8.665
+ $Y=1.485 $X2=8.81 $Y2=1.62
r92 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.725
+ $Y=1.485 $X2=7.87 $Y2=1.96
r93 1 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=6.805
+ $Y=1.485 $X2=6.93 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_27_47# 1 2 3 4 5 16 22 23 24 28 30 34
+ 40
c77 23 0 1.98558e-19 $X=2.2 $Y=0.725
r78 32 34 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.015 $Y=0.725
+ $X2=4.015 $Y2=0.39
r79 31 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.265 $Y=0.815
+ $X2=3.075 $Y2=0.815
r80 30 32 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=3.825 $Y=0.815
+ $X2=4.015 $Y2=0.725
r81 30 31 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.825 $Y=0.815
+ $X2=3.265 $Y2=0.815
r82 26 40 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.075 $Y=0.725
+ $X2=3.075 $Y2=0.815
r83 26 28 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.075 $Y=0.725
+ $X2=3.075 $Y2=0.39
r84 25 39 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.325 $Y=0.815
+ $X2=2.2 $Y2=0.815
r85 24 40 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=0.815
+ $X2=3.075 $Y2=0.815
r86 24 25 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=2.885 $Y=0.815
+ $X2=2.325 $Y2=0.815
r87 23 39 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.2 $Y=0.725 $X2=2.2
+ $Y2=0.815
r88 22 37 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=2.2 $Y=0.475 $X2=2.2
+ $Y2=0.365
r89 22 23 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=2.2 $Y=0.475 $X2=2.2
+ $Y2=0.725
r90 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=0.28 $Y=0.365
+ $X2=1.22 $Y2=0.365
r91 16 37 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=2.075 $Y=0.365
+ $X2=2.2 $Y2=0.365
r92 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=2.075 $Y=0.365
+ $X2=1.22 $Y2=0.365
r93 5 34 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.39
r94 4 28 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.39
r95 3 39 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.73
r96 3 37 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r97 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.39
r98 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 56 57 59 60 61 89 90 95
r151 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r152 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r153 86 87 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r154 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r155 83 84 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r156 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r157 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r158 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=8.05
+ $Y2=0
r159 77 78 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r160 75 78 0.916224 $w=4.8e-07 $l=3.22e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=7.13 $Y2=0
r161 74 77 210.075 $w=1.68e-07 $l=3.22e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=7.13
+ $Y2=0
r162 74 75 2.325 $w=1.7e-07 $l=6.8e-07 $layer=mcon $count=4 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r163 72 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r164 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r165 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r166 69 95 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=0.23
+ $Y2=0
r167 68 69 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r168 64 68 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r169 64 95 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r170 61 95 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r171 59 86 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=9.89 $Y2=0
r172 59 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.135 $Y=0
+ $X2=10.22 $Y2=0
r173 58 89 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=10.305 $Y=0
+ $X2=10.81 $Y2=0
r174 58 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.305 $Y=0
+ $X2=10.22 $Y2=0
r175 56 83 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=9.195 $Y=0
+ $X2=8.97 $Y2=0
r176 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.195 $Y=0 $X2=9.28
+ $Y2=0
r177 55 86 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.365 $Y=0
+ $X2=9.89 $Y2=0
r178 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.365 $Y=0 $X2=9.28
+ $Y2=0
r179 53 80 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.255 $Y=0
+ $X2=8.05 $Y2=0
r180 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.255 $Y=0 $X2=8.34
+ $Y2=0
r181 52 83 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=8.425 $Y=0
+ $X2=8.97 $Y2=0
r182 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=0 $X2=8.34
+ $Y2=0
r183 50 77 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.13 $Y2=0
r184 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.315 $Y=0 $X2=7.4
+ $Y2=0
r185 49 80 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=7.485 $Y=0 $X2=8.05
+ $Y2=0
r186 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.485 $Y=0 $X2=7.4
+ $Y2=0
r187 47 71 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.45
+ $Y2=0
r188 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.57
+ $Y2=0
r189 46 74 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.655 $Y=0
+ $X2=3.91 $Y2=0
r190 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.57
+ $Y2=0
r191 44 68 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r192 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.63
+ $Y2=0
r193 43 71 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=3.45 $Y2=0
r194 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.63
+ $Y2=0
r195 39 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=0.085
+ $X2=10.22 $Y2=0
r196 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.22 $Y=0.085
+ $X2=10.22 $Y2=0.39
r197 35 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0
r198 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.28 $Y=0.085
+ $X2=9.28 $Y2=0.39
r199 31 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0
r200 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.34 $Y=0.085
+ $X2=8.34 $Y2=0.39
r201 27 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.4 $Y=0.085 $X2=7.4
+ $Y2=0
r202 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.4 $Y=0.085
+ $X2=7.4 $Y2=0.39
r203 23 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r204 23 25 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.39
r205 19 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r206 19 21 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.39
r207 6 41 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=10.035
+ $Y=0.235 $X2=10.22 $Y2=0.39
r208 5 37 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=9.095
+ $Y=0.235 $X2=9.28 $Y2=0.39
r209 4 33 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.155
+ $Y=0.235 $X2=8.34 $Y2=0.39
r210 3 29 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.215
+ $Y=0.235 $X2=7.4 $Y2=0.39
r211 2 25 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.39
r212 1 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_4%A_887_47# 1 2 3 4 5 6 7 24 26 27 33 34
+ 35 38 40 44 46 50 52 56 58 59 60
c122 58 0 2.97897e-20 $X=7.845 $Y=0.815
r123 54 56 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.665 $Y=0.725
+ $X2=10.665 $Y2=0.39
r124 53 60 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=9.915 $Y=0.815
+ $X2=9.725 $Y2=0.815
r125 52 54 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=10.475 $Y=0.815
+ $X2=10.665 $Y2=0.725
r126 52 53 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=10.475 $Y=0.815
+ $X2=9.915 $Y2=0.815
r127 48 60 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=9.725 $Y=0.725
+ $X2=9.725 $Y2=0.815
r128 48 50 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.725 $Y=0.725
+ $X2=9.725 $Y2=0.39
r129 47 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.975 $Y=0.815
+ $X2=8.785 $Y2=0.815
r130 46 60 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=9.535 $Y=0.815
+ $X2=9.725 $Y2=0.815
r131 46 47 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=9.535 $Y=0.815
+ $X2=8.975 $Y2=0.815
r132 42 59 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=8.785 $Y=0.725
+ $X2=8.785 $Y2=0.815
r133 42 44 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.785 $Y=0.725
+ $X2=8.785 $Y2=0.39
r134 41 58 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=8.035 $Y=0.815
+ $X2=7.845 $Y2=0.815
r135 40 59 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.595 $Y=0.815
+ $X2=8.785 $Y2=0.815
r136 40 41 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.595 $Y=0.815
+ $X2=8.035 $Y2=0.815
r137 36 58 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.845 $Y=0.725
+ $X2=7.845 $Y2=0.815
r138 36 38 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.845 $Y=0.725
+ $X2=7.845 $Y2=0.39
r139 34 58 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=7.655 $Y=0.82
+ $X2=7.845 $Y2=0.815
r140 34 35 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=7.655 $Y=0.82
+ $X2=7.145 $Y2=0.82
r141 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.06 $Y=0.735
+ $X2=7.145 $Y2=0.82
r142 32 33 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.06 $Y=0.475
+ $X2=7.06 $Y2=0.735
r143 29 31 74.9088 $w=2.18e-07 $l=1.43e-06 $layer=LI1_cond $X=5.5 $Y=0.365
+ $X2=6.93 $Y2=0.365
r144 27 29 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=4.645 $Y=0.365
+ $X2=5.5 $Y2=0.365
r145 26 32 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.975 $Y=0.365
+ $X2=7.06 $Y2=0.475
r146 26 31 2.35727 $w=2.18e-07 $l=4.5e-08 $layer=LI1_cond $X=6.975 $Y=0.365
+ $X2=6.93 $Y2=0.365
r147 22 27 6.88292 $w=2.2e-07 $l=1.49432e-07 $layer=LI1_cond $X=4.552 $Y=0.475
+ $X2=4.645 $Y2=0.365
r148 22 24 6.29484 $w=1.83e-07 $l=1.05e-07 $layer=LI1_cond $X=4.552 $Y=0.475
+ $X2=4.552 $Y2=0.58
r149 7 56 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=10.555
+ $Y=0.235 $X2=10.69 $Y2=0.39
r150 6 50 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=9.565
+ $Y=0.235 $X2=9.75 $Y2=0.39
r151 5 44 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=8.675
+ $Y=0.235 $X2=8.81 $Y2=0.39
r152 4 38 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.685
+ $Y=0.235 $X2=7.87 $Y2=0.39
r153 3 31 91 $w=1.7e-07 $l=6.98212e-07 $layer=licon1_NDIFF $count=2 $X=6.305
+ $Y=0.235 $X2=6.93 $Y2=0.39
r154 2 29 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.315
+ $Y=0.235 $X2=5.5 $Y2=0.39
r155 1 24 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.235 $X2=4.56 $Y2=0.58
.ends

