* NGSPICE file created from sky130_fd_sc_hdll__mux2_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__mux2_1 A0 A1 S VGND VNB VPB VPWR X
M1000 a_245_47# S VGND VNB nshort w=420000u l=150000u
+  ad=1.512e+11p pd=1.56e+06u as=4.745e+11p ps=4.06e+06u
M1001 VGND a_657_21# a_499_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=3.318e+11p ps=2.42e+06u
M1002 a_79_21# A0 a_243_374# VPB phighvt w=420000u l=180000u
+  ad=4.515e+11p pd=2.99e+06u as=1.743e+11p ps=1.67e+06u
M1003 a_613_374# A1 a_79_21# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=0p ps=0u
M1004 a_79_21# A1 a_245_47# VNB nshort w=420000u l=150000u
+  ad=2.562e+11p pd=2.06e+06u as=0p ps=0u
M1005 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=4.926e+11p pd=4.44e+06u as=2.7e+11p ps=2.54e+06u
M1006 VPWR a_657_21# a_613_374# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_499_47# A0 a_79_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_657_21# S VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1009 a_243_374# S VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1011 a_657_21# S VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
.ends

