* File: sky130_fd_sc_hdll__clkbuf_2.spice
* Created: Thu Aug 27 19:01:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_2.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.1323 PD=0.745 PS=1.47 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1000_d N_A_27_47#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06825 AS=0.0777 PD=0.745 PS=0.79 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_A_27_47#_M1003_g N_X_M1001_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.0777 PD=1.36 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1725 AS=0.275 PD=1.345 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1002_d N_A_27_47#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1725 AS=0.145 PD=1.345 PS=1.29 NRD=10.8153 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_27_47#_M1005_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_8 X X PROBETYPE=1
pX8_noxref noxref_9 X X PROBETYPE=1
pX9_noxref noxref_10 X X PROBETYPE=1
pX10_noxref noxref_11 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__clkbuf_2.pxi.spice"
*
.ends
*
*
