# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkinv_12
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  9.200000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  3.996000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 7.925000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  3.290400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 8.655000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 8.655000 1.630000 ;
        RECT 0.595000 1.630000 0.865000 2.465000 ;
        RECT 1.535000 1.630000 1.805000 2.465000 ;
        RECT 2.005000 0.255000 2.275000 0.695000 ;
        RECT 2.475000 1.630000 2.745000 2.465000 ;
        RECT 2.945000 0.255000 3.215000 0.695000 ;
        RECT 3.415000 1.630000 3.685000 2.465000 ;
        RECT 3.885000 0.255000 4.155000 0.695000 ;
        RECT 4.355000 1.630000 4.625000 2.465000 ;
        RECT 4.825000 0.255000 5.095000 0.695000 ;
        RECT 5.295000 1.630000 5.565000 2.465000 ;
        RECT 5.765000 0.255000 6.035000 0.695000 ;
        RECT 6.235000 1.630000 6.505000 2.465000 ;
        RECT 6.705000 0.255000 6.975000 0.695000 ;
        RECT 7.175000 1.630000 7.445000 2.465000 ;
        RECT 8.100000 0.865000 8.655000 1.460000 ;
        RECT 8.115000 1.630000 8.385000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.095000  1.800000 0.425000 2.635000 ;
      RECT 1.035000  1.800000 1.365000 2.635000 ;
      RECT 1.165000  0.085000 1.835000 0.525000 ;
      RECT 1.975000  1.800000 2.305000 2.635000 ;
      RECT 2.445000  0.085000 2.775000 0.525000 ;
      RECT 2.915000  1.800000 3.245000 2.635000 ;
      RECT 3.385000  0.085000 3.715000 0.525000 ;
      RECT 3.855000  1.800000 4.185000 2.635000 ;
      RECT 4.325000  0.085000 4.655000 0.525000 ;
      RECT 4.795000  1.800000 5.125000 2.635000 ;
      RECT 5.265000  0.085000 5.595000 0.525000 ;
      RECT 5.735000  1.800000 6.065000 2.635000 ;
      RECT 6.205000  0.085000 6.535000 0.525000 ;
      RECT 6.675000  1.800000 7.005000 2.635000 ;
      RECT 7.145000  0.085000 7.815000 0.525000 ;
      RECT 7.615000  1.800000 7.945000 2.635000 ;
      RECT 8.555000  1.800000 8.885000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkinv_12
