* File: sky130_fd_sc_hdll__dlxtn_2.pex.spice
* Created: Wed Sep  2 08:30:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%GATE_N 4 5 7 8 10 13 19 20 24 26
c41 19 0 2.67999e-20 $X=0.23 $Y=1.19
c42 13 0 2.71124e-20 $X=0.52 $Y=0.805
r43 24 27 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.4
r44 24 26 48.2986 $w=2.75e-07 $l=1.65e-07 $layer=POLY_cond $X=0.242 $Y=1.235
+ $X2=0.242 $Y2=1.07
r45 19 20 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.207 $Y=1.19
+ $X2=0.207 $Y2=1.53
r46 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r47 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r48 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r49 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r50 5 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r51 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r52 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r53 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r54 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r55 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%A_27_47# 1 2 8 9 11 14 18 19 21 24 28 29
+ 30 38 39 42 45 47 52 54 56 57 60 63 64 69 72 78
c166 19 0 4.94193e-20 $X=3.605 $Y=1.99
c167 8 0 2.67999e-20 $X=0.965 $Y=1.64
r168 68 69 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r169 64 78 6.77715 $w=3.38e-07 $l=1.15e-07 $layer=LI1_cond $X=3.34 $Y=1.53
+ $X2=3.34 $Y2=1.415
r170 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.26 $Y=1.53
+ $X2=3.26 $Y2=1.53
r171 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.745 $Y=1.53
+ $X2=0.745 $Y2=1.53
r172 57 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.89 $Y=1.53
+ $X2=0.745 $Y2=1.53
r173 56 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.115 $Y=1.53
+ $X2=3.26 $Y2=1.53
r174 56 57 2.75371 $w=1.4e-07 $l=2.225e-06 $layer=MET1_cond $X=3.115 $Y=1.53
+ $X2=0.89 $Y2=1.53
r175 52 72 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.025 $Y=0.87
+ $X2=3.025 $Y2=0.705
r176 51 54 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=3 $Y=0.87
+ $X2=3.255 $Y2=0.87
r177 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=0.87
+ $X2=3 $Y2=0.87
r178 49 60 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.745 $Y=1.795
+ $X2=0.745 $Y2=1.53
r179 48 60 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.745 $Y=1.4
+ $X2=0.745 $Y2=1.53
r180 46 68 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r181 45 48 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=1.235
+ $X2=0.775 $Y2=1.4
r182 45 47 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=1.235
+ $X2=0.775 $Y2=1.07
r183 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r184 39 75 27.028 $w=3.21e-07 $l=1.8e-07 $layer=POLY_cond $X=3.425 $Y=1.797
+ $X2=3.605 $Y2=1.797
r185 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r186 36 64 1.86425 $w=3.38e-07 $l=5.5e-08 $layer=LI1_cond $X=3.34 $Y=1.585
+ $X2=3.34 $Y2=1.53
r187 36 38 5.25378 $w=3.38e-07 $l=1.55e-07 $layer=LI1_cond $X=3.34 $Y=1.585
+ $X2=3.34 $Y2=1.74
r188 34 54 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=0.87
r189 34 78 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=3.255 $Y=1.035
+ $X2=3.255 $Y2=1.415
r190 32 47 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.745 $Y=0.805
+ $X2=0.745 $Y2=1.07
r191 31 42 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r192 30 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.745 $Y2=1.795
r193 30 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r194 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.745 $Y2=0.805
r195 28 29 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r196 22 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r197 22 24 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r198 19 75 16.2883 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.605 $Y=1.99
+ $X2=3.605 $Y2=1.797
r199 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.605 $Y=1.99
+ $X2=3.605 $Y2=2.275
r200 18 72 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.99 $Y=0.415
+ $X2=2.99 $Y2=0.705
r201 12 69 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r202 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r203 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r204 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r205 7 68 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r206 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r207 2 42 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r208 1 24 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%D 2 3 5 8 10 14 17
c43 14 0 1.07893e-19 $X=1.725 $Y=1.04
r44 16 17 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.04
+ $X2=1.98 $Y2=1.04
r45 13 16 40.2181 $w=3.3e-07 $l=2.3e-07 $layer=POLY_cond $X=1.725 $Y=1.04
+ $X2=1.955 $Y2=1.04
r46 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.04 $X2=1.725 $Y2=1.04
r47 10 14 4.06745 $w=4.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.677 $Y=1.19
+ $X2=1.677 $Y2=1.04
r48 6 17 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=0.875
+ $X2=1.98 $Y2=1.04
r49 6 8 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=1.98 $Y=0.875 $X2=1.98
+ $Y2=0.445
r50 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r52 1 16 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.04
r53 1 2 154.183 $w=2e-07 $l=4.65e-07 $layer=POLY_cond $X=1.955 $Y=1.205
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%A_319_47# 1 2 8 9 11 14 17 19 21 22 23 24
+ 26 33 35
c89 33 0 1.07893e-19 $X=2.405 $Y=0.93
c90 19 0 7.13094e-20 $X=2.12 $Y=0.7
r91 33 36 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.93
+ $X2=2.43 $Y2=1.095
r92 33 35 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=2.43 $Y=0.93
+ $X2=2.43 $Y2=0.765
r93 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=0.93 $X2=2.405 $Y2=0.93
r94 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.72 $Y=0.51
+ $X2=1.72 $Y2=0.7
r95 23 32 8.96999 $w=3.41e-07 $l=2.18746e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.33 $Y2=0.93
r96 23 24 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.205 $Y=1.095
+ $X2=2.205 $Y2=1.495
r97 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=2.205 $Y2=1.495
r98 21 22 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=2.12 $Y=1.58
+ $X2=1.885 $Y2=1.58
r99 20 28 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.805 $Y=0.7
+ $X2=1.72 $Y2=0.7
r100 19 32 8.22874 $w=3.41e-07 $l=3.18119e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=2.33 $Y2=0.93
r101 19 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.12 $Y=0.7
+ $X2=1.805 $Y2=0.7
r102 15 22 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.885 $Y2=1.58
r103 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r104 14 35 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.45 $Y=0.445
+ $X2=2.45 $Y2=0.765
r105 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r106 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r107 8 36 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r108 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r109 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%A_211_363# 1 2 7 8 9 11 12 16 20 22 24 25
+ 28 31 37
c111 37 0 4.94193e-20 $X=2.87 $Y=1.52
c112 8 0 1.86795e-19 $X=2.95 $Y=1.89
r113 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.52 $X2=2.87 $Y2=1.52
r114 34 36 33.8246 $w=2.85e-07 $l=2e-07 $layer=POLY_cond $X=2.892 $Y=1.32
+ $X2=2.892 $Y2=1.52
r115 32 37 14.1528 $w=2.83e-07 $l=3.5e-07 $layer=LI1_cond $X=2.812 $Y=1.87
+ $X2=2.812 $Y2=1.52
r116 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.755 $Y=1.87
+ $X2=2.755 $Y2=1.87
r117 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.255 $Y=1.87
+ $X2=1.255 $Y2=1.87
r118 25 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.4 $Y=1.87
+ $X2=1.255 $Y2=1.87
r119 24 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.61 $Y=1.87
+ $X2=2.755 $Y2=1.87
r120 24 25 1.49752 $w=1.4e-07 $l=1.21e-06 $layer=MET1_cond $X=2.61 $Y=1.87
+ $X2=1.4 $Y2=1.87
r121 22 28 3.73904 $w=2.23e-07 $l=7.3e-08 $layer=LI1_cond $X=1.227 $Y=1.797
+ $X2=1.227 $Y2=1.87
r122 22 23 6.45221 $w=2.23e-07 $l=1.12e-07 $layer=LI1_cond $X=1.227 $Y=1.797
+ $X2=1.227 $Y2=1.685
r123 20 23 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=1.2 $Y=0.51
+ $X2=1.2 $Y2=1.685
r124 14 16 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.515 $Y=1.245
+ $X2=3.515 $Y2=0.415
r125 13 34 17.7656 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=3.05 $Y=1.32
+ $X2=2.892 $Y2=1.32
r126 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.44 $Y=1.32
+ $X2=3.515 $Y2=1.245
r127 12 13 199.979 $w=1.5e-07 $l=3.9e-07 $layer=POLY_cond $X=3.44 $Y=1.32
+ $X2=3.05 $Y2=1.32
r128 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99
+ $X2=2.95 $Y2=2.275
r129 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r130 7 36 32.2493 $w=2.85e-07 $l=1.9182e-07 $layer=POLY_cond $X=2.95 $Y=1.685
+ $X2=2.892 $Y2=1.52
r131 7 8 67.9733 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=2.95 $Y=1.685 $X2=2.95
+ $Y2=1.89
r132 2 28 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r133 1 20 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%A_783_21# 1 2 9 11 13 14 16 17 19 20 22 23
+ 25 26 33 37 40 42 45 48 50 51 56
r92 56 57 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=5.945 $Y=1.202
+ $X2=5.97 $Y2=1.202
r93 55 56 57.0452 $w=3.76e-07 $l=4.45e-07 $layer=POLY_cond $X=5.5 $Y=1.202
+ $X2=5.945 $Y2=1.202
r94 54 55 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.202
+ $X2=5.5 $Y2=1.202
r95 46 54 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=5.45 $Y=1.202
+ $X2=5.475 $Y2=1.202
r96 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=1.16 $X2=5.45 $Y2=1.16
r97 43 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.905 $Y=1.16
+ $X2=4.82 $Y2=1.16
r98 43 45 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.905 $Y=1.16
+ $X2=5.45 $Y2=1.16
r99 42 50 7.80489 $w=1.95e-07 $l=1.77059e-07 $layer=LI1_cond $X=4.82 $Y=1.535
+ $X2=4.795 $Y2=1.7
r100 41 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=1.325
+ $X2=4.82 $Y2=1.16
r101 41 42 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.82 $Y=1.325
+ $X2=4.82 $Y2=1.535
r102 40 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=1.16
r103 40 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.82 $Y=0.995
+ $X2=4.82 $Y2=0.825
r104 35 50 7.80489 $w=1.95e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=1.865
+ $X2=4.795 $Y2=1.7
r105 35 37 21.2154 $w=2.18e-07 $l=4.05e-07 $layer=LI1_cond $X=4.795 $Y=1.865
+ $X2=4.795 $Y2=2.27
r106 31 48 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=4.795 $Y=0.715
+ $X2=4.795 $Y2=0.825
r107 31 33 7.07181 $w=2.18e-07 $l=1.35e-07 $layer=LI1_cond $X=4.795 $Y=0.715
+ $X2=4.795 $Y2=0.58
r108 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.27
+ $Y=1.7 $X2=4.27 $Y2=1.7
r109 26 50 0.463323 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.685 $Y=1.7
+ $X2=4.795 $Y2=1.7
r110 26 28 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=4.685 $Y=1.7
+ $X2=4.27 $Y2=1.7
r111 23 57 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=1.202
r112 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.97 $Y=0.995
+ $X2=5.97 $Y2=0.56
r113 20 56 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.202
r114 20 22 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.985
r115 17 55 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.5 $Y=0.995
+ $X2=5.5 $Y2=1.202
r116 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.5 $Y=0.995
+ $X2=5.5 $Y2=0.56
r117 14 54 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.202
r118 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.475 $Y=1.41
+ $X2=5.475 $Y2=1.985
r119 11 29 49.5109 $w=4.1e-07 $l=3.55176e-07 $layer=POLY_cond $X=4.015 $Y=1.99
+ $X2=4.16 $Y2=1.7
r120 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.015 $Y=1.99
+ $X2=4.015 $Y2=2.275
r121 7 29 39.7867 $w=4.1e-07 $l=2.38642e-07 $layer=POLY_cond $X=3.99 $Y=1.535
+ $X2=4.16 $Y2=1.7
r122 7 9 558.915 $w=1.5e-07 $l=1.09e-06 $layer=POLY_cond $X=3.99 $Y=1.535
+ $X2=3.99 $Y2=0.445
r123 2 50 600 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.485 $X2=4.77 $Y2=1.755
r124 2 37 600 $w=1.7e-07 $l=8.45192e-07 $layer=licon1_PDIFF $count=1 $X=4.645
+ $Y=1.485 $X2=4.77 $Y2=2.27
r125 1 33 182 $w=1.7e-07 $l=4.02679e-07 $layer=licon1_NDIFF $count=1 $X=4.645
+ $Y=0.235 $X2=4.77 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%A_608_413# 1 2 7 9 10 12 13 14 15 19 24 25
+ 26 29
c80 25 0 1.7336e-19 $X=3.86 $Y=1.325
c81 14 0 1.25081e-19 $X=5.005 $Y=1.202
r82 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.46
+ $Y=1.16 $X2=4.46 $Y2=1.16
r83 27 29 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=3.945 $Y=1.16
+ $X2=4.46 $Y2=1.16
r84 25 27 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.86 $Y=1.325
+ $X2=3.785 $Y2=1.16
r85 25 26 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.86 $Y=1.325
+ $X2=3.86 $Y2=2.255
r86 24 27 9.34553 $w=2.47e-07 $l=1.98997e-07 $layer=LI1_cond $X=3.71 $Y=0.995
+ $X2=3.785 $Y2=1.16
r87 23 24 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.71 $Y=0.535
+ $X2=3.71 $Y2=0.995
r88 19 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.775 $Y=2.34
+ $X2=3.86 $Y2=2.255
r89 19 21 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.775 $Y=2.34
+ $X2=3.31 $Y2=2.34
r90 15 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.625 $Y=0.45
+ $X2=3.71 $Y2=0.535
r91 15 17 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=3.625 $Y=0.45
+ $X2=3.25 $Y2=0.45
r92 13 30 77.8133 $w=3.3e-07 $l=4.45e-07 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=4.46 $Y2=1.16
r93 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.905 $Y=1.16
+ $X2=5.005 $Y2=1.202
r94 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.005 $Y2=1.202
r95 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.03 $Y=0.995
+ $X2=5.03 $Y2=0.56
r96 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.202
r97 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.005 $Y=1.41
+ $X2=5.005 $Y2=1.985
r98 2 21 600 $w=1.7e-07 $l=3.87137e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.31 $Y2=2.34
r99 1 17 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=3.065
+ $Y=0.235 $X2=3.25 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%VPWR 1 2 3 4 5 18 22 26 30 32 34 37 38 39
+ 41 53 60 65 71 74 77 81
c95 22 0 1.86795e-19 $X=2.19 $Y=2
r96 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r97 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r99 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r100 69 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r101 69 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r102 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r103 66 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.405 $Y=2.72
+ $X2=5.27 $Y2=2.72
r104 66 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=2.72
+ $X2=5.75 $Y2=2.72
r105 65 80 4.04153 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=6.267 $Y2=2.72
r106 65 68 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r107 64 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r108 64 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r109 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r110 61 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.315 $Y2=2.72
r111 61 63 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=4.465 $Y=2.72
+ $X2=4.83 $Y2=2.72
r112 60 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=5.27 $Y2=2.72
r113 60 63 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=2.72
+ $X2=4.83 $Y2=2.72
r114 59 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r116 56 59 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r117 55 58 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r118 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r119 53 74 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=4.315 $Y2=2.72
r120 53 58 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r121 52 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r123 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 49 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 48 51 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 48 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r127 46 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r128 46 48 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 41 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r130 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r131 39 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 39 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r133 37 51 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r134 37 38 8.33247 $w=1.7e-07 $l=1.57e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.262 $Y2=2.72
r135 36 55 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.53 $Y2=2.72
r136 36 38 8.33247 $w=1.7e-07 $l=1.58e-07 $layer=LI1_cond $X=2.42 $Y=2.72
+ $X2=2.262 $Y2=2.72
r137 32 80 3.10164 $w=2.5e-07 $l=1.05924e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.267 $Y2=2.72
r138 32 34 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2
r139 28 77 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=2.72
r140 28 30 38.4148 $w=2.68e-07 $l=9e-07 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=1.735
r141 24 74 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.315 $Y=2.635
+ $X2=4.315 $Y2=2.72
r142 24 26 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=4.315 $Y=2.635
+ $X2=4.315 $Y2=2.3
r143 20 38 0.751525 $w=3.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2.72
r144 20 22 23.2318 $w=3.13e-07 $l=6.35e-07 $layer=LI1_cond $X=2.262 $Y=2.635
+ $X2=2.262 $Y2=2
r145 16 71 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r146 16 18 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r147 5 34 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=2
r148 4 30 300 $w=1.7e-07 $l=3.14245e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=1.485 $X2=5.24 $Y2=1.735
r149 3 26 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=4.105
+ $Y=2.065 $X2=4.25 $Y2=2.3
r150 2 22 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r151 1 18 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%Q 1 2 8 11 12 13 14 15 16
c28 16 0 1.25081e-19 $X=6.21 $Y=1.19
r29 16 32 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=6.21 $Y=1.16
+ $X2=5.825 $Y2=1.16
r30 14 15 15.1637 $w=2.83e-07 $l=3.75e-07 $layer=LI1_cond $X=5.767 $Y=1.835
+ $X2=5.767 $Y2=2.21
r31 13 31 14.599 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=5.767 $Y=0.51
+ $X2=5.767 $Y2=0.825
r32 11 14 8.00645 $w=2.83e-07 $l=1.98e-07 $layer=LI1_cond $X=5.767 $Y=1.637
+ $X2=5.767 $Y2=1.835
r33 11 12 7.60349 $w=2.83e-07 $l=1.42e-07 $layer=LI1_cond $X=5.767 $Y=1.637
+ $X2=5.767 $Y2=1.495
r34 9 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.16
r35 9 12 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.495
r36 8 32 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.825 $Y=0.995
+ $X2=5.825 $Y2=1.16
r37 8 31 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=5.825 $Y=0.995
+ $X2=5.825 $Y2=0.825
r38 2 14 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.835
r39 1 13 182 $w=1.7e-07 $l=4.0694e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.58
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLXTN_2%VGND 1 2 3 4 5 18 22 24 26 29 30 31 33 38
+ 50 54 61 68 74 78
c95 78 0 2.71124e-20 $X=6.21 $Y=0
c96 2 0 7.13094e-20 $X=2.055 $Y=0.235
r97 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r98 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r99 68 71 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.165 $Y=0 $X2=2.165
+ $Y2=0.36
r100 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r101 61 64 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r102 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r103 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r104 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=5.29
+ $Y2=0
r105 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r106 55 74 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.405 $Y=0 $X2=5.27
+ $Y2=0
r107 55 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=5.405 $Y=0 $X2=5.75
+ $Y2=0
r108 54 77 4.14883 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=0
+ $X2=6.267 $Y2=0
r109 54 57 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.75
+ $Y2=0
r110 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r111 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r112 50 74 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.135 $Y=0 $X2=5.27
+ $Y2=0
r113 50 52 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.135 $Y=0
+ $X2=4.83 $Y2=0
r114 49 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r115 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r116 46 49 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r117 46 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r118 45 48 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r119 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r120 43 68 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.165
+ $Y2=0
r121 43 45 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r122 42 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r123 42 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r124 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r125 39 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r126 39 41 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.61 $Y2=0
r127 38 68 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.975 $Y=0 $X2=2.165
+ $Y2=0
r128 38 41 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=0
+ $X2=1.61 $Y2=0
r129 33 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r130 33 35 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r131 31 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r132 31 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r133 29 48 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=0
+ $X2=3.91 $Y2=0
r134 29 30 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.225
+ $Y2=0
r135 28 52 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=4.415 $Y=0
+ $X2=4.83 $Y2=0
r136 28 30 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.415 $Y=0 $X2=4.225
+ $Y2=0
r137 24 77 3.06338 $w=2.6e-07 $l=1.03899e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.267 $Y2=0
r138 24 26 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.225 $Y=0.085
+ $X2=6.225 $Y2=0.38
r139 20 74 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0
r140 20 22 19.8476 $w=2.68e-07 $l=4.65e-07 $layer=LI1_cond $X=5.27 $Y=0.085
+ $X2=5.27 $Y2=0.55
r141 16 30 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0
r142 16 18 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0.445
r143 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.38
r144 4 22 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=5.105
+ $Y=0.235 $X2=5.24 $Y2=0.55
r145 3 18 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=4.065
+ $Y=0.235 $X2=4.25 $Y2=0.445
r146 2 71 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r147 1 64 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

