* File: sky130_fd_sc_hdll__sdfsbp_1.pex.spice
* Created: Thu Aug 27 19:26:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%SCD 1 2 3 5 6 8 13 14
c35 13 0 1.17581e-19 $X=0.23 $Y=0.85
c36 6 0 3.51615e-20 $X=0.495 $Y=1.77
r37 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r38 14 19 15.2287 $w=2.78e-07 $l=3.7e-07 $layer=LI1_cond $X=0.225 $Y=1.53
+ $X2=0.225 $Y2=1.16
r39 13 19 12.7592 $w=2.78e-07 $l=3.1e-07 $layer=LI1_cond $X=0.225 $Y=0.85
+ $X2=0.225 $Y2=1.16
r40 6 9 89.734 $w=1.5e-07 $l=1.75e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.32 $Y2=1.695
r41 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r42 3 18 87.8413 $w=2.62e-07 $l=4.96377e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.327 $Y2=1.16
r43 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r44 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.32 $Y=1.62 $X2=0.32
+ $Y2=1.695
r45 1 18 39.0894 $w=2.62e-07 $l=1.68464e-07 $layer=POLY_cond $X=0.32 $Y=1.325
+ $X2=0.327 $Y2=1.16
r46 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.32 $Y=1.325
+ $X2=0.32 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%SCE 3 6 7 9 11 12 14 17 19 20 22 25 30 33
+ 34 38 48
c104 22 0 1.07953e-19 $X=2.73 $Y=1.19
c105 7 0 2.34944e-19 $X=0.965 $Y=1.77
r106 38 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.715 $Y=1.19
+ $X2=0.715 $Y2=1.19
r107 33 36 37.7183 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.767 $Y=1.16
+ $X2=2.767 $Y2=1.325
r108 33 35 46.255 $w=3.35e-07 $l=1.65e-07 $layer=POLY_cond $X=2.767 $Y=1.16
+ $X2=2.767 $Y2=0.995
r109 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r110 30 31 7.25418 $w=2.99e-07 $l=4.5e-08 $layer=POLY_cond $X=0.92 $Y=1.245
+ $X2=0.965 $Y2=1.245
r111 28 30 23.3746 $w=2.99e-07 $l=1.45e-07 $layer=POLY_cond $X=0.775 $Y=1.245
+ $X2=0.92 $Y2=1.245
r112 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.775
+ $Y=1.245 $X2=0.775 $Y2=1.245
r113 25 48 0.00320802 $w=2.3e-07 $l=5e-09 $layer=MET1_cond $X=0.69 $Y=1.19
+ $X2=0.695 $Y2=1.19
r114 22 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.73 $Y=1.19
+ $X2=2.73 $Y2=1.19
r115 20 48 0.128299 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=0.86 $Y=1.19
+ $X2=0.695 $Y2=1.19
r116 19 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=2.73 $Y2=1.19
r117 19 20 2.1349 $w=1.4e-07 $l=1.725e-06 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=0.86 $Y2=1.19
r118 17 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.86 $Y=0.445
+ $X2=2.86 $Y2=0.995
r119 12 14 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.835 $Y=1.77
+ $X2=2.835 $Y2=2.165
r120 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.835 $Y=1.67 $X2=2.835
+ $Y2=1.77
r121 11 36 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=2.835 $Y=1.67
+ $X2=2.835 $Y2=1.325
r122 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.77
+ $X2=0.965 $Y2=2.165
r123 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.67 $X2=0.965
+ $Y2=1.77
r124 5 31 12.2124 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.245
r125 5 6 86.2101 $w=2e-07 $l=2.6e-07 $layer=POLY_cond $X=0.965 $Y=1.41 $X2=0.965
+ $Y2=1.67
r126 1 30 18.89 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.92 $Y=1.08 $X2=0.92
+ $Y2=1.245
r127 1 3 325.606 $w=1.5e-07 $l=6.35e-07 $layer=POLY_cond $X=0.92 $Y=1.08
+ $X2=0.92 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%D 2 3 5 8 9 10 14 16
c46 9 0 8.70679e-20 $X=1.14 $Y=0.85
r47 14 17 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=0.93
+ $X2=1.34 $Y2=1.095
r48 14 16 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.34 $Y=0.93
+ $X2=1.34 $Y2=0.765
r49 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.34
+ $Y=0.93 $X2=1.34 $Y2=0.93
r50 10 15 17.5055 $w=3.93e-07 $l=6e-07 $layer=LI1_cond $X=1.227 $Y=1.53
+ $X2=1.227 $Y2=0.93
r51 9 15 2.33406 $w=3.93e-07 $l=8e-08 $layer=LI1_cond $X=1.227 $Y=0.85 $X2=1.227
+ $Y2=0.93
r52 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.4 $Y=0.445 $X2=1.4
+ $Y2=0.765
r53 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.375 $Y=1.77
+ $X2=1.375 $Y2=2.165
r54 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.375 $Y=1.67 $X2=1.375
+ $Y2=1.77
r55 2 17 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=1.375 $Y=1.67
+ $X2=1.375 $Y2=1.095
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_349_21# 1 2 9 12 13 15 19 20 21 23 33
+ 35
c76 20 0 1.59069e-19 $X=2.15 $Y=1.16
r77 37 39 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.82 $Y=1.16
+ $X2=1.845 $Y2=1.16
r78 33 35 0.841466 $w=3.13e-07 $l=2.3e-08 $layer=LI1_cond $X=2.577 $Y=1.927
+ $X2=2.6 $Y2=1.927
r79 21 23 12.4283 $w=2.53e-07 $l=2.75e-07 $layer=LI1_cond $X=2.587 $Y=0.715
+ $X2=2.587 $Y2=0.44
r80 20 39 53.3327 $w=3.3e-07 $l=3.05e-07 $layer=POLY_cond $X=2.15 $Y=1.16
+ $X2=1.845 $Y2=1.16
r81 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r82 17 33 12.622 $w=3.13e-07 $l=3.45e-07 $layer=LI1_cond $X=2.232 $Y=1.927
+ $X2=2.577 $Y2=1.927
r83 17 19 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.232 $Y=1.77
+ $X2=2.232 $Y2=1.16
r84 16 21 20.7225 $w=1.88e-07 $l=3.55e-07 $layer=LI1_cond $X=2.232 $Y=0.81
+ $X2=2.587 $Y2=0.81
r85 16 19 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.232 $Y=0.905
+ $X2=2.232 $Y2=1.16
r86 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.845 $Y=1.77
+ $X2=1.845 $Y2=2.165
r87 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.845 $Y=1.67 $X2=1.845
+ $Y2=1.77
r88 11 39 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.16
r89 11 12 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.67
r90 7 37 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.82 $Y2=1.16
r91 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.445
r92 2 35 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.845 $X2=2.6 $Y2=1.99
r93 1 23 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.235 $X2=2.63 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%CLK 7 8 10 13 15 16 17 18 22 23 24 26
c72 23 0 3.24882e-20 $X=3.68 $Y=1.255
c73 16 0 9.66133e-20 $X=3.795 $Y=1.77
c74 13 0 1.11374e-19 $X=3.88 $Y=0.805
r75 23 26 15.6478 $w=4.6e-07 $l=7.3675e-07 $layer=LI1_cond $X=3.485 $Y=1.255
+ $X2=3.155 $Y2=1.845
r76 22 25 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.42
r77 22 24 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.09
r78 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.255 $X2=3.68 $Y2=1.255
r79 18 23 1.72391 $w=4.6e-07 $l=6.5e-08 $layer=LI1_cond $X=3.485 $Y=1.19
+ $X2=3.485 $Y2=1.255
r80 17 26 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=1.845
+ $X2=3.155 $Y2=1.845
r81 15 16 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.795 $Y=1.62
+ $X2=3.795 $Y2=1.77
r82 15 25 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.74 $Y=1.62 $X2=3.74
+ $Y2=1.42
r83 11 13 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.74 $Y=0.805
+ $X2=3.88 $Y2=0.805
r84 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.805
r85 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.445
r86 7 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=1.77
r87 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=0.805
r88 1 24 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_693_369# 1 2 8 9 11 12 14 17 19 21 22
+ 24 26 27 29 32 34 37 41 43 44 45 46 48 50 51 55 56 57 58 61 64 65 66 67 68 77
+ 81 85 91
c293 91 0 6.89134e-20 $X=9.81 $Y=1.08
c294 85 0 1.8066e-19 $X=5.73 $Y=1.74
c295 81 0 3.24882e-20 $X=4.235 $Y=1.09
c296 77 0 2.03002e-19 $X=8.29 $Y=1.87
c297 50 0 9.66133e-20 $X=4.21 $Y=1.255
c298 27 0 1.31062e-19 $X=8.585 $Y=1.57
r299 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.74 $X2=5.73 $Y2=1.74
r300 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.29 $Y=1.87
+ $X2=8.29 $Y2=1.87
r301 74 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.69 $Y=1.87
+ $X2=5.69 $Y2=1.87
r302 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.21 $Y=1.87
+ $X2=4.21 $Y2=1.87
r303 68 74 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.885 $Y=1.87
+ $X2=5.69 $Y2=1.87
r304 67 77 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.145 $Y=1.87
+ $X2=8.29 $Y2=1.87
r305 67 68 2.79702 $w=1.4e-07 $l=2.26e-06 $layer=MET1_cond $X=8.145 $Y=1.87
+ $X2=5.885 $Y2=1.87
r306 66 70 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=4.405 $Y=1.87
+ $X2=4.21 $Y2=1.87
r307 65 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=5.69 $Y2=1.87
r308 65 66 1.41089 $w=1.4e-07 $l=1.14e-06 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=4.405 $Y2=1.87
r309 64 78 6.37042 $w=4.58e-07 $l=2.45e-07 $layer=LI1_cond $X=8.535 $Y=1.725
+ $X2=8.29 $Y2=1.725
r310 62 91 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=9.7 $Y=1.08
+ $X2=9.81 $Y2=1.08
r311 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.7
+ $Y=1.08 $X2=9.7 $Y2=1.08
r312 59 61 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=9.75 $Y=0.895
+ $X2=9.75 $Y2=1.08
r313 57 59 7.06569 $w=2e-07 $l=1.83303e-07 $layer=LI1_cond $X=9.61 $Y=0.795
+ $X2=9.75 $Y2=0.895
r314 57 58 47.4136 $w=1.98e-07 $l=8.55e-07 $layer=LI1_cond $X=9.61 $Y=0.795
+ $X2=8.755 $Y2=0.795
r315 56 88 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.645 $Y=1.16
+ $X2=8.645 $Y2=1.325
r316 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.62
+ $Y=1.16 $X2=8.62 $Y2=1.16
r317 53 64 7.98384 $w=4.6e-07 $l=2.79643e-07 $layer=LI1_cond $X=8.645 $Y=1.495
+ $X2=8.535 $Y2=1.725
r318 53 55 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=8.645 $Y=1.495
+ $X2=8.645 $Y2=1.16
r319 52 58 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=8.645 $Y=0.895
+ $X2=8.755 $Y2=0.795
r320 52 55 13.8817 $w=2.18e-07 $l=2.65e-07 $layer=LI1_cond $X=8.645 $Y=0.895
+ $X2=8.645 $Y2=1.16
r321 51 82 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.42
r322 51 81 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.09
r323 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.255 $X2=4.21 $Y2=1.255
r324 48 71 2.91016 $w=2.6e-07 $l=9e-08 $layer=LI1_cond $X=4.165 $Y=1.775
+ $X2=4.165 $Y2=1.865
r325 48 50 23.0489 $w=2.58e-07 $l=5.2e-07 $layer=LI1_cond $X=4.165 $Y=1.775
+ $X2=4.165 $Y2=1.255
r326 47 50 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.165 $Y=0.885
+ $X2=4.165 $Y2=1.255
r327 45 47 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=4.165 $Y2=0.885
r328 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=3.705 $Y2=0.8
r329 43 71 4.20357 $w=1.8e-07 $l=1.3e-07 $layer=LI1_cond $X=4.035 $Y=1.865
+ $X2=4.165 $Y2=1.865
r330 43 44 22.1818 $w=1.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=1.865
+ $X2=3.675 $Y2=1.865
r331 39 46 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.705 $Y2=0.8
r332 39 41 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.612 $Y2=0.44
r333 35 44 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.59 $Y=1.955
+ $X2=3.675 $Y2=1.865
r334 35 37 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=3.59 $Y=1.955
+ $X2=3.59 $Y2=2.16
r335 30 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.81 $Y=0.915
+ $X2=9.81 $Y2=1.08
r336 30 32 241 $w=1.5e-07 $l=4.7e-07 $layer=POLY_cond $X=9.81 $Y=0.915 $X2=9.81
+ $Y2=0.445
r337 27 29 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.585 $Y=1.57
+ $X2=8.585 $Y2=2.065
r338 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.585 $Y=1.47 $X2=8.585
+ $Y2=1.57
r339 26 88 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.585 $Y=1.47
+ $X2=8.585 $Y2=1.325
r340 22 84 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=1.74
r341 22 24 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=2.275
r342 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.34 $Y=0.73
+ $X2=5.34 $Y2=0.445
r343 18 34 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.395 $Y=0.805
+ $X2=4.32 $Y2=0.805
r344 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=5.34 $Y2=0.73
r345 17 18 446.106 $w=1.5e-07 $l=8.7e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=4.395 $Y2=0.805
r346 15 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=0.88
+ $X2=4.32 $Y2=0.805
r347 15 81 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.32 $Y=0.88
+ $X2=4.32 $Y2=1.09
r348 12 34 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.32 $Y=0.73
+ $X2=4.32 $Y2=0.805
r349 12 14 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.32 $Y=0.73
+ $X2=4.32 $Y2=0.445
r350 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.295 $Y=1.77
+ $X2=4.295 $Y2=2.165
r351 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.295 $Y=1.67 $X2=4.295
+ $Y2=1.77
r352 8 82 82.8943 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.295 $Y=1.67
+ $X2=4.295 $Y2=1.42
r353 2 37 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.845 $X2=3.59 $Y2=2.16
r354 1 41 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.495
+ $Y=0.235 $X2=3.62 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_877_369# 1 2 8 9 11 12 13 15 18 22 24
+ 26 32 33 36 39 40 43 46 47 54 63
c183 63 0 8.42613e-20 $X=4.677 $Y=1.09
c184 47 0 9.89235e-21 $X=9.31 $Y=1.19
c185 43 0 1.3308e-19 $X=4.67 $Y=1.19
c186 18 0 8.99086e-20 $X=5.81 $Y=0.445
c187 11 0 2.89743e-19 $X=5.195 $Y=1.915
c188 9 0 1.70908e-19 $X=5.735 $Y=1.165
c189 8 0 1.8066e-19 $X=4.965 $Y=1.84
r190 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.305
+ $Y=1.74 $X2=9.305 $Y2=1.74
r191 53 54 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.255
+ $X2=5.04 $Y2=1.255
r192 50 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.755 $Y=1.255
+ $X2=4.965 $Y2=1.255
r193 47 57 22.6373 $w=2.78e-07 $l=5.5e-07 $layer=LI1_cond $X=9.255 $Y=1.19
+ $X2=9.255 $Y2=1.74
r194 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.31 $Y=1.19
+ $X2=9.31 $Y2=1.19
r195 43 64 8.46186 $w=3.23e-07 $l=2.3e-07 $layer=LI1_cond $X=4.677 $Y=1.19
+ $X2=4.677 $Y2=1.42
r196 43 63 6.15528 $w=3.23e-07 $l=1e-07 $layer=LI1_cond $X=4.677 $Y=1.19
+ $X2=4.677 $Y2=1.09
r197 43 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.255 $X2=4.755 $Y2=1.255
r198 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.67 $Y=1.19
+ $X2=4.67 $Y2=1.19
r199 40 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.815 $Y=1.19
+ $X2=4.67 $Y2=1.19
r200 39 46 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=9.115 $Y=1.19
+ $X2=9.31 $Y2=1.19
r201 39 40 5.32177 $w=1.4e-07 $l=4.3e-06 $layer=MET1_cond $X=9.115 $Y=1.19
+ $X2=4.815 $Y2=1.19
r202 38 63 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=4.6 $Y=0.585
+ $X2=4.6 $Y2=1.09
r203 36 38 9.16686 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=4.572 $Y=0.42
+ $X2=4.572 $Y2=0.585
r204 33 64 29.9635 $w=2.73e-07 $l=7.15e-07 $layer=LI1_cond $X=4.652 $Y=2.135
+ $X2=4.652 $Y2=1.42
r205 32 33 6.01906 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.617 $Y=2.3
+ $X2=4.617 $Y2=2.135
r206 24 56 46.294 $w=3.33e-07 $l=2.65989e-07 $layer=POLY_cond $X=9.26 $Y=1.99
+ $X2=9.227 $Y2=1.74
r207 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.26 $Y=1.99
+ $X2=9.26 $Y2=2.275
r208 20 56 38.6212 $w=3.33e-07 $l=2.23226e-07 $layer=POLY_cond $X=9.09 $Y=1.575
+ $X2=9.227 $Y2=1.74
r209 20 22 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.09 $Y=1.575
+ $X2=9.09 $Y2=0.555
r210 16 18 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.81 $Y=1.09
+ $X2=5.81 $Y2=0.445
r211 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.285 $Y=1.99
+ $X2=5.285 $Y2=2.275
r212 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.285 $Y2=1.99
r213 11 12 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.04 $Y2=1.915
r214 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.81 $Y2=1.09
r215 9 54 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.04 $Y2=1.165
r216 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.965 $Y=1.84
+ $X2=5.04 $Y2=1.915
r217 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.255
r218 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.84
r219 2 32 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.845 $X2=4.53 $Y2=2.3
r220 1 36 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.235 $X2=4.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_1219_21# 1 2 9 12 13 15 18 21 23 24 27
+ 31 33 42
c95 33 0 4.24205e-20 $X=6.267 $Y=0.72
r96 37 42 12.2196 $w=2.7e-07 $l=5.5e-08 $layer=POLY_cond $X=6.26 $Y=0.93
+ $X2=6.315 $Y2=0.93
r97 37 39 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=6.26 $Y=0.93 $X2=6.17
+ $Y2=0.93
r98 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.26
+ $Y=0.93 $X2=6.26 $Y2=0.93
r99 33 36 5.83164 $w=4.13e-07 $l=2.1e-07 $layer=LI1_cond $X=6.267 $Y=0.72
+ $X2=6.267 $Y2=0.93
r100 29 31 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.232 $Y=2.105
+ $X2=7.232 $Y2=2.285
r101 25 27 4.64695 $w=3.08e-07 $l=1.25e-07 $layer=LI1_cond $X=6.93 $Y=0.635
+ $X2=6.93 $Y2=0.51
r102 23 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.1 $Y=2.02
+ $X2=7.232 $Y2=2.105
r103 23 24 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=7.1 $Y=2.02
+ $X2=6.595 $Y2=2.02
r104 22 33 6.00275 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.475 $Y=0.72
+ $X2=6.267 $Y2=0.72
r105 21 25 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=6.775 $Y=0.72
+ $X2=6.93 $Y2=0.635
r106 21 22 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=6.775 $Y=0.72
+ $X2=6.475 $Y2=0.72
r107 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.51
+ $Y=1.74 $X2=6.51 $Y2=1.74
r108 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.595 $Y2=2.02
r109 16 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.51 $Y2=1.74
r110 13 19 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.43 $Y2=1.74
r111 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.315 $Y2=2.275
r112 12 19 31.7097 $w=3.82e-07 $l=2.14942e-07 $layer=POLY_cond $X=6.315 $Y=1.575
+ $X2=6.43 $Y2=1.74
r113 11 42 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=6.315 $Y=1.065
+ $X2=6.315 $Y2=0.93
r114 11 12 169.104 $w=2e-07 $l=5.1e-07 $layer=POLY_cond $X=6.315 $Y=1.065
+ $X2=6.315 $Y2=1.575
r115 7 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.17 $Y=0.795
+ $X2=6.17 $Y2=0.93
r116 7 9 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.17 $Y=0.795
+ $X2=6.17 $Y2=0.445
r117 2 31 600 $w=1.7e-07 $l=2.91033e-07 $layer=licon1_PDIFF $count=1 $X=7.045
+ $Y=2.065 $X2=7.21 $Y2=2.285
r118 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.825
+ $Y=0.235 $X2=6.95 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_1075_413# 1 2 8 10 11 13 14 16 18 19 21
+ 24 27 31 33 38 43 47 48 50 51 52 57 60
c159 10 0 4.24205e-20 $X=6.96 $Y=1.095
r160 56 57 1.11087 $w=2.7e-07 $l=5e-09 $layer=POLY_cond $X=6.955 $Y=1.23
+ $X2=6.96 $Y2=1.23
r161 51 61 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.16
+ $X2=8.115 $Y2=1.325
r162 51 60 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.115 $Y=1.16
+ $X2=8.115 $Y2=0.995
r163 50 52 4.87734 $w=3.48e-07 $l=1.4e-07 $layer=LI1_cond $X=8.09 $Y=1.15
+ $X2=7.95 $Y2=1.15
r164 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=1.16 $X2=8.09 $Y2=1.16
r165 48 52 38.991 $w=2.98e-07 $l=1.015e-06 $layer=LI1_cond $X=6.935 $Y=1.125
+ $X2=7.95 $Y2=1.125
r166 46 56 23.3282 $w=2.7e-07 $l=1.05e-07 $layer=POLY_cond $X=6.85 $Y=1.23
+ $X2=6.955 $Y2=1.23
r167 45 48 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.85 $Y=1.185
+ $X2=6.935 $Y2=1.185
r168 45 47 6.95306 $w=4.18e-07 $l=1e-07 $layer=LI1_cond $X=6.85 $Y=1.185
+ $X2=6.75 $Y2=1.185
r169 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.23 $X2=6.85 $Y2=1.23
r170 40 43 3.80956 $w=1.7e-07 $l=8.46434e-07 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=5.4 $Y2=1.225
r171 40 47 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=6.75 $Y2=1.31
r172 37 43 2.88756 $w=3.3e-07 $l=8.005e-07 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=5.4 $Y2=1.225
r173 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=6.12 $Y2=2.135
r174 33 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=6.12 $Y2=2.135
r175 33 35 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=5.52 $Y2=2.3
r176 29 43 2.88756 $w=3.3e-07 $l=2.45e-07 $layer=LI1_cond $X=5.645 $Y=1.225
+ $X2=5.4 $Y2=1.225
r177 29 31 19.6499 $w=4.88e-07 $l=8.05e-07 $layer=LI1_cond $X=5.645 $Y=1.225
+ $X2=5.645 $Y2=0.42
r178 24 60 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.2 $Y=0.555
+ $X2=8.2 $Y2=0.995
r179 19 21 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.17 $Y=1.57
+ $X2=8.17 $Y2=2.065
r180 18 19 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.17 $Y=1.47 $X2=8.17
+ $Y2=1.57
r181 18 61 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.17 $Y=1.47
+ $X2=8.17 $Y2=1.325
r182 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.805
r183 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.445
r184 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.955 $Y=1.99
+ $X2=6.955 $Y2=2.275
r185 10 57 11.0446 $w=1.9e-07 $l=1.35e-07 $layer=POLY_cond $X=6.96 $Y=1.095
+ $X2=6.96 $Y2=1.23
r186 9 27 153.83 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=6.96 $Y=0.805 $X2=7.26
+ $Y2=0.805
r187 9 10 77.3358 $w=1.9e-07 $l=2.15e-07 $layer=POLY_cond $X=6.96 $Y=0.88
+ $X2=6.96 $Y2=1.095
r188 8 11 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.955 $Y=1.89 $X2=6.955
+ $Y2=1.99
r189 7 56 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=6.955 $Y=1.365
+ $X2=6.955 $Y2=1.23
r190 7 8 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=6.955 $Y=1.365
+ $X2=6.955 $Y2=1.89
r191 2 35 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.065 $X2=5.52 $Y2=2.3
r192 1 31 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%SET_B 2 3 5 8 10 12 15 18 22 26 27 29 30
+ 32 33 35 42 53
c146 42 0 4.99305e-20 $X=7.53 $Y=1.53
c147 29 0 1.31062e-19 $X=9.675 $Y=1.53
c148 18 0 2.59025e-20 $X=7.567 $Y=1.365
c149 10 0 8.83008e-20 $X=10.495 $Y=1.99
c150 3 0 1.53071e-19 $X=7.54 $Y=1.99
r151 39 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.45
+ $Y=1.68 $X2=7.45 $Y2=1.68
r152 35 53 0.0545364 $w=2.3e-07 $l=8.5e-08 $layer=MET1_cond $X=7.53 $Y=1.53
+ $X2=7.615 $Y2=1.53
r153 35 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.53 $Y=1.53
+ $X2=7.53 $Y2=1.53
r154 33 48 3.98117 $w=2.73e-07 $l=9.5e-08 $layer=LI1_cond $X=9.822 $Y=1.53
+ $X2=9.822 $Y2=1.625
r155 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.82 $Y=1.53
+ $X2=9.82 $Y2=1.53
r156 30 53 0.0930106 $w=2.3e-07 $l=1.1e-07 $layer=MET1_cond $X=7.725 $Y=1.53
+ $X2=7.615 $Y2=1.53
r157 29 32 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.675 $Y=1.53
+ $X2=9.82 $Y2=1.53
r158 29 30 2.41336 $w=1.4e-07 $l=1.95e-06 $layer=MET1_cond $X=9.675 $Y=1.53
+ $X2=7.725 $Y2=1.53
r159 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.85
+ $Y=1.61 $X2=10.85 $Y2=1.61
r160 24 48 2.60351 $w=2e-07 $l=1.38e-07 $layer=LI1_cond $X=9.96 $Y=1.625
+ $X2=9.822 $Y2=1.625
r161 24 26 49.3545 $w=1.98e-07 $l=8.9e-07 $layer=LI1_cond $X=9.96 $Y=1.625
+ $X2=10.85 $Y2=1.625
r162 22 27 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=10.875 $Y=1.605
+ $X2=10.875 $Y2=1.61
r163 22 23 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=10.875 $Y=1.605
+ $X2=10.875 $Y2=1.445
r164 21 27 40.5733 $w=3.2e-07 $l=2.25e-07 $layer=POLY_cond $X=10.875 $Y=1.835
+ $X2=10.875 $Y2=1.61
r165 17 18 72.2668 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=7.567 $Y=1.16
+ $X2=7.567 $Y2=1.365
r166 15 23 512.766 $w=1.5e-07 $l=1e-06 $layer=POLY_cond $X=10.96 $Y=0.445
+ $X2=10.96 $Y2=1.445
r167 10 21 121.298 $w=1.51e-07 $l=3.8e-07 $layer=POLY_cond $X=10.495 $Y=1.912
+ $X2=10.875 $Y2=1.912
r168 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.495 $Y=1.99
+ $X2=10.495 $Y2=2.275
r169 8 17 366.628 $w=1.5e-07 $l=7.15e-07 $layer=POLY_cond $X=7.62 $Y=0.445
+ $X2=7.62 $Y2=1.16
r170 3 39 55.7735 $w=3.21e-07 $l=3.51255e-07 $layer=POLY_cond $X=7.54 $Y=1.99
+ $X2=7.452 $Y2=1.68
r171 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.54 $Y=1.99
+ $X2=7.54 $Y2=2.275
r172 2 39 31.5854 $w=3.21e-07 $l=2.04316e-07 $layer=POLY_cond $X=7.54 $Y=1.515
+ $X2=7.452 $Y2=1.68
r173 2 18 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.54 $Y=1.515 $X2=7.54
+ $Y2=1.365
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_1930_295# 1 2 8 9 11 12 13 16 19 22 23
+ 25 26 29 32 36 38
c108 26 0 6.89134e-20 $X=10.365 $Y=1.27
c109 9 0 9.89235e-21 $X=9.75 $Y=1.99
r110 34 36 3.23493 $w=2.83e-07 $l=8e-08 $layer=LI1_cond $X=11.775 $Y=0.397
+ $X2=11.855 $Y2=0.397
r111 32 38 4.14756 $w=2.2e-07 $l=1.03078e-07 $layer=LI1_cond $X=11.855 $Y=1.185
+ $X2=11.815 $Y2=1.27
r112 31 36 3.4259 $w=1.8e-07 $l=1.43e-07 $layer=LI1_cond $X=11.855 $Y=0.54
+ $X2=11.855 $Y2=0.397
r113 31 32 39.7424 $w=1.78e-07 $l=6.45e-07 $layer=LI1_cond $X=11.855 $Y=0.54
+ $X2=11.855 $Y2=1.185
r114 27 38 4.14756 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=11.815 $Y=1.355
+ $X2=11.815 $Y2=1.27
r115 27 29 41.222 $w=2.58e-07 $l=9.3e-07 $layer=LI1_cond $X=11.815 $Y=1.355
+ $X2=11.815 $Y2=2.285
r116 25 38 2.28545 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.685 $Y=1.27
+ $X2=11.815 $Y2=1.27
r117 25 26 86.1176 $w=1.68e-07 $l=1.32e-06 $layer=LI1_cond $X=11.685 $Y=1.27
+ $X2=10.365 $Y2=1.27
r118 23 41 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.255 $Y=1.02
+ $X2=10.255 $Y2=1.185
r119 23 40 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.255 $Y=1.02
+ $X2=10.255 $Y2=0.855
r120 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.23
+ $Y=1.02 $X2=10.23 $Y2=1.02
r121 20 26 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=10.252 $Y=1.185
+ $X2=10.365 $Y2=1.27
r122 20 22 8.45125 $w=2.23e-07 $l=1.65e-07 $layer=LI1_cond $X=10.252 $Y=1.185
+ $X2=10.252 $Y2=1.02
r123 19 41 96.1574 $w=2e-07 $l=2.9e-07 $layer=POLY_cond $X=10.195 $Y=1.475
+ $X2=10.195 $Y2=1.185
r124 16 40 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.17 $Y=0.445
+ $X2=10.17 $Y2=0.855
r125 12 19 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=10.095 $Y=1.55
+ $X2=10.195 $Y2=1.475
r126 12 13 125.628 $w=1.5e-07 $l=2.45e-07 $layer=POLY_cond $X=10.095 $Y=1.55
+ $X2=9.85 $Y2=1.55
r127 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.75 $Y=1.99
+ $X2=9.75 $Y2=2.275
r128 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.75 $Y=1.89 $X2=9.75
+ $Y2=1.99
r129 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=9.75 $Y=1.625
+ $X2=9.85 $Y2=1.55
r130 7 8 87.868 $w=2e-07 $l=2.65e-07 $layer=POLY_cond $X=9.75 $Y=1.625 $X2=9.75
+ $Y2=1.89
r131 2 29 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=11.625
+ $Y=2.065 $X2=11.77 $Y2=2.285
r132 1 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=11.64
+ $Y=0.235 $X2=11.775 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_1735_329# 1 2 3 11 12 14 17 18 20 22 23
+ 25 26 29 30 32 35 37 38 39 43 47 50 53 55 57 58 60 64 67 71 73
c172 67 0 4.09687e-20 $X=9.65 $Y=1.98
c173 64 0 1.93782e-19 $X=11.38 $Y=1.69
r174 74 75 23.2317 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.442 $Y=1.16
+ $X2=11.442 $Y2=1.325
r175 64 65 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.38
+ $Y=1.69 $X2=11.38 $Y2=1.69
r176 62 64 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=11.355 $Y=1.895
+ $X2=11.355 $Y2=1.69
r177 61 71 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=10.86 $Y=1.98
+ $X2=10.752 $Y2=1.98
r178 60 62 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=11.245 $Y=1.98
+ $X2=11.355 $Y2=1.895
r179 60 61 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=11.245 $Y=1.98
+ $X2=10.86 $Y2=1.98
r180 58 74 32.3836 $w=3.95e-07 $l=2.3e-07 $layer=POLY_cond $X=11.442 $Y=0.93
+ $X2=11.442 $Y2=1.16
r181 58 73 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=11.442 $Y=0.93
+ $X2=11.442 $Y2=0.765
r182 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.38
+ $Y=0.93 $X2=11.38 $Y2=0.93
r183 55 57 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.775 $Y=0.93
+ $X2=11.38 $Y2=0.93
r184 51 71 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.752 $Y=2.065
+ $X2=10.752 $Y2=1.98
r185 51 53 11.7924 $w=2.13e-07 $l=2.2e-07 $layer=LI1_cond $X=10.752 $Y=2.065
+ $X2=10.752 $Y2=2.285
r186 50 55 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.69 $Y=0.845
+ $X2=10.775 $Y2=0.93
r187 49 50 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=10.69 $Y=0.445
+ $X2=10.69 $Y2=0.845
r188 48 67 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.735 $Y=1.98
+ $X2=9.65 $Y2=1.98
r189 47 71 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=10.645 $Y=1.98
+ $X2=10.752 $Y2=1.98
r190 47 48 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=10.645 $Y=1.98
+ $X2=9.735 $Y2=1.98
r191 43 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.605 $Y=0.36
+ $X2=10.69 $Y2=0.445
r192 43 45 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=10.605 $Y=0.36
+ $X2=9.375 $Y2=0.36
r193 39 67 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=9.65 $Y=2.292
+ $X2=9.65 $Y2=1.98
r194 39 41 20.6408 $w=3.33e-07 $l=6e-07 $layer=LI1_cond $X=9.565 $Y=2.292
+ $X2=8.965 $Y2=2.292
r195 33 38 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=13.545 $Y=0.995
+ $X2=13.52 $Y2=1.16
r196 33 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=13.545 $Y=0.995
+ $X2=13.545 $Y2=0.445
r197 30 32 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=13.52 $Y=1.7
+ $X2=13.52 $Y2=2.095
r198 29 30 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=13.52 $Y=1.6 $X2=13.52
+ $Y2=1.7
r199 28 38 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=13.52 $Y=1.325
+ $X2=13.52 $Y2=1.16
r200 28 29 91.1837 $w=2e-07 $l=2.75e-07 $layer=POLY_cond $X=13.52 $Y=1.325
+ $X2=13.52 $Y2=1.6
r201 27 37 4.88773 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=12.63 $Y=1.16
+ $X2=12.53 $Y2=1.202
r202 26 38 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=13.42 $Y=1.16
+ $X2=13.52 $Y2=1.16
r203 26 27 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=13.42 $Y=1.16
+ $X2=12.63 $Y2=1.16
r204 23 37 21.2562 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.53 $Y=1.41
+ $X2=12.53 $Y2=1.202
r205 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.53 $Y=1.41
+ $X2=12.53 $Y2=1.985
r206 20 37 21.2562 $w=1.5e-07 $l=2.19144e-07 $layer=POLY_cond $X=12.505 $Y=0.995
+ $X2=12.53 $Y2=1.202
r207 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.505 $Y=0.995
+ $X2=12.505 $Y2=0.56
r208 19 74 7.07907 $w=3.3e-07 $l=1.98e-07 $layer=POLY_cond $X=11.64 $Y=1.16
+ $X2=11.442 $Y2=1.16
r209 18 37 4.88773 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=12.43 $Y=1.16
+ $X2=12.53 $Y2=1.202
r210 18 19 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=12.43 $Y=1.16
+ $X2=11.64 $Y2=1.16
r211 17 73 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.565 $Y=0.445
+ $X2=11.565 $Y2=0.765
r212 12 65 54.406 $w=3.19e-07 $l=3.44238e-07 $layer=POLY_cond $X=11.535 $Y=1.99
+ $X2=11.44 $Y2=1.69
r213 12 14 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.535 $Y=1.99
+ $X2=11.535 $Y2=2.275
r214 11 65 2.97574 $w=3.9e-07 $l=1e-08 $layer=POLY_cond $X=11.44 $Y=1.68
+ $X2=11.44 $Y2=1.69
r215 11 75 50.6243 $w=3.9e-07 $l=3.55e-07 $layer=POLY_cond $X=11.44 $Y=1.68
+ $X2=11.44 $Y2=1.325
r216 3 53 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=10.585
+ $Y=2.065 $X2=10.73 $Y2=2.285
r217 2 41 600 $w=1.7e-07 $l=7.76579e-07 $layer=licon1_PDIFF $count=1 $X=8.675
+ $Y=1.645 $X2=8.965 $Y2=2.29
r218 1 45 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=9.165
+ $Y=0.235 $X2=9.375 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_2632_47# 1 2 7 9 10 12 15 19 23 26
r45 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.965
+ $Y=1.16 $X2=13.965 $Y2=1.16
r46 21 26 0.221902 $w=3.3e-07 $l=1.05e-07 $layer=LI1_cond $X=13.37 $Y=1.16
+ $X2=13.265 $Y2=1.16
r47 21 23 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=13.37 $Y=1.16
+ $X2=13.965 $Y2=1.16
r48 17 26 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=13.265 $Y=1.325
+ $X2=13.265 $Y2=1.16
r49 17 19 31.9524 $w=2.08e-07 $l=6.05e-07 $layer=LI1_cond $X=13.265 $Y=1.325
+ $X2=13.265 $Y2=1.93
r50 13 26 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=13.265 $Y=0.995
+ $X2=13.265 $Y2=1.16
r51 13 15 29.3117 $w=2.08e-07 $l=5.55e-07 $layer=LI1_cond $X=13.265 $Y=0.995
+ $X2=13.265 $Y2=0.44
r52 10 24 38.6072 $w=2.91e-07 $l=2.02287e-07 $layer=POLY_cond $X=14.07 $Y=0.995
+ $X2=13.987 $Y2=1.16
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.07 $Y=0.995
+ $X2=14.07 $Y2=0.56
r54 7 24 48.3784 $w=2.91e-07 $l=2.77489e-07 $layer=POLY_cond $X=14.045 $Y=1.41
+ $X2=13.987 $Y2=1.16
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.045 $Y=1.41
+ $X2=14.045 $Y2=1.985
r56 2 19 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=13.16
+ $Y=1.775 $X2=13.285 $Y2=1.93
r57 1 15 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=13.16
+ $Y=0.235 $X2=13.285 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_27_369# 1 2 7 10 11 13 14 16
r52 14 16 46.2121 $w=2.08e-07 $l=8.75e-07 $layer=LI1_cond $X=1.205 $Y=2.36
+ $X2=2.08 $Y2=2.36
r53 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.12 $Y=2.255
+ $X2=1.205 $Y2=2.36
r54 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.12 $Y=2.025
+ $X2=1.12 $Y2=2.255
r55 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.035 $Y=1.935
+ $X2=1.12 $Y2=2.025
r56 10 11 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=1.035 $Y=1.935
+ $X2=0.345 $Y2=1.935
r57 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r58 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r59 2 16 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.845 $X2=2.08 $Y2=2.34
r60 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%VPWR 1 2 3 4 5 6 7 8 9 30 34 36 40 42 43
+ 46 50 52 56 62 67 69 70 72 73 74 76 81 86 105 117 118 121 124 127 134 139 141
+ 144 148
c214 118 0 1.67702e-19 $X=14.49 $Y=2.72
r215 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r216 142 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=12.19 $Y2=2.72
r217 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r218 137 139 11.292 $w=6.78e-07 $l=2e-07 $layer=LI1_cond $X=8.51 $Y=2.465
+ $X2=8.71 $Y2=2.465
r219 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r220 134 135 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r221 130 131 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r222 127 130 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=2.36
+ $X2=4.035 $Y2=2.72
r223 125 131 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r224 124 125 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r225 121 122 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r226 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r227 115 118 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.49 $Y2=2.72
r228 114 115 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r229 112 115 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.57 $Y2=2.72
r230 112 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r231 111 114 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.65 $Y=2.72
+ $X2=13.57 $Y2=2.72
r232 111 112 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r233 109 144 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=12.38 $Y=2.72
+ $X2=12.275 $Y2=2.72
r234 109 111 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.38 $Y=2.72
+ $X2=12.65 $Y2=2.72
r235 108 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r236 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r237 105 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.135 $Y=2.72
+ $X2=11.3 $Y2=2.72
r238 105 107 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=11.135 $Y=2.72
+ $X2=10.81 $Y2=2.72
r239 104 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r240 103 104 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r241 101 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r242 101 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r243 100 103 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r244 100 139 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=8.71 $Y2=2.72
r245 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r246 97 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r247 97 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r248 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r249 94 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.775 $Y=2.72
+ $X2=6.61 $Y2=2.72
r250 94 96 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=6.775 $Y=2.72
+ $X2=7.59 $Y2=2.72
r251 93 135 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r252 92 93 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r253 90 93 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r254 90 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r255 89 92 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r256 89 90 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r257 87 130 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.035 $Y2=2.72
r258 87 89 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.37 $Y2=2.72
r259 86 134 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.445 $Y=2.72
+ $X2=6.61 $Y2=2.72
r260 86 92 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.445 $Y=2.72
+ $X2=6.21 $Y2=2.72
r261 85 125 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r262 85 122 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r263 84 85 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r264 82 121 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.665 $Y2=2.72
r265 82 84 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r266 81 124 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=3.11 $Y2=2.72
r267 81 84 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=1.15 $Y2=2.72
r268 78 148 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r269 76 121 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.665 $Y2=2.72
r270 76 78 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r271 74 122 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r272 74 148 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r273 72 114 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=13.725 $Y=2.72
+ $X2=13.57 $Y2=2.72
r274 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.725 $Y=2.72
+ $X2=13.81 $Y2=2.72
r275 71 117 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=13.895 $Y=2.72
+ $X2=14.49 $Y2=2.72
r276 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.895 $Y=2.72
+ $X2=13.81 $Y2=2.72
r277 69 103 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=9.89 $Y2=2.72
r278 69 70 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.045 $Y=2.72
+ $X2=10.235 $Y2=2.72
r279 68 107 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=10.425 $Y=2.72
+ $X2=10.81 $Y2=2.72
r280 68 70 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.425 $Y=2.72
+ $X2=10.235 $Y2=2.72
r281 67 96 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=7.655 $Y=2.72
+ $X2=7.59 $Y2=2.72
r282 66 67 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.82 $Y=2.465
+ $X2=7.655 $Y2=2.465
r283 60 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.81 $Y=2.635
+ $X2=13.81 $Y2=2.72
r284 60 62 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=13.81 $Y=2.635
+ $X2=13.81 $Y2=1.9
r285 56 59 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=12.275 $Y=1.66
+ $X2=12.275 $Y2=2.34
r286 54 144 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=12.275 $Y=2.635
+ $X2=12.275 $Y2=2.72
r287 54 59 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=12.275 $Y=2.635
+ $X2=12.275 $Y2=2.34
r288 53 141 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.465 $Y=2.72
+ $X2=11.3 $Y2=2.72
r289 52 144 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=12.17 $Y=2.72
+ $X2=12.275 $Y2=2.72
r290 52 53 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=12.17 $Y=2.72
+ $X2=11.465 $Y2=2.72
r291 48 141 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.3 $Y=2.635
+ $X2=11.3 $Y2=2.72
r292 48 50 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=11.3 $Y=2.635
+ $X2=11.3 $Y2=2.34
r293 44 70 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.235 $Y=2.635
+ $X2=10.235 $Y2=2.72
r294 44 46 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=10.235 $Y=2.635
+ $X2=10.235 $Y2=2.36
r295 43 66 3.07814 $w=6.78e-07 $l=1.75e-07 $layer=LI1_cond $X=7.995 $Y=2.465
+ $X2=7.82 $Y2=2.465
r296 42 137 2.46251 $w=6.78e-07 $l=1.4e-07 $layer=LI1_cond $X=8.37 $Y=2.465
+ $X2=8.51 $Y2=2.465
r297 42 43 6.59602 $w=6.78e-07 $l=3.75e-07 $layer=LI1_cond $X=8.37 $Y=2.465
+ $X2=7.995 $Y2=2.465
r298 38 134 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.61 $Y=2.635
+ $X2=6.61 $Y2=2.72
r299 38 40 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.61 $Y=2.635
+ $X2=6.61 $Y2=2.36
r300 37 124 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.28 $Y=2.72
+ $X2=3.11 $Y2=2.72
r301 36 130 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=4.035 $Y2=2.72
r302 36 37 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=3.28 $Y2=2.72
r303 32 124 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=2.635
+ $X2=3.11 $Y2=2.72
r304 32 34 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.11 $Y=2.635
+ $X2=3.11 $Y2=2.34
r305 28 121 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.665 $Y=2.635
+ $X2=0.665 $Y2=2.72
r306 28 30 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=0.665 $Y=2.635
+ $X2=0.665 $Y2=2.36
r307 9 62 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=13.61
+ $Y=1.775 $X2=13.81 $Y2=1.9
r308 8 59 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=12.17
+ $Y=1.485 $X2=12.295 $Y2=2.34
r309 8 56 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=12.17
+ $Y=1.485 $X2=12.295 $Y2=1.66
r310 7 50 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=11.175
+ $Y=2.065 $X2=11.3 $Y2=2.34
r311 6 46 600 $w=1.7e-07 $l=4.96034e-07 $layer=licon1_PDIFF $count=1 $X=9.84
+ $Y=2.065 $X2=10.21 $Y2=2.36
r312 5 66 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=7.63
+ $Y=2.065 $X2=7.82 $Y2=2.36
r313 4 40 600 $w=1.7e-07 $l=3.84057e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=2.065 $X2=6.61 $Y2=2.36
r314 3 127 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.845 $X2=4.06 $Y2=2.36
r315 2 34 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.845 $X2=3.07 $Y2=2.34
r316 1 30 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%A_199_47# 1 2 3 4 13 19 21 23 29 33 36 37
+ 40 43 44
c126 43 0 4.73361e-19 $X=5.095 $Y=1.53
c127 37 0 1.59069e-19 $X=1.955 $Y=1.53
c128 29 0 1.6927e-19 $X=1.75 $Y=1.87
c129 19 0 8.99086e-20 $X=5.08 $Y=0.42
r130 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.095 $Y=1.53
+ $X2=5.095 $Y2=1.53
r131 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.76 $Y=1.53
+ $X2=1.76 $Y2=1.53
r132 37 39 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=1.955 $Y=1.53
+ $X2=1.76 $Y2=1.53
r133 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=5.095 $Y2=1.53
r134 36 37 3.70668 $w=1.4e-07 $l=2.995e-06 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=1.955 $Y2=1.53
r135 35 44 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.095 $Y=1.59
+ $X2=5.095 $Y2=1.53
r136 33 44 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.095 $Y=0.92
+ $X2=5.095 $Y2=1.53
r137 31 40 56.622 $w=1.88e-07 $l=9.7e-07 $layer=LI1_cond $X=1.75 $Y=0.56
+ $X2=1.75 $Y2=1.53
r138 29 40 19.8469 $w=1.88e-07 $l=3.4e-07 $layer=LI1_cond $X=1.75 $Y=1.87
+ $X2=1.75 $Y2=1.53
r139 26 29 7.57428 $w=2.03e-07 $l=1.4e-07 $layer=LI1_cond $X=1.61 $Y=1.972
+ $X2=1.75 $Y2=1.972
r140 21 35 6.3875 $w=2.18e-07 $l=1.1e-07 $layer=LI1_cond $X=5.07 $Y=1.7 $X2=5.07
+ $Y2=1.59
r141 21 23 31.4303 $w=2.18e-07 $l=6e-07 $layer=LI1_cond $X=5.07 $Y=1.7 $X2=5.07
+ $Y2=2.3
r142 17 33 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.017 $Y=0.758
+ $X2=5.017 $Y2=0.92
r143 17 19 11.9854 $w=3.23e-07 $l=3.38e-07 $layer=LI1_cond $X=5.017 $Y=0.758
+ $X2=5.017 $Y2=0.42
r144 13 31 7.1467 $w=2.8e-07 $l=1.81384e-07 $layer=LI1_cond $X=1.655 $Y=0.42
+ $X2=1.75 $Y2=0.56
r145 13 15 19.1388 $w=2.78e-07 $l=4.65e-07 $layer=LI1_cond $X=1.655 $Y=0.42
+ $X2=1.19 $Y2=0.42
r146 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=2.065 $X2=5.05 $Y2=2.3
r147 3 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=1.845 $X2=1.61 $Y2=1.97
r148 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.08 $Y2=0.42
r149 1 15 182 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_NDIFF $count=1 $X=0.995
+ $Y=0.235 $X2=1.19 $Y2=0.405
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%Q_N 1 2 7 8 9 10 11 12 20
r19 12 37 3.79093 $w=3.78e-07 $l=1.25e-07 $layer=LI1_cond $X=12.74 $Y=2.21
+ $X2=12.74 $Y2=2.335
r20 11 12 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=12.74 $Y=1.87
+ $X2=12.74 $Y2=2.21
r21 11 31 6.5204 $w=3.78e-07 $l=2.15e-07 $layer=LI1_cond $X=12.74 $Y=1.87
+ $X2=12.74 $Y2=1.655
r22 10 31 3.79093 $w=3.78e-07 $l=1.25e-07 $layer=LI1_cond $X=12.74 $Y=1.53
+ $X2=12.74 $Y2=1.655
r23 9 10 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=12.74 $Y=1.19
+ $X2=12.74 $Y2=1.53
r24 8 9 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=12.74 $Y=0.85
+ $X2=12.74 $Y2=1.19
r25 7 8 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=12.74 $Y=0.51
+ $X2=12.74 $Y2=0.85
r26 7 20 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=12.74 $Y=0.51
+ $X2=12.74 $Y2=0.38
r27 2 37 400 $w=1.7e-07 $l=9.19647e-07 $layer=licon1_PDIFF $count=1 $X=12.62
+ $Y=1.485 $X2=12.765 $Y2=2.335
r28 2 31 400 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=12.62
+ $Y=1.485 $X2=12.765 $Y2=1.655
r29 1 20 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=12.58
+ $Y=0.235 $X2=12.765 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%Q 1 2 7 8 9 10 11 12 24 38 45
r20 45 46 2.34364 $w=5.58e-07 $l=3.5e-08 $layer=LI1_cond $X=14.345 $Y=1.53
+ $X2=14.345 $Y2=1.495
r21 29 49 2.45623 $w=5.58e-07 $l=1.15e-07 $layer=LI1_cond $X=14.345 $Y=1.775
+ $X2=14.345 $Y2=1.66
r22 24 43 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=14.447 $Y=0.85
+ $X2=14.447 $Y2=0.825
r23 12 35 2.77661 $w=5.58e-07 $l=1.3e-07 $layer=LI1_cond $X=14.345 $Y=2.21
+ $X2=14.345 $Y2=2.34
r24 11 12 7.2619 $w=5.58e-07 $l=3.4e-07 $layer=LI1_cond $X=14.345 $Y=1.87
+ $X2=14.345 $Y2=2.21
r25 11 29 2.02906 $w=5.58e-07 $l=9.5e-08 $layer=LI1_cond $X=14.345 $Y=1.87
+ $X2=14.345 $Y2=1.775
r26 10 49 2.24265 $w=5.58e-07 $l=1.05e-07 $layer=LI1_cond $X=14.345 $Y=1.555
+ $X2=14.345 $Y2=1.66
r27 10 45 0.533964 $w=5.58e-07 $l=2.5e-08 $layer=LI1_cond $X=14.345 $Y=1.555
+ $X2=14.345 $Y2=1.53
r28 10 46 0.81158 $w=3.53e-07 $l=2.5e-08 $layer=LI1_cond $X=14.447 $Y=1.47
+ $X2=14.447 $Y2=1.495
r29 9 10 9.08969 $w=3.53e-07 $l=2.8e-07 $layer=LI1_cond $X=14.447 $Y=1.19
+ $X2=14.447 $Y2=1.47
r30 8 43 2.23684 $w=5.58e-07 $l=3e-08 $layer=LI1_cond $X=14.345 $Y=0.795
+ $X2=14.345 $Y2=0.825
r31 8 9 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=14.447 $Y=0.88
+ $X2=14.447 $Y2=1.19
r32 8 24 0.973895 $w=3.53e-07 $l=3e-08 $layer=LI1_cond $X=14.447 $Y=0.88
+ $X2=14.447 $Y2=0.85
r33 7 8 6.08718 $w=5.58e-07 $l=2.85e-07 $layer=LI1_cond $X=14.345 $Y=0.51
+ $X2=14.345 $Y2=0.795
r34 7 38 2.34944 $w=5.58e-07 $l=1.1e-07 $layer=LI1_cond $X=14.345 $Y=0.51
+ $X2=14.345 $Y2=0.4
r35 2 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.135
+ $Y=1.485 $X2=14.28 $Y2=1.66
r36 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.135
+ $Y=1.485 $X2=14.28 $Y2=2.34
r37 1 38 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=14.145
+ $Y=0.235 $X2=14.28 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSBP_1%VGND 1 2 3 4 5 6 7 8 9 28 30 34 36 40 44
+ 48 50 54 58 61 62 64 65 66 68 77 89 102 103 109 112 124 130 132 135 139
c183 130 0 2.59025e-20 $X=8.275 $Y=0.302
c184 103 0 2.71124e-20 $X=14.49 $Y=0
r185 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r186 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.27 $Y=0
+ $X2=12.19 $Y2=0
r187 132 133 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r188 128 130 12.2054 $w=7.73e-07 $l=2.25e-07 $layer=LI1_cond $X=8.05 $Y=0.302
+ $X2=8.275 $Y2=0.302
r189 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r190 126 128 2.62366 $w=7.73e-07 $l=1.7e-07 $layer=LI1_cond $X=7.88 $Y=0.302
+ $X2=8.05 $Y2=0.302
r191 123 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.05 $Y2=0
r192 122 126 4.47565 $w=7.73e-07 $l=2.9e-07 $layer=LI1_cond $X=7.59 $Y=0.302
+ $X2=7.88 $Y2=0.302
r193 122 124 9.5046 $w=7.73e-07 $l=5e-08 $layer=LI1_cond $X=7.59 $Y=0.302
+ $X2=7.54 $Y2=0.302
r194 122 123 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r195 112 113 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r196 110 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r197 109 110 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r198 106 139 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r199 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r200 100 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.49 $Y2=0
r201 99 100 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r202 97 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r203 97 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r204 96 99 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r205 96 97 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r206 94 135 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=12.38 $Y=0
+ $X2=12.275 $Y2=0
r207 94 96 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=12.38 $Y=0 $X2=12.65
+ $Y2=0
r208 93 133 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=11.27 $Y2=0
r209 93 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r210 92 130 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=8.51 $Y=0
+ $X2=8.275 $Y2=0
r211 92 93 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r212 89 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0
+ $X2=11.305 $Y2=0
r213 89 92 176.802 $w=1.68e-07 $l=2.71e-06 $layer=LI1_cond $X=11.22 $Y=0
+ $X2=8.51 $Y2=0
r214 88 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r215 88 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=6.21 $Y2=0
r216 87 124 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=7.54
+ $Y2=0
r217 87 88 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r218 85 87 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.67
+ $Y2=0
r219 83 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r220 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r221 80 83 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r222 79 82 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r223 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r224 77 119 8.49551 $w=5.33e-07 $l=3.8e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.327 $Y2=0.38
r225 77 85 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.595 $Y2=0
r226 77 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r227 77 82 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=5.75
+ $Y2=0
r228 76 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r229 76 113 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=2.99 $Y2=0
r230 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r231 73 112 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.11
+ $Y2=0
r232 73 75 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.28 $Y=0 $X2=3.91
+ $Y2=0
r233 72 110 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r234 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r235 69 106 4.96256 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=0
+ $X2=0.215 $Y2=0
r236 69 71 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.69
+ $Y2=0
r237 68 109 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.115
+ $Y2=0
r238 68 71 87.0963 $w=1.68e-07 $l=1.335e-06 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=0.69 $Y2=0
r239 66 72 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r240 66 139 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r241 64 99 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=13.69 $Y=0
+ $X2=13.57 $Y2=0
r242 64 65 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=13.69 $Y=0
+ $X2=13.792 $Y2=0
r243 63 102 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=13.895 $Y=0
+ $X2=14.49 $Y2=0
r244 63 65 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=13.895 $Y=0
+ $X2=13.792 $Y2=0
r245 61 75 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.93 $Y=0 $X2=3.91
+ $Y2=0
r246 61 62 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=3.93 $Y=0 $X2=4.085
+ $Y2=0
r247 60 79 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.37
+ $Y2=0
r248 60 62 8.23795 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=4.24 $Y=0 $X2=4.085
+ $Y2=0
r249 56 65 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=13.792 $Y=0.085
+ $X2=13.792 $Y2=0
r250 56 58 18.6652 $w=2.03e-07 $l=3.45e-07 $layer=LI1_cond $X=13.792 $Y=0.085
+ $X2=13.792 $Y2=0.43
r251 52 135 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=12.275 $Y=0.085
+ $X2=12.275 $Y2=0
r252 52 54 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=12.275 $Y=0.085
+ $X2=12.275 $Y2=0.38
r253 51 132 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.39 $Y=0
+ $X2=11.305 $Y2=0
r254 50 135 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=12.17 $Y=0
+ $X2=12.275 $Y2=0
r255 50 51 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=12.17 $Y=0
+ $X2=11.39 $Y2=0
r256 46 132 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.305 $Y=0.085
+ $X2=11.305 $Y2=0
r257 46 48 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.305 $Y=0.085
+ $X2=11.305 $Y2=0.36
r258 42 62 0.701276 $w=3.1e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r259 42 44 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.36
r260 38 112 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0
r261 38 40 9.99914 $w=3.38e-07 $l=2.95e-07 $layer=LI1_cond $X=3.11 $Y=0.085
+ $X2=3.11 $Y2=0.38
r262 37 109 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.115
+ $Y2=0
r263 36 112 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.11
+ $Y2=0
r264 36 37 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.94 $Y=0
+ $X2=2.205 $Y2=0
r265 32 109 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0
r266 32 34 18.1768 $w=1.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.115 $Y=0.085
+ $X2=2.115 $Y2=0.38
r267 28 106 2.93137 $w=3.45e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.215 $Y2=0
r268 28 30 11.5244 $w=3.43e-07 $l=3.45e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.43
r269 9 58 182 $w=1.7e-07 $l=2.73998e-07 $layer=licon1_NDIFF $count=1 $X=13.62
+ $Y=0.235 $X2=13.81 $Y2=0.43
r270 8 54 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=12.17
+ $Y=0.235 $X2=12.295 $Y2=0.38
r271 7 48 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.235 $X2=11.305 $Y2=0.36
r272 6 126 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.695
+ $Y=0.235 $X2=7.88 $Y2=0.36
r273 5 119 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.245
+ $Y=0.235 $X2=6.43 $Y2=0.38
r274 4 44 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.36
r275 3 40 182 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=1 $X=2.935
+ $Y=0.235 $X2=3.1 $Y2=0.38
r276 2 34 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.11 $Y2=0.38
r277 1 30 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

