* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 a_530_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_334_297# A0 a_424_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND a_424_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_27_47# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VPWR a_424_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND a_27_47# a_226_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 X a_424_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 X a_424_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_424_297# A1 a_530_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_334_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND a_424_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR a_27_47# a_222_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_27_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 X a_424_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_226_47# A0 a_424_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VPWR a_424_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 X a_424_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_424_297# A1 a_222_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
