* File: sky130_fd_sc_hdll__and2b_1.spice
* Created: Wed Sep  2 08:21:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and2b_1.pex.spice"
.subckt sky130_fd_sc_hdll__and2b_1  VNB VPB A_N B VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1006 N_A_27_413#_M1006_d N_A_N_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 A_327_47# N_A_27_413#_M1003_g N_A_225_413#_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0609 AS=0.1302 PD=0.71 PS=1.46 NRD=25.704 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_B_M1001_g A_327_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0922822 AS=0.0609 PD=0.816449 PS=0.71 NRD=18.564 NRS=25.704 M=1 R=2.8
+ SA=75000.7 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_X_M1004_d N_A_225_413#_M1004_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.195 AS=0.142818 PD=1.9 PS=1.26355 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_413#_M1000_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0756 AS=0.1134 PD=0.78 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1002 N_A_225_413#_M1002_d N_A_27_413#_M1002_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0651 AS=0.0756 PD=0.73 PS=0.78 NRD=7.0329 NRS=35.1645 M=1
+ R=2.33333 SA=90000.7 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_B_M1007_g N_A_225_413#_M1002_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.145225 AS=0.0651 PD=1.0707 PS=0.73 NRD=25.7873 NRS=7.0329 M=1 R=2.33333
+ SA=90001.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1005 N_X_M1005_d N_A_225_413#_M1005_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.31 AS=0.345775 PD=2.62 PS=2.5493 NRD=8.8453 NRS=18.715 M=1 R=5.55556
+ SA=90001 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX9_noxref noxref_11 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and2b_1.pxi.spice"
*
.ends
*
*
