* File: sky130_fd_sc_hdll__mux2i_4.spice
* Created: Wed Sep  2 08:35:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2i_4.pex.spice"
.subckt sky130_fd_sc_hdll__mux2i_4  VNB VPB A0 A1 S Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1010 N_A_109_47#_M1010_d N_A0_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1012 N_A_109_47#_M1010_d N_A0_M1012_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1025 N_A_109_47#_M1025_d N_A0_M1025_g N_Y_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1032 N_A_109_47#_M1025_d N_A0_M1032_g N_Y_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1032_s N_A1_M1013_g N_A_485_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1019 N_Y_M1019_d N_A1_M1019_g N_A_485_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1026 N_Y_M1019_d N_A1_M1026_g N_A_485_47#_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1027 N_Y_M1027_d N_A1_M1027_g N_A_485_47#_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_S_M1006_g N_A_485_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_S_M1008_g N_A_485_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1008_d N_S_M1016_g N_A_485_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1024_d N_S_M1024_g N_A_485_47#_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1024_d N_A_1311_21#_M1001_g N_A_109_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.1 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_1311_21#_M1004_g N_A_109_47#_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75002.5 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1004_d N_A_1311_21#_M1021_g N_A_109_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.138125 PD=0.97 PS=1.075 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75003 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1028 N_VGND_M1028_d N_A_1311_21#_M1028_g N_A_109_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.118625 AS=0.138125 PD=1.015 PS=1.075 NRD=7.38 NRS=18.456 M=1
+ R=4.33333 SA=75003.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1029 N_A_1311_21#_M1029_d N_S_M1029_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.118625 PD=1.82 PS=1.015 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_Y_M1002_d N_A0_M1002_g N_A_117_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1015_d N_A0_M1015_g N_A_117_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1022 N_Y_M1015_d N_A0_M1022_g N_A_117_297#_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1030 N_Y_M1030_d N_A0_M1030_g N_A_117_297#_M1022_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1030_d N_A1_M1000_g N_A_493_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g N_A_493_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1007_d N_A1_M1011_g N_A_493_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1017 N_Y_M1017_d N_A1_M1017_g N_A_493_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_117_297#_M1005_d N_S_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004 A=0.18 P=2.36 MULT=1
MM1009 N_A_117_297#_M1005_d N_S_M1009_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003.6 A=0.18 P=2.36 MULT=1
MM1020 N_A_117_297#_M1020_d N_S_M1020_g N_VPWR_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1031 N_A_117_297#_M1020_d N_S_M1031_g N_VPWR_M1031_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1031_s N_A_1311_21#_M1003_g N_A_493_297#_M1003_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.1 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_A_1311_21#_M1014_g N_A_493_297#_M1003_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.5 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1014_d N_A_1311_21#_M1018_g N_A_493_297#_M1018_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.1725 PD=1.29 PS=1.345 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1023_d N_A_1311_21#_M1023_g N_A_493_297#_M1018_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.1675 AS=0.1725 PD=1.335 PS=1.345 NRD=9.8303 NRS=11.8003 M=1
+ R=5.55556 SA=90003.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1033 N_A_1311_21#_M1033_d N_S_M1033_g N_VPWR_M1023_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.1675 PD=2.54 PS=1.335 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004 SB=90000.2 A=0.18 P=2.36 MULT=1
DX34_noxref VNB VPB NWDIODE A=15.3759 P=22.37
*
.include "sky130_fd_sc_hdll__mux2i_4.pxi.spice"
*
.ends
*
*
