* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__einvn_2 A TE_B VGND VNB VPB VPWR Z
M1000 VPWR TE_B a_222_309# VPB phighvt w=940000u l=180000u
+  ad=5.526e+11p pd=4.99e+06u as=5.626e+11p ps=5.04e+06u
M1001 VPWR TE_B a_27_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1002 a_222_309# TE_B VPWR VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_234_47# A Z VNB nshort w=650000u l=150000u
+  ad=6.5975e+11p pd=5.93e+06u as=2.08e+11p ps=1.94e+06u
M1004 VGND TE_B a_27_47# VNB nshort w=420000u l=150000u
+  ad=2.847e+11p pd=3.2e+06u as=1.302e+11p ps=1.46e+06u
M1005 a_234_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_27_47# a_234_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 Z A a_222_309# VPB phighvt w=1e+06u l=180000u
+  ad=5.6e+11p pd=5.12e+06u as=0p ps=0u
M1008 Z A a_234_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_222_309# A Z VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
