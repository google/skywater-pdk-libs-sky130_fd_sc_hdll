* NGSPICE file created from sky130_fd_sc_hdll__o21a_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
M1000 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6e+11p pd=5.2e+06u as=1.76e+12p ps=1.352e+07u
M1001 a_80_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=6.5e+11p pd=5.3e+06u as=0p ps=0u
M1002 X a_80_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_525_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=8.84e+11p pd=7.92e+06u as=1.0075e+12p ps=9.6e+06u
M1004 a_80_21# A2 a_826_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.5e+11p ps=2.5e+06u
M1005 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1006 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND A2 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR A1 a_1008_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=3e+11p ps=2.6e+06u
M1009 X a_80_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR B1 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_525_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_525_47# B1 a_80_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.755e+11p ps=1.84e+06u
M1014 a_826_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_80_21# B1 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_525_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_80_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_80_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_1008_297# A2 a_80_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

