# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o211ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o211ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.400000 1.075000 1.560000 1.330000 ;
        RECT 1.015000 1.330000 1.560000 1.515000 ;
        RECT 1.015000 1.515000 4.030000 1.685000 ;
        RECT 3.700000 0.995000 4.030000 1.515000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.855000 1.075000 3.530000 1.345000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.200000 0.995000 5.525000 1.410000 ;
        RECT 4.710000 1.410000 5.525000 1.515000 ;
        RECT 4.710000 1.515000 7.800000 1.685000 ;
        RECT 7.580000 0.995000 7.800000 1.515000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.970000 1.075000 7.140000 1.345000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  0.832000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.740000 0.085000 ;
        RECT 0.525000  0.085000 0.905000 0.445000 ;
        RECT 1.535000  0.085000 1.865000 0.455000 ;
        RECT 2.445000  0.085000 2.825000 0.445000 ;
        RECT 3.405000  0.085000 3.785000 0.445000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.480000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.740000 2.805000 ;
        RECT 0.090000 1.665000 0.385000 2.635000 ;
        RECT 1.005000 2.275000 1.385000 2.635000 ;
        RECT 4.015000 2.195000 4.285000 2.635000 ;
        RECT 4.885000 2.275000 5.265000 2.635000 ;
        RECT 5.830000 2.275000 6.210000 2.635000 ;
        RECT 6.770000 2.275000 7.155000 2.635000 ;
        RECT 8.155000 2.275000 8.485000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.218500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 1.855000 8.480000 2.025000 ;
        RECT 1.955000 2.025000 3.820000 2.105000 ;
        RECT 4.495000 2.025000 8.480000 2.105000 ;
        RECT 5.830000 0.270000 7.485000 0.450000 ;
        RECT 7.265000 0.450000 7.485000 0.655000 ;
        RECT 7.265000 0.655000 8.160000 0.825000 ;
        RECT 7.980000 0.825000 8.160000 1.340000 ;
        RECT 7.980000 1.340000 8.480000 1.855000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.155000 0.535000 0.355000 0.625000 ;
      RECT 0.155000 0.625000 4.235000 0.795000 ;
      RECT 0.155000 0.795000 3.480000 0.905000 ;
      RECT 0.605000 1.860000 0.825000 1.935000 ;
      RECT 0.605000 1.935000 1.785000 2.105000 ;
      RECT 0.605000 2.105000 0.825000 2.190000 ;
      RECT 1.125000 0.425000 1.340000 0.625000 ;
      RECT 1.605000 2.105000 1.785000 2.275000 ;
      RECT 1.605000 2.275000 3.785000 2.465000 ;
      RECT 4.005000 0.255000 5.470000 0.455000 ;
      RECT 4.005000 0.455000 4.235000 0.625000 ;
      RECT 4.405000 0.635000 6.870000 0.815000 ;
      RECT 7.730000 0.310000 8.490000 0.480000 ;
      RECT 8.320000 0.480000 8.490000 0.595000 ;
    LAYER mcon ;
      RECT 1.170000 0.425000 1.340000 0.595000 ;
      RECT 8.320000 0.425000 8.490000 0.595000 ;
    LAYER met1 ;
      RECT 1.110000 0.395000 1.400000 0.440000 ;
      RECT 1.110000 0.440000 8.550000 0.580000 ;
      RECT 1.110000 0.580000 1.400000 0.625000 ;
      RECT 8.260000 0.395000 8.550000 0.440000 ;
      RECT 8.260000 0.580000 8.550000 0.625000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o211ai_4
