# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and3_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and3_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.995000 0.875000 1.340000 ;
        RECT 0.115000 1.340000 0.330000 2.335000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.045000 0.745000 1.355000 1.340000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.995000 2.050000 1.325000 ;
    END
  END C
  PIN VGND
    ANTENNADIFFAREA  0.708500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  1.435000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  1.061500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.650000 0.515000 2.840000 0.615000 ;
        RECT 2.650000 0.615000 4.490000 0.845000 ;
        RECT 2.650000 1.535000 4.490000 1.760000 ;
        RECT 2.650000 1.760000 2.840000 2.465000 ;
        RECT 3.610000 0.255000 3.800000 0.615000 ;
        RECT 3.610000 1.760000 4.490000 1.765000 ;
        RECT 3.610000 1.765000 3.800000 2.465000 ;
        RECT 4.210000 0.845000 4.490000 1.535000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.465000  0.255000 1.825000 0.445000 ;
      RECT 0.465000  0.445000 0.800000 0.805000 ;
      RECT 0.500000  1.580000 2.430000 1.750000 ;
      RECT 0.500000  1.750000 0.680000 2.465000 ;
      RECT 0.895000  1.935000 1.395000 2.635000 ;
      RECT 1.620000  1.750000 1.800000 2.465000 ;
      RECT 1.635000  0.445000 1.825000 0.615000 ;
      RECT 1.635000  0.615000 2.430000 0.805000 ;
      RECT 2.055000  0.085000 2.385000 0.445000 ;
      RECT 2.060000  1.935000 2.390000 2.635000 ;
      RECT 2.220000  0.805000 2.430000 1.020000 ;
      RECT 2.220000  1.020000 3.905000 1.355000 ;
      RECT 2.220000  1.355000 2.430000 1.580000 ;
      RECT 3.010000  0.085000 3.390000 0.445000 ;
      RECT 3.010000  1.935000 3.390000 2.635000 ;
      RECT 3.970000  0.085000 4.350000 0.445000 ;
      RECT 3.970000  1.935000 4.350000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and3_4
END LIBRARY
