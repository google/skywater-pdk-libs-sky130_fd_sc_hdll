* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2oi_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
M1000 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.99e+12p pd=1.798e+07u as=1.74e+12p ps=1.548e+07u
M1001 VGND A1_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=2.067e+12p pd=1.806e+07u as=8.97e+11p ps=7.96e+06u
M1002 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_831_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_27_297# a_831_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1005 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_831_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=8.97e+11p ps=7.96e+06u
M1007 a_831_21# A2_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=1.43e+12p ps=1.286e+07u
M1008 Y a_831_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y a_831_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.995e+11p ps=7.66e+06u
M1012 VGND B1 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VPWR A1_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_109_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_831_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_1259_297# A2_N a_831_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_831_21# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND A1_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1259_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_831_21# A2_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_27_297# a_831_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 a_831_21# A1_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VGND A2_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_27_297# B2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1027 VPWR A1_N a_1259_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_1259_297# A1_N VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1029 Y a_831_21# a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 Y B2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_109_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_109_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 Y B2 a_109_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1035 Y a_831_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_1259_297# A2_N a_831_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_831_21# A2_N VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_109_47# B1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND A2_N a_831_21# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
