* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and3b_2 A_N B C VGND VNB VPB VPWR X
M1000 a_117_311# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.176e+11p pd=1.4e+06u as=6.936e+11p ps=5.94e+06u
M1001 a_317_53# a_117_311# a_225_311# VNB nshort w=420000u l=150000u
+  ad=1.344e+11p pd=1.48e+06u as=1.218e+11p ps=1.42e+06u
M1002 a_117_311# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=9.409e+11p ps=8.31e+06u
M1003 a_225_311# B VPWR VPB phighvt w=420000u l=180000u
+  ad=2.7055e+11p pd=3.05e+06u as=0p ps=0u
M1004 VPWR C a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_225_311# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1006 X a_225_311# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR a_117_311# a_225_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_225_311# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1009 a_411_53# B a_317_53# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=0p ps=0u
M1010 VGND C a_411_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_225_311# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
