* File: sky130_fd_sc_hdll__inv_2.pex.spice
* Created: Wed Sep  2 08:33:04 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_2%A 1 3 4 6 7 9 10 12 13 20
r35 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.975 $Y=1.202
+ $X2=1 $Y2=1.202
r36 19 20 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=0.53 $Y=1.202
+ $X2=0.975 $Y2=1.202
r37 18 19 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.505 $Y=1.202
+ $X2=0.53 $Y2=1.202
r38 16 18 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=0.27 $Y=1.202
+ $X2=0.505 $Y2=1.202
r39 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r40 10 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=1.202
r41 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1 $Y=0.995 $X2=1
+ $Y2=0.56
r42 7 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.202
r43 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
r44 4 19 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.53 $Y=0.995
+ $X2=0.53 $Y2=1.202
r45 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.53 $Y=0.995 $X2=0.53
+ $Y2=0.56
r46 1 18 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.202
r47 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_2%VPWR 1 2 7 9 13 17 21 25 26 32
r22 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r23 26 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r24 25 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r25 23 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.23 $Y2=2.72
r26 23 25 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 21 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r28 21 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r29 17 20 35.9134 $w=2.08e-07 $l=6.8e-07 $layer=LI1_cond $X=1.23 $Y=1.66
+ $X2=1.23 $Y2=2.34
r30 15 32 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r31 15 20 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.34
r32 14 29 3.83185 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=2.72
+ $X2=0.177 $Y2=2.72
r33 13 32 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.125 $Y=2.72
+ $X2=1.23 $Y2=2.72
r34 13 14 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.125 $Y=2.72
+ $X2=0.355 $Y2=2.72
r35 9 12 34.0722 $w=2.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.24 $Y=1.66 $X2=0.24
+ $Y2=2.34
r36 7 29 3.18603 $w=2.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.177 $Y2=2.72
r37 7 12 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=2.635
+ $X2=0.24 $Y2=2.34
r38 2 20 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.485 $X2=1.21 $Y2=2.34
r39 2 17 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.485 $X2=1.21 $Y2=1.66
r40 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=2.34
r41 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_2%Y 1 2 9 13 15 16 17 31 34
r24 34 35 1.90772 $w=3.78e-07 $l=4.5e-08 $layer=LI1_cond $X=0.715 $Y=1.53
+ $X2=0.715 $Y2=1.485
r25 31 32 1.60444 $w=3.78e-07 $l=3.5e-08 $layer=LI1_cond $X=0.715 $Y=0.85
+ $X2=0.715 $Y2=0.885
r26 17 38 3.33602 $w=3.78e-07 $l=1.1e-07 $layer=LI1_cond $X=0.715 $Y=1.55
+ $X2=0.715 $Y2=1.66
r27 17 34 0.606549 $w=3.78e-07 $l=2e-08 $layer=LI1_cond $X=0.715 $Y=1.55
+ $X2=0.715 $Y2=1.53
r28 17 35 0.768295 $w=2.98e-07 $l=2e-08 $layer=LI1_cond $X=0.755 $Y=1.465
+ $X2=0.755 $Y2=1.485
r29 16 17 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=0.755 $Y=1.19
+ $X2=0.755 $Y2=1.465
r30 15 31 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=0.715 $Y=0.825
+ $X2=0.715 $Y2=0.85
r31 15 16 10.7561 $w=2.98e-07 $l=2.8e-07 $layer=LI1_cond $X=0.755 $Y=0.91
+ $X2=0.755 $Y2=1.19
r32 15 32 0.960369 $w=2.98e-07 $l=2.5e-08 $layer=LI1_cond $X=0.755 $Y=0.91
+ $X2=0.755 $Y2=0.885
r33 11 38 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.715 $Y=1.675
+ $X2=0.715 $Y2=1.66
r34 11 13 20.1678 $w=3.78e-07 $l=6.65e-07 $layer=LI1_cond $X=0.715 $Y=1.675
+ $X2=0.715 $Y2=2.34
r35 7 15 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=0.715 $Y=0.695
+ $X2=0.715 $Y2=0.825
r36 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.715 $Y=0.695
+ $X2=0.715 $Y2=0.38
r37 2 38 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=1.66
r38 2 13 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=1.485 $X2=0.74 $Y2=2.34
r39 1 9 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=0.605
+ $Y=0.235 $X2=0.74 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_2%VGND 1 2 7 9 11 15 17 21 22 28
r22 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r23 22 29 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r24 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r25 19 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.23
+ $Y2=0
r26 19 21 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=1.335 $Y=0 $X2=1.61
+ $Y2=0
r27 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r28 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r29 13 28 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r30 13 15 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.38
r31 12 25 3.83185 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r32 11 28 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=1.23
+ $Y2=0
r33 11 12 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.125 $Y=0 $X2=0.355
+ $Y2=0
r34 7 25 3.18603 $w=2.3e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.177 $Y2=0
r35 7 9 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.24 $Y=0.085
+ $X2=0.24 $Y2=0.38
r36 2 15 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.21 $Y2=0.38
r37 1 9 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.38
.ends

