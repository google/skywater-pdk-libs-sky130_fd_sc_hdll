* File: sky130_fd_sc_hdll__o21ba_4.pex.spice
* Created: Wed Sep  2 08:44:00 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%B1_N 1 3 4 6 7 8 14
r36 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r37 8 14 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=0.77 $Y=1.53
+ $X2=0.77 $Y2=1.285
r38 7 14 4.22511 $w=2.08e-07 $l=8e-08 $layer=LI1_cond $X=0.69 $Y=1.18 $X2=0.77
+ $Y2=1.18
r39 7 13 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.69 $Y=1.18 $X2=0.59
+ $Y2=1.18
r40 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=0.64 $Y=0.995
+ $X2=0.615 $Y2=1.16
r41 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.64 $Y=0.995 $X2=0.64
+ $Y2=0.56
r42 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=0.615 $Y=1.41
+ $X2=0.615 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.615 $Y=1.41
+ $X2=0.615 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A_197_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 40 41 42 45 47 48 49 51 53 56 59 69
c162 69 0 1.33641e-19 $X=2.495 $Y=1.202
c163 47 0 8.46699e-20 $X=3.84 $Y=0.895
c164 42 0 1.24542e-19 $X=2.815 $Y=0.77
c165 28 0 1.73969e-19 $X=2.495 $Y=1.41
r166 69 70 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.495 $Y=1.202
+ $X2=2.52 $Y2=1.202
r167 66 67 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2 $Y=1.202
+ $X2=2.025 $Y2=1.202
r168 65 66 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.555 $Y=1.202
+ $X2=2 $Y2=1.202
r169 64 65 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.53 $Y=1.202
+ $X2=1.555 $Y2=1.202
r170 63 64 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.085 $Y=1.202
+ $X2=1.53 $Y2=1.202
r171 62 63 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.06 $Y=1.202
+ $X2=1.085 $Y2=1.202
r172 51 61 3.19664 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=4.707 $Y=1.795
+ $X2=4.707 $Y2=1.96
r173 51 53 8.23174 $w=2.43e-07 $l=1.75e-07 $layer=LI1_cond $X=4.707 $Y=1.795
+ $X2=4.707 $Y2=1.62
r174 50 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.935 $Y=1.88
+ $X2=3.84 $Y2=1.88
r175 49 61 3.91346 $w=1.7e-07 $l=1.56984e-07 $layer=LI1_cond $X=4.585 $Y=1.88
+ $X2=4.707 $Y2=1.96
r176 49 50 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=4.585 $Y=1.88
+ $X2=3.935 $Y2=1.88
r177 48 59 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.84 $Y=1.795
+ $X2=3.84 $Y2=1.88
r178 47 58 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=3.84 $Y=0.895
+ $X2=3.84 $Y2=0.77
r179 47 48 52.5359 $w=1.88e-07 $l=9e-07 $layer=LI1_cond $X=3.84 $Y=0.895
+ $X2=3.84 $Y2=1.795
r180 46 56 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.285 $Y=1.88
+ $X2=3.2 $Y2=1.88
r181 45 59 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.745 $Y=1.88
+ $X2=3.84 $Y2=1.88
r182 45 46 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.745 $Y=1.88
+ $X2=3.285 $Y2=1.88
r183 41 58 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=3.745 $Y=0.77
+ $X2=3.84 $Y2=0.77
r184 41 42 42.8709 $w=2.48e-07 $l=9.3e-07 $layer=LI1_cond $X=3.745 $Y=0.77
+ $X2=2.815 $Y2=0.77
r185 39 42 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.73 $Y=0.895
+ $X2=2.815 $Y2=0.77
r186 39 40 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.73 $Y=0.895
+ $X2=2.73 $Y2=1.08
r187 37 69 8.42204 $w=3.72e-07 $l=6.5e-08 $layer=POLY_cond $X=2.43 $Y=1.202
+ $X2=2.495 $Y2=1.202
r188 37 67 52.4758 $w=3.72e-07 $l=4.05e-07 $layer=POLY_cond $X=2.43 $Y=1.202
+ $X2=2.025 $Y2=1.202
r189 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.43
+ $Y=1.165 $X2=2.43 $Y2=1.165
r190 34 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=1.165
+ $X2=2.73 $Y2=1.08
r191 34 36 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.645 $Y=1.165
+ $X2=2.43 $Y2=1.165
r192 31 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=1.202
r193 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.52 $Y=0.995
+ $X2=2.52 $Y2=0.56
r194 28 69 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=1.202
r195 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=1.985
r196 25 67 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.025 $Y=1.41
+ $X2=2.025 $Y2=1.202
r197 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.025 $Y=1.41
+ $X2=2.025 $Y2=1.985
r198 22 66 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2 $Y=0.995 $X2=2
+ $Y2=1.202
r199 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2 $Y=0.995 $X2=2
+ $Y2=0.56
r200 19 65 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.555 $Y=1.41
+ $X2=1.555 $Y2=1.202
r201 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.555 $Y=1.41
+ $X2=1.555 $Y2=1.985
r202 16 64 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=1.202
r203 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.53 $Y=0.995
+ $X2=1.53 $Y2=0.56
r204 13 63 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.085 $Y=1.41
+ $X2=1.085 $Y2=1.202
r205 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.085 $Y=1.41
+ $X2=1.085 $Y2=1.985
r206 10 62 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.06 $Y=0.995
+ $X2=1.06 $Y2=1.202
r207 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.06 $Y=0.995
+ $X2=1.06 $Y2=0.56
r208 3 61 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.71 $Y2=1.96
r209 3 53 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.565
+ $Y=1.485 $X2=4.71 $Y2=1.62
r210 2 56 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.055
+ $Y=1.485 $X2=3.2 $Y2=1.96
r211 1 58 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.77 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A_27_297# 1 2 7 9 10 12 13 15 16 18 22 25
+ 27 30 32 34 38 39 41 49 55
c108 49 0 1.33641e-19 $X=3.27 $Y=1.16
c109 32 0 1.73969e-19 $X=3.095 $Y=1.445
c110 7 0 1.54638e-19 $X=2.965 $Y=1.41
r111 55 56 63.2793 $w=3.58e-07 $l=4.7e-07 $layer=POLY_cond $X=3.51 $Y=1.202
+ $X2=3.98 $Y2=1.202
r112 54 55 10.0978 $w=3.58e-07 $l=7.5e-08 $layer=POLY_cond $X=3.435 $Y=1.202
+ $X2=3.51 $Y2=1.202
r113 50 54 22.2151 $w=3.58e-07 $l=1.65e-07 $layer=POLY_cond $X=3.27 $Y=1.202
+ $X2=3.435 $Y2=1.202
r114 50 52 41.0642 $w=3.58e-07 $l=3.05e-07 $layer=POLY_cond $X=3.27 $Y=1.202
+ $X2=2.965 $Y2=1.202
r115 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.27
+ $Y=1.16 $X2=3.27 $Y2=1.16
r116 38 39 8.48848 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.26 $Y=1.62
+ $X2=0.26 $Y2=1.455
r117 36 39 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=0.17 $Y=0.855
+ $X2=0.17 $Y2=1.455
r118 34 36 17.0806 $w=4.58e-07 $l=4.65e-07 $layer=LI1_cond $X=0.315 $Y=0.39
+ $X2=0.315 $Y2=0.855
r119 32 42 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=3.095 $Y=1.53
+ $X2=2.73 $Y2=1.53
r120 31 49 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.095 $Y=1.16
+ $X2=3.27 $Y2=1.16
r121 31 32 10.4768 $w=2.18e-07 $l=2e-07 $layer=LI1_cond $X=3.095 $Y=1.245
+ $X2=3.095 $Y2=1.445
r122 29 42 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=1.615
+ $X2=2.73 $Y2=1.53
r123 29 30 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=2.73 $Y=1.615
+ $X2=2.73 $Y2=1.875
r124 28 41 4.03347 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.435 $Y=1.96
+ $X2=0.26 $Y2=1.96
r125 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.645 $Y=1.96
+ $X2=2.73 $Y2=1.875
r126 27 28 144.182 $w=1.68e-07 $l=2.21e-06 $layer=LI1_cond $X=2.645 $Y=1.96
+ $X2=0.435 $Y2=1.96
r127 23 41 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=1.96
r128 23 25 8.39637 $w=3.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.26 $Y=2.045
+ $X2=0.26 $Y2=2.3
r129 22 41 2.73602 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=1.875
+ $X2=0.26 $Y2=1.96
r130 21 38 0.329269 $w=3.48e-07 $l=1e-08 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=1.62
r131 21 22 8.0671 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=1.875
r132 16 56 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=1.202
r133 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.98 $Y=0.995
+ $X2=3.98 $Y2=0.56
r134 13 55 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.202
r135 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r136 10 54 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.202
r137 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.435 $Y=1.41
+ $X2=3.435 $Y2=1.985
r138 7 52 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.202
r139 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.965 $Y=1.41
+ $X2=2.965 $Y2=1.985
r140 2 41 600 $w=1.7e-07 $l=5.72495e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=1.96
r141 2 38 600 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=1.62
r142 2 25 600 $w=1.7e-07 $l=9.16215e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.35 $Y2=2.3
r143 1 34 91 $w=1.7e-07 $l=2.35053e-07 $layer=licon1_NDIFF $count=2 $X=0.21
+ $Y=0.235 $X2=0.38 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A2 1 3 4 6 7 9 10 12 13 20 23
c54 20 0 1.21795e-19 $X=4.945 $Y=1.202
c55 1 0 8.46699e-20 $X=4.45 $Y=0.995
r56 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.945 $Y=1.202
+ $X2=4.97 $Y2=1.202
r57 19 23 18.8545 $w=1.98e-07 $l=3.4e-07 $layer=LI1_cond $X=4.71 $Y=1.175
+ $X2=4.37 $Y2=1.175
r58 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.71 $Y=1.202
+ $X2=4.945 $Y2=1.202
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.71
+ $Y=1.16 $X2=4.71 $Y2=1.16
r60 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.475 $Y=1.202
+ $X2=4.71 $Y2=1.202
r61 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.45 $Y=1.202
+ $X2=4.475 $Y2=1.202
r62 13 19 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=4.82 $Y=1.175 $X2=4.71
+ $Y2=1.175
r63 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.97 $Y=0.995
+ $X2=4.97 $Y2=1.202
r64 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.97 $Y=0.995
+ $X2=4.97 $Y2=0.56
r65 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.945 $Y=1.41
+ $X2=4.945 $Y2=1.202
r66 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.945 $Y=1.41
+ $X2=4.945 $Y2=1.985
r67 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.202
r68 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.475 $Y=1.41
+ $X2=4.475 $Y2=1.985
r69 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.45 $Y=0.995
+ $X2=4.45 $Y2=1.202
r70 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.45 $Y=0.995 $X2=4.45
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A1 1 3 4 6 7 9 10 12 13 20 25
c38 13 0 1.21795e-19 $X=5.755 $Y=1.105
r39 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.885 $Y=1.202
+ $X2=5.91 $Y2=1.202
r40 19 25 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=5.705 $Y=1.175
+ $X2=5.825 $Y2=1.175
r41 18 20 22.8316 $w=3.8e-07 $l=1.8e-07 $layer=POLY_cond $X=5.705 $Y=1.202
+ $X2=5.885 $Y2=1.202
r42 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.705
+ $Y=1.16 $X2=5.705 $Y2=1.16
r43 16 18 36.7842 $w=3.8e-07 $l=2.9e-07 $layer=POLY_cond $X=5.415 $Y=1.202
+ $X2=5.705 $Y2=1.202
r44 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.39 $Y=1.202
+ $X2=5.415 $Y2=1.202
r45 13 25 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=5.84 $Y=1.175
+ $X2=5.825 $Y2=1.175
r46 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.91 $Y=0.995
+ $X2=5.91 $Y2=1.202
r47 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.91 $Y=0.995
+ $X2=5.91 $Y2=0.56
r48 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.885 $Y=1.41
+ $X2=5.885 $Y2=1.202
r49 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.885 $Y=1.41
+ $X2=5.885 $Y2=1.985
r50 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.415 $Y=1.41
+ $X2=5.415 $Y2=1.202
r51 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.415 $Y=1.41
+ $X2=5.415 $Y2=1.985
r52 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.39 $Y=0.995
+ $X2=5.39 $Y2=1.202
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.39 $Y=0.995 $X2=5.39
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%VPWR 1 2 3 4 5 20 22 26 28 32 36 40 43 44
+ 46 47 48 61 62 65 68 71
r108 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r109 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r111 66 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r112 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r114 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r115 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r116 56 59 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r117 55 58 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r118 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 53 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r120 53 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r121 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r122 50 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.895 $Y=2.72
+ $X2=2.705 $Y2=2.72
r123 50 52 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.895 $Y=2.72
+ $X2=3.45 $Y2=2.72
r124 48 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r125 46 58 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=5.435 $Y=2.72
+ $X2=5.29 $Y2=2.72
r126 46 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.435 $Y=2.72
+ $X2=5.625 $Y2=2.72
r127 45 61 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=6.21 $Y2=2.72
r128 45 47 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=5.625 $Y2=2.72
r129 43 52 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.55 $Y=2.72 $X2=3.45
+ $Y2=2.72
r130 43 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.55 $Y=2.72
+ $X2=3.675 $Y2=2.72
r131 42 55 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.8 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 42 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.8 $Y=2.72
+ $X2=3.675 $Y2=2.72
r133 38 47 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.625 $Y=2.635
+ $X2=5.625 $Y2=2.72
r134 38 40 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=5.625 $Y=2.635
+ $X2=5.625 $Y2=2
r135 34 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=2.635
+ $X2=3.675 $Y2=2.72
r136 34 36 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.675 $Y=2.635
+ $X2=3.675 $Y2=2.3
r137 30 71 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.705 $Y=2.635
+ $X2=2.705 $Y2=2.72
r138 30 32 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.705 $Y=2.635
+ $X2=2.705 $Y2=2.3
r139 29 68 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.955 $Y=2.72
+ $X2=1.765 $Y2=2.72
r140 28 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=2.705 $Y2=2.72
r141 28 29 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=1.955 $Y2=2.72
r142 24 68 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.765 $Y=2.635
+ $X2=1.765 $Y2=2.72
r143 24 26 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.765 $Y=2.635
+ $X2=1.765 $Y2=2.3
r144 23 65 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.015 $Y=2.72
+ $X2=0.825 $Y2=2.72
r145 22 68 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.575 $Y=2.72
+ $X2=1.765 $Y2=2.72
r146 22 23 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.575 $Y=2.72
+ $X2=1.015 $Y2=2.72
r147 18 65 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.825 $Y=2.635
+ $X2=0.825 $Y2=2.72
r148 18 20 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.825 $Y=2.635
+ $X2=0.825 $Y2=2.3
r149 5 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.505
+ $Y=1.485 $X2=5.65 $Y2=2
r150 4 36 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.525
+ $Y=1.485 $X2=3.67 $Y2=2.3
r151 3 32 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.485 $X2=2.73 $Y2=2.3
r152 2 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.645
+ $Y=1.485 $X2=1.79 $Y2=2.3
r153 1 20 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.705
+ $Y=1.485 $X2=0.85 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%X 1 2 3 4 15 18 19 23 25 29 32
c57 25 0 1.74983e-19 $X=1.43 $Y=0.817
c58 23 0 1.54638e-19 $X=2.26 $Y=1.62
r59 29 32 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=2.21 $Y=0.51 $X2=2.21
+ $Y2=0.39
r60 28 29 7.50834 $w=3.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.21 $Y=0.725
+ $X2=2.21 $Y2=0.51
r61 21 27 5.44553 $w=2.6e-07 $l=2.75e-07 $layer=LI1_cond $X=1.705 $Y=1.575
+ $X2=1.43 $Y2=1.575
r62 21 23 24.6002 $w=2.58e-07 $l=5.55e-07 $layer=LI1_cond $X=1.705 $Y=1.575
+ $X2=2.26 $Y2=1.575
r63 20 25 4.58449 $w=1.85e-07 $l=2.75e-07 $layer=LI1_cond $X=1.705 $Y=0.817
+ $X2=1.43 $Y2=0.817
r64 19 28 7.54394 $w=1.85e-07 $l=2.05925e-07 $layer=LI1_cond $X=2.045 $Y=0.817
+ $X2=2.21 $Y2=0.725
r65 19 20 20.3833 $w=1.83e-07 $l=3.4e-07 $layer=LI1_cond $X=2.045 $Y=0.817
+ $X2=1.705 $Y2=0.817
r66 18 27 2.57425 $w=5.5e-07 $l=1.3e-07 $layer=LI1_cond $X=1.43 $Y=1.445
+ $X2=1.43 $Y2=1.575
r67 17 25 2.39439 $w=4.4e-07 $l=9.3e-08 $layer=LI1_cond $X=1.43 $Y=0.91 $X2=1.43
+ $Y2=0.817
r68 17 18 11.6346 $w=5.48e-07 $l=5.35e-07 $layer=LI1_cond $X=1.43 $Y=0.91
+ $X2=1.43 $Y2=1.445
r69 13 25 2.39439 $w=4.4e-07 $l=1.49064e-07 $layer=LI1_cond $X=1.32 $Y=0.725
+ $X2=1.43 $Y2=0.817
r70 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.32 $Y=0.725
+ $X2=1.32 $Y2=0.39
r71 4 23 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.115
+ $Y=1.485 $X2=2.26 $Y2=1.62
r72 3 27 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.175
+ $Y=1.485 $X2=1.32 $Y2=1.62
r73 2 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.075
+ $Y=0.235 $X2=2.21 $Y2=0.39
r74 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.135
+ $Y=0.235 $X2=1.32 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A_823_297# 1 2 3 10 12 13 14 16 18 21
r39 16 29 3.02719 $w=2.75e-07 $l=1.05e-07 $layer=LI1_cond $X=6.172 $Y=1.665
+ $X2=6.172 $Y2=1.56
r40 16 18 26.611 $w=2.73e-07 $l=6.35e-07 $layer=LI1_cond $X=6.172 $Y=1.665
+ $X2=6.172 $Y2=2.3
r41 15 25 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.265 $Y=1.56
+ $X2=5.18 $Y2=1.56
r42 14 29 3.94976 $w=2.1e-07 $l=1.37e-07 $layer=LI1_cond $X=6.035 $Y=1.56
+ $X2=6.172 $Y2=1.56
r43 14 15 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=6.035 $Y=1.56
+ $X2=5.265 $Y2=1.56
r44 13 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.18 $Y=2.295
+ $X2=5.18 $Y2=2.38
r45 12 25 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.18 $Y=1.665
+ $X2=5.18 $Y2=1.56
r46 12 13 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=5.18 $Y=1.665
+ $X2=5.18 $Y2=2.295
r47 11 21 3.86198 $w=1.7e-07 $l=1.80624e-07 $layer=LI1_cond $X=4.325 $Y=2.38
+ $X2=4.18 $Y2=2.3
r48 10 27 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=2.38
+ $X2=5.18 $Y2=2.38
r49 10 11 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.095 $Y=2.38
+ $X2=4.325 $Y2=2.38
r50 3 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.485 $X2=6.12 $Y2=1.62
r51 3 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.975
+ $Y=1.485 $X2=6.12 $Y2=2.3
r52 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=1.485 $X2=5.18 $Y2=2.3
r53 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.035
+ $Y=1.485 $X2=5.18 $Y2=1.62
r54 1 21 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=4.115
+ $Y=1.485 $X2=4.24 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 49 50 51 73 74
r108 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r109 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r110 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r111 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r112 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r113 65 68 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=4.37 $Y2=0
r114 64 67 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.37
+ $Y2=0
r115 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r116 62 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r117 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r118 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r119 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r120 55 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r121 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r122 51 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r123 49 70 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=5.29 $Y2=0
r124 49 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.65
+ $Y2=0
r125 48 73 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=6.21 $Y2=0
r126 48 50 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.65
+ $Y2=0
r127 46 67 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.625 $Y=0
+ $X2=4.37 $Y2=0
r128 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.71
+ $Y2=0
r129 45 70 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=5.29 $Y2=0
r130 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.71
+ $Y2=0
r131 43 61 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.53
+ $Y2=0
r132 43 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.73
+ $Y2=0
r133 42 64 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.99
+ $Y2=0
r134 42 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.73
+ $Y2=0
r135 40 58 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.61
+ $Y2=0
r136 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=0 $X2=1.79
+ $Y2=0
r137 39 61 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.875 $Y=0
+ $X2=2.53 $Y2=0
r138 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.875 $Y=0 $X2=1.79
+ $Y2=0
r139 37 54 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.69
+ $Y2=0
r140 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.765 $Y=0 $X2=0.85
+ $Y2=0
r141 36 58 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=0.935 $Y=0
+ $X2=1.61 $Y2=0
r142 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0 $X2=0.85
+ $Y2=0
r143 32 50 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.65 $Y=0.085
+ $X2=5.65 $Y2=0
r144 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.65 $Y=0.085
+ $X2=5.65 $Y2=0.39
r145 28 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=0.085
+ $X2=4.71 $Y2=0
r146 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.71 $Y=0.085
+ $X2=4.71 $Y2=0.39
r147 24 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.73 $Y=0.085
+ $X2=2.73 $Y2=0
r148 24 26 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.73 $Y=0.085
+ $X2=2.73 $Y2=0.39
r149 20 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0
r150 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.79 $Y=0.085
+ $X2=1.79 $Y2=0.39
r151 16 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.85 $Y=0.085
+ $X2=0.85 $Y2=0
r152 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.85 $Y=0.085
+ $X2=0.85 $Y2=0.39
r153 5 34 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.235 $X2=5.65 $Y2=0.39
r154 4 30 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.525
+ $Y=0.235 $X2=4.71 $Y2=0.39
r155 3 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.595
+ $Y=0.235 $X2=2.73 $Y2=0.39
r156 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.605
+ $Y=0.235 $X2=1.79 $Y2=0.39
r157 1 18 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=0.715
+ $Y=0.235 $X2=0.85 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_4%A_635_47# 1 2 3 4 13 17 18 19 23 25 29 35
r67 27 29 9.53255 $w=4.03e-07 $l=3.35e-07 $layer=LI1_cond $X=6.107 $Y=0.725
+ $X2=6.107 $Y2=0.39
r68 26 35 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.345 $Y=0.815
+ $X2=5.155 $Y2=0.815
r69 25 27 8.21845 $w=1.8e-07 $l=2.42866e-07 $layer=LI1_cond $X=5.905 $Y=0.815
+ $X2=6.107 $Y2=0.725
r70 25 26 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.905 $Y=0.815
+ $X2=5.345 $Y2=0.815
r71 21 35 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.155 $Y=0.725
+ $X2=5.155 $Y2=0.815
r72 21 23 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.155 $Y=0.725
+ $X2=5.155 $Y2=0.39
r73 20 34 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.405 $Y=0.815
+ $X2=4.28 $Y2=0.815
r74 19 35 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.965 $Y=0.815
+ $X2=5.155 $Y2=0.815
r75 19 20 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.965 $Y=0.815
+ $X2=4.405 $Y2=0.815
r76 18 34 2.95288 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=4.28 $Y=0.725 $X2=4.28
+ $Y2=0.815
r77 17 32 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=4.28 $Y=0.475
+ $X2=4.28 $Y2=0.365
r78 17 18 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.28 $Y=0.475
+ $X2=4.28 $Y2=0.725
r79 13 32 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=4.155 $Y=0.365
+ $X2=4.28 $Y2=0.365
r80 13 15 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=4.155 $Y=0.365
+ $X2=3.3 $Y2=0.365
r81 4 29 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.985
+ $Y=0.235 $X2=6.12 $Y2=0.39
r82 3 23 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.045
+ $Y=0.235 $X2=5.18 $Y2=0.39
r83 2 34 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.24 $Y2=0.73
r84 2 32 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.055
+ $Y=0.235 $X2=4.24 $Y2=0.39
r85 1 15 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.175
+ $Y=0.235 $X2=3.3 $Y2=0.39
.ends

