# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21o_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.340000 1.010000 4.965000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.010000 4.170000 1.275000 ;
        RECT 3.945000 1.275000 4.170000 1.510000 ;
        RECT 3.945000 1.510000 5.435000 1.680000 ;
        RECT 5.135000 1.055000 5.600000 1.290000 ;
        RECT 5.135000 1.290000 5.435000 1.510000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.500000 0.995000 2.905000 1.525000 ;
    END
  END B1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.615000 1.885000 0.785000 ;
        RECT 0.145000 0.785000 0.680000 1.585000 ;
        RECT 0.145000 1.585000 1.885000 1.755000 ;
        RECT 0.675000 1.755000 0.845000 2.185000 ;
        RECT 1.635000 1.755000 1.885000 2.185000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.105000  0.085000 0.445000 0.445000 ;
      RECT 0.115000  1.935000 0.445000 2.635000 ;
      RECT 0.850000  0.995000 2.300000 1.325000 ;
      RECT 1.025000  0.085000 1.405000 0.445000 ;
      RECT 1.025000  1.935000 1.405000 2.635000 ;
      RECT 2.065000  1.515000 2.315000 2.635000 ;
      RECT 2.110000  0.085000 2.885000 0.445000 ;
      RECT 2.130000  0.615000 3.295000 0.670000 ;
      RECT 2.130000  0.670000 4.765000 0.785000 ;
      RECT 2.130000  0.785000 2.300000 0.995000 ;
      RECT 2.655000  1.695000 2.825000 2.295000 ;
      RECT 2.655000  2.295000 3.765000 2.465000 ;
      RECT 3.125000  0.255000 3.295000 0.615000 ;
      RECT 3.125000  0.785000 4.765000 0.840000 ;
      RECT 3.125000  0.840000 3.295000 2.125000 ;
      RECT 3.555000  0.085000 3.885000 0.445000 ;
      RECT 3.585000  1.445000 3.765000 1.850000 ;
      RECT 3.585000  1.850000 5.860000 2.020000 ;
      RECT 3.585000  2.020000 3.765000 2.295000 ;
      RECT 3.935000  2.275000 4.315000 2.635000 ;
      RECT 4.485000  0.405000 4.765000 0.670000 ;
      RECT 4.535000  2.020000 4.705000 2.465000 ;
      RECT 4.875000  2.275000 5.255000 2.635000 ;
      RECT 5.445000  0.085000 5.725000 0.885000 ;
      RECT 5.530000  2.020000 5.860000 2.395000 ;
      RECT 5.605000  1.460000 5.860000 1.850000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_4
END LIBRARY
