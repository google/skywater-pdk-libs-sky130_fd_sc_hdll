* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_16 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_27_47# A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_117_297# a_973_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_597_297# A0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_27_47# A1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_973_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_119_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_973_297# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_27_47# A0 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_117_297# A1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_597_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_119_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_27_47# A1 a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_1163_47# a_973_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# A0 a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR a_973_297# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_27_47# A0 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_117_297# a_973_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_27_47# A0 a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 a_119_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 VPWR S a_973_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 a_27_47# A1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 VGND a_973_297# a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 a_1163_47# a_973_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 a_597_297# A0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X45 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 VGND S a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X48 a_1163_47# A0 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 a_119_47# A1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 VPWR S a_597_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 VGND a_973_297# a_1163_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X52 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X53 a_117_297# A1 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 VGND S a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X55 a_1163_47# A0 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X59 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X60 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X61 VPWR a_973_297# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X62 VGND S a_973_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X63 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X64 a_597_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X67 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
