* NGSPICE file created from sky130_fd_sc_hdll__o22ai_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
M1000 Y A2 a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u
M1001 VPWR B1 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=5.16e+06u as=8.7e+11p ps=7.74e+06u
M1002 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.2415e+12p pd=1.032e+07u as=4.81e+11p ps=4.08e+06u
M1003 a_27_297# B2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 Y B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=4.81e+11p pd=4.08e+06u as=0p ps=0u
M1007 a_27_47# B2 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_515_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND A2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR A1 a_515_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_27_297# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 Y B2 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_27_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_515_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

