* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__mux2_8 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_870_297# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_1420_297# a_1369_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VPWR S a_1369_199# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND S a_872_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X6 VGND a_1369_199# a_1422_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X7 a_79_21# A0 a_1422_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR S a_870_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_872_47# A1 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X13 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_1422_47# a_1369_199# VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X16 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_79_21# A0 a_870_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_79_21# A1 a_1420_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_870_297# A0 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_1420_297# A1 a_79_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VPWR a_79_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_79_21# A1 a_872_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X26 a_872_47# S VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X27 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VGND a_79_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND S a_1369_199# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_1422_47# A0 a_79_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 VPWR a_1369_199# a_1420_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 X a_79_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 X a_79_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
