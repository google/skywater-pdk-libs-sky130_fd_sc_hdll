# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o21ba_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.350000 1.075000 3.895000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.645000 1.075000 3.180000 1.285000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.825000 1.325000 ;
        RECT 0.605000 1.325000 0.825000 1.695000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.571700 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.995000 0.295000 1.380000 0.465000 ;
        RECT 0.995000 0.465000 1.235000 1.495000 ;
        RECT 0.995000 1.495000 1.455000 1.695000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.085000  0.430000 0.345000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.495000 ;
      RECT 0.085000  1.495000 0.395000 1.865000 ;
      RECT 0.085000  1.865000 2.085000 2.035000 ;
      RECT 0.520000  2.205000 0.960000 2.635000 ;
      RECT 0.645000  0.085000 0.825000 0.825000 ;
      RECT 1.405000  0.655000 2.470000 0.825000 ;
      RECT 1.405000  0.825000 1.575000 1.325000 ;
      RECT 1.520000  2.205000 2.380000 2.635000 ;
      RECT 1.560000  0.085000 1.925000 0.465000 ;
      RECT 1.915000  0.995000 2.085000 1.865000 ;
      RECT 2.140000  0.255000 2.470000 0.655000 ;
      RECT 2.255000  0.825000 2.470000 1.455000 ;
      RECT 2.255000  1.455000 2.925000 2.035000 ;
      RECT 2.600000  2.035000 2.925000 2.465000 ;
      RECT 2.695000  0.365000 2.945000 0.735000 ;
      RECT 2.695000  0.735000 3.890000 0.905000 ;
      RECT 3.165000  0.085000 3.335000 0.555000 ;
      RECT 3.450000  1.875000 3.830000 2.635000 ;
      RECT 3.555000  0.270000 3.890000 0.735000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_2
END LIBRARY
