* File: sky130_fd_sc_hdll__and2_1.pex.spice
* Created: Wed Sep  2 08:21:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2_1%A 2 3 5 8 10 12 19 22 28
r33 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.16
+ $X2=0.54 $Y2=1.16
r34 16 28 10.833 $w=2.48e-07 $l=2.35e-07 $layer=LI1_cond $X=0.295 $Y=1.2
+ $X2=0.53 $Y2=1.2
r35 15 18 38.4695 $w=3.3e-07 $l=2.2e-07 $layer=POLY_cond $X=0.295 $Y=1.16
+ $X2=0.515 $Y2=1.16
r36 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.295
+ $Y=1.16 $X2=0.295 $Y2=1.16
r37 12 28 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=0.555 $Y=1.2
+ $X2=0.53 $Y2=1.2
r38 10 16 0.829759 $w=2.48e-07 $l=1.8e-08 $layer=LI1_cond $X=0.277 $Y=1.2
+ $X2=0.295 $Y2=1.2
r39 10 22 2.16659 $w=2.48e-07 $l=4.7e-08 $layer=LI1_cond $X=0.277 $Y=1.2
+ $X2=0.23 $Y2=1.2
r40 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.16
r41 6 8 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.585
r42 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.515 $Y=1.78
+ $X2=0.515 $Y2=2.065
r43 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.515 $Y=1.68 $X2=0.515
+ $Y2=1.78
r44 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.515 $Y=1.325
+ $X2=0.515 $Y2=1.16
r45 1 2 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.515 $Y=1.325 $X2=0.515
+ $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_1%B 3 6 7 9 10 13
r41 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.16
+ $X2=1.045 $Y2=1.325
r42 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.045 $Y=1.16
+ $X2=1.045 $Y2=0.995
r43 10 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.05
+ $Y=1.16 $X2=1.05 $Y2=1.16
r44 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.985 $Y=1.78
+ $X2=0.985 $Y2=2.065
r45 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.78
r46 6 16 117.71 $w=2e-07 $l=3.55e-07 $layer=POLY_cond $X=0.985 $Y=1.68 $X2=0.985
+ $Y2=1.325
r47 3 15 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=0.96 $Y=0.585
+ $X2=0.96 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_1%A_27_75# 1 2 7 9 10 12 15 17 18 21 23 24 25
+ 26
r74 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.575
+ $Y=1.16 $X2=1.575 $Y2=1.16
r75 27 29 19.8605 $w=2.15e-07 $l=3.5e-07 $layer=LI1_cond $X=1.532 $Y=0.81
+ $X2=1.532 $Y2=1.16
r76 25 29 9.93147 $w=2.15e-07 $l=1.84811e-07 $layer=LI1_cond $X=1.49 $Y=1.325
+ $X2=1.532 $Y2=1.16
r77 25 26 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.49 $Y=1.325
+ $X2=1.49 $Y2=1.575
r78 23 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.405 $Y=1.66
+ $X2=1.49 $Y2=1.575
r79 23 24 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=1.405 $Y=1.66
+ $X2=0.925 $Y2=1.66
r80 19 24 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.775 $Y=1.745
+ $X2=0.925 $Y2=1.66
r81 19 21 14.7897 $w=2.98e-07 $l=3.85e-07 $layer=LI1_cond $X=0.775 $Y=1.745
+ $X2=0.775 $Y2=2.13
r82 17 27 1.45963 $w=1.9e-07 $l=1.27e-07 $layer=LI1_cond $X=1.405 $Y=0.81
+ $X2=1.532 $Y2=0.81
r83 17 18 55.4545 $w=1.88e-07 $l=9.5e-07 $layer=LI1_cond $X=1.405 $Y=0.81
+ $X2=0.455 $Y2=0.81
r84 13 18 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.455 $Y2=0.81
r85 13 15 6.80989 $w=3.28e-07 $l=1.95e-07 $layer=LI1_cond $X=0.29 $Y=0.715
+ $X2=0.29 $Y2=0.52
r86 10 30 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.54 $Y=1.41
+ $X2=1.575 $Y2=1.16
r87 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.54 $Y=1.41
+ $X2=1.54 $Y2=1.985
r88 7 30 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.515 $Y=0.995
+ $X2=1.575 $Y2=1.16
r89 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.515 $Y=0.995
+ $X2=1.515 $Y2=0.56
r90 2 21 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.855 $X2=0.75 $Y2=2.13
r91 1 15 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.375 $X2=0.28 $Y2=0.52
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_1%VPWR 1 2 7 9 11 15 17 21 22 28
r28 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 22 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r31 19 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=1.26 $Y2=2.72
r32 19 21 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=2.07 $Y2=2.72
r33 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r34 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r35 13 28 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=2.635
+ $X2=1.26 $Y2=2.72
r36 13 15 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=1.26 $Y=2.635
+ $X2=1.26 $Y2=2
r37 12 25 4.25667 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r38 11 28 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=1.26 $Y2=2.72
r39 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.405 $Y2=2.72
r40 7 25 3.10338 $w=2.8e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.202 $Y2=2.72
r41 7 9 20.7851 $w=2.78e-07 $l=5.05e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=2.13
r42 2 15 300 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=2 $X=1.075
+ $Y=1.855 $X2=1.26 $Y2=2
r43 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.855 $X2=0.28 $Y2=2.13
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_1%X 1 2 7 10 11 12 13 14 15 24 35
r22 35 40 1.75796 $w=2.93e-07 $l=4.5e-08 $layer=LI1_cond $X=2.007 $Y=1.87
+ $X2=2.007 $Y2=1.915
r23 15 42 5.69442 $w=4.23e-07 $l=2.1e-07 $layer=LI1_cond $X=1.942 $Y=2.21
+ $X2=1.942 $Y2=2
r24 14 42 1.76256 $w=4.23e-07 $l=6.5e-08 $layer=LI1_cond $X=1.942 $Y=1.935
+ $X2=1.942 $Y2=2
r25 14 40 1.63189 $w=4.23e-07 $l=2e-08 $layer=LI1_cond $X=1.942 $Y=1.935
+ $X2=1.942 $Y2=1.915
r26 14 35 0.781317 $w=2.93e-07 $l=2e-08 $layer=LI1_cond $X=2.007 $Y=1.85
+ $X2=2.007 $Y2=1.87
r27 13 14 12.5011 $w=2.93e-07 $l=3.2e-07 $layer=LI1_cond $X=2.007 $Y=1.53
+ $X2=2.007 $Y2=1.85
r28 12 13 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.007 $Y=1.19
+ $X2=2.007 $Y2=1.53
r29 11 12 13.2824 $w=2.93e-07 $l=3.4e-07 $layer=LI1_cond $X=2.007 $Y=0.85
+ $X2=2.007 $Y2=1.19
r30 10 24 3.38522 $w=2.95e-07 $l=1.45e-07 $layer=LI1_cond $X=2.007 $Y=0.4
+ $X2=2.007 $Y2=0.545
r31 10 11 10.9384 $w=2.93e-07 $l=2.8e-07 $layer=LI1_cond $X=2.007 $Y=0.57
+ $X2=2.007 $Y2=0.85
r32 10 24 0.976647 $w=2.93e-07 $l=2.5e-08 $layer=LI1_cond $X=2.007 $Y=0.57
+ $X2=2.007 $Y2=0.545
r33 7 10 3.43192 $w=2.9e-07 $l=1.47e-07 $layer=LI1_cond $X=1.86 $Y=0.4 $X2=2.007
+ $Y2=0.4
r34 7 9 2.10345 $w=2.9e-07 $l=5e-08 $layer=LI1_cond $X=1.86 $Y=0.4 $X2=1.81
+ $Y2=0.4
r35 2 42 300 $w=1.7e-07 $l=6.39863e-07 $layer=licon1_PDIFF $count=2 $X=1.63
+ $Y=1.485 $X2=1.91 $Y2=2
r36 1 9 182 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.235 $X2=1.81 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_1%VGND 1 6 8 10 17 18 21
r29 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r30 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r31 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r32 15 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=1.23
+ $Y2=0
r33 15 17 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.355 $Y=0 $X2=2.07
+ $Y2=0
r34 10 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=1.23
+ $Y2=0
r35 10 12 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=1.105 $Y=0 $X2=0.23
+ $Y2=0
r36 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r37 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r38 4 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0
r39 4 6 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.085
+ $X2=1.23 $Y2=0.38
r40 1 6 182 $w=1.7e-07 $l=2.37487e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.375 $X2=1.27 $Y2=0.38
.ends

