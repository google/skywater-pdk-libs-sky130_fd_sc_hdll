* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand2b_1 A_N B VGND VNB VPB VPWR Y
M1000 VPWR A_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=5.757e+11p pd=5.25e+06u as=1.134e+11p ps=1.38e+06u
M1001 VPWR a_27_93# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 VGND A_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=2.33e+11p pd=2.07e+06u as=1.302e+11p ps=1.46e+06u
M1003 Y B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 Y a_27_93# a_226_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=1.755e+11p ps=1.84e+06u
M1005 a_226_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
