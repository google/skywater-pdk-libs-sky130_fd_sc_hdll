* NGSPICE file created from sky130_fd_sc_hdll__nand4bb_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__nand4bb_2 A_N B_N C D VGND VNB VPB VPWR Y
M1000 a_211_413# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.974e+11p pd=1.78e+06u as=3.424e+11p ps=3.42e+06u
M1001 Y C VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=2.0218e+12p ps=1.522e+07u
M1002 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_361_47# a_211_413# Y VNB nshort w=650000u l=150000u
+  ad=5.785e+11p pd=5.68e+06u as=2.08e+11p ps=1.94e+06u
M1004 Y a_211_413# a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR D Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_841_47# D VGND VNB nshort w=650000u l=150000u
+  ad=5.59e+11p pd=5.62e+06u as=0p ps=0u
M1007 Y a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND D a_841_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_211_413# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_841_47# C a_641_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1012 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1013 a_211_413# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=2.016e+11p pd=1.8e+06u as=0p ps=0u
M1014 Y a_211_413# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 a_361_47# a_27_47# a_641_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_27_47# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_641_47# a_27_47# a_361_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_641_47# C a_841_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

