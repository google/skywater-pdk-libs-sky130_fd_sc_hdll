* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or3b_1 A B C_N VGND VNB VPB VPWR X
M1000 a_225_53# B VGND VNB nshort w=420000u l=150000u
+  ad=2.835e+11p pd=3.03e+06u as=4.787e+11p ps=4.92e+06u
M1001 VGND A a_225_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 VGND a_117_297# a_225_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_117_297# C_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=4.241e+11p ps=4.1e+06u
M1004 VPWR A a_399_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.407e+11p ps=1.51e+06u
M1005 a_399_297# B a_315_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.008e+11p ps=1.32e+06u
M1006 a_117_297# C_N VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1007 a_315_297# a_117_297# a_225_53# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1008 X a_225_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.85e+11p pd=2.57e+06u as=0p ps=0u
M1009 X a_225_53# VGND VNB nshort w=650000u l=150000u
+  ad=1.7875e+11p pd=1.85e+06u as=0p ps=0u
.ends
