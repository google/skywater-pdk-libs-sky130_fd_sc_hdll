* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfxbp_2 CLK D SCD SCE VGND VNB VPB VPWR Q Q_N
X0 a_1117_47# a_1179_183# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 VPWR a_1653_315# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VPWR a_1001_47# a_1179_183# VPB sky130_fd_pr__pfet_01v8_hvt w=750000u l=180000u
X3 a_1653_315# a_1464_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1111_413# a_1179_183# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 a_1558_413# a_1653_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 Q a_1653_315# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND a_1001_47# a_1179_183# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X8 a_1615_47# a_1653_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X10 a_698_369# SCD VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X11 a_604_369# a_211_363# a_1001_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X12 VGND a_2234_47# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_1001_47# a_27_47# a_1111_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X14 a_319_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VGND a_319_47# a_529_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_1653_315# a_1464_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 a_1464_413# a_211_363# a_1558_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X19 a_2234_47# a_1653_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_1179_183# a_27_47# a_1464_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X21 a_604_369# SCE a_717_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X22 a_604_369# a_27_47# a_1001_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 a_1179_183# a_211_363# a_1464_413# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X24 Q a_1653_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 VPWR SCE a_503_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X26 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_529_47# D a_604_369# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 Q_N a_2234_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X30 a_717_47# SCD VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_1464_413# a_27_47# a_1615_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X32 a_604_369# a_319_47# a_698_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X33 a_1001_47# a_211_363# a_1117_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X34 a_2234_47# a_1653_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X35 a_503_369# D a_604_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X36 Q_N a_2234_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_319_47# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X38 VPWR a_2234_47# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VGND a_1653_315# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
