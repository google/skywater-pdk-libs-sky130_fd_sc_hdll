* File: sky130_fd_sc_hdll__o32ai_2.pex.spice
* Created: Wed Sep  2 08:47:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%B2 1 3 4 6 7 9 10 12 13 14 22 29
c38 29 0 1.58116e-19 $X=0.695 $Y=1.19
r39 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r40 20 22 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.73 $Y=1.202
+ $X2=0.965 $Y2=1.202
r41 20 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.73
+ $Y=1.16 $X2=0.73 $Y2=1.16
r42 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.73 $Y2=1.202
r43 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r44 14 29 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.2 $X2=0.695
+ $Y2=1.2
r45 13 14 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=0.235 $Y=1.2
+ $X2=0.69 $Y2=1.2
r46 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r47 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r48 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r49 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r50 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r51 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r52 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r53 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%B1 1 3 4 6 7 9 10 12 13 14 22 25
c52 22 0 1.58116e-19 $X=1.905 $Y=1.202
c53 14 0 9.67856e-20 $X=1.615 $Y=1.19
r54 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r55 20 22 42.4921 $w=3.8e-07 $l=3.35e-07 $layer=POLY_cond $X=1.57 $Y=1.202
+ $X2=1.905 $Y2=1.202
r56 18 20 17.1237 $w=3.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.57 $Y2=1.202
r57 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r58 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.16 $X2=1.57 $Y2=1.16
r59 13 14 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=1.17 $Y=1.2 $X2=1.57
+ $Y2=1.2
r60 13 25 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=1.17 $Y=1.2
+ $X2=1.155 $Y2=1.2
r61 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r62 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r63 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r64 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r65 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r66 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r67 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r68 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995 $X2=1.41
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A3 3 5 6 7 9 10 12 13 15 16 21 22 25
c57 6 0 1.02109e-19 $X=2.425 $Y=1.19
c58 3 0 9.67856e-20 $X=2.35 $Y=0.56
r59 22 23 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=3.44 $Y=1.202
+ $X2=3.475 $Y2=1.202
r60 20 22 30.4421 $w=3.8e-07 $l=2.4e-07 $layer=POLY_cond $X=3.2 $Y=1.202
+ $X2=3.44 $Y2=1.202
r61 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.2
+ $Y=1.16 $X2=3.2 $Y2=1.16
r62 18 20 24.7342 $w=3.8e-07 $l=1.95e-07 $layer=POLY_cond $X=3.005 $Y=1.202
+ $X2=3.2 $Y2=1.202
r63 16 21 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=3.005 $Y=1.2
+ $X2=3.2 $Y2=1.2
r64 16 25 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=3.005 $Y=1.2
+ $X2=2.985 $Y2=1.2
r65 13 23 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.475 $Y=1.41
+ $X2=3.475 $Y2=1.202
r66 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.475 $Y=1.41
+ $X2=3.475 $Y2=1.985
r67 10 22 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=1.202
r68 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.44 $Y=0.995
+ $X2=3.44 $Y2=0.56
r69 7 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.202
r70 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.985
r71 5 18 30.9734 $w=3.8e-07 $l=1.0583e-07 $layer=POLY_cond $X=2.905 $Y=1.19
+ $X2=3.005 $Y2=1.202
r72 5 6 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=2.905 $Y=1.19
+ $X2=2.425 $Y2=1.19
r73 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.35 $Y=1.115
+ $X2=2.425 $Y2=1.19
r74 1 3 284.585 $w=1.5e-07 $l=5.55e-07 $layer=POLY_cond $X=2.35 $Y=1.115
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A2 1 3 4 6 7 9 10 12 13 14 22 30
r46 22 23 4.4867 $w=3.76e-07 $l=3.5e-08 $layer=POLY_cond $X=4.38 $Y=1.202
+ $X2=4.415 $Y2=1.202
r47 20 22 30.766 $w=3.76e-07 $l=2.4e-07 $layer=POLY_cond $X=4.14 $Y=1.202
+ $X2=4.38 $Y2=1.202
r48 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.14
+ $Y=1.16 $X2=4.14 $Y2=1.16
r49 18 20 24.9973 $w=3.76e-07 $l=1.95e-07 $layer=POLY_cond $X=3.945 $Y=1.202
+ $X2=4.14 $Y2=1.202
r50 17 18 10.8963 $w=3.76e-07 $l=8.5e-08 $layer=POLY_cond $X=3.86 $Y=1.202
+ $X2=3.945 $Y2=1.202
r51 14 30 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=4.37 $Y=1.2 $X2=4.375
+ $Y2=1.2
r52 14 21 10.6025 $w=2.48e-07 $l=2.3e-07 $layer=LI1_cond $X=4.37 $Y=1.2 $X2=4.14
+ $Y2=1.2
r53 13 21 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.915 $Y=1.2
+ $X2=4.14 $Y2=1.2
r54 10 23 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.415 $Y=1.41
+ $X2=4.415 $Y2=1.202
r55 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.415 $Y=1.41
+ $X2=4.415 $Y2=1.985
r56 7 22 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=1.202
r57 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.38 $Y=0.995 $X2=4.38
+ $Y2=0.56
r58 4 18 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.945 $Y=1.41
+ $X2=3.945 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.945 $Y=1.41
+ $X2=3.945 $Y2=1.985
r60 1 17 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995 $X2=3.86
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A1 1 3 4 6 7 9 10 12 13 14 15 24 29 33
r39 24 25 13.496 $w=3.75e-07 $l=1.05e-07 $layer=POLY_cond $X=5.79 $Y=1.202
+ $X2=5.895 $Y2=1.202
r40 23 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.59 $Y=1.2
+ $X2=5.295 $Y2=1.2
r41 22 24 25.7067 $w=3.75e-07 $l=2e-07 $layer=POLY_cond $X=5.59 $Y=1.202
+ $X2=5.79 $Y2=1.202
r42 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.59
+ $Y=1.16 $X2=5.59 $Y2=1.16
r43 20 22 21.208 $w=3.75e-07 $l=1.65e-07 $layer=POLY_cond $X=5.425 $Y=1.202
+ $X2=5.59 $Y2=1.202
r44 19 20 13.496 $w=3.75e-07 $l=1.05e-07 $layer=POLY_cond $X=5.32 $Y=1.202
+ $X2=5.425 $Y2=1.202
r45 15 33 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=6.21 $Y=1.2
+ $X2=5.755 $Y2=1.2
r46 14 33 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=5.735 $Y=1.2
+ $X2=5.755 $Y2=1.2
r47 14 23 6.68417 $w=2.48e-07 $l=1.45e-07 $layer=LI1_cond $X=5.735 $Y=1.2
+ $X2=5.59 $Y2=1.2
r48 13 29 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=5.285 $Y=1.2
+ $X2=5.295 $Y2=1.2
r49 10 25 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.895 $Y=1.41
+ $X2=5.895 $Y2=1.202
r50 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.895 $Y=1.41
+ $X2=5.895 $Y2=1.985
r51 7 24 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=1.202
r52 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.79 $Y=0.995 $X2=5.79
+ $Y2=0.56
r53 4 20 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.425 $Y=1.41
+ $X2=5.425 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.425 $Y=1.41
+ $X2=5.425 $Y2=1.985
r55 1 19 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995 $X2=5.32
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_297# 1 2 3 10 12 14 16 17 18 27
c45 27 0 1.02109e-19 $X=2.14 $Y=2
c46 3 0 3.98522e-20 $X=1.995 $Y=1.485
r47 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.365 $Y=1.92
+ $X2=1.24 $Y2=1.92
r48 18 27 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.925 $Y=1.92
+ $X2=2.115 $Y2=1.92
r49 18 19 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=1.92
+ $X2=1.365 $Y2=1.92
r50 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.24 $Y=2.005
+ $X2=1.24 $Y2=1.92
r51 16 17 13.3683 $w=2.48e-07 $l=2.9e-07 $layer=LI1_cond $X=1.24 $Y=2.005
+ $X2=1.24 $Y2=2.295
r52 15 23 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=2.38
+ $X2=0.217 $Y2=2.38
r53 14 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.115 $Y=2.38
+ $X2=1.24 $Y2=2.295
r54 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.38
+ $X2=0.345 $Y2=2.38
r55 10 23 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.217 $Y=2.295
+ $X2=0.217 $Y2=2.38
r56 10 12 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.217 $Y=2.295
+ $X2=0.217 $Y2=1.66
r57 3 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r58 2 25 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r59 1 23 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r60 1 12 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%Y 1 2 3 4 13 21 23 28 31 32 33
c78 33 0 1.01631e-19 $X=2.075 $Y=1.53
r79 33 39 1.35792 $w=3.85e-07 $l=8.5e-08 $layer=LI1_cond $X=2.177 $Y=1.58
+ $X2=2.177 $Y2=1.495
r80 33 39 0.74834 $w=3.83e-07 $l=2.5e-08 $layer=LI1_cond $X=2.177 $Y=1.47
+ $X2=2.177 $Y2=1.495
r81 33 38 5.17851 $w=3.83e-07 $l=1.73e-07 $layer=LI1_cond $X=2.177 $Y=1.47
+ $X2=2.177 $Y2=1.297
r82 32 38 3.20289 $w=3.83e-07 $l=1.07e-07 $layer=LI1_cond $X=2.177 $Y=1.19
+ $X2=2.177 $Y2=1.297
r83 29 32 6.44568 $w=4.28e-07 $l=2e-07 $layer=LI1_cond $X=2.115 $Y=0.905
+ $X2=2.115 $Y2=1.105
r84 24 33 9.56655 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=2.37 $Y=1.58
+ $X2=2.177 $Y2=1.58
r85 23 31 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.025 $Y=1.58
+ $X2=3.215 $Y2=1.58
r86 23 24 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=3.025 $Y=1.58
+ $X2=2.37 $Y2=1.58
r87 22 28 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r88 21 33 9.56655 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=1.985 $Y=1.58
+ $X2=2.177 $Y2=1.58
r89 21 22 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.985 $Y=1.58
+ $X2=0.895 $Y2=1.58
r90 15 18 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.73 $Y=0.78
+ $X2=1.67 $Y2=0.78
r91 13 29 6.8199 $w=2.5e-07 $l=1.82071e-07 $layer=LI1_cond $X=1.985 $Y=0.78
+ $X2=2.115 $Y2=0.905
r92 13 18 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=1.985 $Y=0.78
+ $X2=1.67 $Y2=0.78
r93 4 31 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=3.095
+ $Y=1.485 $X2=3.24 $Y2=1.66
r94 3 28 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r95 2 18 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.74
r96 1 15 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%VPWR 1 2 3 12 16 18 20 25 26 27 29 41 46
+ 50
r81 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r82 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r83 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r84 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r85 41 49 3.7175 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=6.242 $Y2=2.72
r86 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=5.75 $Y2=2.72
r87 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r88 39 40 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r89 37 40 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r90 37 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r91 36 39 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r92 36 37 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 34 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=1.67 $Y2=2.72
r94 34 36 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=2.07 $Y2=2.72
r95 29 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=1.67 $Y2=2.72
r96 29 31 88.4011 $w=1.68e-07 $l=1.355e-06 $layer=LI1_cond $X=1.585 $Y=2.72
+ $X2=0.23 $Y2=2.72
r97 27 47 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r98 27 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 25 39 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=5.07 $Y=2.72
+ $X2=4.83 $Y2=2.72
r100 25 26 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.07 $Y=2.72
+ $X2=5.172 $Y2=2.72
r101 24 43 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 24 26 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=5.275 $Y=2.72
+ $X2=5.172 $Y2=2.72
r103 20 23 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=6.155 $Y=1.66
+ $X2=6.155 $Y2=2.34
r104 18 49 3.24574 $w=2.2e-07 $l=1.22327e-07 $layer=LI1_cond $X=6.155 $Y=2.635
+ $X2=6.242 $Y2=2.72
r105 18 23 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=6.155 $Y=2.635
+ $X2=6.155 $Y2=2.34
r106 14 26 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.172 $Y=2.635
+ $X2=5.172 $Y2=2.72
r107 14 16 34.3548 $w=2.03e-07 $l=6.35e-07 $layer=LI1_cond $X=5.172 $Y=2.635
+ $X2=5.172 $Y2=2
r108 10 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r109 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.34
r110 3 23 400 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=1.485 $X2=6.15 $Y2=2.34
r111 3 20 400 $w=1.7e-07 $l=2.43926e-07 $layer=licon1_PDIFF $count=1 $X=5.985
+ $Y=1.485 $X2=6.15 $Y2=1.66
r112 2 16 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=5.065
+ $Y=1.485 $X2=5.19 $Y2=2
r113 1 12 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A_525_297# 1 2 3 10 12 14 18 20 22 24 29
r42 22 31 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=4.71 $Y=2.255
+ $X2=4.71 $Y2=2.35
r43 22 24 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.71 $Y=2.255
+ $X2=4.71 $Y2=2
r44 21 29 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.795 $Y=2.35
+ $X2=3.71 $Y2=2.35
r45 20 31 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=2.35
+ $X2=4.71 $Y2=2.35
r46 20 21 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=4.585 $Y=2.35
+ $X2=3.795 $Y2=2.35
r47 16 29 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.71 $Y=2.255
+ $X2=3.71 $Y2=2.35
r48 16 18 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=3.71 $Y=2.255
+ $X2=3.71 $Y2=1.66
r49 15 27 3.96742 $w=1.9e-07 $l=1.25e-07 $layer=LI1_cond $X=2.835 $Y=2.35
+ $X2=2.71 $Y2=2.35
r50 14 29 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.625 $Y=2.35
+ $X2=3.71 $Y2=2.35
r51 14 15 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=3.625 $Y=2.35
+ $X2=2.835 $Y2=2.35
r52 10 27 3.01524 $w=2.5e-07 $l=9.5e-08 $layer=LI1_cond $X=2.71 $Y=2.255
+ $X2=2.71 $Y2=2.35
r53 10 12 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=2.71 $Y=2.255
+ $X2=2.71 $Y2=2
r54 3 31 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.485 $X2=4.67 $Y2=2.34
r55 3 24 600 $w=1.7e-07 $l=5.91777e-07 $layer=licon1_PDIFF $count=1 $X=4.505
+ $Y=1.485 $X2=4.67 $Y2=2
r56 2 29 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.565
+ $Y=1.485 $X2=3.71 $Y2=2.34
r57 2 18 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=3.565
+ $Y=1.485 $X2=3.71 $Y2=1.66
r58 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=1.485 $X2=2.75 $Y2=2.34
r59 1 12 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=2.625
+ $Y=1.485 $X2=2.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A_807_297# 1 2 9 11 13 16
r33 11 18 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.66 $Y=1.665 $X2=5.66
+ $Y2=1.58
r34 11 13 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.66 $Y=1.665
+ $X2=5.66 $Y2=2.34
r35 10 16 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.345 $Y=1.58
+ $X2=4.18 $Y2=1.58
r36 9 18 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.495 $Y=1.58
+ $X2=5.66 $Y2=1.58
r37 9 10 75.0267 $w=1.68e-07 $l=1.15e-06 $layer=LI1_cond $X=5.495 $Y=1.58
+ $X2=4.345 $Y2=1.58
r38 2 18 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=1.485 $X2=5.66 $Y2=1.66
r39 2 13 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.515
+ $Y=1.485 $X2=5.66 $Y2=2.34
r40 1 16 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=4.035
+ $Y=1.485 $X2=4.18 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%A_27_47# 1 2 3 4 5 6 19 21 23 30 31 32 35
+ 39 43 47 50 51
r93 49 51 9.67895 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.01 $Y=0.58
+ $X2=5.175 $Y2=0.58
r94 49 50 15.9354 $w=6.48e-07 $l=5.05e-07 $layer=LI1_cond $X=5.01 $Y=0.58
+ $X2=4.505 $Y2=0.58
r95 41 43 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.14 $Y=0.715
+ $X2=6.14 $Y2=0.38
r96 39 41 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=5.975 $Y=0.81
+ $X2=6.14 $Y2=0.715
r97 39 51 46.6986 $w=1.88e-07 $l=8e-07 $layer=LI1_cond $X=5.975 $Y=0.81
+ $X2=5.175 $Y2=0.81
r98 38 47 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.815 $Y=0.81
+ $X2=3.625 $Y2=0.81
r99 38 50 40.2775 $w=1.88e-07 $l=6.9e-07 $layer=LI1_cond $X=3.815 $Y=0.81
+ $X2=4.505 $Y2=0.81
r100 33 47 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.625 $Y=0.715
+ $X2=3.625 $Y2=0.81
r101 33 35 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.625 $Y=0.715
+ $X2=3.625 $Y2=0.38
r102 31 47 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.435 $Y=0.81
+ $X2=3.625 $Y2=0.81
r103 31 32 45.5311 $w=1.88e-07 $l=7.8e-07 $layer=LI1_cond $X=3.435 $Y=0.81
+ $X2=2.655 $Y2=0.81
r104 30 32 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.57 $Y=0.715
+ $X2=2.655 $Y2=0.81
r105 29 30 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.57 $Y=0.485
+ $X2=2.57 $Y2=0.715
r106 26 28 47.0998 $w=2.28e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=0.37
+ $X2=2.14 $Y2=0.37
r107 24 46 3.603 $w=2.3e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=0.217 $Y2=0.37
r108 24 26 42.8408 $w=2.28e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=0.37
+ $X2=1.2 $Y2=0.37
r109 23 29 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.485 $Y=0.37
+ $X2=2.57 $Y2=0.485
r110 23 28 17.2866 $w=2.28e-07 $l=3.45e-07 $layer=LI1_cond $X=2.485 $Y=0.37
+ $X2=2.14 $Y2=0.37
r111 19 46 3.23707 $w=2.55e-07 $l=1.15e-07 $layer=LI1_cond $X=0.217 $Y=0.485
+ $X2=0.217 $Y2=0.37
r112 19 21 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.217 $Y=0.485
+ $X2=0.217 $Y2=0.74
r113 6 43 91 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.235 $X2=6.14 $Y2=0.38
r114 5 49 45.5 $w=1.7e-07 $l=6.23298e-07 $layer=licon1_NDIFF $count=4 $X=4.455
+ $Y=0.235 $X2=5.01 $Y2=0.38
r115 4 35 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.515
+ $Y=0.235 $X2=3.65 $Y2=0.38
r116 3 28 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r117 2 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r118 1 46 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r119 1 21 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_2%VGND 1 2 3 12 16 20 23 24 26 27 28 30 49
+ 50 53
r79 53 54 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r80 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r81 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r82 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r83 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r84 43 46 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r85 43 44 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r86 41 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r87 41 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r88 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r89 38 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.06
+ $Y2=0
r90 38 40 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.25 $Y=0 $X2=3.91
+ $Y2=0
r91 37 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r92 36 37 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r93 32 36 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r94 30 53 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.06
+ $Y2=0
r95 30 36 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=2.53
+ $Y2=0
r96 28 37 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r97 28 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r98 26 46 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.29
+ $Y2=0
r99 26 27 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.355 $Y=0 $X2=5.545
+ $Y2=0
r100 25 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=6.21 $Y2=0
r101 25 27 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.545
+ $Y2=0
r102 23 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.035 $Y=0
+ $X2=3.91 $Y2=0
r103 23 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0 $X2=4.12
+ $Y2=0
r104 22 43 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.205 $Y=0
+ $X2=4.37 $Y2=0
r105 22 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.205 $Y=0 $X2=4.12
+ $Y2=0
r106 18 27 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.545 $Y=0.085
+ $X2=5.545 $Y2=0
r107 18 20 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.545 $Y=0.085
+ $X2=5.545 $Y2=0.38
r108 14 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.12 $Y=0.085
+ $X2=4.12 $Y2=0
r109 14 16 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.12 $Y=0.085
+ $X2=4.12 $Y2=0.38
r110 10 53 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.06 $Y2=0
r111 10 12 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.06 $Y=0.085
+ $X2=3.06 $Y2=0.38
r112 3 20 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.58 $Y2=0.38
r113 2 16 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.12 $Y2=0.38
r114 1 12 182 $w=1.7e-07 $l=6.78638e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=3.035 $Y2=0.38
.ends

