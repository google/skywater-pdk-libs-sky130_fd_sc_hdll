* NGSPICE file created from sky130_fd_sc_hdll__o21ai_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
M1000 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=1.2e+12p pd=1.04e+07u as=1.2e+12p ps=1.04e+07u
M1001 a_32_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=1.4625e+12p pd=1.36e+07u as=8.515e+11p ps=7.82e+06u
M1002 a_32_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.49e+12p pd=1.298e+07u as=0p ps=0u
M1004 a_123_297# A2 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_32_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND A2 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND A2 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Y B1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=4.615e+11p pd=4.02e+06u as=0p ps=0u
M1012 a_32_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y A2 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND A1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 Y B1 a_32_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 Y B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_32_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_32_47# B1 Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 a_123_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 VPWR A1 a_123_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

