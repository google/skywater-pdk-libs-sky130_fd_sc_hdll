* File: sky130_fd_sc_hdll__sdfsbp_2.pxi.spice
* Created: Wed Sep  2 08:51:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%SCD N_SCD_c_294_n N_SCD_c_298_n N_SCD_c_295_n
+ N_SCD_M1038_g N_SCD_c_299_n N_SCD_M1007_g SCD SCD
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%SCD
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%SCE N_SCE_M1028_g N_SCE_c_336_n N_SCE_c_337_n
+ N_SCE_M1036_g N_SCE_c_338_n N_SCE_c_339_n N_SCE_M1011_g N_SCE_M1004_g
+ N_SCE_c_331_n N_SCE_c_350_n N_SCE_c_374_p SCE N_SCE_c_332_n N_SCE_c_333_n
+ N_SCE_c_334_n N_SCE_c_335_n SCE PM_SKY130_FD_SC_HDLL__SDFSBP_2%SCE
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%D N_D_c_433_n N_D_c_438_n N_D_M1040_g
+ N_D_M1032_g D D N_D_c_435_n N_D_c_436_n PM_SKY130_FD_SC_HDLL__SDFSBP_2%D
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_349_21# N_A_349_21#_M1004_s
+ N_A_349_21#_M1011_s N_A_349_21#_M1000_g N_A_349_21#_c_484_n
+ N_A_349_21#_c_485_n N_A_349_21#_M1022_g N_A_349_21#_c_480_n
+ N_A_349_21#_c_481_n N_A_349_21#_c_482_n N_A_349_21#_c_483_n
+ N_A_349_21#_c_488_n N_A_349_21#_c_489_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_349_21#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%CLK N_CLK_M1044_g N_CLK_c_555_n N_CLK_M1017_g
+ N_CLK_c_556_n N_CLK_c_560_n N_CLK_c_561_n CLK CLK N_CLK_c_557_n N_CLK_c_558_n
+ N_CLK_c_559_n N_CLK_c_564_n CLK PM_SKY130_FD_SC_HDLL__SDFSBP_2%CLK
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_693_369# N_A_693_369#_M1017_s
+ N_A_693_369#_M1044_s N_A_693_369#_c_644_n N_A_693_369#_c_645_n
+ N_A_693_369#_M1027_g N_A_693_369#_c_627_n N_A_693_369#_M1018_g
+ N_A_693_369#_c_628_n N_A_693_369#_c_629_n N_A_693_369#_M1031_g
+ N_A_693_369#_c_646_n N_A_693_369#_M1041_g N_A_693_369#_c_647_n
+ N_A_693_369#_c_648_n N_A_693_369#_M1012_g N_A_693_369#_M1045_g
+ N_A_693_369#_c_631_n N_A_693_369#_c_661_n N_A_693_369#_c_632_n
+ N_A_693_369#_c_649_n N_A_693_369#_c_650_n N_A_693_369#_c_633_n
+ N_A_693_369#_c_634_n N_A_693_369#_c_726_p N_A_693_369#_c_635_n
+ N_A_693_369#_c_636_n N_A_693_369#_c_637_n N_A_693_369#_c_638_n
+ N_A_693_369#_c_639_n N_A_693_369#_c_640_n N_A_693_369#_c_641_n
+ N_A_693_369#_c_655_n N_A_693_369#_c_656_n N_A_693_369#_c_657_n
+ N_A_693_369#_c_658_n N_A_693_369#_c_659_n N_A_693_369#_c_776_p
+ N_A_693_369#_c_642_n N_A_693_369#_c_660_n N_A_693_369#_c_643_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_693_369#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_877_369# N_A_877_369#_M1018_d
+ N_A_877_369#_M1027_d N_A_877_369#_c_930_n N_A_877_369#_c_920_n
+ N_A_877_369#_c_931_n N_A_877_369#_c_932_n N_A_877_369#_c_933_n
+ N_A_877_369#_M1003_g N_A_877_369#_M1024_g N_A_877_369#_M1005_g
+ N_A_877_369#_c_935_n N_A_877_369#_M1009_g N_A_877_369#_c_936_n
+ N_A_877_369#_c_937_n N_A_877_369#_c_976_n N_A_877_369#_c_923_n
+ N_A_877_369#_c_924_n N_A_877_369#_c_925_n N_A_877_369#_c_926_n
+ N_A_877_369#_c_927_n N_A_877_369#_c_928_n N_A_877_369#_c_929_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_877_369#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1219_21# N_A_1219_21#_M1021_s
+ N_A_1219_21#_M1008_d N_A_1219_21#_M1029_g N_A_1219_21#_c_1104_n
+ N_A_1219_21#_c_1110_n N_A_1219_21#_M1042_g N_A_1219_21#_c_1111_n
+ N_A_1219_21#_c_1105_n N_A_1219_21#_c_1112_n N_A_1219_21#_c_1113_n
+ N_A_1219_21#_c_1106_n N_A_1219_21#_c_1167_p N_A_1219_21#_c_1107_n
+ N_A_1219_21#_c_1108_n PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1219_21#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1075_413# N_A_1075_413#_M1031_d
+ N_A_1075_413#_M1003_d N_A_1075_413#_c_1210_n N_A_1075_413#_c_1198_n
+ N_A_1075_413#_c_1211_n N_A_1075_413#_M1008_g N_A_1075_413#_c_1199_n
+ N_A_1075_413#_M1021_g N_A_1075_413#_c_1212_n N_A_1075_413#_c_1213_n
+ N_A_1075_413#_M1035_g N_A_1075_413#_M1010_g N_A_1075_413#_c_1200_n
+ N_A_1075_413#_c_1201_n N_A_1075_413#_c_1230_n N_A_1075_413#_c_1214_n
+ N_A_1075_413#_c_1202_n N_A_1075_413#_c_1203_n N_A_1075_413#_c_1204_n
+ N_A_1075_413#_c_1205_n N_A_1075_413#_c_1206_n N_A_1075_413#_c_1207_n
+ N_A_1075_413#_c_1208_n N_A_1075_413#_c_1209_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1075_413#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%SET_B N_SET_B_c_1360_n N_SET_B_c_1361_n
+ N_SET_B_M1023_g N_SET_B_M1025_g N_SET_B_c_1362_n N_SET_B_M1013_g
+ N_SET_B_M1043_g N_SET_B_c_1359_n N_SET_B_c_1365_n N_SET_B_c_1366_n
+ N_SET_B_c_1367_n N_SET_B_c_1368_n N_SET_B_c_1369_n N_SET_B_c_1370_n
+ N_SET_B_c_1371_n SET_B N_SET_B_c_1372_n SET_B
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%SET_B
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1930_295# N_A_1930_295#_M1001_d
+ N_A_1930_295#_M1002_d N_A_1930_295#_c_1510_n N_A_1930_295#_c_1511_n
+ N_A_1930_295#_M1020_g N_A_1930_295#_c_1512_n N_A_1930_295#_c_1513_n
+ N_A_1930_295#_M1039_g N_A_1930_295#_c_1504_n N_A_1930_295#_c_1505_n
+ N_A_1930_295#_c_1506_n N_A_1930_295#_c_1507_n N_A_1930_295#_c_1516_n
+ N_A_1930_295#_c_1517_n N_A_1930_295#_c_1508_n N_A_1930_295#_c_1509_n
+ N_A_1930_295#_c_1518_n PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1930_295#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1735_329# N_A_1735_329#_M1005_d
+ N_A_1735_329#_M1012_d N_A_1735_329#_M1013_d N_A_1735_329#_c_1623_n
+ N_A_1735_329#_c_1624_n N_A_1735_329#_M1002_g N_A_1735_329#_M1001_g
+ N_A_1735_329#_c_1611_n N_A_1735_329#_c_1612_n N_A_1735_329#_M1015_g
+ N_A_1735_329#_c_1626_n N_A_1735_329#_M1019_g N_A_1735_329#_c_1613_n
+ N_A_1735_329#_M1030_g N_A_1735_329#_c_1627_n N_A_1735_329#_M1037_g
+ N_A_1735_329#_c_1614_n N_A_1735_329#_c_1615_n N_A_1735_329#_c_1630_n
+ N_A_1735_329#_c_1631_n N_A_1735_329#_M1016_g N_A_1735_329#_M1033_g
+ N_A_1735_329#_c_1617_n N_A_1735_329#_c_1640_n N_A_1735_329#_c_1641_n
+ N_A_1735_329#_c_1633_n N_A_1735_329#_c_1618_n N_A_1735_329#_c_1634_n
+ N_A_1735_329#_c_1619_n N_A_1735_329#_c_1620_n N_A_1735_329#_c_1621_n
+ N_A_1735_329#_c_1636_n N_A_1735_329#_c_1667_n N_A_1735_329#_c_1637_n
+ N_A_1735_329#_c_1675_n N_A_1735_329#_c_1622_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_1735_329#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_2739_47# N_A_2739_47#_M1033_s
+ N_A_2739_47#_M1016_s N_A_2739_47#_c_1800_n N_A_2739_47#_M1014_g
+ N_A_2739_47#_c_1795_n N_A_2739_47#_M1006_g N_A_2739_47#_c_1801_n
+ N_A_2739_47#_M1026_g N_A_2739_47#_c_1796_n N_A_2739_47#_M1034_g
+ N_A_2739_47#_c_1797_n N_A_2739_47#_c_1802_n N_A_2739_47#_c_1798_n
+ N_A_2739_47#_c_1816_n N_A_2739_47#_c_1799_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_2739_47#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_27_369# N_A_27_369#_M1007_s
+ N_A_27_369#_M1022_d N_A_27_369#_c_1855_n N_A_27_369#_c_1856_n
+ N_A_27_369#_c_1857_n N_A_27_369#_c_1864_n N_A_27_369#_c_1871_n
+ N_A_27_369#_c_1858_n PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_27_369#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%VPWR N_VPWR_M1007_d N_VPWR_M1011_d
+ N_VPWR_M1044_d N_VPWR_M1042_d N_VPWR_M1023_d N_VPWR_M1020_d N_VPWR_M1002_s
+ N_VPWR_M1019_d N_VPWR_M1037_d N_VPWR_M1016_d N_VPWR_M1026_d N_VPWR_c_1908_n
+ N_VPWR_c_1909_n N_VPWR_c_1910_n N_VPWR_c_1911_n N_VPWR_c_1912_n
+ N_VPWR_c_1913_n N_VPWR_c_1914_n N_VPWR_c_1915_n N_VPWR_c_1916_n
+ N_VPWR_c_1917_n N_VPWR_c_1918_n N_VPWR_c_1919_n N_VPWR_c_1920_n
+ N_VPWR_c_1921_n N_VPWR_c_1922_n N_VPWR_c_1923_n N_VPWR_c_1924_n
+ N_VPWR_c_1925_n N_VPWR_c_1926_n N_VPWR_c_1927_n N_VPWR_c_1928_n VPWR
+ N_VPWR_c_1929_n N_VPWR_c_1930_n N_VPWR_c_1931_n N_VPWR_c_1932_n
+ N_VPWR_c_1933_n N_VPWR_c_1934_n N_VPWR_c_1935_n N_VPWR_c_1936_n
+ N_VPWR_c_1937_n N_VPWR_c_1938_n N_VPWR_c_1939_n N_VPWR_c_1940_n
+ N_VPWR_c_1907_n VPWR PM_SKY130_FD_SC_HDLL__SDFSBP_2%VPWR
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_199_47# N_A_199_47#_M1028_d
+ N_A_199_47#_M1031_s N_A_199_47#_M1040_d N_A_199_47#_M1003_s
+ N_A_199_47#_c_2154_n N_A_199_47#_c_2143_n N_A_199_47#_c_2147_n
+ N_A_199_47#_c_2148_n N_A_199_47#_c_2157_n N_A_199_47#_c_2144_n
+ N_A_199_47#_c_2149_n N_A_199_47#_c_2150_n N_A_199_47#_c_2145_n
+ N_A_199_47#_c_2152_n N_A_199_47#_c_2146_n
+ PM_SKY130_FD_SC_HDLL__SDFSBP_2%A_199_47#
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%Q_N N_Q_N_M1015_s N_Q_N_M1019_s Q_N Q_N Q_N Q_N
+ Q_N Q_N N_Q_N_c_2279_n PM_SKY130_FD_SC_HDLL__SDFSBP_2%Q_N
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%Q N_Q_M1006_d N_Q_M1014_s Q Q Q Q Q Q Q
+ N_Q_c_2305_n Q PM_SKY130_FD_SC_HDLL__SDFSBP_2%Q
x_PM_SKY130_FD_SC_HDLL__SDFSBP_2%VGND N_VGND_M1038_s N_VGND_M1000_d
+ N_VGND_M1004_d N_VGND_M1017_d N_VGND_M1029_d N_VGND_M1025_d N_VGND_M1043_d
+ N_VGND_M1015_d N_VGND_M1030_d N_VGND_M1033_d N_VGND_M1034_s N_VGND_c_2317_n
+ N_VGND_c_2318_n N_VGND_c_2319_n N_VGND_c_2320_n N_VGND_c_2321_n
+ N_VGND_c_2322_n N_VGND_c_2323_n N_VGND_c_2324_n N_VGND_c_2325_n
+ N_VGND_c_2326_n N_VGND_c_2327_n N_VGND_c_2328_n N_VGND_c_2329_n
+ N_VGND_c_2330_n N_VGND_c_2331_n N_VGND_c_2332_n N_VGND_c_2333_n
+ N_VGND_c_2334_n N_VGND_c_2335_n VGND N_VGND_c_2336_n N_VGND_c_2337_n
+ N_VGND_c_2338_n N_VGND_c_2339_n N_VGND_c_2340_n N_VGND_c_2341_n
+ N_VGND_c_2342_n N_VGND_c_2343_n N_VGND_c_2344_n N_VGND_c_2345_n
+ N_VGND_c_2346_n VGND PM_SKY130_FD_SC_HDLL__SDFSBP_2%VGND
cc_1 VNB N_SCD_c_294_n 0.0611035f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.325
cc_2 VNB N_SCD_c_295_n 0.0186791f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_3 VNB SCD 0.0211184f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_4 VNB N_SCE_M1028_g 0.0328557f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.73
cc_5 VNB N_SCE_M1004_g 0.040964f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_6 VNB N_SCE_c_331_n 0.00686301f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_7 VNB N_SCE_c_332_n 0.022827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_SCE_c_333_n 0.0305635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_SCE_c_334_n 0.00345895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_SCE_c_335_n 0.00950707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_D_c_433_n 0.0102691f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.62
cc_12 VNB D 0.00527061f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_13 VNB N_D_c_435_n 0.0244402f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_14 VNB N_D_c_436_n 0.0170109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_349_21#_M1000_g 0.0310156f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_16 VNB N_A_349_21#_c_480_n 0.00445814f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_17 VNB N_A_349_21#_c_481_n 0.0435879f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=0.85
cc_18 VNB N_A_349_21#_c_482_n 0.015063f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_349_21#_c_483_n 0.00723186f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.16
cc_20 VNB N_CLK_c_555_n 0.017386f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_21 VNB N_CLK_c_556_n 0.0189011f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_22 VNB N_CLK_c_557_n 0.0170927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_CLK_c_558_n 0.018041f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.16
cc_24 VNB N_CLK_c_559_n 0.0169683f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.53
cc_25 VNB N_A_693_369#_c_627_n 0.0175643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_693_369#_c_628_n 0.0568461f $X=-0.19 $Y=-0.24 $X2=0.327 $Y2=1.16
cc_27 VNB N_A_693_369#_c_629_n 0.0174152f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_28 VNB N_A_693_369#_M1045_g 0.0243943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_693_369#_c_631_n 0.00444385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_693_369#_c_632_n 0.00137399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_693_369#_c_633_n 0.00761502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_693_369#_c_634_n 0.00370284f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_693_369#_c_635_n 0.0034525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_693_369#_c_636_n 0.0185312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_693_369#_c_637_n 0.0020228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_693_369#_c_638_n 0.0294047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_693_369#_c_639_n 0.0114808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_693_369#_c_640_n 2.43863e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_693_369#_c_641_n 0.00446849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_693_369#_c_642_n 0.011579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_693_369#_c_643_n 0.0326406f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_877_369#_c_920_n 0.0484121f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_43 VNB N_A_877_369#_M1024_g 0.0313379f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_44 VNB N_A_877_369#_M1005_g 0.0378327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_877_369#_c_923_n 0.019416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_877_369#_c_924_n 0.00204181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_877_369#_c_925_n 0.00332704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_877_369#_c_926_n 0.00447837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_877_369#_c_927_n 0.00272906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_877_369#_c_928_n 0.0173258f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_877_369#_c_929_n 0.00482291f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_1219_21#_M1029_g 0.0185139f $X=-0.19 $Y=-0.24 $X2=0.32 $Y2=1.695
cc_53 VNB N_A_1219_21#_c_1104_n 0.0135546f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1219_21#_c_1105_n 0.0072695f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1219_21#_c_1106_n 0.00485794f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1219_21#_c_1107_n 0.00281667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1219_21#_c_1108_n 0.031422f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1075_413#_c_1198_n 0.0134372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1075_413#_c_1199_n 0.0169531f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_60 VNB N_A_1075_413#_c_1200_n 0.0296707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1075_413#_c_1201_n 0.00696624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1075_413#_c_1202_n 0.00499843f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_A_1075_413#_c_1203_n 0.00176087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_A_1075_413#_c_1204_n 0.00237739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_A_1075_413#_c_1205_n 0.00718886f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_A_1075_413#_c_1206_n 0.0224114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_A_1075_413#_c_1207_n 0.0198052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_A_1075_413#_c_1208_n 0.020101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_A_1075_413#_c_1209_n 0.0200017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_SET_B_M1025_g 0.03768f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.165
cc_71 VNB N_SET_B_M1043_g 0.0487505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_SET_B_c_1359_n 0.0115466f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_73 VNB N_A_1930_295#_M1039_g 0.0239654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB N_A_1930_295#_c_1504_n 0.00837455f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_75 VNB N_A_1930_295#_c_1505_n 0.00149329f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_1930_295#_c_1506_n 0.0333096f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.16
cc_77 VNB N_A_1930_295#_c_1507_n 0.012176f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_A_1930_295#_c_1508_n 0.00793643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_A_1930_295#_c_1509_n 0.00312622f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_A_1735_329#_c_1611_n 0.0476297f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_81 VNB N_A_1735_329#_c_1612_n 0.019902f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=0.85
cc_82 VNB N_A_1735_329#_c_1613_n 0.0202814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_A_1735_329#_c_1614_n 0.0555202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_A_1735_329#_c_1615_n 0.0260454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_A_1735_329#_M1033_g 0.0326111f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_A_1735_329#_c_1617_n 0.00971673f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_A_1735_329#_c_1618_n 0.00460174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_1735_329#_c_1619_n 0.00332814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_1735_329#_c_1620_n 0.00806916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_A_1735_329#_c_1621_n 0.0429734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_A_1735_329#_c_1622_n 0.0209837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_A_2739_47#_c_1795_n 0.0176056f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_A_2739_47#_c_1796_n 0.0219834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_A_2739_47#_c_1797_n 0.00715705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_A_2739_47#_c_1798_n 0.00194757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_A_2739_47#_c_1799_n 0.0554028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VPWR_c_1907_n 0.649277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_A_199_47#_c_2143_n 0.00565332f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_99 VNB N_A_199_47#_c_2144_n 0.00132503f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_A_199_47#_c_2145_n 0.00436412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_A_199_47#_c_2146_n 0.00350897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB Q 0.00108985f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.53
cc_103 VNB N_VGND_c_2317_n 0.0102501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_2318_n 0.0172739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_2319_n 0.00479834f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_2320_n 0.0199154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_2321_n 0.00925188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_2322_n 0.00264923f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_2323_n 0.00469188f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_2324_n 0.0210126f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_2325_n 0.00709087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_2326_n 0.0145246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_2327_n 0.00356736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_2328_n 0.0112855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_2329_n 0.0343045f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_2330_n 0.0169909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_2331_n 0.0047213f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_2332_n 0.0220745f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_VGND_c_2333_n 0.00557808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_VGND_c_2334_n 0.0153065f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_VGND_c_2335_n 0.00625144f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_VGND_c_2336_n 0.0418631f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_VGND_c_2337_n 0.0623478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_VGND_c_2338_n 0.0755482f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_VGND_c_2339_n 0.0210195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_VGND_c_2340_n 0.00343497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_VGND_c_2341_n 0.00651182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_VGND_c_2342_n 0.0252938f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_VGND_c_2343_n 0.016038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_VGND_c_2344_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_VGND_c_2345_n 0.00403782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_VGND_c_2346_n 0.733196f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VPB N_SCD_c_294_n 0.00539454f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.325
cc_134 VPB N_SCD_c_298_n 0.0197136f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.62
cc_135 VPB N_SCD_c_299_n 0.049218f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_136 VPB SCD 0.0150047f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_137 VPB N_SCE_c_336_n 0.0141631f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.77
cc_138 VPB N_SCE_c_337_n 0.0221025f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_139 VPB N_SCE_c_338_n 0.0263105f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_140 VPB N_SCE_c_339_n 0.0305056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_SCE_c_332_n 0.0134912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_SCE_c_333_n 0.00526365f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_SCE_c_334_n 0.00431909f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_SCE_c_335_n 0.00618619f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_D_c_433_n 0.018242f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.62
cc_146 VPB N_D_c_438_n 0.0222486f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_147 VPB D 0.00243874f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.695
cc_148 VPB N_A_349_21#_c_484_n 0.0220272f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_349_21#_c_485_n 0.0251734f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_150 VPB N_A_349_21#_c_480_n 0.0105451f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_151 VPB N_A_349_21#_c_481_n 0.0141049f $X=-0.19 $Y=1.305 $X2=0.225 $Y2=0.85
cc_152 VPB N_A_349_21#_c_488_n 0.00405142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_349_21#_c_489_n 0.0117185f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_CLK_c_560_n 0.0122703f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_CLK_c_561_n 0.0358246f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_CLK_c_557_n 0.0107383f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_CLK_c_558_n 0.0172631f $X=-0.19 $Y=1.305 $X2=0.225 $Y2=1.16
cc_158 VPB N_CLK_c_564_n 0.00254669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_693_369#_c_644_n 0.0149524f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_160 VPB N_A_693_369#_c_645_n 0.0250798f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.695
cc_161 VPB N_A_693_369#_c_646_n 0.0571331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_A_693_369#_c_647_n 0.00755818f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_693_369#_c_648_n 0.0202963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_693_369#_c_649_n 0.00152611f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_693_369#_c_650_n 0.00168159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_693_369#_c_635_n 0.00340077f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_A_693_369#_c_636_n 0.0107444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_A_693_369#_c_637_n 0.00132283f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_A_693_369#_c_638_n 0.0051338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_A_693_369#_c_655_n 0.0041777f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_A_693_369#_c_656_n 0.00689926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_693_369#_c_657_n 4.12566e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_A_693_369#_c_658_n 0.00751057f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_A_693_369#_c_659_n 0.00220179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_A_693_369#_c_660_n 0.00224501f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_A_877_369#_c_930_n 0.0246271f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_177 VPB N_A_877_369#_c_931_n 0.0201586f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_178 VPB N_A_877_369#_c_932_n 0.0106624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_A_877_369#_c_933_n 0.0193133f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_180 VPB N_A_877_369#_M1005_g 0.0159604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_A_877_369#_c_935_n 0.0634698f $X=-0.19 $Y=1.305 $X2=0.225 $Y2=1.53
cc_182 VPB N_A_877_369#_c_936_n 0.0048654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_A_877_369#_c_937_n 0.00969938f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_A_877_369#_c_925_n 0.0012792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_A_877_369#_c_926_n 3.90977e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_877_369#_c_927_n 0.00759351f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_A_877_369#_c_928_n 0.0170356f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_A_1219_21#_c_1104_n 0.0179577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_A_1219_21#_c_1110_n 0.0632234f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_190 VPB N_A_1219_21#_c_1111_n 0.00179081f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_191 VPB N_A_1219_21#_c_1112_n 0.00592289f $X=-0.19 $Y=1.305 $X2=0.225
+ $Y2=1.16
cc_192 VPB N_A_1219_21#_c_1113_n 7.95296e-19 $X=-0.19 $Y=1.305 $X2=0.225
+ $Y2=1.53
cc_193 VPB N_A_1075_413#_c_1210_n 0.030077f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.165
cc_194 VPB N_A_1075_413#_c_1211_n 0.0238391f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_195 VPB N_A_1075_413#_c_1212_n 0.00875029f $X=-0.19 $Y=1.305 $X2=0.26
+ $Y2=1.16
cc_196 VPB N_A_1075_413#_c_1213_n 0.0207135f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_197 VPB N_A_1075_413#_c_1214_n 0.0161187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_A_1075_413#_c_1202_n 0.00609637f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_A_1075_413#_c_1203_n 0.00282717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1075_413#_c_1204_n 0.00137632f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_A_1075_413#_c_1205_n 0.00100061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_A_1075_413#_c_1206_n 0.00401989f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_A_1075_413#_c_1208_n 0.00937693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_SET_B_c_1360_n 0.00902906f $X=-0.19 $Y=1.305 $X2=0.32 $Y2=1.62
cc_205 VPB N_SET_B_c_1361_n 0.0618594f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.73
cc_206 VPB N_SET_B_c_1362_n 0.0583889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_SET_B_M1043_g 0.00785288f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_SET_B_c_1359_n 0.00566645f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_209 VPB N_SET_B_c_1365_n 0.0151814f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_SET_B_c_1366_n 0.0119596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_SET_B_c_1367_n 0.01954f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_SET_B_c_1368_n 0.015713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_SET_B_c_1369_n 0.00201394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_SET_B_c_1370_n 0.00562445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_SET_B_c_1371_n 0.00390488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_SET_B_c_1372_n 0.00832064f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_A_1930_295#_c_1510_n 0.0195441f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.165
cc_218 VPB N_A_1930_295#_c_1511_n 0.0237364f $X=-0.19 $Y=1.305 $X2=0.32
+ $Y2=1.695
cc_219 VPB N_A_1930_295#_c_1512_n 0.0315412f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_A_1930_295#_c_1513_n 0.00816498f $X=-0.19 $Y=1.305 $X2=0.15
+ $Y2=0.765
cc_221 VPB N_A_1930_295#_c_1504_n 0.0146843f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_222 VPB N_A_1930_295#_c_1507_n 0.00838362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_A_1930_295#_c_1516_n 6.44545e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_A_1930_295#_c_1517_n 0.0205401f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_A_1930_295#_c_1518_n 3.56731e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_A_1735_329#_c_1623_n 0.0287274f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_227 VPB N_A_1735_329#_c_1624_n 0.0506654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_A_1735_329#_c_1611_n 0.0297022f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_229 VPB N_A_1735_329#_c_1626_n 0.0193293f $X=-0.19 $Y=1.305 $X2=0.225
+ $Y2=1.16
cc_230 VPB N_A_1735_329#_c_1627_n 0.0195239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_A_1735_329#_c_1614_n 0.0337413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_A_1735_329#_c_1615_n 0.0217262f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_A_1735_329#_c_1630_n 0.0178894f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_A_1735_329#_c_1631_n 0.0294934f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_A_1735_329#_c_1617_n 6.17389e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB N_A_1735_329#_c_1633_n 0.0112061f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_A_1735_329#_c_1634_n 0.00434434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_A_1735_329#_c_1621_n 0.00118414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_A_1735_329#_c_1636_n 0.00743639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_A_1735_329#_c_1637_n 0.00232516f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_A_2739_47#_c_1800_n 0.0168206f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=2.165
cc_242 VPB N_A_2739_47#_c_1801_n 0.0207521f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_243 VPB N_A_2739_47#_c_1802_n 0.0124243f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_A_2739_47#_c_1798_n 0.00246016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_A_2739_47#_c_1799_n 0.0278658f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_A_27_369#_c_1855_n 0.0170416f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.165
cc_247 VPB N_A_27_369#_c_1856_n 8.25607e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_A_27_369#_c_1857_n 0.00945086f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.695
cc_249 VPB N_A_27_369#_c_1858_n 0.00263317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_VPWR_c_1908_n 0.00243094f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_VPWR_c_1909_n 0.00982329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_VPWR_c_1910_n 0.0155023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_VPWR_c_1911_n 0.0056301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_VPWR_c_1912_n 0.0049533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_VPWR_c_1913_n 0.00925213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_VPWR_c_1914_n 0.00315146f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_VPWR_c_1915_n 0.0059826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_VPWR_c_1916_n 0.0188969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_VPWR_c_1917_n 0.00697695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_VPWR_c_1918_n 0.0181682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_VPWR_c_1919_n 0.00380756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_VPWR_c_1920_n 0.0112596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_VPWR_c_1921_n 0.0477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_VPWR_c_1922_n 0.0240263f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_VPWR_c_1923_n 0.0321741f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_VPWR_c_1924_n 0.00609289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_VPWR_c_1925_n 0.0220745f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_VPWR_c_1926_n 0.00555219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_VPWR_c_1927_n 0.0153065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_VPWR_c_1928_n 0.00628472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_VPWR_c_1929_n 0.0143786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 VPB N_VPWR_c_1930_n 0.0516265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_273 VPB N_VPWR_c_1931_n 0.0567553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_274 VPB N_VPWR_c_1932_n 0.0174067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_275 VPB N_VPWR_c_1933_n 0.0209859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_276 VPB N_VPWR_c_1934_n 0.00426174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_277 VPB N_VPWR_c_1935_n 0.00651315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_278 VPB N_VPWR_c_1936_n 0.00546385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_279 VPB N_VPWR_c_1937_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_280 VPB N_VPWR_c_1938_n 0.00644418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_281 VPB N_VPWR_c_1939_n 0.00513206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_282 VPB N_VPWR_c_1940_n 0.00401193f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_283 VPB N_VPWR_c_1907_n 0.0845131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_284 VPB N_A_199_47#_c_2147_n 9.1992e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_285 VPB N_A_199_47#_c_2148_n 0.00241998f $X=-0.19 $Y=1.305 $X2=0.225 $Y2=1.16
cc_286 VPB N_A_199_47#_c_2149_n 0.0331926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_287 VPB N_A_199_47#_c_2150_n 0.00325906f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_288 VPB N_A_199_47#_c_2145_n 0.00362768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_289 VPB N_A_199_47#_c_2152_n 0.00776824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_290 VPB N_A_199_47#_c_2146_n 0.00386902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_291 VPB Q 0.00119084f $X=-0.19 $Y=1.305 $X2=0.225 $Y2=1.53
cc_292 N_SCD_c_294_n N_SCE_M1028_g 0.00412822f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_293 N_SCD_c_295_n N_SCE_M1028_g 0.0324759f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_294 SCD N_SCE_M1028_g 2.38515e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_295 N_SCD_c_298_n N_SCE_c_336_n 0.00344219f $X=0.32 $Y=1.62 $X2=0 $Y2=0
cc_296 N_SCD_c_299_n N_SCE_c_336_n 0.00779034f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_297 N_SCD_c_299_n N_SCE_c_337_n 0.0232684f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_298 SCD N_SCE_c_350_n 0.00154533f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_299 N_SCD_c_294_n N_SCE_c_332_n 0.0165133f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_300 SCD N_SCE_c_332_n 3.37737e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_301 N_SCD_c_294_n N_SCE_c_335_n 0.00653076f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_302 N_SCD_c_299_n N_SCE_c_335_n 0.00324317f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_303 SCD N_SCE_c_335_n 0.0647404f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_304 N_SCD_c_299_n N_A_27_369#_c_1855_n 0.00843386f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_305 N_SCD_c_299_n N_A_27_369#_c_1856_n 0.0155652f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_306 N_SCD_c_294_n N_A_27_369#_c_1857_n 5.05332e-19 $X=0.32 $Y=1.325 $X2=0
+ $Y2=0
cc_307 N_SCD_c_299_n N_A_27_369#_c_1857_n 0.00303881f $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_308 SCD N_A_27_369#_c_1857_n 0.0232839f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_309 N_SCD_c_299_n N_A_27_369#_c_1864_n 7.29534e-19 $X=0.495 $Y=1.77 $X2=0
+ $Y2=0
cc_310 N_SCD_c_299_n N_VPWR_c_1908_n 0.0115093f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_311 N_SCD_c_299_n N_VPWR_c_1929_n 0.00317293f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_312 N_SCD_c_299_n N_VPWR_c_1907_n 0.0048112f $X=0.495 $Y=1.77 $X2=0 $Y2=0
cc_313 N_SCD_c_295_n N_A_199_47#_c_2154_n 8.18391e-19 $X=0.47 $Y=0.73 $X2=0
+ $Y2=0
cc_314 N_SCD_c_294_n N_VGND_c_2318_n 0.00470012f $X=0.32 $Y=1.325 $X2=0 $Y2=0
cc_315 N_SCD_c_295_n N_VGND_c_2318_n 0.0144114f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_316 SCD N_VGND_c_2318_n 0.0231483f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_317 N_SCD_c_295_n N_VGND_c_2336_n 0.00447018f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_318 N_SCD_c_295_n N_VGND_c_2346_n 0.00776376f $X=0.47 $Y=0.73 $X2=0 $Y2=0
cc_319 SCD N_VGND_c_2346_n 0.00108189f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_320 N_SCE_c_331_n N_D_c_433_n 0.00233005f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_321 N_SCE_c_332_n N_D_c_433_n 0.0243839f $X=0.92 $Y=1.245 $X2=0 $Y2=0
cc_322 N_SCE_c_335_n N_D_c_433_n 2.84464e-19 $X=0.715 $Y=1.19 $X2=0 $Y2=0
cc_323 N_SCE_c_336_n N_D_c_438_n 0.016356f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_324 N_SCE_c_337_n N_D_c_438_n 0.0474155f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_325 N_SCE_M1028_g D 0.00353673f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_326 N_SCE_c_336_n D 0.00546242f $X=0.965 $Y=1.67 $X2=0 $Y2=0
cc_327 N_SCE_c_337_n D 4.10161e-19 $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_328 N_SCE_c_331_n D 0.0296879f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_329 N_SCE_c_350_n D 7.09436e-19 $X=0.86 $Y=1.19 $X2=0 $Y2=0
cc_330 N_SCE_c_332_n D 0.0045233f $X=0.92 $Y=1.245 $X2=0 $Y2=0
cc_331 N_SCE_c_335_n D 0.0695562f $X=0.715 $Y=1.19 $X2=0 $Y2=0
cc_332 N_SCE_M1028_g N_D_c_435_n 0.0192745f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_333 N_SCE_c_335_n N_D_c_435_n 2.52763e-19 $X=0.715 $Y=1.19 $X2=0 $Y2=0
cc_334 N_SCE_M1028_g N_D_c_436_n 0.0120539f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_335 N_SCE_c_338_n N_A_349_21#_c_480_n 0.00698607f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_336 N_SCE_M1004_g N_A_349_21#_c_480_n 0.00264967f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_337 N_SCE_c_331_n N_A_349_21#_c_480_n 0.0173777f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_338 N_SCE_c_374_p N_A_349_21#_c_480_n 6.89964e-19 $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_339 N_SCE_c_333_n N_A_349_21#_c_480_n 0.00255221f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_340 N_SCE_c_334_n N_A_349_21#_c_480_n 0.0364712f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_341 N_SCE_c_331_n N_A_349_21#_c_481_n 0.00893887f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_342 N_SCE_c_333_n N_A_349_21#_c_481_n 0.0167318f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_343 N_SCE_c_334_n N_A_349_21#_c_481_n 6.66667e-19 $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_344 N_SCE_M1004_g N_A_349_21#_c_482_n 0.00850096f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_345 N_SCE_c_331_n N_A_349_21#_c_482_n 0.00905152f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_346 N_SCE_c_374_p N_A_349_21#_c_482_n 0.00100397f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_347 N_SCE_c_333_n N_A_349_21#_c_482_n 0.0028405f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_348 N_SCE_c_334_n N_A_349_21#_c_482_n 0.00946334f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_349 N_SCE_M1004_g N_A_349_21#_c_483_n 0.00604711f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_350 N_SCE_c_339_n N_A_349_21#_c_488_n 0.0080547f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_351 N_SCE_c_339_n N_A_349_21#_c_489_n 0.00522959f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_352 N_SCE_c_333_n N_A_349_21#_c_489_n 3.7662e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_353 N_SCE_c_334_n N_A_349_21#_c_489_n 0.00610545f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_354 N_SCE_c_333_n N_CLK_c_557_n 0.00434241f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_355 N_SCE_c_334_n N_CLK_c_557_n 6.64246e-19 $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_356 N_SCE_c_338_n N_CLK_c_558_n 0.00539997f $X=2.835 $Y=1.67 $X2=0 $Y2=0
cc_357 N_SCE_c_374_p N_CLK_c_558_n 0.00158915f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_358 N_SCE_c_333_n N_CLK_c_558_n 0.00338404f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_359 N_SCE_c_334_n N_CLK_c_558_n 0.0336849f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_360 N_SCE_c_339_n N_CLK_c_564_n 0.0123265f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_361 N_SCE_c_334_n N_CLK_c_564_n 0.00589458f $X=2.735 $Y=1.16 $X2=0 $Y2=0
cc_362 N_SCE_c_339_n N_A_693_369#_c_661_n 0.00418407f $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_363 N_SCE_M1004_g N_A_693_369#_c_632_n 0.0037991f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_SCE_c_339_n N_A_693_369#_c_650_n 6.23463e-19 $X=2.835 $Y=1.77 $X2=0
+ $Y2=0
cc_365 N_SCE_M1004_g N_A_693_369#_c_634_n 0.00453904f $X=2.86 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_SCE_c_337_n N_A_27_369#_c_1856_n 0.0141586f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_367 N_SCE_c_331_n N_A_27_369#_c_1856_n 0.00493245f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_368 N_SCE_c_350_n N_A_27_369#_c_1856_n 0.00104372f $X=0.86 $Y=1.19 $X2=0
+ $Y2=0
cc_369 N_SCE_c_332_n N_A_27_369#_c_1856_n 8.01447e-19 $X=0.92 $Y=1.245 $X2=0
+ $Y2=0
cc_370 N_SCE_c_335_n N_A_27_369#_c_1856_n 0.0214161f $X=0.715 $Y=1.19 $X2=0
+ $Y2=0
cc_371 N_SCE_c_337_n N_A_27_369#_c_1864_n 0.00505317f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_372 N_SCE_c_337_n N_A_27_369#_c_1871_n 0.00471403f $X=0.965 $Y=1.77 $X2=0
+ $Y2=0
cc_373 N_SCE_c_337_n N_VPWR_c_1908_n 0.0042885f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_374 N_SCE_c_339_n N_VPWR_c_1909_n 0.0050341f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_375 N_SCE_c_337_n N_VPWR_c_1930_n 0.0051032f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_376 N_SCE_c_339_n N_VPWR_c_1930_n 0.00635181f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_377 N_SCE_c_337_n N_VPWR_c_1907_n 0.00666674f $X=0.965 $Y=1.77 $X2=0 $Y2=0
cc_378 N_SCE_c_339_n N_VPWR_c_1907_n 0.0129491f $X=2.835 $Y=1.77 $X2=0 $Y2=0
cc_379 N_SCE_M1028_g N_A_199_47#_c_2154_n 0.00552246f $X=0.92 $Y=0.445 $X2=0
+ $Y2=0
cc_380 N_SCE_c_331_n N_A_199_47#_c_2154_n 0.0104741f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_381 N_SCE_c_331_n N_A_199_47#_c_2157_n 0.00565156f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_382 N_SCE_c_338_n N_A_199_47#_c_2149_n 0.00717356f $X=2.835 $Y=1.67 $X2=0
+ $Y2=0
cc_383 N_SCE_c_331_n N_A_199_47#_c_2149_n 0.0490896f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_384 N_SCE_c_374_p N_A_199_47#_c_2149_n 0.0249445f $X=2.73 $Y=1.19 $X2=0 $Y2=0
cc_385 N_SCE_c_334_n N_A_199_47#_c_2149_n 0.0169978f $X=2.735 $Y=1.16 $X2=0
+ $Y2=0
cc_386 N_SCE_c_331_n N_A_199_47#_c_2150_n 0.0305807f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_387 N_SCE_c_331_n N_A_199_47#_c_2145_n 0.0189564f $X=2.585 $Y=1.19 $X2=0
+ $Y2=0
cc_388 N_SCE_M1028_g N_VGND_c_2318_n 0.00226101f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_389 N_SCE_M1004_g N_VGND_c_2319_n 0.00245709f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_390 N_SCE_c_331_n N_VGND_c_2319_n 0.00127321f $X=2.585 $Y=1.19 $X2=0 $Y2=0
cc_391 N_SCE_M1004_g N_VGND_c_2320_n 0.00585385f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_392 N_SCE_M1004_g N_VGND_c_2321_n 0.00496436f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_393 N_SCE_M1028_g N_VGND_c_2336_n 0.00555741f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_394 N_SCE_M1028_g N_VGND_c_2346_n 0.0098437f $X=0.92 $Y=0.445 $X2=0 $Y2=0
cc_395 N_SCE_M1004_g N_VGND_c_2346_n 0.0132032f $X=2.86 $Y=0.445 $X2=0 $Y2=0
cc_396 N_SCE_c_335_n N_VGND_c_2346_n 0.0128517f $X=0.715 $Y=1.19 $X2=0 $Y2=0
cc_397 D N_A_349_21#_M1000_g 0.00101694f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_398 N_D_c_436_n N_A_349_21#_M1000_g 0.018979f $X=1.34 $Y=0.765 $X2=0 $Y2=0
cc_399 N_D_c_433_n N_A_349_21#_c_484_n 0.018979f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_400 N_D_c_438_n N_A_349_21#_c_485_n 0.0424801f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_401 N_D_c_435_n N_A_349_21#_c_481_n 0.018979f $X=1.34 $Y=0.93 $X2=0 $Y2=0
cc_402 N_D_c_438_n N_A_27_369#_c_1856_n 0.00149383f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_403 D N_A_27_369#_c_1856_n 0.0125499f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_404 N_D_c_438_n N_A_27_369#_c_1864_n 0.00438564f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_405 N_D_c_438_n N_A_27_369#_c_1858_n 0.0135943f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_406 D N_A_27_369#_c_1858_n 0.00495298f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_407 N_D_c_438_n N_VPWR_c_1930_n 0.00429453f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_408 N_D_c_438_n N_VPWR_c_1907_n 0.0060009f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_409 D N_A_199_47#_c_2154_n 0.0230444f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_410 N_D_c_435_n N_A_199_47#_c_2154_n 6.89124e-19 $X=1.34 $Y=0.93 $X2=0 $Y2=0
cc_411 N_D_c_436_n N_A_199_47#_c_2154_n 0.0112593f $X=1.34 $Y=0.765 $X2=0 $Y2=0
cc_412 N_D_c_438_n N_A_199_47#_c_2157_n 0.00530414f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_413 D N_A_199_47#_c_2157_n 0.00194167f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_414 N_D_c_433_n N_A_199_47#_c_2150_n 0.00427772f $X=1.375 $Y=1.67 $X2=0 $Y2=0
cc_415 D N_A_199_47#_c_2150_n 0.0073578f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_416 N_D_c_438_n N_A_199_47#_c_2145_n 0.00168939f $X=1.375 $Y=1.77 $X2=0 $Y2=0
cc_417 D N_A_199_47#_c_2145_n 0.0510276f $X=1.08 $Y=0.765 $X2=0 $Y2=0
cc_418 N_D_c_436_n N_A_199_47#_c_2145_n 0.0116756f $X=1.34 $Y=0.765 $X2=0 $Y2=0
cc_419 N_D_c_436_n N_VGND_c_2336_n 0.00363059f $X=1.34 $Y=0.765 $X2=0 $Y2=0
cc_420 N_D_c_436_n N_VGND_c_2346_n 0.00542863f $X=1.34 $Y=0.765 $X2=0 $Y2=0
cc_421 N_A_349_21#_c_480_n N_CLK_c_564_n 0.00191349f $X=2.15 $Y=1.16 $X2=0 $Y2=0
cc_422 N_A_349_21#_c_489_n N_CLK_c_564_n 0.016878f $X=2.6 $Y=1.99 $X2=0 $Y2=0
cc_423 N_A_349_21#_c_489_n N_A_27_369#_M1022_d 0.00558673f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_424 N_A_349_21#_c_485_n N_A_27_369#_c_1858_n 0.0110384f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_425 N_A_349_21#_c_488_n N_A_27_369#_c_1858_n 0.0146603f $X=2.577 $Y=1.927
+ $X2=0 $Y2=0
cc_426 N_A_349_21#_c_489_n N_A_27_369#_c_1858_n 0.0132953f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_427 N_A_349_21#_c_485_n N_VPWR_c_1930_n 0.00429453f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_428 N_A_349_21#_c_488_n N_VPWR_c_1930_n 0.0143696f $X=2.577 $Y=1.927 $X2=0
+ $Y2=0
cc_429 N_A_349_21#_c_489_n N_VPWR_c_1930_n 0.00433681f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_430 N_A_349_21#_M1011_s N_VPWR_c_1907_n 0.00425811f $X=2.475 $Y=1.845 $X2=0
+ $Y2=0
cc_431 N_A_349_21#_c_485_n N_VPWR_c_1907_n 0.00736445f $X=1.845 $Y=1.77 $X2=0
+ $Y2=0
cc_432 N_A_349_21#_c_488_n N_VPWR_c_1907_n 0.00808388f $X=2.577 $Y=1.927 $X2=0
+ $Y2=0
cc_433 N_A_349_21#_c_489_n N_VPWR_c_1907_n 0.00699177f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_434 N_A_349_21#_M1000_g N_A_199_47#_c_2154_n 0.00877574f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_435 N_A_349_21#_c_483_n N_A_199_47#_c_2154_n 4.62381e-19 $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_436 N_A_349_21#_c_485_n N_A_199_47#_c_2157_n 0.00499317f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_437 N_A_349_21#_c_489_n N_A_199_47#_c_2157_n 0.0139951f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_438 N_A_349_21#_c_480_n N_A_199_47#_c_2149_n 0.0184928f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_439 N_A_349_21#_c_481_n N_A_199_47#_c_2149_n 0.00172463f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_440 N_A_349_21#_c_489_n N_A_199_47#_c_2149_n 0.0129846f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_441 N_A_349_21#_c_484_n N_A_199_47#_c_2150_n 0.00546081f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_442 N_A_349_21#_c_480_n N_A_199_47#_c_2150_n 0.00296292f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_443 N_A_349_21#_M1000_g N_A_199_47#_c_2145_n 0.0112054f $X=1.82 $Y=0.445
+ $X2=0 $Y2=0
cc_444 N_A_349_21#_c_484_n N_A_199_47#_c_2145_n 0.0072174f $X=1.845 $Y=1.67
+ $X2=0 $Y2=0
cc_445 N_A_349_21#_c_485_n N_A_199_47#_c_2145_n 0.00500146f $X=1.845 $Y=1.77
+ $X2=0 $Y2=0
cc_446 N_A_349_21#_c_480_n N_A_199_47#_c_2145_n 0.0488018f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_447 N_A_349_21#_c_481_n N_A_199_47#_c_2145_n 0.00926658f $X=2.15 $Y=1.16
+ $X2=0 $Y2=0
cc_448 N_A_349_21#_c_482_n N_A_199_47#_c_2145_n 0.0125538f $X=2.587 $Y=0.715
+ $X2=0 $Y2=0
cc_449 N_A_349_21#_c_483_n N_A_199_47#_c_2145_n 0.00436191f $X=2.63 $Y=0.44
+ $X2=0 $Y2=0
cc_450 N_A_349_21#_c_489_n N_A_199_47#_c_2145_n 0.00653816f $X=2.6 $Y=1.99 $X2=0
+ $Y2=0
cc_451 N_A_349_21#_M1000_g N_VGND_c_2319_n 0.0107253f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_452 N_A_349_21#_c_481_n N_VGND_c_2319_n 0.00128608f $X=2.15 $Y=1.16 $X2=0
+ $Y2=0
cc_453 N_A_349_21#_c_482_n N_VGND_c_2319_n 0.010779f $X=2.587 $Y=0.715 $X2=0
+ $Y2=0
cc_454 N_A_349_21#_c_483_n N_VGND_c_2319_n 0.0166351f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_455 N_A_349_21#_c_482_n N_VGND_c_2320_n 0.00401857f $X=2.587 $Y=0.715 $X2=0
+ $Y2=0
cc_456 N_A_349_21#_c_483_n N_VGND_c_2320_n 0.0173505f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_457 N_A_349_21#_M1000_g N_VGND_c_2336_n 0.00437031f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_458 N_A_349_21#_M1004_s N_VGND_c_2346_n 0.00468725f $X=2.505 $Y=0.235 $X2=0
+ $Y2=0
cc_459 N_A_349_21#_M1000_g N_VGND_c_2346_n 0.00852325f $X=1.82 $Y=0.445 $X2=0
+ $Y2=0
cc_460 N_A_349_21#_c_482_n N_VGND_c_2346_n 0.00745898f $X=2.587 $Y=0.715 $X2=0
+ $Y2=0
cc_461 N_A_349_21#_c_483_n N_VGND_c_2346_n 0.00964668f $X=2.63 $Y=0.44 $X2=0
+ $Y2=0
cc_462 N_CLK_c_560_n N_A_693_369#_c_644_n 0.00590278f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_463 N_CLK_c_561_n N_A_693_369#_c_644_n 0.00655864f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_464 N_CLK_c_558_n N_A_693_369#_c_644_n 2.4441e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_465 N_CLK_c_561_n N_A_693_369#_c_645_n 0.022554f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_466 N_CLK_c_555_n N_A_693_369#_c_627_n 0.00982747f $X=3.88 $Y=0.73 $X2=0
+ $Y2=0
cc_467 N_CLK_c_556_n N_A_693_369#_c_631_n 0.00982747f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_468 N_CLK_c_561_n N_A_693_369#_c_661_n 0.00657215f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_469 N_CLK_c_558_n N_A_693_369#_c_661_n 0.0011771f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_470 N_CLK_c_555_n N_A_693_369#_c_632_n 0.00564782f $X=3.88 $Y=0.73 $X2=0
+ $Y2=0
cc_471 N_CLK_c_561_n N_A_693_369#_c_649_n 0.0171228f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_472 N_CLK_c_558_n N_A_693_369#_c_649_n 0.00788865f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_473 N_CLK_c_561_n N_A_693_369#_c_650_n 3.33569e-19 $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_474 N_CLK_c_557_n N_A_693_369#_c_650_n 6.2151e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_475 N_CLK_c_558_n N_A_693_369#_c_650_n 0.0277101f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_476 N_CLK_c_555_n N_A_693_369#_c_633_n 0.00405994f $X=3.88 $Y=0.73 $X2=0
+ $Y2=0
cc_477 N_CLK_c_556_n N_A_693_369#_c_633_n 0.00866962f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_478 N_CLK_c_558_n N_A_693_369#_c_633_n 0.00798345f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_479 N_CLK_c_559_n N_A_693_369#_c_633_n 0.00151349f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_480 N_CLK_c_556_n N_A_693_369#_c_634_n 0.00402268f $X=3.88 $Y=0.805 $X2=0
+ $Y2=0
cc_481 N_CLK_c_557_n N_A_693_369#_c_634_n 8.52949e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_482 N_CLK_c_558_n N_A_693_369#_c_634_n 0.0161366f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_483 N_CLK_c_559_n N_A_693_369#_c_634_n 5.59955e-19 $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_484 N_CLK_c_560_n N_A_693_369#_c_635_n 6.001e-19 $X=3.795 $Y=1.62 $X2=0 $Y2=0
cc_485 N_CLK_c_561_n N_A_693_369#_c_635_n 0.00368077f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_486 N_CLK_c_558_n N_A_693_369#_c_635_n 0.0341939f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_487 N_CLK_c_559_n N_A_693_369#_c_635_n 0.00565736f $X=3.68 $Y=1.09 $X2=0
+ $Y2=0
cc_488 N_CLK_c_557_n N_A_693_369#_c_636_n 0.0164171f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_489 N_CLK_c_558_n N_A_693_369#_c_636_n 3.92042e-19 $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_490 N_CLK_c_561_n N_A_693_369#_c_657_n 4.94593e-19 $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_491 N_CLK_c_559_n N_A_693_369#_c_642_n 0.0047227f $X=3.68 $Y=1.09 $X2=0 $Y2=0
cc_492 N_CLK_c_558_n N_VPWR_M1011_d 7.09937e-19 $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_493 N_CLK_c_564_n N_VPWR_M1011_d 0.00208896f $X=3.155 $Y=1.845 $X2=0 $Y2=0
cc_494 N_CLK_c_561_n N_VPWR_c_1909_n 0.00416373f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_495 N_CLK_c_558_n N_VPWR_c_1909_n 0.0107374f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_496 N_CLK_c_564_n N_VPWR_c_1909_n 0.0134722f $X=3.155 $Y=1.845 $X2=0 $Y2=0
cc_497 N_CLK_c_561_n N_VPWR_c_1910_n 0.00429282f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_498 N_CLK_c_558_n N_VPWR_c_1910_n 8.87093e-19 $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_499 N_CLK_c_564_n N_VPWR_c_1930_n 0.00101383f $X=3.155 $Y=1.845 $X2=0 $Y2=0
cc_500 N_CLK_c_561_n N_VPWR_c_1936_n 0.011012f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_501 N_CLK_c_561_n N_VPWR_c_1907_n 0.00532542f $X=3.795 $Y=1.77 $X2=0 $Y2=0
cc_502 N_CLK_c_558_n N_VPWR_c_1907_n 0.00207708f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_503 N_CLK_c_564_n N_VPWR_c_1907_n 0.00265567f $X=3.155 $Y=1.845 $X2=0 $Y2=0
cc_504 N_CLK_c_560_n N_A_199_47#_c_2149_n 0.00255456f $X=3.795 $Y=1.62 $X2=0
+ $Y2=0
cc_505 N_CLK_c_561_n N_A_199_47#_c_2149_n 0.00327618f $X=3.795 $Y=1.77 $X2=0
+ $Y2=0
cc_506 N_CLK_c_558_n N_A_199_47#_c_2149_n 0.0462271f $X=3.68 $Y=1.255 $X2=0
+ $Y2=0
cc_507 N_CLK_c_564_n N_A_199_47#_c_2149_n 0.0124022f $X=3.155 $Y=1.845 $X2=0
+ $Y2=0
cc_508 N_CLK_c_555_n N_VGND_c_2321_n 0.0019914f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_509 N_CLK_c_558_n N_VGND_c_2321_n 0.00531942f $X=3.68 $Y=1.255 $X2=0 $Y2=0
cc_510 N_CLK_c_555_n N_VGND_c_2322_n 0.00794414f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_511 N_CLK_c_555_n N_VGND_c_2330_n 0.00362954f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_512 N_CLK_c_556_n N_VGND_c_2330_n 4.55781e-19 $X=3.88 $Y=0.805 $X2=0 $Y2=0
cc_513 N_CLK_c_555_n N_VGND_c_2346_n 0.00567184f $X=3.88 $Y=0.73 $X2=0 $Y2=0
cc_514 N_A_693_369#_c_656_n N_A_877_369#_M1027_d 0.00109658f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_515 N_A_693_369#_c_657_n N_A_877_369#_M1027_d 6.85484e-19 $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_516 N_A_693_369#_c_644_n N_A_877_369#_c_930_n 0.00686143f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_517 N_A_693_369#_c_645_n N_A_877_369#_c_930_n 0.00519819f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_518 N_A_693_369#_c_646_n N_A_877_369#_c_930_n 0.00286715f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_519 N_A_693_369#_c_656_n N_A_877_369#_c_930_n 0.00108936f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_520 N_A_693_369#_c_646_n N_A_877_369#_c_920_n 0.0103538f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_521 N_A_693_369#_c_656_n N_A_877_369#_c_920_n 5.38573e-19 $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_522 N_A_693_369#_c_660_n N_A_877_369#_c_920_n 2.56925e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_523 N_A_693_369#_c_646_n N_A_877_369#_c_931_n 0.00899979f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_524 N_A_693_369#_c_656_n N_A_877_369#_c_931_n 0.00501369f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_525 N_A_693_369#_c_659_n N_A_877_369#_c_931_n 7.59275e-19 $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_526 N_A_693_369#_c_660_n N_A_877_369#_c_931_n 6.19475e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_527 N_A_693_369#_c_656_n N_A_877_369#_c_932_n 0.00170021f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_528 N_A_693_369#_c_646_n N_A_877_369#_c_933_n 0.0111876f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_529 N_A_693_369#_c_629_n N_A_877_369#_M1024_g 0.0157045f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_530 N_A_693_369#_c_647_n N_A_877_369#_M1005_g 0.00875009f $X=8.585 $Y=1.47
+ $X2=0 $Y2=0
cc_531 N_A_693_369#_c_648_n N_A_877_369#_M1005_g 0.00538907f $X=8.585 $Y=1.57
+ $X2=0 $Y2=0
cc_532 N_A_693_369#_M1045_g N_A_877_369#_M1005_g 0.0162509f $X=9.81 $Y=0.445
+ $X2=0 $Y2=0
cc_533 N_A_693_369#_c_637_n N_A_877_369#_M1005_g 0.00561652f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_534 N_A_693_369#_c_638_n N_A_877_369#_M1005_g 0.0214546f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_535 N_A_693_369#_c_639_n N_A_877_369#_M1005_g 0.0169448f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_536 N_A_693_369#_c_641_n N_A_877_369#_M1005_g 0.00134438f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_537 N_A_693_369#_c_655_n N_A_877_369#_M1005_g 0.00176342f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_538 N_A_693_369#_c_643_n N_A_877_369#_M1005_g 0.00987946f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_539 N_A_693_369#_c_648_n N_A_877_369#_c_935_n 0.0205398f $X=8.585 $Y=1.57
+ $X2=0 $Y2=0
cc_540 N_A_693_369#_c_639_n N_A_877_369#_c_935_n 0.00137216f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_541 N_A_693_369#_c_655_n N_A_877_369#_c_935_n 0.00201823f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_542 N_A_693_369#_c_656_n N_A_877_369#_c_936_n 0.00228522f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_543 N_A_693_369#_c_644_n N_A_877_369#_c_937_n 0.00327724f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_544 N_A_693_369#_c_645_n N_A_877_369#_c_937_n 0.00734806f $X=4.295 $Y=1.77
+ $X2=0 $Y2=0
cc_545 N_A_693_369#_c_726_p N_A_877_369#_c_937_n 0.00919493f $X=4.165 $Y=1.775
+ $X2=0 $Y2=0
cc_546 N_A_693_369#_c_656_n N_A_877_369#_c_937_n 0.0194314f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_547 N_A_693_369#_c_657_n N_A_877_369#_c_937_n 0.0036187f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_548 N_A_693_369#_c_628_n N_A_877_369#_c_976_n 0.00114551f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_549 N_A_693_369#_c_628_n N_A_877_369#_c_923_n 0.00138193f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_550 N_A_693_369#_c_637_n N_A_877_369#_c_923_n 0.0210866f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_551 N_A_693_369#_c_638_n N_A_877_369#_c_923_n 0.00420192f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_552 N_A_693_369#_c_639_n N_A_877_369#_c_923_n 0.0147683f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_553 N_A_693_369#_c_655_n N_A_877_369#_c_923_n 0.00223864f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_554 N_A_693_369#_c_656_n N_A_877_369#_c_923_n 0.0141918f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_555 N_A_693_369#_c_658_n N_A_877_369#_c_923_n 0.0621551f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_556 N_A_693_369#_c_659_n N_A_877_369#_c_923_n 0.0147709f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_557 N_A_693_369#_c_660_n N_A_877_369#_c_923_n 8.31647e-19 $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_558 N_A_693_369#_c_628_n N_A_877_369#_c_924_n 0.00178278f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_559 N_A_693_369#_c_635_n N_A_877_369#_c_924_n 0.00153409f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_560 N_A_693_369#_c_628_n N_A_877_369#_c_925_n 0.00171814f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_561 N_A_693_369#_c_636_n N_A_877_369#_c_925_n 0.00327724f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_562 N_A_693_369#_c_637_n N_A_877_369#_c_926_n 0.00195297f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_563 N_A_693_369#_c_638_n N_A_877_369#_c_926_n 4.54037e-19 $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_564 N_A_693_369#_c_639_n N_A_877_369#_c_926_n 0.00503543f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_565 N_A_693_369#_c_641_n N_A_877_369#_c_926_n 0.00565473f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_566 N_A_693_369#_c_643_n N_A_877_369#_c_926_n 0.00358039f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_567 N_A_693_369#_c_647_n N_A_877_369#_c_927_n 3.23748e-19 $X=8.585 $Y=1.47
+ $X2=0 $Y2=0
cc_568 N_A_693_369#_c_648_n N_A_877_369#_c_927_n 8.17584e-19 $X=8.585 $Y=1.57
+ $X2=0 $Y2=0
cc_569 N_A_693_369#_c_637_n N_A_877_369#_c_927_n 0.0136833f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_570 N_A_693_369#_c_638_n N_A_877_369#_c_927_n 8.6434e-19 $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_571 N_A_693_369#_c_639_n N_A_877_369#_c_927_n 0.0176397f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_572 N_A_693_369#_c_641_n N_A_877_369#_c_927_n 0.00858102f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_573 N_A_693_369#_c_655_n N_A_877_369#_c_927_n 0.0180481f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_574 N_A_693_369#_c_643_n N_A_877_369#_c_927_n 0.00131619f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_575 N_A_693_369#_c_628_n N_A_877_369#_c_928_n 0.0525427f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_576 N_A_693_369#_c_635_n N_A_877_369#_c_928_n 2.98087e-19 $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_577 N_A_693_369#_c_636_n N_A_877_369#_c_928_n 0.0187786f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_578 N_A_693_369#_c_627_n N_A_877_369#_c_929_n 0.00444102f $X=4.32 $Y=0.73
+ $X2=0 $Y2=0
cc_579 N_A_693_369#_c_628_n N_A_877_369#_c_929_n 0.0134963f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_580 N_A_693_369#_c_633_n N_A_877_369#_c_929_n 0.010534f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_581 N_A_693_369#_c_635_n N_A_877_369#_c_929_n 0.0523483f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_582 N_A_693_369#_c_642_n N_A_877_369#_c_929_n 0.00327724f $X=4.235 $Y=1.09
+ $X2=0 $Y2=0
cc_583 N_A_693_369#_c_646_n N_A_1219_21#_c_1110_n 0.0334006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_584 N_A_693_369#_c_658_n N_A_1219_21#_c_1110_n 0.00835454f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_585 N_A_693_369#_c_658_n N_A_1219_21#_c_1111_n 0.0111901f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_586 N_A_693_369#_c_655_n N_A_1219_21#_c_1112_n 6.46547e-19 $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_587 N_A_693_369#_c_658_n N_A_1219_21#_c_1112_n 0.0274448f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_588 N_A_693_369#_c_658_n N_A_1219_21#_c_1113_n 0.0032337f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_589 N_A_693_369#_c_658_n N_A_1075_413#_c_1210_n 0.00369378f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_590 N_A_693_369#_c_658_n N_A_1075_413#_c_1211_n 7.16017e-19 $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_591 N_A_693_369#_c_647_n N_A_1075_413#_c_1212_n 0.00764195f $X=8.585 $Y=1.47
+ $X2=0 $Y2=0
cc_592 N_A_693_369#_c_637_n N_A_1075_413#_c_1212_n 0.00114063f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_593 N_A_693_369#_c_648_n N_A_1075_413#_c_1213_n 0.067034f $X=8.585 $Y=1.57
+ $X2=0 $Y2=0
cc_594 N_A_693_369#_c_655_n N_A_1075_413#_c_1213_n 0.0211451f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_595 N_A_693_369#_c_776_p N_A_1075_413#_c_1213_n 0.00160461f $X=8.29 $Y=1.87
+ $X2=0 $Y2=0
cc_596 N_A_693_369#_c_628_n N_A_1075_413#_c_1201_n 0.00479017f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_597 N_A_693_369#_c_629_n N_A_1075_413#_c_1201_n 0.00694463f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_598 N_A_693_369#_c_646_n N_A_1075_413#_c_1230_n 0.0154392f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_599 N_A_693_369#_c_656_n N_A_1075_413#_c_1230_n 0.00374204f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_600 N_A_693_369#_c_658_n N_A_1075_413#_c_1230_n 0.00492445f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_601 N_A_693_369#_c_659_n N_A_1075_413#_c_1230_n 0.00557824f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_602 N_A_693_369#_c_660_n N_A_1075_413#_c_1230_n 0.013294f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_603 N_A_693_369#_c_646_n N_A_1075_413#_c_1214_n 0.00612006f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_604 N_A_693_369#_c_658_n N_A_1075_413#_c_1214_n 0.0152429f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_605 N_A_693_369#_c_659_n N_A_1075_413#_c_1214_n 0.00314702f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_606 N_A_693_369#_c_660_n N_A_1075_413#_c_1214_n 0.0267088f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_607 N_A_693_369#_c_646_n N_A_1075_413#_c_1202_n 0.00314884f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_608 N_A_693_369#_c_656_n N_A_1075_413#_c_1202_n 0.00396196f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_609 N_A_693_369#_c_658_n N_A_1075_413#_c_1202_n 0.00354029f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_610 N_A_693_369#_c_659_n N_A_1075_413#_c_1202_n 0.00343992f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_611 N_A_693_369#_c_660_n N_A_1075_413#_c_1202_n 0.0183007f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_612 N_A_693_369#_c_658_n N_A_1075_413#_c_1203_n 0.00831647f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_613 N_A_693_369#_c_637_n N_A_1075_413#_c_1205_n 0.0260852f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_614 N_A_693_369#_c_638_n N_A_1075_413#_c_1205_n 0.00195155f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_615 N_A_693_369#_c_655_n N_A_1075_413#_c_1205_n 0.0268779f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_616 N_A_693_369#_c_637_n N_A_1075_413#_c_1206_n 3.90905e-19 $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_617 N_A_693_369#_c_638_n N_A_1075_413#_c_1206_n 0.0212873f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_618 N_A_693_369#_c_655_n N_A_1075_413#_c_1206_n 0.00268124f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_619 N_A_693_369#_c_655_n N_A_1075_413#_c_1207_n 0.00210703f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_620 N_A_693_369#_c_658_n N_A_1075_413#_c_1207_n 0.00302221f $X=8.145 $Y=1.87
+ $X2=0 $Y2=0
cc_621 N_A_693_369#_c_637_n N_A_1075_413#_c_1209_n 0.00268604f $X=8.62 $Y=1.16
+ $X2=0 $Y2=0
cc_622 N_A_693_369#_c_640_n N_A_1075_413#_c_1209_n 0.00746519f $X=8.755 $Y=0.795
+ $X2=0 $Y2=0
cc_623 N_A_693_369#_c_655_n N_SET_B_c_1360_n 8.88943e-19 $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_624 N_A_693_369#_c_655_n N_SET_B_c_1361_n 0.00342541f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_625 N_A_693_369#_c_658_n N_SET_B_c_1361_n 0.0105854f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_626 N_A_693_369#_c_647_n N_SET_B_c_1368_n 5.5681e-19 $X=8.585 $Y=1.47 $X2=0
+ $Y2=0
cc_627 N_A_693_369#_c_637_n N_SET_B_c_1368_n 0.00574163f $X=8.62 $Y=1.16 $X2=0
+ $Y2=0
cc_628 N_A_693_369#_c_638_n N_SET_B_c_1368_n 7.93137e-19 $X=8.62 $Y=1.16 $X2=0
+ $Y2=0
cc_629 N_A_693_369#_c_639_n N_SET_B_c_1368_n 0.00555644f $X=9.61 $Y=0.795 $X2=0
+ $Y2=0
cc_630 N_A_693_369#_c_641_n N_SET_B_c_1368_n 0.00193527f $X=9.7 $Y=1.08 $X2=0
+ $Y2=0
cc_631 N_A_693_369#_c_655_n N_SET_B_c_1368_n 0.0317941f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_632 N_A_693_369#_c_658_n N_SET_B_c_1368_n 0.0327067f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_633 N_A_693_369#_c_776_p N_SET_B_c_1368_n 0.0249445f $X=8.29 $Y=1.87 $X2=0
+ $Y2=0
cc_634 N_A_693_369#_c_643_n N_SET_B_c_1368_n 0.00119869f $X=9.81 $Y=1.08 $X2=0
+ $Y2=0
cc_635 N_A_693_369#_c_655_n N_SET_B_c_1369_n 0.0013569f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_636 N_A_693_369#_c_658_n N_SET_B_c_1369_n 0.0305426f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_637 N_A_693_369#_c_641_n N_SET_B_c_1370_n 0.00198942f $X=9.7 $Y=1.08 $X2=0
+ $Y2=0
cc_638 N_A_693_369#_c_641_n N_SET_B_c_1371_n 0.0141719f $X=9.7 $Y=1.08 $X2=0
+ $Y2=0
cc_639 N_A_693_369#_c_643_n N_SET_B_c_1371_n 5.26002e-19 $X=9.81 $Y=1.08 $X2=0
+ $Y2=0
cc_640 N_A_693_369#_c_655_n N_SET_B_c_1372_n 0.0202323f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_641 N_A_693_369#_c_658_n N_SET_B_c_1372_n 0.0116927f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_642 N_A_693_369#_c_641_n N_A_1930_295#_c_1513_n 3.58483e-19 $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_643 N_A_693_369#_c_643_n N_A_1930_295#_c_1513_n 0.0137905f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_644 N_A_693_369#_M1045_g N_A_1930_295#_M1039_g 0.03639f $X=9.81 $Y=0.445
+ $X2=0 $Y2=0
cc_645 N_A_693_369#_c_639_n N_A_1930_295#_M1039_g 0.00438668f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_646 N_A_693_369#_M1045_g N_A_1930_295#_c_1505_n 3.88967e-19 $X=9.81 $Y=0.445
+ $X2=0 $Y2=0
cc_647 N_A_693_369#_c_639_n N_A_1930_295#_c_1505_n 0.00246646f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_648 N_A_693_369#_c_641_n N_A_1930_295#_c_1505_n 0.0164774f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_649 N_A_693_369#_c_641_n N_A_1930_295#_c_1506_n 0.00211855f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_650 N_A_693_369#_c_643_n N_A_1930_295#_c_1506_n 0.03639f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_651 N_A_693_369#_c_641_n N_A_1930_295#_c_1516_n 0.00368955f $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_652 N_A_693_369#_c_639_n N_A_1735_329#_M1005_d 0.00390782f $X=9.61 $Y=0.795
+ $X2=-0.19 $Y2=-0.24
cc_653 N_A_693_369#_c_655_n N_A_1735_329#_M1012_d 0.00467074f $X=8.535 $Y=1.725
+ $X2=0 $Y2=0
cc_654 N_A_693_369#_c_648_n N_A_1735_329#_c_1640_n 0.00139431f $X=8.585 $Y=1.57
+ $X2=0 $Y2=0
cc_655 N_A_693_369#_M1045_g N_A_1735_329#_c_1641_n 0.0109876f $X=9.81 $Y=0.445
+ $X2=0 $Y2=0
cc_656 N_A_693_369#_c_639_n N_A_1735_329#_c_1641_n 0.0328142f $X=9.61 $Y=0.795
+ $X2=0 $Y2=0
cc_657 N_A_693_369#_c_643_n N_A_1735_329#_c_1641_n 5.24431e-19 $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_658 N_A_693_369#_c_641_n N_A_1735_329#_c_1637_n 8.42276e-19 $X=9.7 $Y=1.08
+ $X2=0 $Y2=0
cc_659 N_A_693_369#_c_643_n N_A_1735_329#_c_1637_n 0.00144539f $X=9.81 $Y=1.08
+ $X2=0 $Y2=0
cc_660 N_A_693_369#_c_649_n N_VPWR_M1044_d 8.59632e-19 $X=4.035 $Y=1.865 $X2=0
+ $Y2=0
cc_661 N_A_693_369#_c_726_p N_VPWR_M1044_d 0.00112408f $X=4.165 $Y=1.775 $X2=0
+ $Y2=0
cc_662 N_A_693_369#_c_657_n N_VPWR_M1044_d 0.00140392f $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_663 N_A_693_369#_c_655_n N_VPWR_M1023_d 0.00543586f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_664 N_A_693_369#_c_658_n N_VPWR_M1023_d 0.00122696f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_665 N_A_693_369#_c_661_n N_VPWR_c_1909_n 0.0118222f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_666 N_A_693_369#_c_661_n N_VPWR_c_1910_n 0.00607628f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_667 N_A_693_369#_c_658_n N_VPWR_c_1911_n 0.00119067f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_668 N_A_693_369#_c_776_p N_VPWR_c_1912_n 0.00339415f $X=8.29 $Y=1.87 $X2=0
+ $Y2=0
cc_669 N_A_693_369#_c_655_n N_VPWR_c_1913_n 0.0333891f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_670 N_A_693_369#_c_658_n N_VPWR_c_1913_n 0.00918422f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_671 N_A_693_369#_c_645_n N_VPWR_c_1931_n 0.0062441f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_672 N_A_693_369#_c_646_n N_VPWR_c_1931_n 0.00429453f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_673 N_A_693_369#_c_645_n N_VPWR_c_1936_n 0.00817812f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_674 N_A_693_369#_c_661_n N_VPWR_c_1936_n 0.00373276f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_675 N_A_693_369#_c_649_n N_VPWR_c_1936_n 0.00556421f $X=4.035 $Y=1.865 $X2=0
+ $Y2=0
cc_676 N_A_693_369#_c_726_p N_VPWR_c_1936_n 0.005601f $X=4.165 $Y=1.775 $X2=0
+ $Y2=0
cc_677 N_A_693_369#_c_657_n N_VPWR_c_1936_n 0.00180068f $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_678 N_A_693_369#_c_648_n N_VPWR_c_1938_n 0.0230452f $X=8.585 $Y=1.57 $X2=0
+ $Y2=0
cc_679 N_A_693_369#_c_655_n N_VPWR_c_1938_n 0.0110409f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_680 N_A_693_369#_M1044_s N_VPWR_c_1907_n 0.00405031f $X=3.465 $Y=1.845 $X2=0
+ $Y2=0
cc_681 N_A_693_369#_c_645_n N_VPWR_c_1907_n 0.0065951f $X=4.295 $Y=1.77 $X2=0
+ $Y2=0
cc_682 N_A_693_369#_c_646_n N_VPWR_c_1907_n 0.00620168f $X=5.755 $Y=1.99 $X2=0
+ $Y2=0
cc_683 N_A_693_369#_c_661_n N_VPWR_c_1907_n 0.00593257f $X=3.59 $Y=2.16 $X2=0
+ $Y2=0
cc_684 N_A_693_369#_c_649_n N_VPWR_c_1907_n 0.00631759f $X=4.035 $Y=1.865 $X2=0
+ $Y2=0
cc_685 N_A_693_369#_c_726_p N_VPWR_c_1907_n 0.00130914f $X=4.165 $Y=1.775 $X2=0
+ $Y2=0
cc_686 N_A_693_369#_c_655_n N_VPWR_c_1907_n 0.00372941f $X=8.535 $Y=1.725 $X2=0
+ $Y2=0
cc_687 N_A_693_369#_c_656_n N_VPWR_c_1907_n 0.0554324f $X=5.545 $Y=1.87 $X2=0
+ $Y2=0
cc_688 N_A_693_369#_c_657_n N_VPWR_c_1907_n 0.0177757f $X=4.405 $Y=1.87 $X2=0
+ $Y2=0
cc_689 N_A_693_369#_c_658_n N_VPWR_c_1907_n 0.103409f $X=8.145 $Y=1.87 $X2=0
+ $Y2=0
cc_690 N_A_693_369#_c_659_n N_VPWR_c_1907_n 0.018311f $X=5.885 $Y=1.87 $X2=0
+ $Y2=0
cc_691 N_A_693_369#_c_776_p N_VPWR_c_1907_n 0.0143696f $X=8.29 $Y=1.87 $X2=0
+ $Y2=0
cc_692 N_A_693_369#_c_628_n N_A_199_47#_c_2143_n 0.0087293f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_693 N_A_693_369#_c_629_n N_A_199_47#_c_2143_n 0.00393123f $X=5.34 $Y=0.73
+ $X2=0 $Y2=0
cc_694 N_A_693_369#_c_646_n N_A_199_47#_c_2148_n 3.68983e-19 $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_695 N_A_693_369#_c_656_n N_A_199_47#_c_2148_n 0.0165286f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_696 N_A_693_369#_c_659_n N_A_199_47#_c_2148_n 0.00274637f $X=5.885 $Y=1.87
+ $X2=0 $Y2=0
cc_697 N_A_693_369#_c_628_n N_A_199_47#_c_2144_n 0.00917259f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_698 N_A_693_369#_c_644_n N_A_199_47#_c_2149_n 0.00641873f $X=4.295 $Y=1.67
+ $X2=0 $Y2=0
cc_699 N_A_693_369#_c_628_n N_A_199_47#_c_2149_n 0.0024753f $X=5.265 $Y=0.805
+ $X2=0 $Y2=0
cc_700 N_A_693_369#_c_649_n N_A_199_47#_c_2149_n 0.012588f $X=4.035 $Y=1.865
+ $X2=0 $Y2=0
cc_701 N_A_693_369#_c_650_n N_A_199_47#_c_2149_n 0.00440477f $X=3.675 $Y=1.865
+ $X2=0 $Y2=0
cc_702 N_A_693_369#_c_633_n N_A_199_47#_c_2149_n 0.00714467f $X=4.035 $Y=0.8
+ $X2=0 $Y2=0
cc_703 N_A_693_369#_c_634_n N_A_199_47#_c_2149_n 7.06126e-19 $X=3.705 $Y=0.8
+ $X2=0 $Y2=0
cc_704 N_A_693_369#_c_635_n N_A_199_47#_c_2149_n 0.0226415f $X=4.21 $Y=1.255
+ $X2=0 $Y2=0
cc_705 N_A_693_369#_c_656_n N_A_199_47#_c_2149_n 0.0426897f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_706 N_A_693_369#_c_657_n N_A_199_47#_c_2149_n 0.030156f $X=4.405 $Y=1.87
+ $X2=0 $Y2=0
cc_707 N_A_693_369#_c_646_n N_A_199_47#_c_2152_n 0.00118188f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_708 N_A_693_369#_c_656_n N_A_199_47#_c_2152_n 0.0256821f $X=5.545 $Y=1.87
+ $X2=0 $Y2=0
cc_709 N_A_693_369#_c_660_n N_A_199_47#_c_2152_n 0.00187515f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_710 N_A_693_369#_c_646_n N_A_199_47#_c_2146_n 0.00245294f $X=5.755 $Y=1.99
+ $X2=0 $Y2=0
cc_711 N_A_693_369#_c_660_n N_A_199_47#_c_2146_n 0.0103393f $X=5.73 $Y=1.74
+ $X2=0 $Y2=0
cc_712 N_A_693_369#_c_655_n A_1652_329# 5.60832e-19 $X=8.535 $Y=1.725 $X2=-0.19
+ $Y2=-0.24
cc_713 N_A_693_369#_c_776_p A_1652_329# 0.00169225f $X=8.29 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_714 N_A_693_369#_c_632_n N_VGND_c_2321_n 0.0184201f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_715 N_A_693_369#_c_627_n N_VGND_c_2322_n 0.00315208f $X=4.32 $Y=0.73 $X2=0
+ $Y2=0
cc_716 N_A_693_369#_c_632_n N_VGND_c_2322_n 0.017284f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_717 N_A_693_369#_c_633_n N_VGND_c_2322_n 0.0211484f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_718 N_A_693_369#_c_636_n N_VGND_c_2322_n 5.1204e-19 $X=4.21 $Y=1.255 $X2=0
+ $Y2=0
cc_719 N_A_693_369#_c_632_n N_VGND_c_2330_n 0.0127969f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_720 N_A_693_369#_c_633_n N_VGND_c_2330_n 0.00324829f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_721 N_A_693_369#_c_627_n N_VGND_c_2337_n 0.00535706f $X=4.32 $Y=0.73 $X2=0
+ $Y2=0
cc_722 N_A_693_369#_c_628_n N_VGND_c_2337_n 0.00396629f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_723 N_A_693_369#_c_629_n N_VGND_c_2337_n 0.00564131f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_724 N_A_693_369#_c_633_n N_VGND_c_2337_n 8.32209e-19 $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_725 N_A_693_369#_M1045_g N_VGND_c_2338_n 0.00362032f $X=9.81 $Y=0.445 $X2=0
+ $Y2=0
cc_726 N_A_693_369#_c_639_n N_VGND_c_2338_n 0.00572424f $X=9.61 $Y=0.795 $X2=0
+ $Y2=0
cc_727 N_A_693_369#_c_640_n N_VGND_c_2338_n 0.00375056f $X=8.755 $Y=0.795 $X2=0
+ $Y2=0
cc_728 N_A_693_369#_M1017_s N_VGND_c_2346_n 0.00388795f $X=3.495 $Y=0.235 $X2=0
+ $Y2=0
cc_729 N_A_693_369#_c_627_n N_VGND_c_2346_n 0.0102775f $X=4.32 $Y=0.73 $X2=0
+ $Y2=0
cc_730 N_A_693_369#_c_628_n N_VGND_c_2346_n 0.00372099f $X=5.265 $Y=0.805 $X2=0
+ $Y2=0
cc_731 N_A_693_369#_c_629_n N_VGND_c_2346_n 0.0116506f $X=5.34 $Y=0.73 $X2=0
+ $Y2=0
cc_732 N_A_693_369#_M1045_g N_VGND_c_2346_n 0.00575709f $X=9.81 $Y=0.445 $X2=0
+ $Y2=0
cc_733 N_A_693_369#_c_632_n N_VGND_c_2346_n 0.00703355f $X=3.62 $Y=0.44 $X2=0
+ $Y2=0
cc_734 N_A_693_369#_c_633_n N_VGND_c_2346_n 0.00794826f $X=4.035 $Y=0.8 $X2=0
+ $Y2=0
cc_735 N_A_693_369#_c_639_n N_VGND_c_2346_n 0.0114601f $X=9.61 $Y=0.795 $X2=0
+ $Y2=0
cc_736 N_A_693_369#_c_640_n N_VGND_c_2346_n 0.00633305f $X=8.755 $Y=0.795 $X2=0
+ $Y2=0
cc_737 N_A_693_369#_c_639_n A_1655_47# 0.00430463f $X=9.61 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_738 N_A_693_369#_c_640_n A_1655_47# 0.00840217f $X=8.755 $Y=0.795 $X2=-0.19
+ $Y2=-0.24
cc_739 N_A_877_369#_M1024_g N_A_1219_21#_M1029_g 0.0611333f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_740 N_A_877_369#_M1024_g N_A_1219_21#_c_1104_n 0.00658605f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_741 N_A_877_369#_c_923_n N_A_1219_21#_c_1104_n 0.00298371f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_742 N_A_877_369#_c_923_n N_A_1219_21#_c_1111_n 5.84337e-19 $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_743 N_A_877_369#_c_923_n N_A_1219_21#_c_1105_n 0.00838091f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_744 N_A_877_369#_M1024_g N_A_1219_21#_c_1107_n 0.00123852f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_745 N_A_877_369#_c_923_n N_A_1219_21#_c_1107_n 0.0108029f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_746 N_A_877_369#_c_923_n N_A_1219_21#_c_1108_n 0.00455149f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_747 N_A_877_369#_c_920_n N_A_1075_413#_c_1201_n 0.0159502f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_748 N_A_877_369#_M1024_g N_A_1075_413#_c_1201_n 0.0218559f $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_749 N_A_877_369#_c_923_n N_A_1075_413#_c_1201_n 0.0362886f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_750 N_A_877_369#_c_920_n N_A_1075_413#_c_1202_n 0.006731f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_751 N_A_877_369#_c_923_n N_A_1075_413#_c_1202_n 0.024704f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_752 N_A_877_369#_c_928_n N_A_1075_413#_c_1202_n 3.66329e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_753 N_A_877_369#_c_923_n N_A_1075_413#_c_1203_n 0.017023f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_754 N_A_877_369#_c_923_n N_A_1075_413#_c_1204_n 0.0118734f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_755 N_A_877_369#_c_923_n N_A_1075_413#_c_1205_n 0.0197335f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_756 N_A_877_369#_c_923_n N_A_1075_413#_c_1207_n 0.0486664f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_757 N_A_877_369#_c_923_n N_A_1075_413#_c_1208_n 0.00125052f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_758 N_A_877_369#_M1005_g N_SET_B_c_1368_n 0.00159382f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_759 N_A_877_369#_c_935_n N_SET_B_c_1368_n 0.00253162f $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_760 N_A_877_369#_c_923_n N_SET_B_c_1368_n 0.110022f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_761 N_A_877_369#_c_926_n N_SET_B_c_1368_n 0.0298544f $X=9.31 $Y=1.19 $X2=0
+ $Y2=0
cc_762 N_A_877_369#_c_927_n N_SET_B_c_1368_n 0.0174459f $X=9.31 $Y=1.19 $X2=0
+ $Y2=0
cc_763 N_A_877_369#_c_923_n N_SET_B_c_1369_n 0.0307796f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_764 N_A_877_369#_c_935_n N_SET_B_c_1370_n 2.51444e-19 $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_765 N_A_877_369#_c_927_n N_SET_B_c_1370_n 0.00223542f $X=9.31 $Y=1.19 $X2=0
+ $Y2=0
cc_766 N_A_877_369#_M1005_g N_SET_B_c_1371_n 3.42341e-19 $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_767 N_A_877_369#_c_935_n N_SET_B_c_1371_n 5.73214e-19 $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_768 N_A_877_369#_c_927_n N_SET_B_c_1371_n 0.0125602f $X=9.31 $Y=1.19 $X2=0
+ $Y2=0
cc_769 N_A_877_369#_c_923_n N_SET_B_c_1372_n 0.00151535f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_770 N_A_877_369#_c_935_n N_A_1930_295#_c_1511_n 0.0284781f $X=9.26 $Y=1.99
+ $X2=0 $Y2=0
cc_771 N_A_877_369#_M1005_g N_A_1930_295#_c_1513_n 0.00237322f $X=9.09 $Y=0.555
+ $X2=0 $Y2=0
cc_772 N_A_877_369#_c_935_n N_A_1930_295#_c_1513_n 0.0212602f $X=9.26 $Y=1.99
+ $X2=0 $Y2=0
cc_773 N_A_877_369#_c_927_n N_A_1930_295#_c_1513_n 0.00217613f $X=9.31 $Y=1.19
+ $X2=0 $Y2=0
cc_774 N_A_877_369#_c_926_n N_A_1930_295#_c_1504_n 0.00120279f $X=9.31 $Y=1.19
+ $X2=0 $Y2=0
cc_775 N_A_877_369#_c_935_n N_A_1735_329#_c_1640_n 0.0230466f $X=9.26 $Y=1.99
+ $X2=0 $Y2=0
cc_776 N_A_877_369#_c_927_n N_A_1735_329#_c_1640_n 0.0134287f $X=9.31 $Y=1.19
+ $X2=0 $Y2=0
cc_777 N_A_877_369#_M1005_g N_A_1735_329#_c_1641_n 0.0109504f $X=9.09 $Y=0.555
+ $X2=0 $Y2=0
cc_778 N_A_877_369#_c_935_n N_A_1735_329#_c_1637_n 0.00478932f $X=9.26 $Y=1.99
+ $X2=0 $Y2=0
cc_779 N_A_877_369#_c_927_n N_A_1735_329#_c_1637_n 7.42195e-19 $X=9.31 $Y=1.19
+ $X2=0 $Y2=0
cc_780 N_A_877_369#_c_935_n N_VPWR_c_1923_n 0.00430708f $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_781 N_A_877_369#_c_931_n N_VPWR_c_1931_n 4.12218e-19 $X=5.195 $Y=1.915 $X2=0
+ $Y2=0
cc_782 N_A_877_369#_c_932_n N_VPWR_c_1931_n 0.00197478f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_783 N_A_877_369#_c_933_n N_VPWR_c_1931_n 0.00702461f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_784 N_A_877_369#_c_936_n N_VPWR_c_1931_n 0.0240597f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_785 N_A_877_369#_c_936_n N_VPWR_c_1936_n 0.0122663f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_786 N_A_877_369#_c_935_n N_VPWR_c_1938_n 0.00165817f $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_787 N_A_877_369#_M1027_d N_VPWR_c_1907_n 0.00224652f $X=4.385 $Y=1.845 $X2=0
+ $Y2=0
cc_788 N_A_877_369#_c_932_n N_VPWR_c_1907_n 0.00145806f $X=5.04 $Y=1.915 $X2=0
+ $Y2=0
cc_789 N_A_877_369#_c_933_n N_VPWR_c_1907_n 0.00872443f $X=5.285 $Y=1.99 $X2=0
+ $Y2=0
cc_790 N_A_877_369#_c_935_n N_VPWR_c_1907_n 0.00663314f $X=9.26 $Y=1.99 $X2=0
+ $Y2=0
cc_791 N_A_877_369#_c_936_n N_VPWR_c_1907_n 0.00624504f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_792 N_A_877_369#_c_976_n N_A_199_47#_c_2143_n 0.0256938f $X=4.56 $Y=0.42
+ $X2=0 $Y2=0
cc_793 N_A_877_369#_c_930_n N_A_199_47#_c_2147_n 0.00360345f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_794 N_A_877_369#_c_937_n N_A_199_47#_c_2147_n 0.0330959f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_795 N_A_877_369#_c_923_n N_A_199_47#_c_2147_n 2.97542e-19 $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_796 N_A_877_369#_c_930_n N_A_199_47#_c_2148_n 0.0023952f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_797 N_A_877_369#_c_931_n N_A_199_47#_c_2148_n 0.00940265f $X=5.195 $Y=1.915
+ $X2=0 $Y2=0
cc_798 N_A_877_369#_c_932_n N_A_199_47#_c_2148_n 0.00350075f $X=5.04 $Y=1.915
+ $X2=0 $Y2=0
cc_799 N_A_877_369#_c_933_n N_A_199_47#_c_2148_n 0.00399253f $X=5.285 $Y=1.99
+ $X2=0 $Y2=0
cc_800 N_A_877_369#_c_936_n N_A_199_47#_c_2148_n 0.0330959f $X=4.53 $Y=2.3 $X2=0
+ $Y2=0
cc_801 N_A_877_369#_M1024_g N_A_199_47#_c_2144_n 7.40209e-19 $X=5.81 $Y=0.445
+ $X2=0 $Y2=0
cc_802 N_A_877_369#_c_923_n N_A_199_47#_c_2144_n 0.00642819f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_803 N_A_877_369#_c_928_n N_A_199_47#_c_2144_n 0.00351906f $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_804 N_A_877_369#_c_929_n N_A_199_47#_c_2144_n 0.0256938f $X=4.677 $Y=1.09
+ $X2=0 $Y2=0
cc_805 N_A_877_369#_c_930_n N_A_199_47#_c_2149_n 0.00243542f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_806 N_A_877_369#_c_937_n N_A_199_47#_c_2149_n 0.0159202f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_807 N_A_877_369#_c_923_n N_A_199_47#_c_2149_n 0.010881f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_808 N_A_877_369#_c_924_n N_A_199_47#_c_2149_n 0.025062f $X=4.815 $Y=1.19
+ $X2=0 $Y2=0
cc_809 N_A_877_369#_c_925_n N_A_199_47#_c_2149_n 0.00146838f $X=4.67 $Y=1.19
+ $X2=0 $Y2=0
cc_810 N_A_877_369#_c_928_n N_A_199_47#_c_2149_n 8.48997e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_811 N_A_877_369#_c_930_n N_A_199_47#_c_2152_n 7.80938e-19 $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_812 N_A_877_369#_c_937_n N_A_199_47#_c_2152_n 0.00216296f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_813 N_A_877_369#_c_923_n N_A_199_47#_c_2152_n 0.0260798f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_814 N_A_877_369#_c_928_n N_A_199_47#_c_2152_n 4.63662e-19 $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_815 N_A_877_369#_c_930_n N_A_199_47#_c_2146_n 0.00416664f $X=4.965 $Y=1.84
+ $X2=0 $Y2=0
cc_816 N_A_877_369#_c_920_n N_A_199_47#_c_2146_n 0.007561f $X=5.735 $Y=1.165
+ $X2=0 $Y2=0
cc_817 N_A_877_369#_c_937_n N_A_199_47#_c_2146_n 0.00868311f $X=4.617 $Y=2.135
+ $X2=0 $Y2=0
cc_818 N_A_877_369#_c_923_n N_A_199_47#_c_2146_n 0.0123027f $X=9.115 $Y=1.19
+ $X2=0 $Y2=0
cc_819 N_A_877_369#_c_924_n N_A_199_47#_c_2146_n 9.4569e-19 $X=4.815 $Y=1.19
+ $X2=0 $Y2=0
cc_820 N_A_877_369#_c_925_n N_A_199_47#_c_2146_n 0.0221582f $X=4.67 $Y=1.19
+ $X2=0 $Y2=0
cc_821 N_A_877_369#_c_928_n N_A_199_47#_c_2146_n 0.00622411f $X=5.04 $Y=1.255
+ $X2=0 $Y2=0
cc_822 N_A_877_369#_c_929_n N_A_199_47#_c_2146_n 0.00790273f $X=4.677 $Y=1.09
+ $X2=0 $Y2=0
cc_823 N_A_877_369#_M1024_g N_VGND_c_2337_n 0.00594529f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_824 N_A_877_369#_c_976_n N_VGND_c_2337_n 0.0154902f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_825 N_A_877_369#_M1005_g N_VGND_c_2338_n 0.00431327f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_826 N_A_877_369#_c_923_n N_VGND_c_2343_n 0.00453482f $X=9.115 $Y=1.19 $X2=0
+ $Y2=0
cc_827 N_A_877_369#_M1018_d N_VGND_c_2346_n 0.00458762f $X=4.395 $Y=0.235 $X2=0
+ $Y2=0
cc_828 N_A_877_369#_M1024_g N_VGND_c_2346_n 0.00523587f $X=5.81 $Y=0.445 $X2=0
+ $Y2=0
cc_829 N_A_877_369#_M1005_g N_VGND_c_2346_n 0.00799794f $X=9.09 $Y=0.555 $X2=0
+ $Y2=0
cc_830 N_A_877_369#_c_976_n N_VGND_c_2346_n 0.0085511f $X=4.56 $Y=0.42 $X2=0
+ $Y2=0
cc_831 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1210_n 0.00620188f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_832 N_A_1219_21#_c_1110_n N_A_1075_413#_c_1210_n 0.0219469f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_833 N_A_1219_21#_c_1111_n N_A_1075_413#_c_1210_n 0.00189088f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_834 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1198_n 6.33239e-19 $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_835 N_A_1219_21#_c_1110_n N_A_1075_413#_c_1211_n 0.0157421f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_836 N_A_1219_21#_c_1111_n N_A_1075_413#_c_1211_n 4.34901e-19 $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_837 N_A_1219_21#_c_1112_n N_A_1075_413#_c_1211_n 0.0157459f $X=7.1 $Y=2.02
+ $X2=0 $Y2=0
cc_838 N_A_1219_21#_c_1105_n N_A_1075_413#_c_1199_n 0.00317995f $X=6.775 $Y=0.72
+ $X2=0 $Y2=0
cc_839 N_A_1219_21#_c_1106_n N_A_1075_413#_c_1199_n 0.0095302f $X=6.95 $Y=0.51
+ $X2=0 $Y2=0
cc_840 N_A_1219_21#_M1029_g N_A_1075_413#_c_1200_n 8.20955e-19 $X=6.17 $Y=0.445
+ $X2=0 $Y2=0
cc_841 N_A_1219_21#_c_1105_n N_A_1075_413#_c_1200_n 0.0119696f $X=6.775 $Y=0.72
+ $X2=0 $Y2=0
cc_842 N_A_1219_21#_c_1107_n N_A_1075_413#_c_1200_n 0.00113481f $X=6.267 $Y=0.72
+ $X2=0 $Y2=0
cc_843 N_A_1219_21#_c_1108_n N_A_1075_413#_c_1200_n 0.0088694f $X=6.315 $Y=0.93
+ $X2=0 $Y2=0
cc_844 N_A_1219_21#_M1029_g N_A_1075_413#_c_1201_n 0.00118237f $X=6.17 $Y=0.445
+ $X2=0 $Y2=0
cc_845 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1201_n 0.00265367f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_846 N_A_1219_21#_c_1107_n N_A_1075_413#_c_1201_n 0.0313291f $X=6.267 $Y=0.72
+ $X2=0 $Y2=0
cc_847 N_A_1219_21#_c_1108_n N_A_1075_413#_c_1201_n 0.00121327f $X=6.315 $Y=0.93
+ $X2=0 $Y2=0
cc_848 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1214_n 0.0114963f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_849 N_A_1219_21#_c_1110_n N_A_1075_413#_c_1214_n 0.00116159f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_850 N_A_1219_21#_c_1111_n N_A_1075_413#_c_1214_n 0.0201747f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_851 N_A_1219_21#_c_1113_n N_A_1075_413#_c_1214_n 0.00880623f $X=6.595 $Y=2.02
+ $X2=0 $Y2=0
cc_852 N_A_1219_21#_c_1107_n N_A_1075_413#_c_1202_n 0.00784248f $X=6.267 $Y=0.72
+ $X2=0 $Y2=0
cc_853 N_A_1219_21#_c_1108_n N_A_1075_413#_c_1202_n 0.00297153f $X=6.315 $Y=0.93
+ $X2=0 $Y2=0
cc_854 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1203_n 0.0150073f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_855 N_A_1219_21#_c_1110_n N_A_1075_413#_c_1203_n 0.00260846f $X=6.315 $Y=1.99
+ $X2=0 $Y2=0
cc_856 N_A_1219_21#_c_1111_n N_A_1075_413#_c_1203_n 0.0109804f $X=6.51 $Y=1.74
+ $X2=0 $Y2=0
cc_857 N_A_1219_21#_c_1105_n N_A_1075_413#_c_1203_n 0.00671458f $X=6.775 $Y=0.72
+ $X2=0 $Y2=0
cc_858 N_A_1219_21#_c_1112_n N_A_1075_413#_c_1203_n 0.00617396f $X=7.1 $Y=2.02
+ $X2=0 $Y2=0
cc_859 N_A_1219_21#_c_1107_n N_A_1075_413#_c_1203_n 0.0134066f $X=6.267 $Y=0.72
+ $X2=0 $Y2=0
cc_860 N_A_1219_21#_c_1108_n N_A_1075_413#_c_1203_n 7.94205e-19 $X=6.315 $Y=0.93
+ $X2=0 $Y2=0
cc_861 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1204_n 0.00185156f $X=6.315
+ $Y=1.575 $X2=0 $Y2=0
cc_862 N_A_1219_21#_c_1105_n N_A_1075_413#_c_1204_n 0.0255064f $X=6.775 $Y=0.72
+ $X2=0 $Y2=0
cc_863 N_A_1219_21#_c_1107_n N_A_1075_413#_c_1204_n 0.00233448f $X=6.267 $Y=0.72
+ $X2=0 $Y2=0
cc_864 N_A_1219_21#_c_1108_n N_A_1075_413#_c_1204_n 0.00163596f $X=6.315 $Y=0.93
+ $X2=0 $Y2=0
cc_865 N_A_1219_21#_c_1112_n N_A_1075_413#_c_1207_n 0.00336414f $X=7.1 $Y=2.02
+ $X2=0 $Y2=0
cc_866 N_A_1219_21#_c_1104_n N_A_1075_413#_c_1208_n 0.0135332f $X=6.315 $Y=1.575
+ $X2=0 $Y2=0
cc_867 N_A_1219_21#_c_1105_n N_A_1075_413#_c_1208_n 0.00200711f $X=6.775 $Y=0.72
+ $X2=0 $Y2=0
cc_868 N_A_1219_21#_c_1112_n N_A_1075_413#_c_1208_n 6.59136e-19 $X=7.1 $Y=2.02
+ $X2=0 $Y2=0
cc_869 N_A_1219_21#_c_1112_n N_SET_B_c_1361_n 0.0071054f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_870 N_A_1219_21#_c_1167_p N_SET_B_c_1361_n 0.00388525f $X=7.21 $Y=2.285 $X2=0
+ $Y2=0
cc_871 N_A_1219_21#_c_1105_n N_SET_B_M1025_g 2.94061e-19 $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_872 N_A_1219_21#_c_1111_n N_SET_B_c_1372_n 0.00579563f $X=6.51 $Y=1.74 $X2=0
+ $Y2=0
cc_873 N_A_1219_21#_c_1112_n N_SET_B_c_1372_n 0.0117875f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_874 N_A_1219_21#_c_1112_n N_VPWR_M1042_d 0.00245852f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_875 N_A_1219_21#_c_1113_n N_VPWR_M1042_d 0.00153636f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_876 N_A_1219_21#_c_1110_n N_VPWR_c_1911_n 0.0054598f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_877 N_A_1219_21#_c_1112_n N_VPWR_c_1911_n 0.0125888f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_878 N_A_1219_21#_c_1113_n N_VPWR_c_1911_n 0.0102436f $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_879 N_A_1219_21#_c_1112_n N_VPWR_c_1922_n 0.00482933f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_880 N_A_1219_21#_c_1167_p N_VPWR_c_1922_n 0.0165035f $X=7.21 $Y=2.285 $X2=0
+ $Y2=0
cc_881 N_A_1219_21#_c_1110_n N_VPWR_c_1931_n 0.00743866f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_882 N_A_1219_21#_M1008_d N_VPWR_c_1907_n 0.00326382f $X=7.045 $Y=2.065 $X2=0
+ $Y2=0
cc_883 N_A_1219_21#_c_1110_n N_VPWR_c_1907_n 0.00840629f $X=6.315 $Y=1.99 $X2=0
+ $Y2=0
cc_884 N_A_1219_21#_c_1112_n N_VPWR_c_1907_n 0.0041491f $X=7.1 $Y=2.02 $X2=0
+ $Y2=0
cc_885 N_A_1219_21#_c_1113_n N_VPWR_c_1907_n 7.82982e-19 $X=6.595 $Y=2.02 $X2=0
+ $Y2=0
cc_886 N_A_1219_21#_c_1167_p N_VPWR_c_1907_n 0.0047097f $X=7.21 $Y=2.285 $X2=0
+ $Y2=0
cc_887 N_A_1219_21#_c_1105_n N_VGND_M1029_d 8.64971e-19 $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_888 N_A_1219_21#_c_1107_n N_VGND_M1029_d 0.00185499f $X=6.267 $Y=0.72 $X2=0
+ $Y2=0
cc_889 N_A_1219_21#_M1029_g N_VGND_c_2337_n 0.0134364f $X=6.17 $Y=0.445 $X2=0
+ $Y2=0
cc_890 N_A_1219_21#_c_1105_n N_VGND_c_2337_n 0.00919218f $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_891 N_A_1219_21#_c_1106_n N_VGND_c_2337_n 0.017353f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_892 N_A_1219_21#_c_1107_n N_VGND_c_2337_n 0.0252557f $X=6.267 $Y=0.72 $X2=0
+ $Y2=0
cc_893 N_A_1219_21#_c_1108_n N_VGND_c_2337_n 0.00107872f $X=6.315 $Y=0.93 $X2=0
+ $Y2=0
cc_894 N_A_1219_21#_c_1105_n N_VGND_c_2342_n 0.00328118f $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_895 N_A_1219_21#_c_1106_n N_VGND_c_2342_n 0.0213909f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_896 N_A_1219_21#_c_1105_n N_VGND_c_2343_n 0.0019843f $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_897 N_A_1219_21#_M1021_s N_VGND_c_2346_n 0.00408247f $X=6.825 $Y=0.235 $X2=0
+ $Y2=0
cc_898 N_A_1219_21#_c_1105_n N_VGND_c_2346_n 0.00566344f $X=6.775 $Y=0.72 $X2=0
+ $Y2=0
cc_899 N_A_1219_21#_c_1106_n N_VGND_c_2346_n 0.0117965f $X=6.95 $Y=0.51 $X2=0
+ $Y2=0
cc_900 N_A_1219_21#_c_1107_n N_VGND_c_2346_n 0.00191018f $X=6.267 $Y=0.72 $X2=0
+ $Y2=0
cc_901 N_A_1075_413#_c_1210_n N_SET_B_c_1360_n 0.00568643f $X=6.955 $Y=1.89
+ $X2=0 $Y2=0
cc_902 N_A_1075_413#_c_1212_n N_SET_B_c_1360_n 0.00292325f $X=8.17 $Y=1.47 $X2=0
+ $Y2=0
cc_903 N_A_1075_413#_c_1210_n N_SET_B_c_1361_n 0.0252833f $X=6.955 $Y=1.89 $X2=0
+ $Y2=0
cc_904 N_A_1075_413#_c_1211_n N_SET_B_c_1361_n 0.0110372f $X=6.955 $Y=1.99 $X2=0
+ $Y2=0
cc_905 N_A_1075_413#_c_1213_n N_SET_B_c_1361_n 0.0261173f $X=8.17 $Y=1.57 $X2=0
+ $Y2=0
cc_906 N_A_1075_413#_c_1200_n N_SET_B_c_1361_n 8.54675e-19 $X=7.26 $Y=0.805
+ $X2=0 $Y2=0
cc_907 N_A_1075_413#_c_1207_n N_SET_B_c_1361_n 8.96199e-19 $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_908 N_A_1075_413#_c_1198_n N_SET_B_M1025_g 0.00662033f $X=6.96 $Y=1.095 $X2=0
+ $Y2=0
cc_909 N_A_1075_413#_c_1199_n N_SET_B_M1025_g 0.0486803f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_910 N_A_1075_413#_c_1206_n N_SET_B_M1025_g 0.0162655f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_911 N_A_1075_413#_c_1207_n N_SET_B_M1025_g 0.0106452f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_912 N_A_1075_413#_c_1209_n N_SET_B_M1025_g 0.0208277f $X=8.115 $Y=0.995 $X2=0
+ $Y2=0
cc_913 N_A_1075_413#_c_1212_n N_SET_B_c_1359_n 0.00163967f $X=8.17 $Y=1.47 $X2=0
+ $Y2=0
cc_914 N_A_1075_413#_c_1204_n N_SET_B_c_1359_n 5.81381e-19 $X=6.935 $Y=1.185
+ $X2=0 $Y2=0
cc_915 N_A_1075_413#_c_1205_n N_SET_B_c_1359_n 0.00109872f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_916 N_A_1075_413#_c_1207_n N_SET_B_c_1359_n 0.010681f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_917 N_A_1075_413#_c_1208_n N_SET_B_c_1359_n 0.00568643f $X=6.96 $Y=1.23 $X2=0
+ $Y2=0
cc_918 N_A_1075_413#_c_1212_n N_SET_B_c_1368_n 0.00130585f $X=8.17 $Y=1.47 $X2=0
+ $Y2=0
cc_919 N_A_1075_413#_c_1213_n N_SET_B_c_1368_n 3.54738e-19 $X=8.17 $Y=1.57 $X2=0
+ $Y2=0
cc_920 N_A_1075_413#_c_1205_n N_SET_B_c_1368_n 0.00262589f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_921 N_A_1075_413#_c_1206_n N_SET_B_c_1368_n 0.0018852f $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_922 N_A_1075_413#_c_1207_n N_SET_B_c_1368_n 0.00557137f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_923 N_A_1075_413#_c_1210_n N_SET_B_c_1369_n 4.49976e-19 $X=6.955 $Y=1.89
+ $X2=0 $Y2=0
cc_924 N_A_1075_413#_c_1212_n N_SET_B_c_1369_n 6.78777e-19 $X=8.17 $Y=1.47 $X2=0
+ $Y2=0
cc_925 N_A_1075_413#_c_1207_n N_SET_B_c_1369_n 0.00199134f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_926 N_A_1075_413#_c_1210_n N_SET_B_c_1372_n 0.00585069f $X=6.955 $Y=1.89
+ $X2=0 $Y2=0
cc_927 N_A_1075_413#_c_1212_n N_SET_B_c_1372_n 7.35449e-19 $X=8.17 $Y=1.47 $X2=0
+ $Y2=0
cc_928 N_A_1075_413#_c_1213_n N_SET_B_c_1372_n 6.66787e-19 $X=8.17 $Y=1.57 $X2=0
+ $Y2=0
cc_929 N_A_1075_413#_c_1207_n N_SET_B_c_1372_n 0.0360668f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_930 N_A_1075_413#_c_1211_n N_VPWR_c_1911_n 0.00587549f $X=6.955 $Y=1.99 $X2=0
+ $Y2=0
cc_931 N_A_1075_413#_c_1213_n N_VPWR_c_1912_n 0.0265199f $X=8.17 $Y=1.57 $X2=0
+ $Y2=0
cc_932 N_A_1075_413#_c_1211_n N_VPWR_c_1922_n 0.00512994f $X=6.955 $Y=1.99 $X2=0
+ $Y2=0
cc_933 N_A_1075_413#_c_1230_n N_VPWR_c_1931_n 0.0467357f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_934 N_A_1075_413#_M1003_d N_VPWR_c_1907_n 0.00227362f $X=5.375 $Y=2.065 $X2=0
+ $Y2=0
cc_935 N_A_1075_413#_c_1211_n N_VPWR_c_1907_n 0.0071219f $X=6.955 $Y=1.99 $X2=0
+ $Y2=0
cc_936 N_A_1075_413#_c_1230_n N_VPWR_c_1907_n 0.0130771f $X=6.035 $Y=2.3 $X2=0
+ $Y2=0
cc_937 N_A_1075_413#_c_1201_n N_A_199_47#_c_2143_n 0.0618132f $X=5.55 $Y=0.42
+ $X2=0 $Y2=0
cc_938 N_A_1075_413#_c_1202_n N_A_199_47#_c_2146_n 0.00960767f $X=5.4 $Y=1.225
+ $X2=0 $Y2=0
cc_939 N_A_1075_413#_c_1230_n A_1169_413# 0.00692155f $X=6.035 $Y=2.3 $X2=-0.19
+ $Y2=-0.24
cc_940 N_A_1075_413#_c_1214_n A_1169_413# 0.00130666f $X=6.12 $Y=2.135 $X2=-0.19
+ $Y2=-0.24
cc_941 N_A_1075_413#_c_1199_n N_VGND_c_2337_n 0.00255767f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_942 N_A_1075_413#_c_1201_n N_VGND_c_2337_n 0.029789f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_943 N_A_1075_413#_c_1199_n N_VGND_c_2342_n 0.00585385f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_944 N_A_1075_413#_c_1200_n N_VGND_c_2342_n 0.00213423f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_945 N_A_1075_413#_c_1199_n N_VGND_c_2343_n 0.0035869f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_946 N_A_1075_413#_c_1206_n N_VGND_c_2343_n 9.9419e-19 $X=8.09 $Y=1.16 $X2=0
+ $Y2=0
cc_947 N_A_1075_413#_c_1207_n N_VGND_c_2343_n 0.0353368f $X=7.95 $Y=1.15 $X2=0
+ $Y2=0
cc_948 N_A_1075_413#_c_1209_n N_VGND_c_2343_n 0.0310659f $X=8.115 $Y=0.995 $X2=0
+ $Y2=0
cc_949 N_A_1075_413#_M1031_d N_VGND_c_2346_n 0.0025535f $X=5.415 $Y=0.235 $X2=0
+ $Y2=0
cc_950 N_A_1075_413#_c_1199_n N_VGND_c_2346_n 0.0120541f $X=7.26 $Y=0.73 $X2=0
+ $Y2=0
cc_951 N_A_1075_413#_c_1200_n N_VGND_c_2346_n 0.00217092f $X=7.26 $Y=0.805 $X2=0
+ $Y2=0
cc_952 N_A_1075_413#_c_1201_n N_VGND_c_2346_n 0.0178988f $X=5.55 $Y=0.42 $X2=0
+ $Y2=0
cc_953 N_A_1075_413#_c_1209_n N_VGND_c_2346_n 0.00217582f $X=8.115 $Y=0.995
+ $X2=0 $Y2=0
cc_954 N_SET_B_c_1362_n N_A_1930_295#_c_1510_n 0.0034701f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_955 N_SET_B_c_1366_n N_A_1930_295#_c_1510_n 6.19792e-19 $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_956 N_SET_B_c_1370_n N_A_1930_295#_c_1510_n 2.8888e-19 $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_957 N_SET_B_c_1371_n N_A_1930_295#_c_1510_n 0.00613246f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_958 N_SET_B_c_1362_n N_A_1930_295#_c_1511_n 0.00838032f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_959 N_SET_B_c_1366_n N_A_1930_295#_c_1512_n 0.0192625f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_960 N_SET_B_c_1367_n N_A_1930_295#_c_1512_n 0.00290311f $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_961 N_SET_B_c_1370_n N_A_1930_295#_c_1512_n 0.00214137f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_962 N_SET_B_c_1371_n N_A_1930_295#_c_1512_n 0.00565092f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_963 N_SET_B_c_1368_n N_A_1930_295#_c_1513_n 0.00133058f $X=9.675 $Y=1.53
+ $X2=0 $Y2=0
cc_964 N_SET_B_c_1370_n N_A_1930_295#_c_1513_n 2.32196e-19 $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_965 N_SET_B_c_1371_n N_A_1930_295#_c_1513_n 0.00349541f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_966 N_SET_B_M1043_g N_A_1930_295#_M1039_g 0.0093392f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_967 N_SET_B_M1043_g N_A_1930_295#_c_1504_n 0.00473733f $X=10.96 $Y=0.445
+ $X2=0 $Y2=0
cc_968 N_SET_B_c_1365_n N_A_1930_295#_c_1504_n 0.00290311f $X=10.875 $Y=1.605
+ $X2=0 $Y2=0
cc_969 N_SET_B_c_1370_n N_A_1930_295#_c_1504_n 0.00157836f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_970 N_SET_B_c_1371_n N_A_1930_295#_c_1504_n 0.00203f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_971 N_SET_B_M1043_g N_A_1930_295#_c_1505_n 9.90788e-19 $X=10.96 $Y=0.445
+ $X2=0 $Y2=0
cc_972 N_SET_B_c_1362_n N_A_1930_295#_c_1506_n 2.09583e-19 $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_973 N_SET_B_M1043_g N_A_1930_295#_c_1506_n 0.00802103f $X=10.96 $Y=0.445
+ $X2=0 $Y2=0
cc_974 N_SET_B_c_1366_n N_A_1930_295#_c_1506_n 3.26955e-19 $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_975 N_SET_B_M1043_g N_A_1930_295#_c_1507_n 0.0112032f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_976 N_SET_B_c_1365_n N_A_1930_295#_c_1507_n 0.00463602f $X=10.875 $Y=1.605
+ $X2=0 $Y2=0
cc_977 N_SET_B_c_1366_n N_A_1930_295#_c_1507_n 0.052296f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_978 N_SET_B_c_1366_n N_A_1930_295#_c_1516_n 0.017477f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_979 N_SET_B_c_1365_n N_A_1735_329#_c_1623_n 0.0250342f $X=10.875 $Y=1.605
+ $X2=0 $Y2=0
cc_980 N_SET_B_c_1366_n N_A_1735_329#_c_1623_n 0.00123477f $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_981 N_SET_B_c_1362_n N_A_1735_329#_c_1624_n 0.00306987f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_982 N_SET_B_c_1367_n N_A_1735_329#_c_1624_n 0.0250342f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_983 N_SET_B_c_1368_n N_A_1735_329#_c_1640_n 0.0147965f $X=9.675 $Y=1.53 $X2=0
+ $Y2=0
cc_984 N_SET_B_M1043_g N_A_1735_329#_c_1641_n 0.00263881f $X=10.96 $Y=0.445
+ $X2=0 $Y2=0
cc_985 N_SET_B_c_1362_n N_A_1735_329#_c_1633_n 0.0152108f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_986 N_SET_B_c_1366_n N_A_1735_329#_c_1633_n 0.0512144f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_987 N_SET_B_c_1370_n N_A_1735_329#_c_1633_n 0.0013632f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_988 N_SET_B_c_1371_n N_A_1735_329#_c_1633_n 0.0156012f $X=9.82 $Y=1.53 $X2=0
+ $Y2=0
cc_989 N_SET_B_M1043_g N_A_1735_329#_c_1618_n 0.0090922f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_990 N_SET_B_c_1362_n N_A_1735_329#_c_1634_n 0.00477237f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_991 N_SET_B_M1043_g N_A_1735_329#_c_1620_n 0.0118997f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_992 N_SET_B_M1043_g N_A_1735_329#_c_1621_n 0.0250342f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_993 N_SET_B_c_1362_n N_A_1735_329#_c_1636_n 0.00797317f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_994 N_SET_B_c_1366_n N_A_1735_329#_c_1636_n 0.0150275f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_995 N_SET_B_c_1362_n N_A_1735_329#_c_1667_n 4.52613e-19 $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_996 N_SET_B_c_1365_n N_A_1735_329#_c_1667_n 2.27844e-19 $X=10.875 $Y=1.605
+ $X2=0 $Y2=0
cc_997 N_SET_B_c_1366_n N_A_1735_329#_c_1667_n 0.0162126f $X=10.85 $Y=1.61 $X2=0
+ $Y2=0
cc_998 N_SET_B_c_1367_n N_A_1735_329#_c_1667_n 0.00109766f $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_999 N_SET_B_c_1362_n N_A_1735_329#_c_1637_n 6.07879e-19 $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_1000 N_SET_B_c_1368_n N_A_1735_329#_c_1637_n 0.0037791f $X=9.675 $Y=1.53
+ $X2=0 $Y2=0
cc_1001 N_SET_B_c_1370_n N_A_1735_329#_c_1637_n 6.09285e-19 $X=9.82 $Y=1.53
+ $X2=0 $Y2=0
cc_1002 N_SET_B_c_1371_n N_A_1735_329#_c_1637_n 0.00347269f $X=9.82 $Y=1.53
+ $X2=0 $Y2=0
cc_1003 N_SET_B_c_1362_n N_A_1735_329#_c_1675_n 0.00907673f $X=10.495 $Y=1.99
+ $X2=0 $Y2=0
cc_1004 N_SET_B_c_1366_n N_A_1735_329#_c_1675_n 0.0165572f $X=10.85 $Y=1.61
+ $X2=0 $Y2=0
cc_1005 N_SET_B_M1043_g N_A_1735_329#_c_1622_n 0.0134742f $X=10.96 $Y=0.445
+ $X2=0 $Y2=0
cc_1006 N_SET_B_c_1361_n N_VPWR_c_1913_n 0.00384082f $X=7.54 $Y=1.99 $X2=0 $Y2=0
cc_1007 N_SET_B_c_1372_n N_VPWR_c_1913_n 0.0013983f $X=7.53 $Y=1.53 $X2=0 $Y2=0
cc_1008 N_SET_B_c_1362_n N_VPWR_c_1914_n 0.00959979f $X=10.495 $Y=1.99 $X2=0
+ $Y2=0
cc_1009 N_SET_B_c_1362_n N_VPWR_c_1915_n 0.0028116f $X=10.495 $Y=1.99 $X2=0
+ $Y2=0
cc_1010 N_SET_B_c_1361_n N_VPWR_c_1922_n 0.00743866f $X=7.54 $Y=1.99 $X2=0 $Y2=0
cc_1011 N_SET_B_c_1362_n N_VPWR_c_1932_n 0.00586964f $X=10.495 $Y=1.99 $X2=0
+ $Y2=0
cc_1012 N_SET_B_c_1368_n N_VPWR_c_1938_n 0.00120798f $X=9.675 $Y=1.53 $X2=0
+ $Y2=0
cc_1013 N_SET_B_c_1361_n N_VPWR_c_1907_n 0.00868094f $X=7.54 $Y=1.99 $X2=0 $Y2=0
cc_1014 N_SET_B_c_1362_n N_VPWR_c_1907_n 0.00655278f $X=10.495 $Y=1.99 $X2=0
+ $Y2=0
cc_1015 N_SET_B_M1043_g N_VGND_c_2323_n 0.00577126f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_1016 N_SET_B_M1043_g N_VGND_c_2338_n 0.00585385f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_1017 N_SET_B_M1025_g N_VGND_c_2343_n 0.0187314f $X=7.62 $Y=0.445 $X2=0 $Y2=0
cc_1018 N_SET_B_M1043_g N_VGND_c_2346_n 0.00754935f $X=10.96 $Y=0.445 $X2=0
+ $Y2=0
cc_1019 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1623_n 0.0123735f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1020 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1623_n 0.0202974f $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1021 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1624_n 0.00679817f $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1022 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1611_n 0.00238264f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1023 N_A_1930_295#_c_1508_n N_A_1735_329#_c_1611_n 0.0197873f $X=11.855
+ $Y=1.185 $X2=0 $Y2=0
cc_1024 N_A_1930_295#_c_1509_n N_A_1735_329#_c_1611_n 0.00116113f $X=11.855
+ $Y=0.397 $X2=0 $Y2=0
cc_1025 N_A_1930_295#_c_1518_n N_A_1735_329#_c_1611_n 0.0159459f $X=11.815
+ $Y=1.27 $X2=0 $Y2=0
cc_1026 N_A_1930_295#_c_1508_n N_A_1735_329#_c_1612_n 0.00230619f $X=11.855
+ $Y=1.185 $X2=0 $Y2=0
cc_1027 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1626_n 0.00292762f $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1028 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1615_n 9.41286e-19 $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1029 N_A_1930_295#_c_1518_n N_A_1735_329#_c_1615_n 5.49649e-19 $X=11.815
+ $Y=1.27 $X2=0 $Y2=0
cc_1030 N_A_1930_295#_c_1511_n N_A_1735_329#_c_1640_n 5.33749e-19 $X=9.75
+ $Y=1.99 $X2=0 $Y2=0
cc_1031 N_A_1930_295#_M1039_g N_A_1735_329#_c_1641_n 0.0128291f $X=10.17
+ $Y=0.445 $X2=0 $Y2=0
cc_1032 N_A_1930_295#_c_1505_n N_A_1735_329#_c_1641_n 0.00609647f $X=10.23
+ $Y=1.02 $X2=0 $Y2=0
cc_1033 N_A_1930_295#_c_1506_n N_A_1735_329#_c_1641_n 0.00199588f $X=10.23
+ $Y=1.02 $X2=0 $Y2=0
cc_1034 N_A_1930_295#_c_1511_n N_A_1735_329#_c_1633_n 0.00945937f $X=9.75
+ $Y=1.99 $X2=0 $Y2=0
cc_1035 N_A_1930_295#_c_1512_n N_A_1735_329#_c_1633_n 0.00241624f $X=10.095
+ $Y=1.55 $X2=0 $Y2=0
cc_1036 N_A_1930_295#_M1039_g N_A_1735_329#_c_1618_n 0.00755004f $X=10.17
+ $Y=0.445 $X2=0 $Y2=0
cc_1037 N_A_1930_295#_M1039_g N_A_1735_329#_c_1619_n 2.40752e-19 $X=10.17
+ $Y=0.445 $X2=0 $Y2=0
cc_1038 N_A_1930_295#_c_1505_n N_A_1735_329#_c_1619_n 0.0101679f $X=10.23
+ $Y=1.02 $X2=0 $Y2=0
cc_1039 N_A_1930_295#_c_1506_n N_A_1735_329#_c_1619_n 0.00160145f $X=10.23
+ $Y=1.02 $X2=0 $Y2=0
cc_1040 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1619_n 0.0143582f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1041 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1620_n 0.0545597f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1042 N_A_1930_295#_c_1508_n N_A_1735_329#_c_1620_n 0.011018f $X=11.855
+ $Y=1.185 $X2=0 $Y2=0
cc_1043 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1621_n 0.0135148f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1044 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1636_n 0.00572977f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1045 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1636_n 0.0114977f $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1046 N_A_1930_295#_c_1507_n N_A_1735_329#_c_1667_n 0.0162897f $X=11.685
+ $Y=1.27 $X2=0 $Y2=0
cc_1047 N_A_1930_295#_c_1517_n N_A_1735_329#_c_1667_n 0.0229496f $X=11.77
+ $Y=2.285 $X2=0 $Y2=0
cc_1048 N_A_1930_295#_c_1511_n N_A_1735_329#_c_1637_n 0.0161207f $X=9.75 $Y=1.99
+ $X2=0 $Y2=0
cc_1049 N_A_1930_295#_c_1508_n N_A_1735_329#_c_1622_n 0.0137675f $X=11.855
+ $Y=1.185 $X2=0 $Y2=0
cc_1050 N_A_1930_295#_c_1509_n N_A_1735_329#_c_1622_n 0.00686122f $X=11.855
+ $Y=0.397 $X2=0 $Y2=0
cc_1051 N_A_1930_295#_c_1511_n N_VPWR_c_1914_n 0.00533159f $X=9.75 $Y=1.99 $X2=0
+ $Y2=0
cc_1052 N_A_1930_295#_c_1517_n N_VPWR_c_1915_n 0.0143781f $X=11.77 $Y=2.285
+ $X2=0 $Y2=0
cc_1053 N_A_1930_295#_c_1517_n N_VPWR_c_1916_n 0.0182101f $X=11.77 $Y=2.285
+ $X2=0 $Y2=0
cc_1054 N_A_1930_295#_c_1517_n N_VPWR_c_1917_n 0.0622168f $X=11.77 $Y=2.285
+ $X2=0 $Y2=0
cc_1055 N_A_1930_295#_c_1511_n N_VPWR_c_1923_n 0.00486131f $X=9.75 $Y=1.99 $X2=0
+ $Y2=0
cc_1056 N_A_1930_295#_M1002_d N_VPWR_c_1907_n 0.00404917f $X=11.625 $Y=2.065
+ $X2=0 $Y2=0
cc_1057 N_A_1930_295#_c_1511_n N_VPWR_c_1907_n 0.00719873f $X=9.75 $Y=1.99 $X2=0
+ $Y2=0
cc_1058 N_A_1930_295#_c_1517_n N_VPWR_c_1907_n 0.00993603f $X=11.77 $Y=2.285
+ $X2=0 $Y2=0
cc_1059 N_A_1930_295#_c_1517_n N_Q_N_c_2279_n 0.0038838f $X=11.77 $Y=2.285 $X2=0
+ $Y2=0
cc_1060 N_A_1930_295#_c_1508_n N_Q_N_c_2279_n 0.00803225f $X=11.855 $Y=1.185
+ $X2=0 $Y2=0
cc_1061 N_A_1930_295#_c_1518_n N_Q_N_c_2279_n 0.00493346f $X=11.815 $Y=1.27
+ $X2=0 $Y2=0
cc_1062 N_A_1930_295#_c_1508_n N_VGND_c_2323_n 2.0356e-19 $X=11.855 $Y=1.185
+ $X2=0 $Y2=0
cc_1063 N_A_1930_295#_c_1509_n N_VGND_c_2323_n 0.0212548f $X=11.855 $Y=0.397
+ $X2=0 $Y2=0
cc_1064 N_A_1930_295#_c_1509_n N_VGND_c_2324_n 0.0234105f $X=11.855 $Y=0.397
+ $X2=0 $Y2=0
cc_1065 N_A_1930_295#_c_1508_n N_VGND_c_2325_n 0.0212846f $X=11.855 $Y=1.185
+ $X2=0 $Y2=0
cc_1066 N_A_1930_295#_c_1509_n N_VGND_c_2325_n 0.0186051f $X=11.855 $Y=0.397
+ $X2=0 $Y2=0
cc_1067 N_A_1930_295#_M1039_g N_VGND_c_2338_n 0.00362032f $X=10.17 $Y=0.445
+ $X2=0 $Y2=0
cc_1068 N_A_1930_295#_M1001_d N_VGND_c_2346_n 0.00209344f $X=11.64 $Y=0.235
+ $X2=0 $Y2=0
cc_1069 N_A_1930_295#_M1039_g N_VGND_c_2346_n 0.00585485f $X=10.17 $Y=0.445
+ $X2=0 $Y2=0
cc_1070 N_A_1930_295#_c_1509_n N_VGND_c_2346_n 0.014068f $X=11.855 $Y=0.397
+ $X2=0 $Y2=0
cc_1071 N_A_1735_329#_c_1630_n N_A_2739_47#_c_1800_n 0.0104722f $X=14.055
+ $Y=1.605 $X2=0 $Y2=0
cc_1072 N_A_1735_329#_c_1631_n N_A_2739_47#_c_1800_n 0.00790691f $X=14.055
+ $Y=1.705 $X2=0 $Y2=0
cc_1073 N_A_1735_329#_M1033_g N_A_2739_47#_c_1795_n 0.0205349f $X=14.08 $Y=0.445
+ $X2=0 $Y2=0
cc_1074 N_A_1735_329#_c_1613_n N_A_2739_47#_c_1797_n 0.00297226f $X=12.975
+ $Y=0.995 $X2=0 $Y2=0
cc_1075 N_A_1735_329#_M1033_g N_A_2739_47#_c_1797_n 0.0112396f $X=14.08 $Y=0.445
+ $X2=0 $Y2=0
cc_1076 N_A_1735_329#_c_1627_n N_A_2739_47#_c_1802_n 0.00282932f $X=13 $Y=1.41
+ $X2=0 $Y2=0
cc_1077 N_A_1735_329#_c_1615_n N_A_2739_47#_c_1802_n 0.00189409f $X=13.1 $Y=1.16
+ $X2=0 $Y2=0
cc_1078 N_A_1735_329#_c_1630_n N_A_2739_47#_c_1802_n 0.0142026f $X=14.055
+ $Y=1.605 $X2=0 $Y2=0
cc_1079 N_A_1735_329#_c_1631_n N_A_2739_47#_c_1802_n 0.00449389f $X=14.055
+ $Y=1.705 $X2=0 $Y2=0
cc_1080 N_A_1735_329#_c_1614_n N_A_2739_47#_c_1798_n 0.00559143f $X=13.955
+ $Y=1.16 $X2=0 $Y2=0
cc_1081 N_A_1735_329#_c_1617_n N_A_2739_47#_c_1798_n 0.0233563f $X=14.055
+ $Y=1.16 $X2=0 $Y2=0
cc_1082 N_A_1735_329#_c_1614_n N_A_2739_47#_c_1816_n 0.0319869f $X=13.955
+ $Y=1.16 $X2=0 $Y2=0
cc_1083 N_A_1735_329#_c_1630_n N_A_2739_47#_c_1799_n 0.00322527f $X=14.055
+ $Y=1.605 $X2=0 $Y2=0
cc_1084 N_A_1735_329#_c_1617_n N_A_2739_47#_c_1799_n 0.0216214f $X=14.055
+ $Y=1.16 $X2=0 $Y2=0
cc_1085 N_A_1735_329#_c_1636_n N_VPWR_M1002_s 0.00211122f $X=11.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1086 N_A_1735_329#_c_1633_n N_VPWR_c_1914_n 0.0268245f $X=10.645 $Y=1.98
+ $X2=0 $Y2=0
cc_1087 N_A_1735_329#_c_1634_n N_VPWR_c_1914_n 0.013391f $X=10.73 $Y=2.285 $X2=0
+ $Y2=0
cc_1088 N_A_1735_329#_c_1637_n N_VPWR_c_1914_n 0.0106386f $X=9.65 $Y=1.98 $X2=0
+ $Y2=0
cc_1089 N_A_1735_329#_c_1624_n N_VPWR_c_1915_n 0.0104645f $X=11.535 $Y=1.99
+ $X2=0 $Y2=0
cc_1090 N_A_1735_329#_c_1634_n N_VPWR_c_1915_n 0.0124141f $X=10.73 $Y=2.285
+ $X2=0 $Y2=0
cc_1091 N_A_1735_329#_c_1636_n N_VPWR_c_1915_n 0.0241606f $X=11.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1092 N_A_1735_329#_c_1624_n N_VPWR_c_1916_n 0.00643335f $X=11.535 $Y=1.99
+ $X2=0 $Y2=0
cc_1093 N_A_1735_329#_c_1624_n N_VPWR_c_1917_n 0.00283678f $X=11.535 $Y=1.99
+ $X2=0 $Y2=0
cc_1094 N_A_1735_329#_c_1611_n N_VPWR_c_1917_n 0.00634276f $X=12.43 $Y=1.16
+ $X2=0 $Y2=0
cc_1095 N_A_1735_329#_c_1626_n N_VPWR_c_1917_n 0.00767971f $X=12.53 $Y=1.41
+ $X2=0 $Y2=0
cc_1096 N_A_1735_329#_c_1627_n N_VPWR_c_1918_n 0.0261524f $X=13 $Y=1.41 $X2=0
+ $Y2=0
cc_1097 N_A_1735_329#_c_1614_n N_VPWR_c_1918_n 0.00856698f $X=13.955 $Y=1.16
+ $X2=0 $Y2=0
cc_1098 N_A_1735_329#_c_1631_n N_VPWR_c_1918_n 0.00308982f $X=14.055 $Y=1.705
+ $X2=0 $Y2=0
cc_1099 N_A_1735_329#_c_1631_n N_VPWR_c_1919_n 0.0220967f $X=14.055 $Y=1.705
+ $X2=0 $Y2=0
cc_1100 N_A_1735_329#_c_1640_n N_VPWR_c_1923_n 0.0402948f $X=9.565 $Y=2.292
+ $X2=0 $Y2=0
cc_1101 N_A_1735_329#_c_1633_n N_VPWR_c_1923_n 0.00522413f $X=10.645 $Y=1.98
+ $X2=0 $Y2=0
cc_1102 N_A_1735_329#_c_1637_n N_VPWR_c_1923_n 0.00927152f $X=9.65 $Y=1.98 $X2=0
+ $Y2=0
cc_1103 N_A_1735_329#_c_1626_n N_VPWR_c_1925_n 0.00605302f $X=12.53 $Y=1.41
+ $X2=0 $Y2=0
cc_1104 N_A_1735_329#_c_1627_n N_VPWR_c_1925_n 0.00567349f $X=13 $Y=1.41 $X2=0
+ $Y2=0
cc_1105 N_A_1735_329#_c_1631_n N_VPWR_c_1927_n 0.00427505f $X=14.055 $Y=1.705
+ $X2=0 $Y2=0
cc_1106 N_A_1735_329#_c_1633_n N_VPWR_c_1932_n 0.00353433f $X=10.645 $Y=1.98
+ $X2=0 $Y2=0
cc_1107 N_A_1735_329#_c_1634_n N_VPWR_c_1932_n 0.0134676f $X=10.73 $Y=2.285
+ $X2=0 $Y2=0
cc_1108 N_A_1735_329#_c_1636_n N_VPWR_c_1932_n 0.00480174f $X=11.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1109 N_A_1735_329#_M1012_d N_VPWR_c_1907_n 0.00826962f $X=8.675 $Y=1.645
+ $X2=0 $Y2=0
cc_1110 N_A_1735_329#_M1013_d N_VPWR_c_1907_n 0.00240388f $X=10.585 $Y=2.065
+ $X2=0 $Y2=0
cc_1111 N_A_1735_329#_c_1624_n N_VPWR_c_1907_n 0.012023f $X=11.535 $Y=1.99 $X2=0
+ $Y2=0
cc_1112 N_A_1735_329#_c_1626_n N_VPWR_c_1907_n 0.0114618f $X=12.53 $Y=1.41 $X2=0
+ $Y2=0
cc_1113 N_A_1735_329#_c_1627_n N_VPWR_c_1907_n 0.0107621f $X=13 $Y=1.41 $X2=0
+ $Y2=0
cc_1114 N_A_1735_329#_c_1631_n N_VPWR_c_1907_n 0.00873932f $X=14.055 $Y=1.705
+ $X2=0 $Y2=0
cc_1115 N_A_1735_329#_c_1640_n N_VPWR_c_1907_n 0.0250088f $X=9.565 $Y=2.292
+ $X2=0 $Y2=0
cc_1116 N_A_1735_329#_c_1633_n N_VPWR_c_1907_n 0.0151012f $X=10.645 $Y=1.98
+ $X2=0 $Y2=0
cc_1117 N_A_1735_329#_c_1634_n N_VPWR_c_1907_n 0.00809922f $X=10.73 $Y=2.285
+ $X2=0 $Y2=0
cc_1118 N_A_1735_329#_c_1636_n N_VPWR_c_1907_n 0.00920524f $X=11.245 $Y=1.98
+ $X2=0 $Y2=0
cc_1119 N_A_1735_329#_c_1637_n N_VPWR_c_1907_n 0.00608385f $X=9.65 $Y=1.98 $X2=0
+ $Y2=0
cc_1120 N_A_1735_329#_c_1640_n A_1870_413# 0.00509751f $X=9.565 $Y=2.292
+ $X2=-0.19 $Y2=-0.24
cc_1121 N_A_1735_329#_c_1637_n A_1870_413# 0.00191133f $X=9.65 $Y=1.98 $X2=-0.19
+ $Y2=-0.24
cc_1122 N_A_1735_329#_c_1612_n N_Q_N_c_2279_n 0.0107292f $X=12.505 $Y=0.995
+ $X2=0 $Y2=0
cc_1123 N_A_1735_329#_c_1626_n N_Q_N_c_2279_n 0.0172757f $X=12.53 $Y=1.41 $X2=0
+ $Y2=0
cc_1124 N_A_1735_329#_c_1613_n N_Q_N_c_2279_n 0.0184062f $X=12.975 $Y=0.995
+ $X2=0 $Y2=0
cc_1125 N_A_1735_329#_c_1627_n N_Q_N_c_2279_n 0.0220641f $X=13 $Y=1.41 $X2=0
+ $Y2=0
cc_1126 N_A_1735_329#_c_1615_n N_Q_N_c_2279_n 0.0587962f $X=13.1 $Y=1.16 $X2=0
+ $Y2=0
cc_1127 N_A_1735_329#_c_1641_n N_VGND_c_2323_n 0.00676624f $X=10.605 $Y=0.36
+ $X2=0 $Y2=0
cc_1128 N_A_1735_329#_c_1618_n N_VGND_c_2323_n 0.00354515f $X=10.69 $Y=0.845
+ $X2=0 $Y2=0
cc_1129 N_A_1735_329#_c_1620_n N_VGND_c_2323_n 0.00796254f $X=11.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1130 N_A_1735_329#_c_1621_n N_VGND_c_2323_n 0.00394879f $X=11.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1131 N_A_1735_329#_c_1622_n N_VGND_c_2323_n 0.00377035f $X=11.442 $Y=0.765
+ $X2=0 $Y2=0
cc_1132 N_A_1735_329#_c_1621_n N_VGND_c_2324_n 0.0019796f $X=11.38 $Y=0.93 $X2=0
+ $Y2=0
cc_1133 N_A_1735_329#_c_1622_n N_VGND_c_2324_n 0.00464047f $X=11.442 $Y=0.765
+ $X2=0 $Y2=0
cc_1134 N_A_1735_329#_c_1611_n N_VGND_c_2325_n 0.00537422f $X=12.43 $Y=1.16
+ $X2=0 $Y2=0
cc_1135 N_A_1735_329#_c_1612_n N_VGND_c_2325_n 0.00444548f $X=12.505 $Y=0.995
+ $X2=0 $Y2=0
cc_1136 N_A_1735_329#_c_1622_n N_VGND_c_2325_n 0.00213038f $X=11.442 $Y=0.765
+ $X2=0 $Y2=0
cc_1137 N_A_1735_329#_c_1613_n N_VGND_c_2326_n 0.0170291f $X=12.975 $Y=0.995
+ $X2=0 $Y2=0
cc_1138 N_A_1735_329#_c_1614_n N_VGND_c_2326_n 0.00915844f $X=13.955 $Y=1.16
+ $X2=0 $Y2=0
cc_1139 N_A_1735_329#_M1033_g N_VGND_c_2326_n 0.00251081f $X=14.08 $Y=0.445
+ $X2=0 $Y2=0
cc_1140 N_A_1735_329#_M1033_g N_VGND_c_2327_n 0.0186193f $X=14.08 $Y=0.445 $X2=0
+ $Y2=0
cc_1141 N_A_1735_329#_c_1612_n N_VGND_c_2332_n 0.0054895f $X=12.505 $Y=0.995
+ $X2=0 $Y2=0
cc_1142 N_A_1735_329#_c_1613_n N_VGND_c_2332_n 0.00435091f $X=12.975 $Y=0.995
+ $X2=0 $Y2=0
cc_1143 N_A_1735_329#_M1033_g N_VGND_c_2334_n 0.00271402f $X=14.08 $Y=0.445
+ $X2=0 $Y2=0
cc_1144 N_A_1735_329#_c_1641_n N_VGND_c_2338_n 0.0842904f $X=10.605 $Y=0.36
+ $X2=0 $Y2=0
cc_1145 N_A_1735_329#_M1005_d N_VGND_c_2346_n 0.00463132f $X=9.165 $Y=0.235
+ $X2=0 $Y2=0
cc_1146 N_A_1735_329#_c_1612_n N_VGND_c_2346_n 0.0111395f $X=12.505 $Y=0.995
+ $X2=0 $Y2=0
cc_1147 N_A_1735_329#_c_1613_n N_VGND_c_2346_n 0.00861527f $X=12.975 $Y=0.995
+ $X2=0 $Y2=0
cc_1148 N_A_1735_329#_M1033_g N_VGND_c_2346_n 0.00634617f $X=14.08 $Y=0.445
+ $X2=0 $Y2=0
cc_1149 N_A_1735_329#_c_1641_n N_VGND_c_2346_n 0.0582503f $X=10.605 $Y=0.36
+ $X2=0 $Y2=0
cc_1150 N_A_1735_329#_c_1620_n N_VGND_c_2346_n 0.0193429f $X=11.38 $Y=0.93 $X2=0
+ $Y2=0
cc_1151 N_A_1735_329#_c_1621_n N_VGND_c_2346_n 0.00267073f $X=11.38 $Y=0.93
+ $X2=0 $Y2=0
cc_1152 N_A_1735_329#_c_1622_n N_VGND_c_2346_n 0.007891f $X=11.442 $Y=0.765
+ $X2=0 $Y2=0
cc_1153 N_A_1735_329#_c_1641_n A_1977_47# 0.00460484f $X=10.605 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_1154 N_A_1735_329#_c_1641_n A_2049_47# 0.0189122f $X=10.605 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_1155 N_A_1735_329#_c_1618_n A_2049_47# 0.00722679f $X=10.69 $Y=0.845
+ $X2=-0.19 $Y2=-0.24
cc_1156 N_A_2739_47#_c_1802_n N_VPWR_c_1918_n 0.0647314f $X=13.82 $Y=1.935 $X2=0
+ $Y2=0
cc_1157 N_A_2739_47#_c_1800_n N_VPWR_c_1919_n 0.00398983f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1158 N_A_2739_47#_c_1802_n N_VPWR_c_1919_n 0.0628748f $X=13.82 $Y=1.935 $X2=0
+ $Y2=0
cc_1159 N_A_2739_47#_c_1798_n N_VPWR_c_1919_n 0.0204719f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_1160 N_A_2739_47#_c_1799_n N_VPWR_c_1919_n 0.00226232f $X=15.05 $Y=1.202
+ $X2=0 $Y2=0
cc_1161 N_A_2739_47#_c_1801_n N_VPWR_c_1921_n 0.00741457f $X=15.05 $Y=1.41 $X2=0
+ $Y2=0
cc_1162 N_A_2739_47#_c_1802_n N_VPWR_c_1927_n 0.0131202f $X=13.82 $Y=1.935 $X2=0
+ $Y2=0
cc_1163 N_A_2739_47#_c_1800_n N_VPWR_c_1933_n 0.00702461f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1164 N_A_2739_47#_c_1801_n N_VPWR_c_1933_n 0.00524286f $X=15.05 $Y=1.41 $X2=0
+ $Y2=0
cc_1165 N_A_2739_47#_c_1800_n N_VPWR_c_1907_n 0.0126497f $X=14.58 $Y=1.41 $X2=0
+ $Y2=0
cc_1166 N_A_2739_47#_c_1801_n N_VPWR_c_1907_n 0.00926612f $X=15.05 $Y=1.41 $X2=0
+ $Y2=0
cc_1167 N_A_2739_47#_c_1802_n N_VPWR_c_1907_n 0.00704765f $X=13.82 $Y=1.935
+ $X2=0 $Y2=0
cc_1168 N_A_2739_47#_c_1801_n Q 0.015334f $X=15.05 $Y=1.41 $X2=0 $Y2=0
cc_1169 N_A_2739_47#_c_1800_n Q 8.35015e-19 $X=14.58 $Y=1.41 $X2=0 $Y2=0
cc_1170 N_A_2739_47#_c_1795_n Q 0.00292937f $X=14.605 $Y=0.995 $X2=0 $Y2=0
cc_1171 N_A_2739_47#_c_1801_n Q 0.00495339f $X=15.05 $Y=1.41 $X2=0 $Y2=0
cc_1172 N_A_2739_47#_c_1796_n Q 0.00773979f $X=15.075 $Y=0.995 $X2=0 $Y2=0
cc_1173 N_A_2739_47#_c_1798_n Q 0.021005f $X=14.5 $Y=1.16 $X2=0 $Y2=0
cc_1174 N_A_2739_47#_c_1799_n Q 0.0400426f $X=15.05 $Y=1.202 $X2=0 $Y2=0
cc_1175 N_A_2739_47#_c_1796_n N_Q_c_2305_n 0.0107839f $X=15.075 $Y=0.995 $X2=0
+ $Y2=0
cc_1176 N_A_2739_47#_c_1799_n N_Q_c_2305_n 0.00103509f $X=15.05 $Y=1.202 $X2=0
+ $Y2=0
cc_1177 N_A_2739_47#_c_1801_n Q 0.00528968f $X=15.05 $Y=1.41 $X2=0 $Y2=0
cc_1178 N_A_2739_47#_c_1799_n Q 0.00315148f $X=15.05 $Y=1.202 $X2=0 $Y2=0
cc_1179 N_A_2739_47#_c_1797_n N_VGND_c_2326_n 0.04163f $X=13.82 $Y=0.44 $X2=0
+ $Y2=0
cc_1180 N_A_2739_47#_c_1795_n N_VGND_c_2327_n 0.00631549f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1181 N_A_2739_47#_c_1797_n N_VGND_c_2327_n 0.0432591f $X=13.82 $Y=0.44 $X2=0
+ $Y2=0
cc_1182 N_A_2739_47#_c_1798_n N_VGND_c_2327_n 0.0337889f $X=14.5 $Y=1.16 $X2=0
+ $Y2=0
cc_1183 N_A_2739_47#_c_1799_n N_VGND_c_2327_n 0.00263742f $X=15.05 $Y=1.202
+ $X2=0 $Y2=0
cc_1184 N_A_2739_47#_c_1796_n N_VGND_c_2329_n 0.0066147f $X=15.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1185 N_A_2739_47#_c_1797_n N_VGND_c_2334_n 0.0128687f $X=13.82 $Y=0.44 $X2=0
+ $Y2=0
cc_1186 N_A_2739_47#_c_1795_n N_VGND_c_2339_n 0.00585385f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1187 N_A_2739_47#_c_1796_n N_VGND_c_2339_n 0.00467644f $X=15.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1188 N_A_2739_47#_M1033_s N_VGND_c_2346_n 0.0069454f $X=13.695 $Y=0.235 $X2=0
+ $Y2=0
cc_1189 N_A_2739_47#_c_1795_n N_VGND_c_2346_n 0.0110943f $X=14.605 $Y=0.995
+ $X2=0 $Y2=0
cc_1190 N_A_2739_47#_c_1796_n N_VGND_c_2346_n 0.00898223f $X=15.075 $Y=0.995
+ $X2=0 $Y2=0
cc_1191 N_A_2739_47#_c_1797_n N_VGND_c_2346_n 0.00704765f $X=13.82 $Y=0.44 $X2=0
+ $Y2=0
cc_1192 N_A_27_369#_c_1856_n N_VPWR_M1007_d 0.00338362f $X=1.035 $Y=1.935
+ $X2=-0.19 $Y2=1.305
cc_1193 N_A_27_369#_c_1855_n N_VPWR_c_1908_n 0.0204331f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1194 N_A_27_369#_c_1856_n N_VPWR_c_1908_n 0.0183997f $X=1.035 $Y=1.935 $X2=0
+ $Y2=0
cc_1195 N_A_27_369#_c_1864_n N_VPWR_c_1908_n 0.00358735f $X=1.12 $Y=2.255 $X2=0
+ $Y2=0
cc_1196 N_A_27_369#_c_1871_n N_VPWR_c_1908_n 0.0140744f $X=1.205 $Y=2.36 $X2=0
+ $Y2=0
cc_1197 N_A_27_369#_c_1855_n N_VPWR_c_1929_n 0.0180865f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1198 N_A_27_369#_c_1856_n N_VPWR_c_1929_n 0.00206566f $X=1.035 $Y=1.935 $X2=0
+ $Y2=0
cc_1199 N_A_27_369#_c_1856_n N_VPWR_c_1930_n 0.002804f $X=1.035 $Y=1.935 $X2=0
+ $Y2=0
cc_1200 N_A_27_369#_c_1871_n N_VPWR_c_1930_n 0.00987263f $X=1.205 $Y=2.36 $X2=0
+ $Y2=0
cc_1201 N_A_27_369#_c_1858_n N_VPWR_c_1930_n 0.0595487f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1202 N_A_27_369#_M1007_s N_VPWR_c_1907_n 0.00244672f $X=0.135 $Y=1.845 $X2=0
+ $Y2=0
cc_1203 N_A_27_369#_M1022_d N_VPWR_c_1907_n 0.00217543f $X=1.935 $Y=1.845 $X2=0
+ $Y2=0
cc_1204 N_A_27_369#_c_1855_n N_VPWR_c_1907_n 0.00991202f $X=0.215 $Y=2.025 $X2=0
+ $Y2=0
cc_1205 N_A_27_369#_c_1856_n N_VPWR_c_1907_n 0.010397f $X=1.035 $Y=1.935 $X2=0
+ $Y2=0
cc_1206 N_A_27_369#_c_1871_n N_VPWR_c_1907_n 0.00643973f $X=1.205 $Y=2.36 $X2=0
+ $Y2=0
cc_1207 N_A_27_369#_c_1858_n N_VPWR_c_1907_n 0.0371977f $X=2.08 $Y=2.34 $X2=0
+ $Y2=0
cc_1208 N_A_27_369#_c_1856_n A_211_369# 0.00269538f $X=1.035 $Y=1.935 $X2=-0.19
+ $Y2=1.305
cc_1209 N_A_27_369#_c_1864_n A_211_369# 0.00240059f $X=1.12 $Y=2.255 $X2=-0.19
+ $Y2=1.305
cc_1210 N_A_27_369#_c_1871_n A_211_369# 9.06933e-19 $X=1.205 $Y=2.36 $X2=-0.19
+ $Y2=1.305
cc_1211 N_A_27_369#_c_1858_n A_211_369# 6.40929e-19 $X=2.08 $Y=2.34 $X2=-0.19
+ $Y2=1.305
cc_1212 N_A_27_369#_c_1858_n N_A_199_47#_M1040_d 0.00358545f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1213 N_A_27_369#_c_1856_n N_A_199_47#_c_2157_n 0.0119789f $X=1.035 $Y=1.935
+ $X2=0 $Y2=0
cc_1214 N_A_27_369#_c_1864_n N_A_199_47#_c_2157_n 0.00338342f $X=1.12 $Y=2.255
+ $X2=0 $Y2=0
cc_1215 N_A_27_369#_c_1858_n N_A_199_47#_c_2157_n 0.0215797f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1216 N_A_27_369#_c_1858_n N_A_199_47#_c_2150_n 0.00286711f $X=2.08 $Y=2.34
+ $X2=0 $Y2=0
cc_1217 N_A_27_369#_c_1856_n N_A_199_47#_c_2145_n 9.93859e-19 $X=1.035 $Y=1.935
+ $X2=0 $Y2=0
cc_1218 N_VPWR_c_1907_n A_211_369# 0.00184695f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1219 N_VPWR_c_1907_n N_A_199_47#_M1040_d 0.00232895f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1220 N_VPWR_c_1907_n N_A_199_47#_M1003_s 0.00206785f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1221 N_VPWR_c_1931_n N_A_199_47#_c_2148_n 0.0139015f $X=6.445 $Y=2.72 $X2=0
+ $Y2=0
cc_1222 N_VPWR_c_1907_n N_A_199_47#_c_2148_n 0.00399922f $X=15.41 $Y=2.72 $X2=0
+ $Y2=0
cc_1223 N_VPWR_c_1909_n N_A_199_47#_c_2149_n 5.11867e-19 $X=3.07 $Y=2.34 $X2=0
+ $Y2=0
cc_1224 N_VPWR_c_1907_n A_1169_413# 0.00263276f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1225 N_VPWR_c_1912_n A_1652_329# 5.2056e-19 $X=8.37 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1226 N_VPWR_c_1938_n A_1652_329# 6.507e-19 $X=8.71 $Y=2.465 $X2=-0.19
+ $Y2=-0.24
cc_1227 N_VPWR_c_1907_n A_1870_413# 0.0024832f $X=15.41 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_1228 N_VPWR_c_1907_n N_Q_N_M1019_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1229 N_VPWR_c_1917_n N_Q_N_c_2279_n 0.0735565f $X=12.295 $Y=1.66 $X2=0 $Y2=0
cc_1230 N_VPWR_c_1918_n N_Q_N_c_2279_n 0.0643033f $X=13.3 $Y=1.66 $X2=0 $Y2=0
cc_1231 N_VPWR_c_1925_n N_Q_N_c_2279_n 0.0267874f $X=13.215 $Y=2.72 $X2=0 $Y2=0
cc_1232 N_VPWR_c_1907_n N_Q_N_c_2279_n 0.0162161f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1233 N_VPWR_c_1907_n N_Q_M1014_s 0.0033595f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1234 N_VPWR_c_1933_n Q 0.0213494f $X=15.25 $Y=2.72 $X2=0 $Y2=0
cc_1235 N_VPWR_c_1907_n Q 0.013832f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_1236 N_VPWR_c_1921_n Q 0.0744069f $X=15.335 $Y=1.66 $X2=0 $Y2=0
cc_1237 N_VPWR_c_1917_n N_VGND_c_2325_n 0.00710932f $X=12.295 $Y=1.66 $X2=0
+ $Y2=0
cc_1238 N_VPWR_c_1918_n N_VGND_c_2326_n 0.0102631f $X=13.3 $Y=1.66 $X2=0 $Y2=0
cc_1239 N_VPWR_c_1921_n N_VGND_c_2329_n 0.00938925f $X=15.335 $Y=1.66 $X2=0
+ $Y2=0
cc_1240 N_A_199_47#_c_2154_n N_VGND_c_2318_n 0.00853026f $X=1.655 $Y=0.42 $X2=0
+ $Y2=0
cc_1241 N_A_199_47#_c_2154_n N_VGND_c_2319_n 0.0200007f $X=1.655 $Y=0.42 $X2=0
+ $Y2=0
cc_1242 N_A_199_47#_c_2154_n N_VGND_c_2336_n 0.0432896f $X=1.655 $Y=0.42 $X2=0
+ $Y2=0
cc_1243 N_A_199_47#_c_2143_n N_VGND_c_2337_n 0.0228313f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1244 N_A_199_47#_M1028_d N_VGND_c_2346_n 0.00264864f $X=0.995 $Y=0.235 $X2=0
+ $Y2=0
cc_1245 N_A_199_47#_M1031_s N_VGND_c_2346_n 0.0054218f $X=4.955 $Y=0.235 $X2=0
+ $Y2=0
cc_1246 N_A_199_47#_c_2154_n N_VGND_c_2346_n 0.0310791f $X=1.655 $Y=0.42 $X2=0
+ $Y2=0
cc_1247 N_A_199_47#_c_2143_n N_VGND_c_2346_n 0.0124358f $X=5.08 $Y=0.42 $X2=0
+ $Y2=0
cc_1248 N_A_199_47#_c_2154_n A_295_47# 0.00409661f $X=1.655 $Y=0.42 $X2=-0.19
+ $Y2=-0.24
cc_1249 N_A_199_47#_c_2145_n A_295_47# 0.00111253f $X=1.76 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_1250 N_Q_N_c_2279_n N_VGND_c_2326_n 0.0413385f $X=12.765 $Y=0.38 $X2=0 $Y2=0
cc_1251 N_Q_N_c_2279_n N_VGND_c_2332_n 0.0268516f $X=12.765 $Y=0.38 $X2=0 $Y2=0
cc_1252 N_Q_N_M1015_s N_VGND_c_2346_n 0.0025535f $X=12.58 $Y=0.235 $X2=0 $Y2=0
cc_1253 N_Q_N_c_2279_n N_VGND_c_2346_n 0.0163533f $X=12.765 $Y=0.38 $X2=0 $Y2=0
cc_1254 N_Q_c_2305_n N_VGND_c_2329_n 0.0471812f $X=14.815 $Y=0.44 $X2=0 $Y2=0
cc_1255 N_Q_c_2305_n N_VGND_c_2339_n 0.0204545f $X=14.815 $Y=0.44 $X2=0 $Y2=0
cc_1256 N_Q_M1006_d N_VGND_c_2346_n 0.00330789f $X=14.68 $Y=0.235 $X2=0 $Y2=0
cc_1257 N_Q_c_2305_n N_VGND_c_2346_n 0.0140179f $X=14.815 $Y=0.44 $X2=0 $Y2=0
cc_1258 N_VGND_c_2346_n A_109_47# 0.0042254f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1259 N_VGND_c_2346_n A_295_47# 0.00218006f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1260 N_VGND_c_2346_n A_1177_47# 0.00726675f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1261 N_VGND_c_2346_n A_1467_47# 0.0087201f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1262 N_VGND_c_2346_n A_1655_47# 0.0171719f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1263 N_VGND_c_2346_n A_1977_47# 0.00169327f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
cc_1264 N_VGND_c_2346_n A_2049_47# 0.00594765f $X=15.41 $Y=0 $X2=-0.19 $Y2=-0.24
