# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdfrbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfrbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.72000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 0.975000 0.490000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.160200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.120000 1.355000 3.655000 2.465000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.564000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.860000 0.265000 13.260000 1.695000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.494750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.770000 1.535000 14.205000 2.080000 ;
        RECT 13.780000 0.310000 14.205000 0.825000 ;
        RECT 14.035000 0.825000 14.205000 1.535000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.230000 0.765000  7.810000 1.045000 ;
        RECT 10.600000 1.065000 11.370000 1.275000 ;
        RECT 11.065000 0.635000 11.370000 1.065000 ;
      LAYER mcon ;
        RECT  7.255000 0.765000  7.425000 0.935000 ;
        RECT  7.615000 0.765000  7.785000 0.935000 ;
        RECT 11.175000 0.765000 11.345000 0.935000 ;
      LAYER met1 ;
        RECT  7.145000 0.735000  7.900000 0.780000 ;
        RECT  7.145000 0.780000 11.405000 0.920000 ;
        RECT  7.145000 0.920000  7.900000 0.965000 ;
        RECT 11.115000 0.735000 11.405000 0.780000 ;
        RECT 11.115000 0.920000 11.405000 0.965000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.172800 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.610000 0.710000 4.955000 1.700000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.467400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.585000 1.070000 1.990000 1.335000 ;
        RECT 1.585000 1.335000 2.220000 1.745000 ;
    END
  END SCE
  PIN VGND
    ANTENNADIFFAREA  1.778050 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.720000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  2.035000  0.085000  2.415000 0.560000 ;
        RECT  2.655000  0.085000  3.035000 0.825000 ;
        RECT  5.005000  0.085000  5.350000 0.540000 ;
        RECT  7.690000  0.085000  8.020000 0.545000 ;
        RECT 10.110000  0.085000 10.330000 0.525000 ;
        RECT 12.325000  0.085000 12.655000 0.485000 ;
        RECT 13.440000  0.085000 13.610000 0.825000 ;
        RECT 14.375000  0.085000 14.545000 0.930000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.720000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.269200 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 14.720000 2.805000 ;
        RECT  0.530000 2.135000  0.910000 2.635000 ;
        RECT  2.600000 2.255000  2.930000 2.635000 ;
        RECT  4.855000 2.275000  5.205000 2.635000 ;
        RECT  7.135000 2.355000  7.465000 2.635000 ;
        RECT  8.150000 2.175000  8.570000 2.635000 ;
        RECT 10.415000 2.195000 10.665000 2.635000 ;
        RECT 11.255000 2.255000 11.635000 2.635000 ;
        RECT 12.255000 2.205000 12.715000 2.635000 ;
        RECT 13.270000 2.255000 13.725000 2.635000 ;
        RECT 14.375000 1.495000 14.625000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
        RECT 14.405000 2.635000 14.575000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 14.720000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.090000 1.795000  0.915000 1.965000 ;
      RECT  0.090000 1.965000  0.345000 2.465000 ;
      RECT  0.095000 0.345000  0.345000 0.635000 ;
      RECT  0.095000 0.635000  0.885000 0.805000 ;
      RECT  0.710000 0.805000  0.885000 0.995000 ;
      RECT  0.710000 0.995000  1.025000 1.325000 ;
      RECT  0.710000 1.325000  0.915000 1.795000 ;
      RECT  1.115000 0.345000  1.365000 0.675000 ;
      RECT  1.135000 1.730000  1.365000 2.465000 ;
      RECT  1.195000 0.675000  1.365000 1.730000 ;
      RECT  1.695000 0.395000  1.865000 0.730000 ;
      RECT  1.695000 0.730000  2.435000 0.900000 ;
      RECT  2.110000 1.915000  2.730000 2.085000 ;
      RECT  2.110000 2.085000  2.380000 2.400000 ;
      RECT  2.265000 0.900000  2.435000 0.995000 ;
      RECT  2.265000 0.995000  3.445000 1.165000 ;
      RECT  2.475000 1.165000  3.445000 1.185000 ;
      RECT  2.475000 1.185000  2.730000 1.915000 ;
      RECT  3.275000 0.255000  4.435000 0.425000 ;
      RECT  3.275000 0.425000  3.445000 0.995000 ;
      RECT  3.665000 0.675000  4.045000 1.075000 ;
      RECT  3.870000 1.075000  4.045000 1.935000 ;
      RECT  3.870000 1.935000  5.650000 2.105000 ;
      RECT  3.870000 2.105000  4.040000 2.465000 ;
      RECT  4.265000 0.425000  4.435000 1.685000 ;
      RECT  5.140000 0.715000  5.720000 0.895000 ;
      RECT  5.140000 0.895000  5.310000 1.935000 ;
      RECT  5.480000 1.065000  5.650000 1.395000 ;
      RECT  5.480000 2.105000  5.650000 2.185000 ;
      RECT  5.480000 2.185000  5.850000 2.435000 ;
      RECT  5.550000 0.335000  5.890000 0.505000 ;
      RECT  5.550000 0.505000  5.720000 0.715000 ;
      RECT  5.820000 1.575000  6.120000 1.955000 ;
      RECT  5.900000 0.705000  6.650000 1.035000 ;
      RECT  5.900000 1.035000  6.120000 1.575000 ;
      RECT  6.095000 2.135000  6.460000 2.465000 ;
      RECT  6.110000 0.305000  7.010000 0.475000 ;
      RECT  6.290000 1.215000  8.150000 1.385000 ;
      RECT  6.290000 1.385000  6.460000 2.135000 ;
      RECT  6.680000 1.935000  7.940000 2.105000 ;
      RECT  6.680000 2.105000  6.850000 2.375000 ;
      RECT  6.840000 0.475000  7.010000 1.215000 ;
      RECT  6.960000 1.595000  8.540000 1.765000 ;
      RECT  7.770000 2.105000  7.940000 2.375000 ;
      RECT  7.980000 1.005000  8.150000 1.215000 ;
      RECT  8.230000 0.275000  8.610000 0.445000 ;
      RECT  8.230000 0.445000  8.540000 0.835000 ;
      RECT  8.230000 1.765000  8.540000 1.835000 ;
      RECT  8.230000 1.835000  8.985000 2.005000 ;
      RECT  8.370000 0.835000  8.540000 1.595000 ;
      RECT  8.710000 0.705000  8.970000 1.495000 ;
      RECT  8.710000 1.495000  9.445000 1.660000 ;
      RECT  8.710000 1.660000  9.845000 1.665000 ;
      RECT  8.780000 0.255000  9.890000 0.535000 ;
      RECT  8.815000 2.005000  8.985000 2.465000 ;
      RECT  9.185000 1.665000  9.845000 1.955000 ;
      RECT  9.195000 2.125000 10.215000 2.465000 ;
      RECT  9.235000 0.920000  9.405000 1.325000 ;
      RECT  9.670000 0.535000  9.890000 1.315000 ;
      RECT  9.670000 1.315000 10.285000 1.485000 ;
      RECT 10.040000 1.485000 10.285000 1.575000 ;
      RECT 10.040000 1.575000 11.370000 1.745000 ;
      RECT 10.040000 1.745000 10.215000 2.125000 ;
      RECT 10.150000 0.695000 10.730000 0.865000 ;
      RECT 10.150000 0.865000 10.370000 1.145000 ;
      RECT 10.560000 0.295000 11.730000 0.465000 ;
      RECT 10.560000 0.465000 10.730000 0.695000 ;
      RECT 10.910000 1.915000 11.730000 2.085000 ;
      RECT 10.910000 2.085000 11.080000 2.375000 ;
      RECT 11.560000 0.465000 11.730000 0.995000 ;
      RECT 11.560000 0.995000 12.205000 1.325000 ;
      RECT 11.560000 1.325000 11.730000 1.915000 ;
      RECT 11.900000 0.345000 12.070000 0.655000 ;
      RECT 11.900000 0.655000 12.640000 0.825000 ;
      RECT 11.900000 1.795000 12.640000 1.865000 ;
      RECT 11.900000 1.865000 13.600000 2.035000 ;
      RECT 11.900000 2.035000 12.075000 2.465000 ;
      RECT 12.465000 0.825000 12.640000 1.795000 ;
      RECT 13.430000 0.995000 13.865000 1.325000 ;
      RECT 13.430000 1.325000 13.600000 1.865000 ;
    LAYER mcon ;
      RECT 0.855000 1.105000 1.025000 1.275000 ;
      RECT 1.135000 1.785000 1.305000 1.955000 ;
      RECT 5.480000 1.105000 5.650000 1.275000 ;
      RECT 5.950000 1.785000 6.120000 1.955000 ;
      RECT 9.235000 1.105000 9.405000 1.275000 ;
      RECT 9.565000 1.785000 9.735000 1.955000 ;
    LAYER met1 ;
      RECT 0.795000 1.075000 1.085000 1.120000 ;
      RECT 0.795000 1.120000 9.465000 1.260000 ;
      RECT 0.795000 1.260000 1.085000 1.305000 ;
      RECT 1.070000 1.755000 1.370000 1.800000 ;
      RECT 1.070000 1.800000 9.795000 1.940000 ;
      RECT 1.070000 1.940000 1.370000 1.985000 ;
      RECT 5.420000 1.075000 5.710000 1.120000 ;
      RECT 5.420000 1.260000 5.710000 1.305000 ;
      RECT 5.890000 1.755000 6.180000 1.800000 ;
      RECT 5.890000 1.940000 6.180000 1.985000 ;
      RECT 9.155000 1.075000 9.465000 1.120000 ;
      RECT 9.155000 1.260000 9.465000 1.305000 ;
      RECT 9.500000 1.755000 9.795000 1.800000 ;
      RECT 9.500000 1.940000 9.795000 1.985000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfrbp_2
