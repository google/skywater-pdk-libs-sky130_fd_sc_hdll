* NGSPICE file created from sky130_fd_sc_hdll__clkbuf_6.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkbuf_6 A VGND VNB VPB VPWR X
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=1.41e+12p pd=1.282e+07u as=8.7e+11p ps=7.74e+06u
M1001 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1002 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND A a_117_297# VNB nshort w=420000u l=150000u
+  ad=7.245e+11p pd=7.65e+06u as=1.134e+11p ps=1.38e+06u
M1005 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=3.423e+11p pd=4.15e+06u as=0p ps=0u
M1006 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_117_297# A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND a_117_297# X VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

