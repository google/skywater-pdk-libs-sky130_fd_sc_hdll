* File: sky130_fd_sc_hdll__o21bai_2.spice
* Created: Thu Aug 27 19:20:03 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21bai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o21bai_2  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1003 N_A_28_297#_M1003_d N_B1_N_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_A_226_47#_M1001_d N_A_28_297#_M1001_g N_Y_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.27625 AS=0.104 PD=2.15 PS=0.97 NRD=29.532 NRS=0 M=1 R=4.33333
+ SA=75000.3 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_226_47#_M1002_d N_A_28_297#_M1002_g N_Y_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1006 N_A_226_47#_M1002_d N_A2_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1012 N_A_226_47#_M1012_d N_A2_M1012_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.8
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1000 N_A_226_47#_M1012_d N_A1_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_A_226_47#_M1008_d N_A1_M1008_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.182 AS=0.12025 PD=1.86 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_VPWR_M1004_d N_B1_N_M1004_g N_A_28_297#_M1004_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=75.1752 NRS=0 M=1
+ R=2.33333 SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1004_d N_A_28_297#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.145 PD=1.90845 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_28_297#_M1009_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1011 N_A_437_297#_M1011_d N_A2_M1011_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_A_437_297#_M1013_d N_A2_M1013_g N_Y_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1007 N_A_437_297#_M1013_d N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_437_297#_M1010_d N_A1_M1010_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_12 B1_N B1_N PROBETYPE=1
pX16_noxref noxref_13 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21bai_2.pxi.spice"
*
.ends
*
*
