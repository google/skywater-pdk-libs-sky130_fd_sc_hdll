* File: sky130_fd_sc_hdll__and2b_4.pxi.spice
* Created: Thu Aug 27 18:57:47 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2B_4%A_33_199# N_A_33_199#_M1006_d
+ N_A_33_199#_M1010_d N_A_33_199#_c_57_n N_A_33_199#_M1005_g N_A_33_199#_c_58_n
+ N_A_33_199#_M1008_g N_A_33_199#_c_62_n N_A_33_199#_c_63_n N_A_33_199#_c_93_p
+ N_A_33_199#_c_59_n N_A_33_199#_c_60_n PM_SKY130_FD_SC_HDLL__AND2B_4%A_33_199#
x_PM_SKY130_FD_SC_HDLL__AND2B_4%B N_B_c_119_n N_B_M1003_g N_B_c_120_n
+ N_B_M1000_g B N_B_c_121_n PM_SKY130_FD_SC_HDLL__AND2B_4%B
x_PM_SKY130_FD_SC_HDLL__AND2B_4%A_27_47# N_A_27_47#_M1008_s N_A_27_47#_M1005_d
+ N_A_27_47#_c_149_n N_A_27_47#_M1002_g N_A_27_47#_c_158_n N_A_27_47#_M1001_g
+ N_A_27_47#_c_150_n N_A_27_47#_M1004_g N_A_27_47#_c_159_n N_A_27_47#_M1007_g
+ N_A_27_47#_c_151_n N_A_27_47#_M1009_g N_A_27_47#_c_160_n N_A_27_47#_M1011_g
+ N_A_27_47#_c_161_n N_A_27_47#_M1013_g N_A_27_47#_c_152_n N_A_27_47#_M1012_g
+ N_A_27_47#_c_153_n N_A_27_47#_c_154_n N_A_27_47#_c_172_n N_A_27_47#_c_173_n
+ N_A_27_47#_c_155_n N_A_27_47#_c_156_n N_A_27_47#_c_163_n N_A_27_47#_c_157_n
+ PM_SKY130_FD_SC_HDLL__AND2B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND2B_4%A_N N_A_N_c_263_n N_A_N_M1010_g N_A_N_c_264_n
+ N_A_N_M1006_g A_N PM_SKY130_FD_SC_HDLL__AND2B_4%A_N
x_PM_SKY130_FD_SC_HDLL__AND2B_4%VPWR N_VPWR_M1005_s N_VPWR_M1000_d
+ N_VPWR_M1007_d N_VPWR_M1013_d N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_296_n
+ N_VPWR_c_297_n N_VPWR_c_298_n N_VPWR_c_299_n N_VPWR_c_300_n VPWR
+ N_VPWR_c_301_n N_VPWR_c_293_n N_VPWR_c_303_n N_VPWR_c_304_n
+ PM_SKY130_FD_SC_HDLL__AND2B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2B_4%X N_X_M1002_s N_X_M1009_s N_X_M1001_s
+ N_X_M1011_s N_X_c_354_n N_X_c_360_n N_X_c_355_n X N_X_c_370_n X
+ PM_SKY130_FD_SC_HDLL__AND2B_4%X
x_PM_SKY130_FD_SC_HDLL__AND2B_4%VGND N_VGND_M1003_d N_VGND_M1004_d
+ N_VGND_M1012_d N_VGND_c_401_n N_VGND_c_402_n N_VGND_c_403_n N_VGND_c_404_n
+ VGND N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n
+ N_VGND_c_409_n PM_SKY130_FD_SC_HDLL__AND2B_4%VGND
cc_1 VNB N_A_33_199#_c_57_n 0.0350476f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_33_199#_c_58_n 0.0216244f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A_33_199#_c_59_n 0.0206663f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.68
cc_4 VNB N_A_33_199#_c_60_n 0.0111949f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_5 VNB N_B_c_119_n 0.0175219f $X=-0.19 $Y=-0.24 $X2=3.63 $Y2=0.465
cc_6 VNB N_B_c_120_n 0.0243247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_121_n 0.00399631f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_8 VNB N_A_27_47#_c_149_n 0.0178199f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_A_27_47#_c_150_n 0.0169022f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.325
cc_10 VNB N_A_27_47#_c_151_n 0.016912f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.68
cc_11 VNB N_A_27_47#_c_152_n 0.0186874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_153_n 0.00980077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_154_n 0.0143075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_155_n 0.00118228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_156_n 0.00185646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_157_n 0.0766183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_N_c_263_n 0.0273411f $X=-0.19 $Y=-0.24 $X2=3.63 $Y2=0.465
cc_18 VNB N_A_N_c_264_n 0.0213062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB A_N 0.00272024f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_20 VNB N_VPWR_c_293_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_401_n 0.00507933f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_22 VNB N_VGND_c_402_n 0.0173771f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.915
cc_23 VNB N_VGND_c_403_n 0.0135958f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=2
cc_24 VNB N_VGND_c_404_n 0.0137344f $X=-0.19 $Y=-0.24 $X2=3.832 $Y2=1.915
cc_25 VNB N_VGND_c_405_n 0.029662f $X=-0.19 $Y=-0.24 $X2=0.34 $Y2=1.16
cc_26 VNB N_VGND_c_406_n 0.0245003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_407_n 0.232568f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_408_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_409_n 0.0053874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_A_33_199#_c_57_n 0.032854f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_31 VPB N_A_33_199#_c_62_n 0.00695362f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.915
cc_32 VPB N_A_33_199#_c_63_n 0.0192746f $X=-0.19 $Y=1.305 $X2=3.725 $Y2=2
cc_33 VPB N_A_33_199#_c_59_n 0.00930852f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.68
cc_34 VPB N_A_33_199#_c_60_n 6.88357e-19 $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_35 VPB N_B_c_120_n 0.0274062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_B_c_121_n 0.00200146f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_37 VPB N_A_27_47#_c_158_n 0.0173633f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_38 VPB N_A_27_47#_c_159_n 0.0160428f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=2
cc_39 VPB N_A_27_47#_c_160_n 0.0157532f $X=-0.19 $Y=1.305 $X2=3.815 $Y2=1.695
cc_40 VPB N_A_27_47#_c_161_n 0.0177229f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_41 VPB N_A_27_47#_c_156_n 0.0031409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_163_n 0.00344008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_157_n 0.0482382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_N_c_263_n 0.0291439f $X=-0.19 $Y=1.305 $X2=3.63 $Y2=0.465
cc_45 VPB A_N 0.00116764f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_46 VPB N_VPWR_c_294_n 0.0102988f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.325
cc_47 VPB N_VPWR_c_295_n 0.0134185f $X=-0.19 $Y=1.305 $X2=3.725 $Y2=2
cc_48 VPB N_VPWR_c_296_n 0.0171055f $X=-0.19 $Y=1.305 $X2=3.832 $Y2=1.915
cc_49 VPB N_VPWR_c_297_n 0.00451311f $X=-0.19 $Y=1.305 $X2=3.832 $Y2=1.695
cc_50 VPB N_VPWR_c_298_n 0.0163056f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.16
cc_51 VPB N_VPWR_c_299_n 0.0167956f $X=-0.19 $Y=1.305 $X2=0.34 $Y2=1.16
cc_52 VPB N_VPWR_c_300_n 0.0132269f $X=-0.19 $Y=1.305 $X2=0.38 $Y2=1.16
cc_53 VPB N_VPWR_c_301_n 0.0239901f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_293_n 0.0538337f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_303_n 0.00631318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_304_n 0.00538144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 N_A_33_199#_c_58_n N_B_c_119_n 0.0384605f $X=0.52 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_58 N_A_33_199#_c_57_n N_B_c_120_n 0.0803275f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_33_199#_c_63_n N_B_c_120_n 0.0139886f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_60 N_A_33_199#_c_60_n N_B_c_120_n 2.24934e-19 $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_33_199#_c_57_n N_B_c_121_n 0.00282251f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_33_199#_c_60_n N_B_c_121_n 0.0253934f $X=0.34 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_33_199#_c_63_n N_A_27_47#_M1005_d 0.00493291f $X=3.725 $Y=2 $X2=0
+ $Y2=0
cc_64 N_A_33_199#_c_63_n N_A_27_47#_c_158_n 0.0164781f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_65 N_A_33_199#_c_63_n N_A_27_47#_c_159_n 0.0131214f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_66 N_A_33_199#_c_63_n N_A_27_47#_c_160_n 0.0133589f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_67 N_A_33_199#_c_63_n N_A_27_47#_c_161_n 0.0163925f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_68 N_A_33_199#_c_57_n N_A_27_47#_c_153_n 0.0059209f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_69 N_A_33_199#_c_60_n N_A_27_47#_c_153_n 0.0178872f $X=0.34 $Y=1.16 $X2=0
+ $Y2=0
cc_70 N_A_33_199#_c_58_n N_A_27_47#_c_172_n 0.0143005f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_71 N_A_33_199#_c_57_n N_A_27_47#_c_173_n 0.00773972f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_72 N_A_33_199#_c_62_n N_A_27_47#_c_173_n 0.018267f $X=0.25 $Y=1.915 $X2=0
+ $Y2=0
cc_73 N_A_33_199#_c_63_n N_A_27_47#_c_173_n 0.0403997f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_74 N_A_33_199#_c_63_n N_A_27_47#_c_156_n 0.012382f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_75 N_A_33_199#_c_63_n N_A_27_47#_c_163_n 0.00471602f $X=3.725 $Y=2 $X2=0
+ $Y2=0
cc_76 N_A_33_199#_c_63_n N_A_27_47#_c_157_n 7.05723e-19 $X=3.725 $Y=2 $X2=0
+ $Y2=0
cc_77 N_A_33_199#_c_63_n N_A_N_c_263_n 0.0144444f $X=3.725 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_33_199#_c_59_n N_A_N_c_263_n 0.00640745f $X=3.81 $Y=0.68 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_33_199#_c_59_n N_A_N_c_264_n 0.016013f $X=3.81 $Y=0.68 $X2=0 $Y2=0
cc_80 N_A_33_199#_c_63_n A_N 0.0249218f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_81 N_A_33_199#_c_59_n A_N 0.0815607f $X=3.81 $Y=0.68 $X2=0 $Y2=0
cc_82 N_A_33_199#_c_62_n N_VPWR_M1005_s 0.0231796f $X=0.25 $Y=1.915 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_33_199#_c_63_n N_VPWR_M1005_s 3.13877e-19 $X=3.725 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_33_199#_c_93_p N_VPWR_M1005_s 0.0100218f $X=0.335 $Y=2 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_33_199#_c_63_n N_VPWR_M1000_d 0.00615695f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_86 N_A_33_199#_c_63_n N_VPWR_M1007_d 0.00359344f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_87 N_A_33_199#_c_63_n N_VPWR_M1013_d 0.00721553f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_88 N_A_33_199#_c_57_n N_VPWR_c_295_n 0.00975695f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_33_199#_c_63_n N_VPWR_c_295_n 0.00227506f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_90 N_A_33_199#_c_93_p N_VPWR_c_295_n 0.0142454f $X=0.335 $Y=2 $X2=0 $Y2=0
cc_91 N_A_33_199#_c_57_n N_VPWR_c_296_n 0.00452725f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_33_199#_c_63_n N_VPWR_c_296_n 0.0100826f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_93 N_A_33_199#_c_63_n N_VPWR_c_297_n 0.019066f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_94 N_A_33_199#_c_63_n N_VPWR_c_298_n 0.00970145f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_95 N_A_33_199#_c_63_n N_VPWR_c_299_n 0.0218583f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_96 N_A_33_199#_c_63_n N_VPWR_c_300_n 0.00861424f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_97 N_A_33_199#_c_63_n N_VPWR_c_301_n 0.0107325f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_98 N_A_33_199#_c_57_n N_VPWR_c_293_n 0.00520867f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_33_199#_c_63_n N_VPWR_c_293_n 0.0700575f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_100 N_A_33_199#_c_93_p N_VPWR_c_293_n 8.51964e-19 $X=0.335 $Y=2 $X2=0 $Y2=0
cc_101 N_A_33_199#_c_63_n N_VPWR_c_304_n 0.0177358f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_102 N_A_33_199#_c_63_n N_X_M1001_s 0.00559492f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_103 N_A_33_199#_c_63_n N_X_M1011_s 0.00477619f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_104 N_A_33_199#_c_63_n N_X_c_354_n 0.0425914f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_105 N_A_33_199#_c_63_n N_X_c_355_n 0.0328136f $X=3.725 $Y=2 $X2=0 $Y2=0
cc_106 N_A_33_199#_c_58_n N_VGND_c_405_n 0.00422112f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_A_33_199#_c_59_n N_VGND_c_406_n 0.00576054f $X=3.81 $Y=0.68 $X2=0 $Y2=0
cc_108 N_A_33_199#_c_58_n N_VGND_c_407_n 0.00665063f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_109 N_A_33_199#_c_59_n N_VGND_c_407_n 0.00708776f $X=3.81 $Y=0.68 $X2=0 $Y2=0
cc_110 N_B_c_119_n N_A_27_47#_c_149_n 0.0195615f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_c_120_n N_A_27_47#_c_158_n 0.0317612f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_119_n N_A_27_47#_c_172_n 0.0130948f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_120_n N_A_27_47#_c_172_n 0.00478288f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_121_n N_A_27_47#_c_172_n 0.0271044f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_115 N_B_c_120_n N_A_27_47#_c_173_n 0.0153421f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B_c_121_n N_A_27_47#_c_173_n 0.0309331f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B_c_119_n N_A_27_47#_c_155_n 0.00381579f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B_c_120_n N_A_27_47#_c_156_n 0.00672893f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B_c_121_n N_A_27_47#_c_156_n 0.0284819f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_c_120_n N_A_27_47#_c_157_n 0.0144946f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B_c_121_n N_A_27_47#_c_157_n 2.81641e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_122 N_B_c_120_n N_VPWR_c_295_n 0.00115542f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B_c_120_n N_VPWR_c_296_n 0.00510113f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_c_120_n N_VPWR_c_297_n 0.00307218f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B_c_120_n N_VPWR_c_293_n 0.00696016f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_126 N_B_c_119_n N_VGND_c_401_n 0.0062316f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_127 N_B_c_119_n N_VGND_c_405_n 0.00422112f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B_c_119_n N_VGND_c_407_n 0.00617105f $X=0.88 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_161_n N_A_N_c_263_n 0.0188572f $X=2.975 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_27_47#_c_157_n N_A_N_c_263_n 0.0247074f $X=2.975 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_131 N_A_27_47#_c_152_n N_A_N_c_264_n 0.0141129f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_161_n A_N 0.00277927f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_152_n A_N 0.00636928f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_173_n N_VPWR_M1000_d 0.00644594f $X=1.245 $Y=1.622 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_156_n N_VPWR_M1000_d 0.00338093f $X=1.455 $Y=1.175 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_158_n N_VPWR_c_297_n 0.00181033f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_27_47#_c_158_n N_VPWR_c_298_n 0.00510113f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_c_159_n N_VPWR_c_298_n 0.00311736f $X=2.035 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_27_47#_c_160_n N_VPWR_c_299_n 0.00112257f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_c_161_n N_VPWR_c_299_n 0.0117289f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_27_47#_c_160_n N_VPWR_c_300_n 0.00453434f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_161_n N_VPWR_c_300_n 0.00311736f $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1005_d N_VPWR_c_293_n 0.00338665f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_c_158_n N_VPWR_c_293_n 0.00693233f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_c_159_n N_VPWR_c_293_n 0.00383364f $X=2.035 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_c_160_n N_VPWR_c_293_n 0.00518254f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_161_n N_VPWR_c_293_n 0.00375605f $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_158_n N_VPWR_c_304_n 0.00115604f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_c_159_n N_VPWR_c_304_n 0.0111217f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_160_n N_VPWR_c_304_n 0.00785399f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_c_161_n N_VPWR_c_304_n 0.00100747f $X=2.975 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_159_n N_X_c_354_n 0.0110852f $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_160_n N_X_c_354_n 0.0048427f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_163_n N_X_c_354_n 0.0344279f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_157_n N_X_c_354_n 0.00963857f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_172_n N_X_c_360_n 0.0123227f $X=1.245 $Y=0.71 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_155_n N_X_c_360_n 0.00115157f $X=1.35 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_163_n N_X_c_360_n 0.0145204f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_157_n N_X_c_360_n 0.00339703f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_160_n N_X_c_355_n 0.00509181f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_161_n N_X_c_355_n 0.00491661f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_150_n X 0.0108646f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_151_n X 0.00676743f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_163_n X 0.018991f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_157_n X 0.00544676f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_151_n N_X_c_370_n 0.00416118f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_152_n N_X_c_370_n 0.00415234f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_150_n X 9.16455e-19 $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_159_n X 7.29709e-19 $X=2.035 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_151_n X 0.0059288f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_160_n X 0.00450101f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_161_n X 0.00299019f $X=2.975 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_152_n X 0.00391765f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_163_n X 0.0205613f $X=1.985 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_157_n X 0.0420653f $X=2.975 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_172_n A_119_47# 0.00271764f $X=1.245 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_27_47#_c_172_n N_VGND_M1003_d 0.0110607f $X=1.245 $Y=0.71 $X2=-0.19
+ $Y2=-0.24
cc_178 N_A_27_47#_c_155_n N_VGND_M1003_d 0.00103313f $X=1.35 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_27_47#_c_149_n N_VGND_c_401_n 0.00321931f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_172_n N_VGND_c_401_n 0.0255338f $X=1.245 $Y=0.71 $X2=0 $Y2=0
cc_181 N_A_27_47#_c_149_n N_VGND_c_402_n 0.00563595f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_150_n N_VGND_c_402_n 0.0033769f $X=1.99 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_172_n N_VGND_c_402_n 8.83096e-19 $X=1.245 $Y=0.71 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_151_n N_VGND_c_403_n 0.00116335f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_152_n N_VGND_c_403_n 0.0149575f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_151_n N_VGND_c_404_n 0.0036573f $X=2.47 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_152_n N_VGND_c_404_n 0.00213258f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_154_n N_VGND_c_405_n 0.0218999f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_172_n N_VGND_c_405_n 0.0096965f $X=1.245 $Y=0.71 $X2=0 $Y2=0
cc_190 N_A_27_47#_M1008_s N_VGND_c_407_n 0.00255893f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_149_n N_VGND_c_407_n 0.0106573f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_150_n N_VGND_c_407_n 0.00410511f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_151_n N_VGND_c_407_n 0.00450312f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_152_n N_VGND_c_407_n 0.00341549f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_154_n N_VGND_c_407_n 0.0127541f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_172_n N_VGND_c_407_n 0.0203275f $X=1.245 $Y=0.71 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_149_n N_VGND_c_409_n 0.00111023f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_150_n N_VGND_c_409_n 0.00882507f $X=1.99 $Y=0.995 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_151_n N_VGND_c_409_n 0.00796296f $X=2.47 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_152_n N_VGND_c_409_n 0.00102739f $X=3 $Y=0.995 $X2=0 $Y2=0
cc_201 A_N N_VPWR_M1013_d 0.00512222f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_202 N_A_N_c_263_n N_VPWR_c_301_n 6.43543e-19 $X=3.53 $Y=1.41 $X2=0 $Y2=0
cc_203 A_N N_X_c_355_n 0.0142199f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_204 N_A_N_c_264_n N_X_c_370_n 2.0294e-19 $X=3.555 $Y=0.995 $X2=0 $Y2=0
cc_205 A_N N_X_c_370_n 0.0135427f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_206 N_A_N_c_263_n X 4.78319e-19 $X=3.53 $Y=1.41 $X2=0 $Y2=0
cc_207 A_N X 0.0478567f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_208 A_N N_VGND_M1012_d 0.00621173f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_209 N_A_N_c_263_n N_VGND_c_403_n 3.1887e-19 $X=3.53 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_N_c_264_n N_VGND_c_403_n 0.00303795f $X=3.555 $Y=0.995 $X2=0 $Y2=0
cc_211 A_N N_VGND_c_403_n 0.0138294f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_212 N_A_N_c_264_n N_VGND_c_406_n 0.00459323f $X=3.555 $Y=0.995 $X2=0 $Y2=0
cc_213 A_N N_VGND_c_406_n 0.00269856f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_214 N_A_N_c_264_n N_VGND_c_407_n 0.00512902f $X=3.555 $Y=0.995 $X2=0 $Y2=0
cc_215 A_N N_VGND_c_407_n 0.00600614f $X=3.365 $Y=1.105 $X2=0 $Y2=0
cc_216 N_VPWR_c_293_n N_X_M1001_s 0.003737f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_217 N_VPWR_c_293_n N_X_M1011_s 0.00338665f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_218 N_VPWR_M1007_d N_X_c_354_n 0.0040425f $X=2.125 $Y=1.485 $X2=0 $Y2=0
cc_219 X N_VGND_M1004_d 0.00557582f $X=2.445 $Y=0.765 $X2=3.62 $Y2=1.485
cc_220 N_X_c_360_n N_VGND_c_402_n 0.00477425f $X=1.77 $Y=0.66 $X2=0.25 $Y2=1.915
cc_221 X N_VGND_c_402_n 0.00259391f $X=2.445 $Y=0.765 $X2=0.25 $Y2=1.915
cc_222 X N_VGND_c_404_n 5.14241e-19 $X=2.445 $Y=0.765 $X2=3.832 $Y2=1.915
cc_223 N_X_c_370_n N_VGND_c_404_n 0.00944884f $X=2.712 $Y=0.825 $X2=3.832
+ $Y2=1.915
cc_224 N_X_M1002_s N_VGND_c_407_n 0.00629831f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_225 N_X_M1009_s N_VGND_c_407_n 0.00435221f $X=2.545 $Y=0.235 $X2=0 $Y2=0
cc_226 N_X_c_360_n N_VGND_c_407_n 0.00607819f $X=1.77 $Y=0.66 $X2=0 $Y2=0
cc_227 X N_VGND_c_407_n 0.00686047f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_228 N_X_c_370_n N_VGND_c_407_n 0.0155137f $X=2.712 $Y=0.825 $X2=0 $Y2=0
cc_229 X N_VGND_c_409_n 0.0199734f $X=2.445 $Y=0.765 $X2=0 $Y2=0
cc_230 A_119_47# N_VGND_c_407_n 0.00239227f $X=0.595 $Y=0.235 $X2=0.425 $Y2=0.71
