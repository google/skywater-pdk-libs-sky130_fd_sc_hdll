* File: sky130_fd_sc_hdll__sdlclkp_1.spice
* Created: Thu Aug 27 19:28:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdlclkp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sdlclkp_1  VNB VPB SCE GATE CLK VPWR GCLK VGND
* 
* VGND	VGND
* GCLK	GCLK
* VPWR	VPWR
* CLK	CLK
* GATE	GATE
* SCE	SCE
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_SCE_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.1302 PD=0.695 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.6 A=0.063 P=1.14 MULT=1
MM1021 N_A_27_47#_M1021_d N_GATE_M1021_g N_VGND_M1015_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0710769 AS=0.05775 PD=0.802308 PS=0.695 NRD=11.424 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75002.2 A=0.063 P=1.14 MULT=1
MM1014 N_A_299_47#_M1014_d N_A_269_21#_M1014_g N_A_27_47#_M1021_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0774 AS=0.0609231 PD=0.79 PS=0.687692 NRD=31.656 NRS=1.656
+ M=1 R=2.4 SA=75001.1 SB=75002 A=0.054 P=1.02 MULT=1
MM1006 A_415_47# N_A_266_243#_M1006_g N_A_299_47#_M1014_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0908308 AS=0.0774 PD=0.853846 PS=0.79 NRD=65.76 NRS=18.324 M=1
+ R=2.4 SA=75001.7 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1011 N_VGND_M1011_d N_A_484_315#_M1011_g A_415_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.102704 AS=0.105969 PD=0.859626 PS=0.996154 NRD=35.712 NRS=56.364 M=1
+ R=2.8 SA=75002.1 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1004 N_A_484_315#_M1004_d N_A_299_47#_M1004_g N_VGND_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.158946 PD=1.82 PS=1.33037 NRD=0 NRS=7.38 M=1 R=4.33333
+ SA=75001.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A_269_21#_M1019_g N_A_266_243#_M1019_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0945 AS=0.1092 PD=0.87 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75000.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_269_21#_M1007_d N_CLK_M1007_g N_VGND_M1019_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0945 PD=1.46 PS=0.87 NRD=12.852 NRS=35.712 M=1 R=2.8 SA=75000.8
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1008 A_1181_47# N_A_484_315#_M1008_g N_A_1089_47#_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0693 AS=0.1302 PD=0.75 PS=1.46 NRD=31.428 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_CLK_M1013_g A_1181_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0889065 AS=0.0693 PD=0.804673 PS=0.75 NRD=0 NRS=31.428 M=1 R=2.8
+ SA=75000.7 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1018 N_GCLK_M1018_d N_A_1089_47#_M1018_g N_VGND_M1013_d VNB NSHORT L=0.15
+ W=0.65 AD=0.18525 AS=0.137593 PD=1.87 PS=1.24533 NRD=3.684 NRS=18.456 M=1
+ R=4.33333 SA=75000.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 A_117_369# N_SCE_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.1728 PD=0.87 PS=1.82 NRD=18.4589 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1003 N_A_27_47#_M1003_d N_GATE_M1003_g A_117_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.122023 AS=0.0736 PD=1.18943 PS=0.87 NRD=18.4589 NRS=18.4589 M=1 R=3.55556
+ SA=90000.6 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1017 N_A_299_47#_M1017_d N_A_266_243#_M1017_g N_A_27_47#_M1003_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0735 AS=0.0800774 PD=0.77 PS=0.780566 NRD=16.4101
+ NRS=2.3443 M=1 R=2.33333 SA=90001.1 SB=90002 A=0.0756 P=1.2 MULT=1
MM1009 A_410_413# N_A_269_21#_M1009_g N_A_299_47#_M1017_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0798 AS=0.0735 PD=0.8 PS=0.77 NRD=63.3158 NRS=16.4101 M=1
+ R=2.33333 SA=90001.6 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_484_315#_M1010_g A_410_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.109821 AS=0.0798 PD=0.902113 PS=0.8 NRD=63.3158 NRS=63.3158 M=1 R=2.33333
+ SA=90002.2 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1000 N_A_484_315#_M1000_d N_A_299_47#_M1000_g N_VPWR_M1010_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.27 AS=0.261479 PD=2.54 PS=2.14789 NRD=0.9653 NRS=21.67 M=1
+ R=5.55556 SA=90001.3 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1020 N_VPWR_M1020_d N_A_269_21#_M1020_g N_A_266_243#_M1020_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.17565 AS=0.1728 PD=1.39 PS=1.82 NRD=67.5316 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90000.8 A=0.1152 P=1.64 MULT=1
MM1002 N_A_269_21#_M1002_d N_CLK_M1002_g N_VPWR_M1020_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.17565 PD=1.82 PS=1.39 NRD=1.5366 NRS=67.5316 M=1
+ R=3.55556 SA=90000.8 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1001 N_A_1089_47#_M1001_d N_A_484_315#_M1001_g N_VPWR_M1001_s VPB PHIGHVT
+ L=0.18 W=0.64 AD=0.096 AS=0.1728 PD=0.94 PS=1.82 NRD=1.5366 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1016 N_VPWR_M1016_d N_CLK_M1016_g N_A_1089_47#_M1001_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.122693 AS=0.096 PD=1.04976 PS=0.94 NRD=10.7562 NRS=4.6098 M=1
+ R=3.55556 SA=90000.7 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1012 N_GCLK_M1012_d N_A_1089_47#_M1012_g N_VPWR_M1016_d VPB PHIGHVT L=0.18 W=1
+ AD=0.295 AS=0.191707 PD=2.59 PS=1.64024 NRD=5.8903 NRS=5.8903 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX22_noxref VNB VPB NWDIODE A=12.4227 P=18.69
c_74 VNB 0 3.23043e-19 $X=0.15 $Y=-0.085
c_138 VPB 0 1.64862e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdlclkp_1.pxi.spice"
*
.ends
*
*
