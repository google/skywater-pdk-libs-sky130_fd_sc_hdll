* File: sky130_fd_sc_hdll__a211oi_2.pxi.spice
* Created: Thu Aug 27 18:51:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__A211OI_2%C1 N_C1_c_79_n N_C1_M1004_g N_C1_c_75_n
+ N_C1_M1012_g N_C1_c_80_n N_C1_M1011_g N_C1_c_76_n N_C1_M1014_g C1 C1
+ N_C1_c_77_n N_C1_c_78_n PM_SKY130_FD_SC_HDLL__A211OI_2%C1
x_PM_SKY130_FD_SC_HDLL__A211OI_2%B1 N_B1_c_116_n N_B1_M1001_g N_B1_c_121_n
+ N_B1_M1005_g N_B1_c_122_n N_B1_M1013_g N_B1_c_117_n N_B1_M1006_g B1 B1 B1
+ N_B1_c_119_n N_B1_c_120_n B1 PM_SKY130_FD_SC_HDLL__A211OI_2%B1
x_PM_SKY130_FD_SC_HDLL__A211OI_2%A1 N_A1_c_166_n N_A1_M1002_g N_A1_c_170_n
+ N_A1_M1003_g N_A1_c_171_n N_A1_M1015_g N_A1_c_167_n N_A1_M1007_g A1 A1
+ N_A1_c_169_n A1 A1 PM_SKY130_FD_SC_HDLL__A211OI_2%A1
x_PM_SKY130_FD_SC_HDLL__A211OI_2%A2 N_A2_c_205_n N_A2_M1009_g N_A2_c_211_n
+ N_A2_M1000_g N_A2_c_212_n N_A2_M1008_g N_A2_c_206_n N_A2_M1010_g A2 A2 A2
+ N_A2_c_209_n A2 N_A2_c_210_n PM_SKY130_FD_SC_HDLL__A211OI_2%A2
x_PM_SKY130_FD_SC_HDLL__A211OI_2%A_37_297# N_A_37_297#_M1004_s
+ N_A_37_297#_M1011_s N_A_37_297#_M1013_s N_A_37_297#_c_248_n
+ N_A_37_297#_c_255_n N_A_37_297#_c_249_n N_A_37_297#_c_259_n
+ N_A_37_297#_c_261_n N_A_37_297#_c_250_n N_A_37_297#_c_251_n
+ N_A_37_297#_c_276_p PM_SKY130_FD_SC_HDLL__A211OI_2%A_37_297#
x_PM_SKY130_FD_SC_HDLL__A211OI_2%Y N_Y_M1012_d N_Y_M1001_d N_Y_M1002_s
+ N_Y_M1004_d N_Y_c_285_n Y Y Y Y Y N_Y_c_295_n Y
+ PM_SKY130_FD_SC_HDLL__A211OI_2%Y
x_PM_SKY130_FD_SC_HDLL__A211OI_2%A_320_297# N_A_320_297#_M1005_d
+ N_A_320_297#_M1003_d N_A_320_297#_M1000_s N_A_320_297#_c_331_n
+ N_A_320_297#_c_370_p N_A_320_297#_c_332_n N_A_320_297#_c_333_n
+ N_A_320_297#_c_371_p N_A_320_297#_c_334_n N_A_320_297#_c_335_n
+ PM_SKY130_FD_SC_HDLL__A211OI_2%A_320_297#
x_PM_SKY130_FD_SC_HDLL__A211OI_2%VPWR N_VPWR_M1003_s N_VPWR_M1015_s
+ N_VPWR_M1008_d N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n
+ N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n N_VPWR_c_388_n
+ N_VPWR_c_389_n VPWR N_VPWR_c_379_n VPWR PM_SKY130_FD_SC_HDLL__A211OI_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A211OI_2%VGND N_VGND_M1012_s N_VGND_M1014_s
+ N_VGND_M1006_s N_VGND_M1009_d N_VGND_c_442_n N_VGND_c_443_n N_VGND_c_444_n
+ N_VGND_c_445_n N_VGND_c_446_n N_VGND_c_447_n N_VGND_c_448_n VGND
+ N_VGND_c_449_n N_VGND_c_450_n N_VGND_c_451_n N_VGND_c_452_n N_VGND_c_453_n
+ VGND PM_SKY130_FD_SC_HDLL__A211OI_2%VGND
x_PM_SKY130_FD_SC_HDLL__A211OI_2%A_525_47# N_A_525_47#_M1002_d
+ N_A_525_47#_M1007_d N_A_525_47#_M1010_s N_A_525_47#_c_513_n
+ N_A_525_47#_c_514_n N_A_525_47#_c_528_n N_A_525_47#_c_515_n
+ PM_SKY130_FD_SC_HDLL__A211OI_2%A_525_47#
cc_1 VNB N_C1_c_75_n 0.0220734f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=0.995
cc_2 VNB N_C1_c_76_n 0.0163511f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_3 VNB N_C1_c_77_n 0.0160237f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_4 VNB N_C1_c_78_n 0.0602555f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.202
cc_5 VNB N_B1_c_116_n 0.0171089f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.41
cc_6 VNB N_B1_c_117_n 0.0218479f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_7 VNB B1 0.00396499f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_c_119_n 0.0486756f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.16
cc_9 VNB N_B1_c_120_n 0.0014706f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.19
cc_10 VNB N_A1_c_166_n 0.0229935f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.41
cc_11 VNB N_A1_c_167_n 0.0173559f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_12 VNB A1 0.0135983f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.445
cc_13 VNB N_A1_c_169_n 0.0421546f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.202
cc_14 VNB N_A2_c_205_n 0.0171406f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.41
cc_15 VNB N_A2_c_206_n 0.0229935f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_16 VNB A2 0.00434725f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.445
cc_17 VNB A2 0.00100822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_209_n 0.043139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_210_n 0.0166807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_285_n 0.00946905f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.202
cc_21 VNB Y 0.00109007f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.202
cc_22 VNB N_VPWR_c_379_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_442_n 0.011635f $X=-0.19 $Y=-0.24 $X2=0.125 $Y2=1.105
cc_24 VNB N_VGND_c_443_n 0.0266241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_444_n 3.38371e-19 $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_26 VNB N_VGND_c_445_n 0.0138317f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.202
cc_27 VNB N_VGND_c_446_n 0.00547462f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_447_n 0.0092224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_448_n 0.0364432f $X=-0.19 $Y=-0.24 $X2=0.252 $Y2=1.53
cc_30 VNB N_VGND_c_449_n 0.0161159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_450_n 0.0212876f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_451_n 0.267118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_452_n 0.00502699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_453_n 0.00576672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_525_47#_c_513_n 0.00254857f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=0.995
cc_36 VNB N_A_525_47#_c_514_n 0.00965734f $X=-0.19 $Y=-0.24 $X2=0.315 $Y2=1.16
cc_37 VNB N_A_525_47#_c_515_n 0.0141126f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.202
cc_38 VPB N_C1_c_79_n 0.0188939f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.41
cc_39 VPB N_C1_c_80_n 0.0161239f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_40 VPB N_C1_c_77_n 0.0148901f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_41 VPB N_C1_c_78_n 0.0312859f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.202
cc_42 VPB N_B1_c_121_n 0.0164342f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=0.995
cc_43 VPB N_B1_c_122_n 0.0204212f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_44 VPB B1 0.00165019f $X=-0.19 $Y=1.305 $X2=0.125 $Y2=1.445
cc_45 VPB N_B1_c_119_n 0.023333f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.16
cc_46 VPB N_A1_c_170_n 0.0204263f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=0.995
cc_47 VPB N_A1_c_171_n 0.0162669f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_48 VPB N_A1_c_169_n 0.0230636f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.202
cc_49 VPB N_A2_c_211_n 0.0162661f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=0.995
cc_50 VPB N_A2_c_212_n 0.0192854f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.41
cc_51 VPB A2 0.0211052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A2_c_209_n 0.0210485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_37_297#_c_248_n 0.0191356f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=0.56
cc_54 VPB N_A_37_297#_c_249_n 0.00746418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_37_297#_c_250_n 0.00246231f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.202
cc_56 VPB N_A_37_297#_c_251_n 0.00474692f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.16
cc_57 VPB Y 9.28314e-19 $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_58 VPB N_A_320_297#_c_331_n 0.0225472f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=0.56
cc_59 VPB N_A_320_297#_c_332_n 0.00577699f $X=-0.19 $Y=1.305 $X2=0.315 $Y2=1.16
cc_60 VPB N_A_320_297#_c_333_n 0.00193259f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_61 VPB N_A_320_297#_c_334_n 0.00180652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_320_297#_c_335_n 0.00163082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_380_n 0.00506779f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=0.56
cc_64 VPB N_VPWR_c_381_n 0.00505418f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_382_n 0.00506779f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.202
cc_66 VPB N_VPWR_c_383_n 0.0650797f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.202
cc_67 VPB N_VPWR_c_384_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.16
cc_68 VPB N_VPWR_c_385_n 0.0206452f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.19
cc_69 VPB N_VPWR_c_386_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_387_n 0.0108943f $X=-0.19 $Y=1.305 $X2=0.252 $Y2=1.53
cc_71 VPB N_VPWR_c_388_n 0.0206452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_389_n 0.0043981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_379_n 0.0621476f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_C1_c_76_n N_B1_c_116_n 0.0220982f $X=1.055 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_75 N_C1_c_80_n N_B1_c_121_n 0.0191741f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_76 N_C1_c_80_n B1 0.00599068f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_77 N_C1_c_78_n B1 0.00316171f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_78 N_C1_c_78_n N_B1_c_119_n 0.0220982f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_79 N_C1_c_78_n N_B1_c_120_n 0.00909282f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_80 N_C1_c_77_n N_A_37_297#_M1004_s 0.00369033f $X=0.315 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_81 N_C1_c_77_n N_A_37_297#_c_248_n 0.0231249f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C1_c_78_n N_A_37_297#_c_248_n 9.3647e-19 $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_83 N_C1_c_79_n N_A_37_297#_c_255_n 0.0125412f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_84 N_C1_c_80_n N_A_37_297#_c_255_n 0.0136838f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_85 N_C1_c_76_n N_Y_c_285_n 0.0125668f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_86 N_C1_c_79_n Y 0.0171663f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_87 N_C1_c_75_n Y 0.0119991f $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_88 N_C1_c_80_n Y 5.95065e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_89 N_C1_c_76_n Y 0.00355601f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_90 N_C1_c_77_n Y 0.0418879f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_91 N_C1_c_78_n Y 0.0317806f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_92 N_C1_c_75_n N_Y_c_295_n 0.00631582f $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_93 N_C1_c_80_n N_A_320_297#_c_334_n 6.96116e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_94 N_C1_c_79_n N_VPWR_c_383_n 0.00431957f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C1_c_80_n N_VPWR_c_383_n 0.00431957f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_96 N_C1_c_79_n N_VPWR_c_379_n 0.00705273f $X=0.55 $Y=1.41 $X2=0 $Y2=0
cc_97 N_C1_c_80_n N_VPWR_c_379_n 0.00614289f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_98 N_C1_c_75_n N_VGND_c_443_n 0.00805774f $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_99 N_C1_c_77_n N_VGND_c_443_n 0.0208132f $X=0.315 $Y=1.16 $X2=0 $Y2=0
cc_100 N_C1_c_78_n N_VGND_c_443_n 0.00168116f $X=1.03 $Y=1.202 $X2=0 $Y2=0
cc_101 N_C1_c_75_n N_VGND_c_444_n 5.29225e-19 $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_102 N_C1_c_76_n N_VGND_c_444_n 0.00977288f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_103 N_C1_c_75_n N_VGND_c_449_n 0.00473044f $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_104 N_C1_c_76_n N_VGND_c_449_n 0.00213283f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C1_c_75_n N_VGND_c_451_n 0.00926759f $X=0.575 $Y=0.995 $X2=0 $Y2=0
cc_106 N_C1_c_76_n N_VGND_c_451_n 0.00289592f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_107 B1 N_A_37_297#_M1011_s 0.00244039f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_108 B1 N_A_37_297#_c_255_n 0.00127477f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_109 B1 N_A_37_297#_c_259_n 0.00952426f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_110 B1 N_A_37_297#_c_259_n 0.00304501f $X=1.655 $Y=1.105 $X2=0 $Y2=0
cc_111 N_B1_c_121_n N_A_37_297#_c_261_n 0.0135559f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B1_c_122_n N_A_37_297#_c_261_n 0.012175f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_116_n N_Y_c_285_n 0.0104488f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_114 N_B1_c_117_n N_Y_c_285_n 0.0143939f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_115 B1 N_Y_c_285_n 0.0396446f $X=1.655 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B1_c_119_n N_Y_c_285_n 0.00468889f $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_117 N_B1_c_120_n N_Y_c_285_n 0.0150107f $X=1.175 $Y=1.285 $X2=0 $Y2=0
cc_118 B1 Y 0.0196438f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_119 N_B1_c_119_n Y 3.38724e-19 $X=1.99 $Y=1.202 $X2=0 $Y2=0
cc_120 N_B1_c_120_n Y 0.0199119f $X=1.175 $Y=1.285 $X2=0 $Y2=0
cc_121 N_B1_c_122_n N_A_320_297#_c_331_n 0.0166106f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_122 B1 N_A_320_297#_c_331_n 0.0013794f $X=1.655 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B1_c_119_n N_A_320_297#_c_331_n 3.63008e-19 $X=1.99 $Y=1.202 $X2=0
+ $Y2=0
cc_124 N_B1_c_121_n N_A_320_297#_c_334_n 0.0125099f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_c_122_n N_A_320_297#_c_334_n 0.0117074f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_126 B1 N_A_320_297#_c_334_n 0.00954721f $X=1.075 $Y=1.445 $X2=0 $Y2=0
cc_127 B1 N_A_320_297#_c_334_n 0.0308488f $X=1.655 $Y=1.105 $X2=0 $Y2=0
cc_128 N_B1_c_119_n N_A_320_297#_c_334_n 0.00777503f $X=1.99 $Y=1.202 $X2=0
+ $Y2=0
cc_129 N_B1_c_122_n N_VPWR_c_380_n 0.00219083f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B1_c_121_n N_VPWR_c_383_n 0.00431957f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_131 N_B1_c_122_n N_VPWR_c_383_n 0.00431957f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B1_c_121_n N_VPWR_c_379_n 0.00614289f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_133 N_B1_c_122_n N_VPWR_c_379_n 0.00737633f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B1_c_116_n N_VGND_c_444_n 0.00856001f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B1_c_117_n N_VGND_c_444_n 0.00112959f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B1_c_116_n N_VGND_c_445_n 0.00355956f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B1_c_117_n N_VGND_c_445_n 0.00213283f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B1_c_116_n N_VGND_c_446_n 0.00125169f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_139 N_B1_c_117_n N_VGND_c_446_n 0.0125705f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_140 N_B1_c_116_n N_VGND_c_451_n 0.0044447f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B1_c_117_n N_VGND_c_451_n 0.0030623f $X=2.015 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_167_n N_A2_c_205_n 0.0221649f $X=3.495 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A1_c_171_n N_A2_c_211_n 0.0224695f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_144 A1 A2 0.0125963f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A1_c_169_n A2 2.9421e-19 $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_146 A1 N_A2_c_209_n 0.00112647f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A1_c_169_n N_A2_c_209_n 0.0221649f $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A1_c_166_n N_Y_c_285_n 0.0117564f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_149 A1 N_Y_c_285_n 0.0356656f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A1_c_169_n N_Y_c_285_n 0.00468889f $X=3.47 $Y=1.202 $X2=0 $Y2=0
cc_151 N_A1_c_170_n N_A_320_297#_c_331_n 0.019037f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_152 A1 N_A_320_297#_c_331_n 0.020833f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_169_n N_A_320_297#_c_331_n 7.48985e-19 $X=3.47 $Y=1.202 $X2=0
+ $Y2=0
cc_154 N_A1_c_171_n N_A_320_297#_c_332_n 0.0166967f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_155 A1 N_A_320_297#_c_332_n 0.0145519f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_169_n N_A_320_297#_c_332_n 7.48985e-19 $X=3.47 $Y=1.202 $X2=0
+ $Y2=0
cc_157 A1 N_A_320_297#_c_335_n 0.0223447f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_158 N_A1_c_169_n N_A_320_297#_c_335_n 0.00688955f $X=3.47 $Y=1.202 $X2=0
+ $Y2=0
cc_159 N_A1_c_170_n N_VPWR_c_380_n 0.00464144f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A1_c_171_n N_VPWR_c_381_n 0.00291222f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A1_c_170_n N_VPWR_c_385_n 0.00702461f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A1_c_171_n N_VPWR_c_385_n 0.00702461f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A1_c_170_n N_VPWR_c_379_n 0.0137545f $X=2.99 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A1_c_171_n N_VPWR_c_379_n 0.0125211f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A1_c_166_n N_VGND_c_446_n 0.00252024f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A1_c_167_n N_VGND_c_447_n 0.00126572f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A1_c_166_n N_VGND_c_448_n 0.00359964f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A1_c_167_n N_VGND_c_448_n 0.00359964f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A1_c_166_n N_VGND_c_451_n 0.00682766f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A1_c_167_n N_VGND_c_451_n 0.00559419f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A1_c_166_n N_A_525_47#_c_513_n 0.00954283f $X=2.965 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A1_c_167_n N_A_525_47#_c_513_n 0.0120706f $X=3.495 $Y=0.995 $X2=0 $Y2=0
cc_173 A1 N_A_525_47#_c_513_n 0.00431881f $X=3.395 $Y=1.105 $X2=0 $Y2=0
cc_174 N_A2_c_211_n N_A_320_297#_c_332_n 0.0170511f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_175 A2 N_A_320_297#_c_332_n 0.0116855f $X=4.685 $Y=1.105 $X2=0 $Y2=0
cc_176 N_A2_c_209_n N_A_320_297#_c_332_n 8.05532e-19 $X=4.43 $Y=1.202 $X2=0
+ $Y2=0
cc_177 N_A2_c_212_n N_A_320_297#_c_333_n 3.88929e-19 $X=4.43 $Y=1.41 $X2=0 $Y2=0
cc_178 A2 N_A_320_297#_c_333_n 0.0223447f $X=4.685 $Y=1.105 $X2=0 $Y2=0
cc_179 A2 N_A_320_297#_c_333_n 0.00522847f $X=4.72 $Y=1.445 $X2=0 $Y2=0
cc_180 N_A2_c_209_n N_A_320_297#_c_333_n 0.00688955f $X=4.43 $Y=1.202 $X2=0
+ $Y2=0
cc_181 A2 N_VPWR_M1008_d 0.00456566f $X=4.72 $Y=1.445 $X2=0 $Y2=0
cc_182 N_A2_c_211_n N_VPWR_c_381_n 0.00291222f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A2_c_212_n N_VPWR_c_382_n 0.00464144f $X=4.43 $Y=1.41 $X2=0 $Y2=0
cc_184 A2 N_VPWR_c_382_n 0.00428501f $X=4.685 $Y=1.105 $X2=0 $Y2=0
cc_185 A2 N_VPWR_c_382_n 0.00840623f $X=4.72 $Y=1.445 $X2=0 $Y2=0
cc_186 N_A2_c_211_n N_VPWR_c_388_n 0.00702461f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A2_c_212_n N_VPWR_c_388_n 0.00702461f $X=4.43 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A2_c_211_n N_VPWR_c_379_n 0.0125211f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A2_c_212_n N_VPWR_c_379_n 0.0134871f $X=4.43 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A2_c_205_n N_VGND_c_447_n 0.00781941f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_206_n N_VGND_c_447_n 0.00323317f $X=4.455 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_205_n N_VGND_c_448_n 0.00354245f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_206_n N_VGND_c_450_n 0.00425094f $X=4.455 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_205_n N_VGND_c_451_n 0.00418343f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_206_n N_VGND_c_451_n 0.00701427f $X=4.455 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_205_n N_A_525_47#_c_514_n 0.0133229f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_206_n N_A_525_47#_c_514_n 0.0141242f $X=4.455 $Y=0.995 $X2=0 $Y2=0
cc_198 A2 N_A_525_47#_c_514_n 0.0504092f $X=4.685 $Y=1.105 $X2=0 $Y2=0
cc_199 N_A2_c_209_n N_A_525_47#_c_514_n 0.0047002f $X=4.43 $Y=1.202 $X2=0 $Y2=0
cc_200 N_A2_c_210_n N_A_525_47#_c_514_n 0.0130672f $X=4.8 $Y=1.285 $X2=0 $Y2=0
cc_201 N_A_37_297#_c_255_n N_Y_M1004_d 0.00376318f $X=1.175 $Y=2.37 $X2=0 $Y2=0
cc_202 N_A_37_297#_c_255_n Y 0.01874f $X=1.175 $Y=2.37 $X2=0 $Y2=0
cc_203 N_A_37_297#_c_261_n N_A_320_297#_M1005_d 0.00383041f $X=2.135 $Y=2.355
+ $X2=-0.19 $Y2=1.305
cc_204 N_A_37_297#_M1013_s N_A_320_297#_c_331_n 0.00327427f $X=2.08 $Y=1.485
+ $X2=0 $Y2=0
cc_205 N_A_37_297#_c_261_n N_A_320_297#_c_331_n 0.00401632f $X=2.135 $Y=2.355
+ $X2=0 $Y2=0
cc_206 N_A_37_297#_c_251_n N_A_320_297#_c_331_n 0.0218566f $X=2.23 $Y=2 $X2=0
+ $Y2=0
cc_207 N_A_37_297#_c_261_n N_A_320_297#_c_334_n 0.018955f $X=2.135 $Y=2.355
+ $X2=0 $Y2=0
cc_208 N_A_37_297#_c_250_n N_VPWR_c_380_n 0.0140848f $X=2.275 $Y=2.255 $X2=0
+ $Y2=0
cc_209 N_A_37_297#_c_251_n N_VPWR_c_380_n 0.0273982f $X=2.23 $Y=2 $X2=0 $Y2=0
cc_210 N_A_37_297#_c_255_n N_VPWR_c_383_n 0.039305f $X=1.175 $Y=2.37 $X2=0 $Y2=0
cc_211 N_A_37_297#_c_249_n N_VPWR_c_383_n 0.0171513f $X=0.405 $Y=2.37 $X2=0
+ $Y2=0
cc_212 N_A_37_297#_c_261_n N_VPWR_c_383_n 0.0396474f $X=2.135 $Y=2.355 $X2=0
+ $Y2=0
cc_213 N_A_37_297#_c_250_n N_VPWR_c_383_n 0.0183943f $X=2.275 $Y=2.255 $X2=0
+ $Y2=0
cc_214 N_A_37_297#_c_276_p N_VPWR_c_383_n 0.0124114f $X=1.27 $Y=2.355 $X2=0
+ $Y2=0
cc_215 N_A_37_297#_M1004_s N_VPWR_c_379_n 0.00221966f $X=0.185 $Y=1.485 $X2=0
+ $Y2=0
cc_216 N_A_37_297#_M1011_s N_VPWR_c_379_n 0.00239679f $X=1.12 $Y=1.485 $X2=0
+ $Y2=0
cc_217 N_A_37_297#_M1013_s N_VPWR_c_379_n 0.00221966f $X=2.08 $Y=1.485 $X2=0
+ $Y2=0
cc_218 N_A_37_297#_c_255_n N_VPWR_c_379_n 0.0267141f $X=1.175 $Y=2.37 $X2=0
+ $Y2=0
cc_219 N_A_37_297#_c_249_n N_VPWR_c_379_n 0.00995095f $X=0.405 $Y=2.37 $X2=0
+ $Y2=0
cc_220 N_A_37_297#_c_261_n N_VPWR_c_379_n 0.0268145f $X=2.135 $Y=2.355 $X2=0
+ $Y2=0
cc_221 N_A_37_297#_c_250_n N_VPWR_c_379_n 0.0106949f $X=2.275 $Y=2.255 $X2=0
+ $Y2=0
cc_222 N_A_37_297#_c_276_p N_VPWR_c_379_n 0.00725819f $X=1.27 $Y=2.355 $X2=0
+ $Y2=0
cc_223 N_Y_c_285_n N_A_320_297#_c_331_n 0.0253539f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_224 N_Y_M1004_d N_VPWR_c_379_n 0.00241318f $X=0.64 $Y=1.485 $X2=0 $Y2=0
cc_225 N_Y_c_285_n N_VGND_M1014_s 0.00357056f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_226 N_Y_c_285_n N_VGND_M1006_s 0.00729184f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_227 Y N_VGND_c_443_n 0.0123602f $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_228 N_Y_c_295_n N_VGND_c_443_n 0.0289134f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_229 N_Y_c_285_n N_VGND_c_444_n 0.0189097f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_230 N_Y_c_295_n N_VGND_c_444_n 0.0171757f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_231 N_Y_c_285_n N_VGND_c_445_n 0.0086905f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_232 N_Y_c_285_n N_VGND_c_446_n 0.0233875f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_233 N_Y_c_285_n N_VGND_c_448_n 0.00335954f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_234 N_Y_c_285_n N_VGND_c_449_n 0.00216426f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_235 N_Y_c_295_n N_VGND_c_449_n 0.0194818f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_236 N_Y_M1012_d N_VGND_c_451_n 0.00301699f $X=0.65 $Y=0.235 $X2=0 $Y2=0
cc_237 N_Y_M1001_d N_VGND_c_451_n 0.00457742f $X=1.56 $Y=0.235 $X2=0 $Y2=0
cc_238 N_Y_M1002_s N_VGND_c_451_n 0.0030567f $X=3.04 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_285_n N_VGND_c_451_n 0.0296938f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_240 Y N_VGND_c_451_n 2.9649e-19 $X=0.585 $Y=0.765 $X2=0 $Y2=0
cc_241 N_Y_c_295_n N_VGND_c_451_n 0.0114508f $X=0.79 $Y=0.42 $X2=0 $Y2=0
cc_242 N_Y_c_285_n N_A_525_47#_M1002_d 0.00708857f $X=3.23 $Y=0.755 $X2=-0.19
+ $Y2=-0.24
cc_243 N_Y_M1002_s N_A_525_47#_c_513_n 0.00548807f $X=3.04 $Y=0.235 $X2=0 $Y2=0
cc_244 N_Y_c_285_n N_A_525_47#_c_513_n 0.0443062f $X=3.23 $Y=0.755 $X2=0 $Y2=0
cc_245 N_A_320_297#_c_331_n N_VPWR_M1003_s 0.00358195f $X=3.095 $Y=1.555
+ $X2=-0.19 $Y2=1.305
cc_246 N_A_320_297#_c_332_n N_VPWR_M1015_s 0.00203544f $X=4.055 $Y=1.555 $X2=0
+ $Y2=0
cc_247 N_A_320_297#_c_331_n N_VPWR_c_380_n 0.0163148f $X=3.095 $Y=1.555 $X2=0
+ $Y2=0
cc_248 N_A_320_297#_c_332_n N_VPWR_c_381_n 0.0146597f $X=4.055 $Y=1.555 $X2=0
+ $Y2=0
cc_249 N_A_320_297#_c_370_p N_VPWR_c_385_n 0.0159891f $X=3.23 $Y=2.3 $X2=0 $Y2=0
cc_250 N_A_320_297#_c_371_p N_VPWR_c_388_n 0.0159891f $X=4.19 $Y=2.3 $X2=0 $Y2=0
cc_251 N_A_320_297#_M1005_d N_VPWR_c_379_n 0.00241318f $X=1.6 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_320_297#_M1003_d N_VPWR_c_379_n 0.00343438f $X=3.08 $Y=1.485 $X2=0
+ $Y2=0
cc_253 N_A_320_297#_M1000_s N_VPWR_c_379_n 0.00343438f $X=4.04 $Y=1.485 $X2=0
+ $Y2=0
cc_254 N_A_320_297#_c_370_p N_VPWR_c_379_n 0.0103212f $X=3.23 $Y=2.3 $X2=0 $Y2=0
cc_255 N_A_320_297#_c_371_p N_VPWR_c_379_n 0.0103212f $X=4.19 $Y=2.3 $X2=0 $Y2=0
cc_256 N_A_320_297#_c_332_n N_A_525_47#_c_514_n 0.00190555f $X=4.055 $Y=1.555
+ $X2=0 $Y2=0
cc_257 N_A_320_297#_c_332_n N_A_525_47#_c_528_n 0.00556674f $X=4.055 $Y=1.555
+ $X2=0 $Y2=0
cc_258 N_VGND_c_451_n N_A_525_47#_M1002_d 0.00213789f $X=4.83 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_259 N_VGND_c_451_n N_A_525_47#_M1007_d 0.00245191f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_260 N_VGND_c_451_n N_A_525_47#_M1010_s 0.00233744f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_261 N_VGND_c_446_n N_A_525_47#_c_513_n 0.0171803f $X=2.23 $Y=0.38 $X2=0 $Y2=0
cc_262 N_VGND_c_448_n N_A_525_47#_c_513_n 0.0671949f $X=3.975 $Y=0 $X2=0 $Y2=0
cc_263 N_VGND_c_451_n N_A_525_47#_c_513_n 0.0437078f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_264 N_VGND_M1009_d N_A_525_47#_c_514_n 0.0054808f $X=4 $Y=0.235 $X2=0 $Y2=0
cc_265 N_VGND_c_447_n N_A_525_47#_c_514_n 0.0212258f $X=4.165 $Y=0 $X2=0 $Y2=0
cc_266 N_VGND_c_448_n N_A_525_47#_c_514_n 0.00261003f $X=3.975 $Y=0 $X2=0 $Y2=0
cc_267 N_VGND_c_450_n N_A_525_47#_c_514_n 0.00327039f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_268 N_VGND_c_451_n N_A_525_47#_c_514_n 0.0120601f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_269 N_VGND_c_450_n N_A_525_47#_c_515_n 0.0162389f $X=4.83 $Y=0 $X2=0 $Y2=0
cc_270 N_VGND_c_451_n N_A_525_47#_c_515_n 0.0094641f $X=4.83 $Y=0 $X2=0 $Y2=0
