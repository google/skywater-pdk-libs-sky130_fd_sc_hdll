* File: sky130_fd_sc_hdll__and3b_2.spice
* Created: Wed Sep  2 08:22:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and3b_2.pex.spice"
.subckt sky130_fd_sc_hdll__and3b_2  VNB VPB A_N B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1000 N_A_117_311#_M1000_d N_A_N_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1176 AS=0.1302 PD=1.4 PS=1.46 NRD=4.284 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 A_317_53# N_A_117_311#_M1001_g N_A_225_311#_M1001_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0672 AS=0.1218 PD=0.74 PS=1.42 NRD=30 NRS=7.14 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1009 A_411_53# N_B_M1009_g A_317_53# VNB NSHORT L=0.15 W=0.42 AD=0.0441
+ AS=0.0672 PD=0.63 PS=0.74 NRD=14.28 NRS=30 M=1 R=2.8 SA=75000.7 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_C_M1010_g A_411_53# VNB NSHORT L=0.15 W=0.42 AD=0.121643
+ AS=0.0441 PD=0.942056 PS=0.63 NRD=62.856 NRS=14.28 M=1 R=2.8 SA=75001
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1010_d N_A_225_311#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.188257 AS=0.104 PD=1.45794 PS=0.97 NRD=9.228 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_225_311#_M1006_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2535 AS=0.104 PD=2.08 PS=0.97 NRD=23.076 NRS=8.304 M=1 R=4.33333
+ SA=75001.7 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_117_311#_M1002_d N_A_N_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1134 PD=1.38 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_A_117_311#_M1007_g N_A_225_311#_M1007_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90002 A=0.0756 P=1.2 MULT=1
MM1003 N_A_225_311#_M1003_d N_B_M1003_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.078575 AS=0.0609 PD=0.835 PS=0.71 NRD=28.1316 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_C_M1004_g N_A_225_311#_M1003_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.078575 PD=0.801549 PS=0.835 NRD=75.1752 NRS=0 M=1 R=2.33333
+ SA=90001 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1004_d N_A_225_311#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.145 PD=1.90845 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.8 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_225_311#_M1011_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.4 AS=0.145 PD=2.8 PS=1.29 NRD=26.5753 NRS=0.9653 M=1 R=5.55556 SA=90001.2
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_13 X X PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and3b_2.pxi.spice"
*
.ends
*
*
