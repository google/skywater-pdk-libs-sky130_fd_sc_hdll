* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4bb_4 A_N B_N C D VGND VNB VPB VPWR Y
X0 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_853_47# C a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND D a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 Y a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_395_47# a_206_47# a_853_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 Y a_27_47# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND D a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_853_47# a_206_47# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1251_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y a_206_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VPWR a_206_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 Y a_27_47# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 a_1251_47# C a_853_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 a_1251_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND B_N a_206_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_1251_47# C a_853_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_395_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 VPWR B_N a_206_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 VPWR a_206_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_395_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 a_853_47# a_206_47# a_395_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 a_395_47# a_206_47# a_853_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X34 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_853_47# C a_1251_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
