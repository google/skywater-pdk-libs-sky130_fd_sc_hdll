* NGSPICE file created from sky130_fd_sc_hdll__o21a_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
M1000 a_79_21# B1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=1.365e+12p ps=8.73e+06u
M1001 X a_79_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.95e+11p pd=2.59e+06u as=0p ps=0u
M1002 a_414_47# B1 a_79_21# VNB nshort w=650000u l=150000u
+  ad=3.8675e+11p pd=3.79e+06u as=2.0475e+11p ps=1.93e+06u
M1003 a_414_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.1825e+11p ps=6.11e+06u
M1004 VGND A2 a_414_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_79_21# VGND VNB nshort w=650000u l=150000u
+  ad=2.1125e+11p pd=1.95e+06u as=0p ps=0u
M1006 VPWR a_79_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_508_297# A2 a_79_21# VPB phighvt w=1e+06u l=180000u
+  ad=5e+11p pd=3e+06u as=0p ps=0u
M1008 VPWR A1 a_508_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VGND a_79_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

