* File: sky130_fd_sc_hdll__mux2_16.pex.spice
* Created: Wed Sep  2 08:34:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39
r88 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.905 $Y2=1.202
r89 37 39 16.8441 $w=3.72e-07 $l=1.3e-07 $layer=POLY_cond $X=1.75 $Y=1.202
+ $X2=1.88 $Y2=1.202
r90 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.75
+ $Y=1.16 $X2=1.75 $Y2=1.16
r91 35 37 37.5753 $w=3.72e-07 $l=2.9e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.75 $Y2=1.202
r92 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r93 33 34 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.435 $Y2=1.202
r94 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r95 30 32 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=0.73 $Y=1.202
+ $X2=0.94 $Y2=1.202
r96 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.73
+ $Y=1.16 $X2=0.73 $Y2=1.16
r97 28 30 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.73 $Y2=1.202
r98 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r99 25 38 27.6586 $w=2.48e-07 $l=6e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=1.75
+ $Y2=1.2
r100 25 31 19.361 $w=2.48e-07 $l=4.2e-07 $layer=LI1_cond $X=1.15 $Y=1.2 $X2=0.73
+ $Y2=1.2
r101 22 40 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r102 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r103 19 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=1.202
r104 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.88 $Y=0.995
+ $X2=1.88 $Y2=0.56
r105 16 35 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r106 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r107 13 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r108 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r109 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r110 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r111 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r112 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=0.56
r113 4 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r114 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r115 1 27 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r116 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%S 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 43 55
r124 55 56 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.245 $Y2=1.202
r125 54 55 54.7135 $w=3.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=5.22 $Y2=1.202
r126 53 54 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r127 52 53 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.775 $Y2=1.202
r128 51 52 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r129 49 51 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=4.11 $Y=1.202
+ $X2=4.28 $Y2=1.202
r130 47 49 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.86 $Y=1.202
+ $X2=4.11 $Y2=1.202
r131 46 47 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r132 45 46 61.227 $w=3.7e-07 $l=4.7e-07 $layer=POLY_cond $X=3.365 $Y=1.202
+ $X2=3.835 $Y2=1.202
r133 44 45 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.365 $Y2=1.202
r134 43 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.11
+ $Y=1.16 $X2=4.11 $Y2=1.16
r135 42 44 32.5676 $w=3.7e-07 $l=2.5e-07 $layer=POLY_cond $X=3.09 $Y=1.202
+ $X2=3.34 $Y2=1.202
r136 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.09
+ $Y=1.16 $X2=3.09 $Y2=1.16
r137 40 42 22.1459 $w=3.7e-07 $l=1.7e-07 $layer=POLY_cond $X=2.92 $Y=1.202
+ $X2=3.09 $Y2=1.202
r138 39 40 3.25676 $w=3.7e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.202
+ $X2=2.92 $Y2=1.202
r139 37 43 0.271111 $w=1.348e-06 $l=3e-08 $layer=LI1_cond $X=3.6 $Y=1.19 $X2=3.6
+ $Y2=1.16
r140 34 56 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.202
r141 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r142 31 55 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r143 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r144 28 54 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r145 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=0.56
r146 25 53 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r147 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r148 22 52 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r149 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r150 19 51 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r151 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r152 16 47 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r153 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r154 13 46 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r155 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r156 10 45 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.202
r157 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r158 7 44 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r159 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r160 4 40 23.9667 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.92 $Y2=1.202
r161 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.92 $Y2=0.56
r162 1 39 19.6139 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.202
r163 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_973_297# 1 2 7 9 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 33 37 46 49 58
r122 58 59 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.1 $Y=1.202
+ $X2=7.125 $Y2=1.202
r123 55 56 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.655 $Y=1.202
+ $X2=6.68 $Y2=1.202
r124 54 55 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.655 $Y2=1.202
r125 53 54 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r126 50 51 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.715 $Y=1.202
+ $X2=5.74 $Y2=1.202
r127 47 58 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=6.93 $Y=1.202
+ $X2=7.1 $Y2=1.202
r128 47 56 32.3925 $w=3.72e-07 $l=2.5e-07 $layer=POLY_cond $X=6.93 $Y=1.202
+ $X2=6.68 $Y2=1.202
r129 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.93
+ $Y=1.16 $X2=6.93 $Y2=1.16
r130 44 53 32.3925 $w=3.72e-07 $l=2.5e-07 $layer=POLY_cond $X=5.91 $Y=1.202
+ $X2=6.16 $Y2=1.202
r131 44 51 22.0269 $w=3.72e-07 $l=1.7e-07 $layer=POLY_cond $X=5.91 $Y=1.202
+ $X2=5.74 $Y2=1.202
r132 43 46 47.0197 $w=2.48e-07 $l=1.02e-06 $layer=LI1_cond $X=5.91 $Y=1.2
+ $X2=6.93 $Y2=1.2
r133 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.91
+ $Y=1.16 $X2=5.91 $Y2=1.16
r134 41 49 2.3589 $w=2.5e-07 $l=1.65e-07 $layer=LI1_cond $X=5.175 $Y=1.2
+ $X2=5.01 $Y2=1.2
r135 41 43 33.8818 $w=2.48e-07 $l=7.35e-07 $layer=LI1_cond $X=5.175 $Y=1.2
+ $X2=5.91 $Y2=1.2
r136 37 39 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=5.01 $Y=1.66
+ $X2=5.01 $Y2=2.34
r137 35 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.01 $Y2=1.2
r138 35 37 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.01 $Y=1.325
+ $X2=5.01 $Y2=1.66
r139 31 49 4.07664 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=5.01 $Y=1.075
+ $X2=5.01 $Y2=1.2
r140 31 33 22.8742 $w=3.28e-07 $l=6.55e-07 $layer=LI1_cond $X=5.01 $Y=1.075
+ $X2=5.01 $Y2=0.42
r141 28 59 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r142 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r143 25 58 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=1.202
r144 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.1 $Y=0.995
+ $X2=7.1 $Y2=0.56
r145 22 56 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=1.202
r146 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.68 $Y=0.995
+ $X2=6.68 $Y2=0.56
r147 19 55 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r148 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r149 16 54 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r150 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r151 13 53 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r152 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r153 10 51 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=1.202
r154 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.74 $Y=0.995
+ $X2=5.74 $Y2=0.56
r155 7 50 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r156 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r157 2 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2.34
r158 2 37 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.66
r159 1 33 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A0 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 38 39
r92 39 40 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.5 $Y=1.202
+ $X2=9.525 $Y2=1.202
r93 37 39 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=9.29 $Y=1.202
+ $X2=9.5 $Y2=1.202
r94 37 38 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.29
+ $Y=1.16 $X2=9.29 $Y2=1.16
r95 35 37 27.2097 $w=3.72e-07 $l=2.1e-07 $layer=POLY_cond $X=9.08 $Y=1.202
+ $X2=9.29 $Y2=1.202
r96 34 35 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=9.055 $Y=1.202
+ $X2=9.08 $Y2=1.202
r97 33 34 60.8979 $w=3.72e-07 $l=4.7e-07 $layer=POLY_cond $X=8.585 $Y=1.202
+ $X2=9.055 $Y2=1.202
r98 32 33 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.56 $Y=1.202
+ $X2=8.585 $Y2=1.202
r99 30 32 37.5753 $w=3.72e-07 $l=2.9e-07 $layer=POLY_cond $X=8.27 $Y=1.202
+ $X2=8.56 $Y2=1.202
r100 30 31 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.27
+ $Y=1.16 $X2=8.27 $Y2=1.16
r101 28 30 16.8441 $w=3.72e-07 $l=1.3e-07 $layer=POLY_cond $X=8.14 $Y=1.202
+ $X2=8.27 $Y2=1.202
r102 27 28 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=8.115 $Y=1.202
+ $X2=8.14 $Y2=1.202
r103 25 38 14.7513 $w=2.48e-07 $l=3.2e-07 $layer=LI1_cond $X=8.97 $Y=1.2
+ $X2=9.29 $Y2=1.2
r104 25 31 32.2684 $w=2.48e-07 $l=7e-07 $layer=LI1_cond $X=8.97 $Y=1.2 $X2=8.27
+ $Y2=1.2
r105 22 40 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.525 $Y=1.41
+ $X2=9.525 $Y2=1.202
r106 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.525 $Y=1.41
+ $X2=9.525 $Y2=1.985
r107 19 39 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=1.202
r108 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.5 $Y=0.995
+ $X2=9.5 $Y2=0.56
r109 16 35 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=1.202
r110 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.08 $Y=0.995
+ $X2=9.08 $Y2=0.56
r111 13 34 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.202
r112 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.055 $Y=1.41
+ $X2=9.055 $Y2=1.985
r113 10 33 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.202
r114 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.585 $Y=1.41
+ $X2=8.585 $Y2=1.985
r115 7 32 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=1.202
r116 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.56 $Y=0.995
+ $X2=8.56 $Y2=0.56
r117 4 28 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=1.202
r118 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.14 $Y=0.995
+ $X2=8.14 $Y2=0.56
r119 1 27 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.202
r120 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.115 $Y=1.41
+ $X2=8.115 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 12 37 39
+ 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61 63 64 66 67 69 70 72 73 75 76 78
+ 79 81 82 84 85 87 88 90 91 93 94 96 97 99 100 102 103 105 106 108 109 111 112
+ 114 115 117 118 120 121 123 124 126 127 129 130 132 135 139 143 145 147 149
+ 151 155 159 161 163 166 168 174 177 180 185 186 187 189 190 197 202 203 204
+ 205 209 212 213 216 219 220 254
c560 219 0 1.96891e-19 $X=9.76 $Y=0.51
c561 213 0 1.96891e-19 $X=0.405 $Y=0.51
r562 254 255 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=17.54 $Y=1.202
+ $X2=17.565 $Y2=1.202
r563 253 254 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=17.12 $Y=1.202
+ $X2=17.54 $Y2=1.202
r564 252 253 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=17.095 $Y=1.202
+ $X2=17.12 $Y2=1.202
r565 249 250 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=16.6 $Y=1.202
+ $X2=16.625 $Y2=1.202
r566 248 249 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=16.18 $Y=1.202
+ $X2=16.6 $Y2=1.202
r567 247 248 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=16.155 $Y=1.202
+ $X2=16.18 $Y2=1.202
r568 246 247 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=15.685 $Y=1.202
+ $X2=16.155 $Y2=1.202
r569 245 246 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.66 $Y=1.202
+ $X2=15.685 $Y2=1.202
r570 244 245 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=15.24 $Y=1.202
+ $X2=15.66 $Y2=1.202
r571 243 244 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=15.215 $Y=1.202
+ $X2=15.24 $Y2=1.202
r572 242 243 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=14.745 $Y=1.202
+ $X2=15.215 $Y2=1.202
r573 241 242 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.72 $Y=1.202
+ $X2=14.745 $Y2=1.202
r574 240 241 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=14.3 $Y=1.202
+ $X2=14.72 $Y2=1.202
r575 239 240 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=14.275 $Y=1.202
+ $X2=14.3 $Y2=1.202
r576 238 239 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=13.805 $Y=1.202
+ $X2=14.275 $Y2=1.202
r577 237 238 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.78 $Y=1.202
+ $X2=13.805 $Y2=1.202
r578 236 237 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=13.36 $Y=1.202
+ $X2=13.78 $Y2=1.202
r579 235 236 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=13.335 $Y=1.202
+ $X2=13.36 $Y2=1.202
r580 234 235 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=12.865 $Y=1.202
+ $X2=13.335 $Y2=1.202
r581 233 234 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.84 $Y=1.202
+ $X2=12.865 $Y2=1.202
r582 232 233 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=12.42 $Y=1.202
+ $X2=12.84 $Y2=1.202
r583 231 232 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=12.395 $Y=1.202
+ $X2=12.42 $Y2=1.202
r584 230 231 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=11.925 $Y=1.202
+ $X2=12.395 $Y2=1.202
r585 229 230 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.9 $Y=1.202
+ $X2=11.925 $Y2=1.202
r586 228 229 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=11.48 $Y=1.202
+ $X2=11.9 $Y2=1.202
r587 227 228 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.455 $Y=1.202
+ $X2=11.48 $Y2=1.202
r588 226 227 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=10.985 $Y=1.202
+ $X2=11.455 $Y2=1.202
r589 225 226 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.96 $Y=1.202
+ $X2=10.985 $Y2=1.202
r590 222 223 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.515 $Y=1.202
+ $X2=10.54 $Y2=1.202
r591 219 220 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.76 $Y=0.51
+ $X2=9.76 $Y2=0.51
r592 216 258 44.177 $w=2.98e-07 $l=1.15e-06 $layer=LI1_cond $X=0.245 $Y=0.51
+ $X2=0.245 $Y2=1.66
r593 215 216 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.26 $Y=0.51
+ $X2=0.26 $Y2=0.51
r594 213 215 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.405 $Y=0.51
+ $X2=0.26 $Y2=0.51
r595 212 219 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.615 $Y=0.51
+ $X2=9.76 $Y2=0.51
r596 212 213 11.3985 $w=1.4e-07 $l=9.21e-06 $layer=MET1_cond $X=9.615 $Y=0.51
+ $X2=0.405 $Y2=0.51
r597 208 220 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=9.775 $Y=1.075
+ $X2=9.775 $Y2=0.51
r598 208 209 4.4274 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.775 $Y=1.075
+ $X2=9.775 $Y2=1.2
r599 205 220 3.26526 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.425
+ $X2=9.775 $Y2=0.51
r600 205 207 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.425
+ $X2=9.775 $Y2=0.34
r601 201 203 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.82 $Y=0.4
+ $X2=8.955 $Y2=0.4
r602 201 202 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=8.82 $Y=0.4
+ $X2=8.685 $Y2=0.4
r603 197 202 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.015 $Y=0.34
+ $X2=8.685 $Y2=0.34
r604 195 197 7.32568 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=7.88 $Y=0.402
+ $X2=8.015 $Y2=0.402
r605 189 190 7.32568 $w=2.93e-07 $l=1.35e-07 $layer=LI1_cond $X=2.14 $Y=0.402
+ $X2=2.005 $Y2=0.402
r606 186 190 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=2.005 $Y2=0.34
r607 184 186 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.4
+ $X2=1.335 $Y2=0.4
r608 184 185 7.32169 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.4
+ $X2=1.065 $Y2=0.4
r609 180 258 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.295
+ $X2=0.245 $Y2=1.66
r610 180 182 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=2.295
+ $X2=0.245 $Y2=2.38
r611 177 216 3.26526 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.51
r612 177 179 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=0.425
+ $X2=0.245 $Y2=0.34
r613 175 252 51.8774 $w=3.67e-07 $l=3.95e-07 $layer=POLY_cond $X=16.7 $Y=1.202
+ $X2=17.095 $Y2=1.202
r614 175 250 9.85014 $w=3.67e-07 $l=7.5e-08 $layer=POLY_cond $X=16.7 $Y=1.202
+ $X2=16.625 $Y2=1.202
r615 174 175 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9 $X=16.7
+ $Y=1.16 $X2=16.7 $Y2=1.16
r616 172 225 49.9074 $w=3.67e-07 $l=3.8e-07 $layer=POLY_cond $X=10.58 $Y=1.202
+ $X2=10.96 $Y2=1.202
r617 172 223 5.25341 $w=3.67e-07 $l=4e-08 $layer=POLY_cond $X=10.58 $Y=1.202
+ $X2=10.54 $Y2=1.202
r618 171 174 282.118 $w=2.48e-07 $l=6.12e-06 $layer=LI1_cond $X=10.58 $Y=1.2
+ $X2=16.7 $Y2=1.2
r619 171 172 15.2926 $w=1.7e-07 $l=1.615e-06 $layer=licon1_POLY $count=9
+ $X=10.58 $Y=1.16 $X2=10.58 $Y2=1.16
r620 169 209 2.0066 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=9.925 $Y=1.2
+ $X2=9.775 $Y2=1.2
r621 169 171 30.194 $w=2.48e-07 $l=6.55e-07 $layer=LI1_cond $X=9.925 $Y=1.2
+ $X2=10.58 $Y2=1.2
r622 166 211 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=2.295
+ $X2=9.775 $Y2=2.38
r623 166 168 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=9.775 $Y=2.295
+ $X2=9.775 $Y2=1.66
r624 165 209 4.4274 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=9.775 $Y=1.325
+ $X2=9.775 $Y2=1.2
r625 165 168 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=9.775 $Y=1.325
+ $X2=9.775 $Y2=1.66
r626 164 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.955 $Y=2.38
+ $X2=8.82 $Y2=2.38
r627 163 211 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.625 $Y=2.38
+ $X2=9.775 $Y2=2.38
r628 163 164 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.625 $Y=2.38
+ $X2=8.955 $Y2=2.38
r629 161 207 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=9.625 $Y=0.34
+ $X2=9.775 $Y2=0.34
r630 161 203 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.625 $Y=0.34
+ $X2=8.955 $Y2=0.34
r631 157 204 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.82 $Y=2.295
+ $X2=8.82 $Y2=2.38
r632 157 159 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.82 $Y=2.295
+ $X2=8.82 $Y2=2
r633 156 199 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=8.015 $Y=2.38
+ $X2=7.865 $Y2=2.38
r634 155 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=8.82 $Y2=2.38
r635 155 156 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.685 $Y=2.38
+ $X2=8.015 $Y2=2.38
r636 149 199 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.295
+ $X2=7.865 $Y2=2.38
r637 149 151 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=7.865 $Y=2.295
+ $X2=7.865 $Y2=1.66
r638 145 193 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.155 $Y2=2.38
r639 145 147 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=2.155 $Y=2.295
+ $X2=2.155 $Y2=1.66
r640 144 187 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.38
+ $X2=1.2 $Y2=2.38
r641 143 193 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.005 $Y=2.38
+ $X2=2.155 $Y2=2.38
r642 143 144 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.38
+ $X2=1.335 $Y2=2.38
r643 137 187 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=2.38
r644 137 139 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=2
r645 136 182 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=2.38
+ $X2=0.245 $Y2=2.38
r646 135 187 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.38
+ $X2=1.2 $Y2=2.38
r647 135 136 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.065 $Y=2.38
+ $X2=0.395 $Y2=2.38
r648 134 179 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=0.34
+ $X2=0.245 $Y2=0.34
r649 134 185 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.395 $Y=0.34
+ $X2=1.065 $Y2=0.34
r650 130 255 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=17.565 $Y=1.41
+ $X2=17.565 $Y2=1.202
r651 130 132 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=17.565 $Y=1.41
+ $X2=17.565 $Y2=1.985
r652 127 254 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=17.54 $Y=0.995
+ $X2=17.54 $Y2=1.202
r653 127 129 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=17.54 $Y=0.995
+ $X2=17.54 $Y2=0.56
r654 124 253 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=17.12 $Y=0.995
+ $X2=17.12 $Y2=1.202
r655 124 126 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=17.12 $Y=0.995
+ $X2=17.12 $Y2=0.56
r656 121 252 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=17.095 $Y=1.41
+ $X2=17.095 $Y2=1.202
r657 121 123 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=17.095 $Y=1.41
+ $X2=17.095 $Y2=1.985
r658 118 250 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=16.625 $Y=1.41
+ $X2=16.625 $Y2=1.202
r659 118 120 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.625 $Y=1.41
+ $X2=16.625 $Y2=1.985
r660 115 249 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=16.6 $Y=0.995
+ $X2=16.6 $Y2=1.202
r661 115 117 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.6 $Y=0.995
+ $X2=16.6 $Y2=0.56
r662 112 248 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=16.18 $Y=0.995
+ $X2=16.18 $Y2=1.202
r663 112 114 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=16.18 $Y=0.995
+ $X2=16.18 $Y2=0.56
r664 109 247 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=16.155 $Y=1.41
+ $X2=16.155 $Y2=1.202
r665 109 111 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.155 $Y=1.41
+ $X2=16.155 $Y2=1.985
r666 106 246 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.685 $Y=1.41
+ $X2=15.685 $Y2=1.202
r667 106 108 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.685 $Y=1.41
+ $X2=15.685 $Y2=1.985
r668 103 245 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.66 $Y=0.995
+ $X2=15.66 $Y2=1.202
r669 103 105 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.66 $Y=0.995
+ $X2=15.66 $Y2=0.56
r670 100 244 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=15.24 $Y=0.995
+ $X2=15.24 $Y2=1.202
r671 100 102 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=15.24 $Y=0.995
+ $X2=15.24 $Y2=0.56
r672 97 243 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=15.215 $Y=1.41
+ $X2=15.215 $Y2=1.202
r673 97 99 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.215 $Y=1.41
+ $X2=15.215 $Y2=1.985
r674 94 242 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.745 $Y=1.41
+ $X2=14.745 $Y2=1.202
r675 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.745 $Y=1.41
+ $X2=14.745 $Y2=1.985
r676 91 241 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.72 $Y=0.995
+ $X2=14.72 $Y2=1.202
r677 91 93 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.72 $Y=0.995
+ $X2=14.72 $Y2=0.56
r678 88 240 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.3 $Y=0.995
+ $X2=14.3 $Y2=1.202
r679 88 90 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.3 $Y=0.995
+ $X2=14.3 $Y2=0.56
r680 85 239 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.275 $Y=1.41
+ $X2=14.275 $Y2=1.202
r681 85 87 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.275 $Y=1.41
+ $X2=14.275 $Y2=1.985
r682 82 238 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.805 $Y=1.41
+ $X2=13.805 $Y2=1.202
r683 82 84 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.805 $Y=1.41
+ $X2=13.805 $Y2=1.985
r684 79 237 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.78 $Y=0.995
+ $X2=13.78 $Y2=1.202
r685 79 81 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.78 $Y=0.995
+ $X2=13.78 $Y2=0.56
r686 76 236 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.36 $Y=0.995
+ $X2=13.36 $Y2=1.202
r687 76 78 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.36 $Y=0.995
+ $X2=13.36 $Y2=0.56
r688 73 235 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.335 $Y=1.41
+ $X2=13.335 $Y2=1.202
r689 73 75 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.335 $Y=1.41
+ $X2=13.335 $Y2=1.985
r690 70 234 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.865 $Y=1.41
+ $X2=12.865 $Y2=1.202
r691 70 72 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.865 $Y=1.41
+ $X2=12.865 $Y2=1.985
r692 67 233 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=1.202
r693 67 69 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.84 $Y=0.995
+ $X2=12.84 $Y2=0.56
r694 64 232 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=12.42 $Y=0.995
+ $X2=12.42 $Y2=1.202
r695 64 66 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=12.42 $Y=0.995
+ $X2=12.42 $Y2=0.56
r696 61 231 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=12.395 $Y=1.41
+ $X2=12.395 $Y2=1.202
r697 61 63 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.395 $Y=1.41
+ $X2=12.395 $Y2=1.985
r698 58 230 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.925 $Y=1.41
+ $X2=11.925 $Y2=1.202
r699 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.925 $Y=1.41
+ $X2=11.925 $Y2=1.985
r700 55 229 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.9 $Y=0.995
+ $X2=11.9 $Y2=1.202
r701 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.9 $Y=0.995
+ $X2=11.9 $Y2=0.56
r702 52 228 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.48 $Y=0.995
+ $X2=11.48 $Y2=1.202
r703 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.48 $Y=0.995
+ $X2=11.48 $Y2=0.56
r704 49 227 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.202
r705 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.985
r706 46 226 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.202
r707 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.985
r708 43 225 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.96 $Y=0.995
+ $X2=10.96 $Y2=1.202
r709 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.96 $Y=0.995
+ $X2=10.96 $Y2=0.56
r710 40 223 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.54 $Y=0.995
+ $X2=10.54 $Y2=1.202
r711 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.54 $Y=0.995
+ $X2=10.54 $Y2=0.56
r712 37 222 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.202
r713 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.985
r714 12 211 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.485 $X2=9.76 $Y2=2.34
r715 12 168 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.615
+ $Y=1.485 $X2=9.76 $Y2=1.66
r716 11 159 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.675
+ $Y=1.485 $X2=8.82 $Y2=2
r717 10 199 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.485 $X2=7.88 $Y2=2.34
r718 10 151 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=7.755
+ $Y=1.485 $X2=7.88 $Y2=1.66
r719 9 193 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.34
r720 9 147 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.66
r721 8 139 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r722 7 258 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r723 7 182 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r724 6 207 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.575
+ $Y=0.235 $X2=9.76 $Y2=0.4
r725 5 201 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.635
+ $Y=0.235 $X2=8.82 $Y2=0.38
r726 4 195 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=7.755
+ $Y=0.235 $X2=7.88 $Y2=0.385
r727 3 189 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.385
r728 2 184 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.38
r729 1 179 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_117_297# 1 2 3 4 13 15 17 20 23 26 29 30
+ 31 32 33 34 37 41 44 46 47
r131 47 59 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=6.89 $Y=1.87
+ $X2=6.89 $Y2=2.34
r132 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.89 $Y=1.87
+ $X2=6.89 $Y2=1.87
r133 44 55 16.4136 $w=3.28e-07 $l=4.7e-07 $layer=LI1_cond $X=5.95 $Y=1.87
+ $X2=5.95 $Y2=2.34
r134 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.95 $Y=1.87
+ $X2=5.95 $Y2=1.87
r135 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.67 $Y=1.87
+ $X2=1.67 $Y2=1.87
r136 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.73 $Y=1.87
+ $X2=0.73 $Y2=1.87
r137 34 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.095 $Y=1.87
+ $X2=5.95 $Y2=1.87
r138 33 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.745 $Y=1.87
+ $X2=6.89 $Y2=1.87
r139 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=6.745 $Y=1.87
+ $X2=6.095 $Y2=1.87
r140 32 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.815 $Y=1.87
+ $X2=1.67 $Y2=1.87
r141 31 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.805 $Y=1.87
+ $X2=5.95 $Y2=1.87
r142 31 32 4.93811 $w=1.4e-07 $l=3.99e-06 $layer=MET1_cond $X=5.805 $Y=1.87
+ $X2=1.815 $Y2=1.87
r143 30 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.875 $Y=1.87
+ $X2=0.73 $Y2=1.87
r144 29 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.525 $Y=1.87
+ $X2=1.67 $Y2=1.87
r145 29 30 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=1.525 $Y=1.87
+ $X2=0.875 $Y2=1.87
r146 26 47 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=6.89 $Y=1.665
+ $X2=6.89 $Y2=1.87
r147 26 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.665
+ $X2=6.89 $Y2=1.58
r148 23 44 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=5.95 $Y=1.665
+ $X2=5.95 $Y2=1.87
r149 23 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.95 $Y=1.665
+ $X2=5.95 $Y2=1.58
r150 20 41 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.87
r151 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r152 17 37 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.87
r153 17 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r154 16 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.115 $Y=1.58
+ $X2=5.95 $Y2=1.58
r155 15 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=1.58
+ $X2=6.89 $Y2=1.58
r156 15 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=6.725 $Y=1.58
+ $X2=6.115 $Y2=1.58
r157 14 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r158 13 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r159 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r160 4 59 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=2.34
r161 4 28 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.66
r162 3 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=2.34
r163 3 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.66
r164 2 22 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r165 1 19 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 48 54 58 64 70 74 80 86 90 94 98 102 106 108 112 114 118 123 124 126 127 129
+ 130 132 133 135 136 138 139 140 142 169 173 178 183 188 193 200 201 204 207
+ 210 213 216 219 222 225 228 232
c301 126 0 1.97192e-19 $X=4.405 $Y=2.72
c302 123 0 1.97192e-19 $X=3.465 $Y=2.72
c303 5 0 1.91318e-19 $X=6.275 $Y=1.485
c304 2 0 1.91318e-19 $X=3.455 $Y=1.485
r305 228 229 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.71 $Y=2.72
+ $X2=17.71 $Y2=2.72
r306 226 229 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.79 $Y=2.72
+ $X2=17.71 $Y2=2.72
r307 225 226 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.79 $Y=2.72
+ $X2=16.79 $Y2=2.72
r308 223 226 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.87 $Y=2.72
+ $X2=16.79 $Y2=2.72
r309 222 223 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=2.72
+ $X2=15.87 $Y2=2.72
r310 219 220 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r311 216 217 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r312 213 214 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r313 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r314 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r315 204 205 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r316 201 229 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=2.72
+ $X2=17.71 $Y2=2.72
r317 200 201 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=2.72
+ $X2=18.17 $Y2=2.72
r318 198 228 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.935 $Y=2.72
+ $X2=17.8 $Y2=2.72
r319 198 200 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=17.935 $Y=2.72
+ $X2=18.17 $Y2=2.72
r320 197 223 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=15.87 $Y2=2.72
r321 197 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=2.72
+ $X2=14.95 $Y2=2.72
r322 196 197 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=2.72
+ $X2=15.41 $Y2=2.72
r323 194 219 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.115 $Y=2.72
+ $X2=14.98 $Y2=2.72
r324 194 196 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.115 $Y=2.72
+ $X2=15.41 $Y2=2.72
r325 193 222 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.785 $Y=2.72
+ $X2=15.92 $Y2=2.72
r326 193 196 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.785 $Y=2.72
+ $X2=15.41 $Y2=2.72
r327 192 220 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r328 192 217 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.03 $Y2=2.72
r329 191 192 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r330 189 216 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.175 $Y=2.72
+ $X2=14.04 $Y2=2.72
r331 189 191 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.175 $Y=2.72
+ $X2=14.49 $Y2=2.72
r332 188 219 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.845 $Y=2.72
+ $X2=14.98 $Y2=2.72
r333 188 191 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.845 $Y=2.72
+ $X2=14.49 $Y2=2.72
r334 187 217 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r335 187 214 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=13.11 $Y2=2.72
r336 186 187 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r337 184 213 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.235 $Y=2.72
+ $X2=13.1 $Y2=2.72
r338 184 186 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.235 $Y=2.72
+ $X2=13.57 $Y2=2.72
r339 183 216 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.905 $Y=2.72
+ $X2=14.04 $Y2=2.72
r340 183 186 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.905 $Y=2.72
+ $X2=13.57 $Y2=2.72
r341 182 214 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r342 182 211 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r343 181 182 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r344 179 210 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.295 $Y=2.72
+ $X2=12.16 $Y2=2.72
r345 179 181 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.295 $Y=2.72
+ $X2=12.65 $Y2=2.72
r346 178 213 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.965 $Y=2.72
+ $X2=13.1 $Y2=2.72
r347 178 181 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.965 $Y=2.72
+ $X2=12.65 $Y2=2.72
r348 177 211 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r349 177 208 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r350 176 177 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r351 174 207 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.355 $Y=2.72
+ $X2=11.22 $Y2=2.72
r352 174 176 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.355 $Y=2.72
+ $X2=11.73 $Y2=2.72
r353 173 210 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=12.16 $Y2=2.72
r354 173 176 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=2.72
+ $X2=11.73 $Y2=2.72
r355 172 208 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r356 171 172 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r357 169 207 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.085 $Y=2.72
+ $X2=11.22 $Y2=2.72
r358 169 171 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.085 $Y=2.72
+ $X2=10.81 $Y2=2.72
r359 168 172 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r360 167 168 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r361 165 168 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r362 164 167 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.89 $Y2=2.72
r363 164 165 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r364 162 165 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r365 161 162 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r366 159 162 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r367 158 159 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r368 156 159 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r369 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r370 153 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r371 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r372 150 153 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r373 150 205 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r374 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r375 147 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=2.66 $Y2=2.72
r376 147 149 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.795 $Y=2.72
+ $X2=3.45 $Y2=2.72
r377 144 232 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r378 142 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.66 $Y2=2.72
r379 142 144 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r380 140 205 0.653023 $w=4.8e-07 $l=2.295e-06 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=2.53 $Y2=2.72
r381 140 232 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r382 138 167 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.145 $Y=2.72
+ $X2=9.89 $Y2=2.72
r383 138 139 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.145 $Y=2.72
+ $X2=10.28 $Y2=2.72
r384 137 171 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.81 $Y2=2.72
r385 137 139 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.415 $Y=2.72
+ $X2=10.28 $Y2=2.72
r386 135 161 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.13 $Y2=2.72
r387 135 136 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.225 $Y=2.72
+ $X2=7.36 $Y2=2.72
r388 134 164 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=7.59 $Y2=2.72
r389 134 136 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.495 $Y=2.72
+ $X2=7.36 $Y2=2.72
r390 132 158 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.21 $Y2=2.72
r391 132 133 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.285 $Y=2.72
+ $X2=6.42 $Y2=2.72
r392 131 161 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=7.13 $Y2=2.72
r393 131 133 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.42 $Y2=2.72
r394 129 155 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r395 129 130 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.48 $Y2=2.72
r396 128 158 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=6.21 $Y2=2.72
r397 128 130 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.48 $Y2=2.72
r398 126 152 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.37 $Y2=2.72
r399 126 127 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.54 $Y2=2.72
r400 125 155 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=5.29 $Y2=2.72
r401 125 127 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=4.54 $Y2=2.72
r402 123 149 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.45 $Y2=2.72
r403 123 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=2.72
+ $X2=3.6 $Y2=2.72
r404 122 152 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=4.37 $Y2=2.72
r405 122 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=2.72
+ $X2=3.6 $Y2=2.72
r406 118 121 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=17.8 $Y=1.66
+ $X2=17.8 $Y2=2.34
r407 116 228 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.8 $Y=2.635
+ $X2=17.8 $Y2=2.72
r408 116 121 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.8 $Y=2.635
+ $X2=17.8 $Y2=2.34
r409 115 225 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.995 $Y=2.72
+ $X2=16.86 $Y2=2.72
r410 114 228 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.665 $Y=2.72
+ $X2=17.8 $Y2=2.72
r411 114 115 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.665 $Y=2.72
+ $X2=16.995 $Y2=2.72
r412 110 225 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.86 $Y=2.635
+ $X2=16.86 $Y2=2.72
r413 110 112 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=16.86 $Y=2.635
+ $X2=16.86 $Y2=2
r414 109 222 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.055 $Y=2.72
+ $X2=15.92 $Y2=2.72
r415 108 225 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.725 $Y=2.72
+ $X2=16.86 $Y2=2.72
r416 108 109 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.725 $Y=2.72
+ $X2=16.055 $Y2=2.72
r417 104 222 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.92 $Y=2.635
+ $X2=15.92 $Y2=2.72
r418 104 106 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=15.92 $Y=2.635
+ $X2=15.92 $Y2=2
r419 100 219 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=2.635
+ $X2=14.98 $Y2=2.72
r420 100 102 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.98 $Y=2.635
+ $X2=14.98 $Y2=2
r421 96 216 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.04 $Y=2.635
+ $X2=14.04 $Y2=2.72
r422 96 98 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=14.04 $Y=2.635
+ $X2=14.04 $Y2=2
r423 92 213 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.1 $Y=2.635
+ $X2=13.1 $Y2=2.72
r424 92 94 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=13.1 $Y=2.635
+ $X2=13.1 $Y2=2
r425 88 210 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.16 $Y=2.635
+ $X2=12.16 $Y2=2.72
r426 88 90 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=12.16 $Y=2.635
+ $X2=12.16 $Y2=2
r427 84 207 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=2.635
+ $X2=11.22 $Y2=2.72
r428 84 86 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=11.22 $Y=2.635
+ $X2=11.22 $Y2=2
r429 80 83 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=10.28 $Y=1.66
+ $X2=10.28 $Y2=2.34
r430 78 139 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.28 $Y2=2.72
r431 78 83 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.28 $Y=2.635
+ $X2=10.28 $Y2=2.34
r432 74 77 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=7.36 $Y=1.66
+ $X2=7.36 $Y2=2.34
r433 72 136 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r434 72 77 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.34
r435 68 133 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r436 68 70 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2
r437 64 67 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.48 $Y=1.66
+ $X2=5.48 $Y2=2.34
r438 62 130 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r439 62 67 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.34
r440 58 61 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.54 $Y=1.66
+ $X2=4.54 $Y2=2.34
r441 56 127 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r442 56 61 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.34
r443 52 124 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2.72
r444 52 54 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.6 $Y=2.635
+ $X2=3.6 $Y2=2
r445 48 51 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.66 $Y=1.66
+ $X2=2.66 $Y2=2.34
r446 46 204 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.72
r447 46 51 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.66 $Y=2.635
+ $X2=2.66 $Y2=2.34
r448 15 121 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=17.655
+ $Y=1.485 $X2=17.8 $Y2=2.34
r449 15 118 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=17.655
+ $Y=1.485 $X2=17.8 $Y2=1.66
r450 14 112 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=16.715
+ $Y=1.485 $X2=16.86 $Y2=2
r451 13 106 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=15.775
+ $Y=1.485 $X2=15.92 $Y2=2
r452 12 102 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=14.835
+ $Y=1.485 $X2=14.98 $Y2=2
r453 11 98 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=13.895
+ $Y=1.485 $X2=14.04 $Y2=2
r454 10 94 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.955
+ $Y=1.485 $X2=13.1 $Y2=2
r455 9 90 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=12.015
+ $Y=1.485 $X2=12.16 $Y2=2
r456 8 86 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.075
+ $Y=1.485 $X2=11.22 $Y2=2
r457 7 83 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.28 $Y2=2.34
r458 7 80 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=10.155
+ $Y=1.485 $X2=10.28 $Y2=1.66
r459 6 77 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=2.34
r460 6 74 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.66
r461 5 70 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2
r462 4 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=2.34
r463 4 64 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.66
r464 3 61 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.34
r465 3 58 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.66
r466 2 54 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2
r467 1 51 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=2.34
r468 1 48 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.66 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_597_297# 1 2 3 4 13 15 17 20 23 26 29 30
+ 31 32 34 35 36 37 38 41 45 48 50 51
c138 32 0 1.97192e-19 $X=4.215 $Y=2.21
c139 31 0 1.91318e-19 $X=7.52 $Y=2.21
c140 30 0 1.97192e-19 $X=3.275 $Y=2.21
c141 29 0 1.91318e-19 $X=3.925 $Y=2.21
r142 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.29 $Y=1.87
+ $X2=9.29 $Y2=1.87
r143 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.35 $Y=1.87
+ $X2=8.35 $Y2=1.87
r144 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.07 $Y=2.21
+ $X2=4.07 $Y2=2.21
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.13 $Y=2.21
+ $X2=3.13 $Y2=2.21
r146 38 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.495 $Y=1.87
+ $X2=8.35 $Y2=1.87
r147 37 50 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.145 $Y=1.87
+ $X2=9.29 $Y2=1.87
r148 37 38 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=9.145 $Y=1.87
+ $X2=8.495 $Y2=1.87
r149 35 47 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.205 $Y=1.87
+ $X2=8.35 $Y2=1.87
r150 35 36 0.674504 $w=1.4e-07 $l=5.45e-07 $layer=MET1_cond $X=8.205 $Y=1.87
+ $X2=7.66 $Y2=1.87
r151 33 36 0.0698411 $w=1.4e-07 $l=9.89949e-08 $layer=MET1_cond $X=7.59 $Y=1.94
+ $X2=7.66 $Y2=1.87
r152 33 34 0.247524 $w=1.4e-07 $l=2e-07 $layer=MET1_cond $X=7.59 $Y=1.94
+ $X2=7.59 $Y2=2.14
r153 32 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.215 $Y=2.21
+ $X2=4.07 $Y2=2.21
r154 31 34 0.0698411 $w=1.4e-07 $l=9.89949e-08 $layer=MET1_cond $X=7.52 $Y=2.21
+ $X2=7.59 $Y2=2.14
r155 31 32 4.09034 $w=1.4e-07 $l=3.305e-06 $layer=MET1_cond $X=7.52 $Y=2.21
+ $X2=4.215 $Y2=2.21
r156 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.275 $Y=2.21
+ $X2=3.13 $Y2=2.21
r157 29 44 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.925 $Y=2.21
+ $X2=4.07 $Y2=2.21
r158 29 30 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=3.925 $Y=2.21
+ $X2=3.275 $Y2=2.21
r159 26 51 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.29 $Y=1.665
+ $X2=9.29 $Y2=1.87
r160 26 28 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.29 $Y=1.665
+ $X2=9.29 $Y2=1.58
r161 23 48 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.35 $Y=1.665
+ $X2=8.35 $Y2=1.87
r162 23 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.35 $Y=1.665
+ $X2=8.35 $Y2=1.58
r163 20 45 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=2.21
r164 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=1.665
+ $X2=4.07 $Y2=1.58
r165 17 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=2.21
r166 17 19 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=1.665
+ $X2=3.13 $Y2=1.58
r167 16 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.515 $Y=1.58
+ $X2=8.35 $Y2=1.58
r168 15 28 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.125 $Y=1.58
+ $X2=9.29 $Y2=1.58
r169 15 16 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.125 $Y=1.58
+ $X2=8.515 $Y2=1.58
r170 14 19 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=1.58
+ $X2=3.13 $Y2=1.58
r171 13 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.905 $Y=1.58
+ $X2=4.07 $Y2=1.58
r172 13 14 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.905 $Y=1.58
+ $X2=3.295 $Y2=1.58
r173 4 28 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=9.145
+ $Y=1.485 $X2=9.29 $Y2=1.66
r174 3 25 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=8.205
+ $Y=1.485 $X2=8.35 $Y2=1.66
r175 2 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2.34
r176 2 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.66
r177 1 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.34
r178 1 19 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 53 55 57 58 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 105 107 111 115
+ 117 119 123 127 129 131 135 139 143 145 146 148 149 151 152 154 155 157 158
+ 160 162 165 166
r299 163 166 8.57305 $w=4.08e-07 $l=3.05e-07 $layer=LI1_cond $X=17.29 $Y=1.495
+ $X2=17.29 $Y2=1.19
r300 163 165 2.59952 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.29 $Y=1.495
+ $X2=17.29 $Y2=1.58
r301 161 166 8.01088 $w=4.08e-07 $l=2.85e-07 $layer=LI1_cond $X=17.29 $Y=0.905
+ $X2=17.29 $Y2=1.19
r302 161 162 2.74001 $w=3.7e-07 $l=9e-08 $layer=LI1_cond $X=17.29 $Y=0.905
+ $X2=17.29 $Y2=0.815
r303 137 165 2.59952 $w=3.7e-07 $l=1.03078e-07 $layer=LI1_cond $X=17.33 $Y=1.665
+ $X2=17.29 $Y2=1.58
r304 137 139 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=17.33 $Y=1.665
+ $X2=17.33 $Y2=2.34
r305 133 162 2.74001 $w=3.7e-07 $l=1.08167e-07 $layer=LI1_cond $X=17.33 $Y=0.725
+ $X2=17.29 $Y2=0.815
r306 133 135 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=17.33 $Y=0.725
+ $X2=17.33 $Y2=0.42
r307 132 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.555 $Y=1.58
+ $X2=16.39 $Y2=1.58
r308 131 165 4.24538 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=17.085 $Y=1.58
+ $X2=17.29 $Y2=1.58
r309 131 132 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=17.085 $Y=1.58
+ $X2=16.555 $Y2=1.58
r310 130 158 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=16.555 $Y=0.815
+ $X2=16.39 $Y2=0.815
r311 129 162 4.02741 $w=1.8e-07 $l=2.05e-07 $layer=LI1_cond $X=17.085 $Y=0.815
+ $X2=17.29 $Y2=0.815
r312 129 130 32.6566 $w=1.78e-07 $l=5.3e-07 $layer=LI1_cond $X=17.085 $Y=0.815
+ $X2=16.555 $Y2=0.815
r313 125 160 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.39 $Y=1.665
+ $X2=16.39 $Y2=1.58
r314 125 127 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=16.39 $Y=1.665
+ $X2=16.39 $Y2=2.34
r315 121 158 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=16.39 $Y=0.725
+ $X2=16.39 $Y2=0.815
r316 121 123 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=16.39 $Y=0.725
+ $X2=16.39 $Y2=0.42
r317 120 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.615 $Y=1.58
+ $X2=15.45 $Y2=1.58
r318 119 160 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.225 $Y=1.58
+ $X2=16.39 $Y2=1.58
r319 119 120 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=16.225 $Y=1.58
+ $X2=15.615 $Y2=1.58
r320 118 155 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.615 $Y=0.815
+ $X2=15.45 $Y2=0.815
r321 117 158 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=16.225 $Y=0.815
+ $X2=16.39 $Y2=0.815
r322 117 118 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=16.225 $Y=0.815
+ $X2=15.615 $Y2=0.815
r323 113 157 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=15.45 $Y=1.665
+ $X2=15.45 $Y2=1.58
r324 113 115 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.45 $Y=1.665
+ $X2=15.45 $Y2=2.34
r325 109 155 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=15.45 $Y=0.725
+ $X2=15.45 $Y2=0.815
r326 109 111 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=15.45 $Y=0.725
+ $X2=15.45 $Y2=0.42
r327 108 154 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.675 $Y=1.58
+ $X2=14.51 $Y2=1.58
r328 107 157 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.285 $Y=1.58
+ $X2=15.45 $Y2=1.58
r329 107 108 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=15.285 $Y=1.58
+ $X2=14.675 $Y2=1.58
r330 106 152 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.675 $Y=0.815
+ $X2=14.51 $Y2=0.815
r331 105 155 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=15.285 $Y=0.815
+ $X2=15.45 $Y2=0.815
r332 105 106 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=15.285 $Y=0.815
+ $X2=14.675 $Y2=0.815
r333 101 154 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=14.51 $Y=1.665
+ $X2=14.51 $Y2=1.58
r334 101 103 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=14.51 $Y=1.665
+ $X2=14.51 $Y2=2.34
r335 97 152 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=14.51 $Y=0.725
+ $X2=14.51 $Y2=0.815
r336 97 99 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=14.51 $Y=0.725
+ $X2=14.51 $Y2=0.42
r337 96 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.735 $Y=1.58
+ $X2=13.57 $Y2=1.58
r338 95 154 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=14.345 $Y=1.58
+ $X2=14.51 $Y2=1.58
r339 95 96 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=14.345 $Y=1.58
+ $X2=13.735 $Y2=1.58
r340 94 149 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.735 $Y=0.815
+ $X2=13.57 $Y2=0.815
r341 93 152 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=14.345 $Y=0.815
+ $X2=14.51 $Y2=0.815
r342 93 94 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=14.345 $Y=0.815
+ $X2=13.735 $Y2=0.815
r343 89 151 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.57 $Y=1.665
+ $X2=13.57 $Y2=1.58
r344 89 91 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=13.57 $Y=1.665
+ $X2=13.57 $Y2=2.34
r345 85 149 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=13.57 $Y=0.725
+ $X2=13.57 $Y2=0.815
r346 85 87 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=13.57 $Y=0.725
+ $X2=13.57 $Y2=0.42
r347 84 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=1.58
+ $X2=12.63 $Y2=1.58
r348 83 151 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=1.58
+ $X2=13.57 $Y2=1.58
r349 83 84 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=13.405 $Y=1.58
+ $X2=12.795 $Y2=1.58
r350 82 146 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.795 $Y=0.815
+ $X2=12.63 $Y2=0.815
r351 81 149 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=0.815
+ $X2=13.57 $Y2=0.815
r352 81 82 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=13.405 $Y=0.815
+ $X2=12.795 $Y2=0.815
r353 77 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.63 $Y=1.665
+ $X2=12.63 $Y2=1.58
r354 77 79 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=12.63 $Y=1.665
+ $X2=12.63 $Y2=2.34
r355 73 146 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=12.63 $Y=0.725
+ $X2=12.63 $Y2=0.815
r356 73 75 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=12.63 $Y=0.725
+ $X2=12.63 $Y2=0.42
r357 72 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.855 $Y=1.58
+ $X2=11.69 $Y2=1.58
r358 71 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=1.58
+ $X2=12.63 $Y2=1.58
r359 71 72 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=12.465 $Y=1.58
+ $X2=11.855 $Y2=1.58
r360 70 143 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.855 $Y=0.815
+ $X2=11.69 $Y2=0.815
r361 69 146 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=12.465 $Y=0.815
+ $X2=12.63 $Y2=0.815
r362 69 70 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=12.465 $Y=0.815
+ $X2=11.855 $Y2=0.815
r363 65 145 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.69 $Y=1.665
+ $X2=11.69 $Y2=1.58
r364 65 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.69 $Y=1.665
+ $X2=11.69 $Y2=2.34
r365 61 143 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=11.69 $Y=0.725
+ $X2=11.69 $Y2=0.815
r366 61 63 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=11.69 $Y=0.725
+ $X2=11.69 $Y2=0.42
r367 60 142 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.915 $Y=1.58
+ $X2=10.75 $Y2=1.58
r368 59 145 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=1.58
+ $X2=11.69 $Y2=1.58
r369 59 60 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=11.525 $Y=1.58
+ $X2=10.915 $Y2=1.58
r370 57 143 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=11.525 $Y=0.815
+ $X2=11.69 $Y2=0.815
r371 57 58 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=11.525 $Y=0.815
+ $X2=10.915 $Y2=0.815
r372 53 142 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.75 $Y2=1.58
r373 53 55 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.75 $Y=1.665
+ $X2=10.75 $Y2=2.34
r374 49 58 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=10.75 $Y=0.725
+ $X2=10.915 $Y2=0.815
r375 49 51 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=10.75 $Y=0.725
+ $X2=10.75 $Y2=0.42
r376 16 165 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=17.185
+ $Y=1.485 $X2=17.33 $Y2=1.66
r377 16 139 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=17.185
+ $Y=1.485 $X2=17.33 $Y2=2.34
r378 15 160 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=16.245
+ $Y=1.485 $X2=16.39 $Y2=1.66
r379 15 127 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=16.245
+ $Y=1.485 $X2=16.39 $Y2=2.34
r380 14 157 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=15.305
+ $Y=1.485 $X2=15.45 $Y2=1.66
r381 14 115 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=15.305
+ $Y=1.485 $X2=15.45 $Y2=2.34
r382 13 154 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=14.365
+ $Y=1.485 $X2=14.51 $Y2=1.66
r383 13 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=14.365
+ $Y=1.485 $X2=14.51 $Y2=2.34
r384 12 151 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=13.425
+ $Y=1.485 $X2=13.57 $Y2=1.66
r385 12 91 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.425
+ $Y=1.485 $X2=13.57 $Y2=2.34
r386 11 148 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.63 $Y2=1.66
r387 11 79 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.485
+ $Y=1.485 $X2=12.63 $Y2=2.34
r388 10 145 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.69 $Y2=1.66
r389 10 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.545
+ $Y=1.485 $X2=11.69 $Y2=2.34
r390 9 142 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.485 $X2=10.75 $Y2=1.66
r391 9 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.605
+ $Y=1.485 $X2=10.75 $Y2=2.34
r392 8 135 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=17.195
+ $Y=0.235 $X2=17.33 $Y2=0.42
r393 7 123 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=16.255
+ $Y=0.235 $X2=16.39 $Y2=0.42
r394 6 111 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=15.315
+ $Y=0.235 $X2=15.45 $Y2=0.42
r395 5 99 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=14.375
+ $Y=0.235 $X2=14.51 $Y2=0.42
r396 4 87 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=13.435
+ $Y=0.235 $X2=13.57 $Y2=0.42
r397 3 75 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=12.495
+ $Y=0.235 $X2=12.63 $Y2=0.42
r398 2 63 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=11.555
+ $Y=0.235 $X2=11.69 $Y2=0.42
r399 1 51 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=10.615
+ $Y=0.235 $X2=10.75 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_119_47# 1 2 3 4 15 19 21 25 30 33 34 35
r83 32 34 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.75
+ $X2=1.835 $Y2=0.75
r84 32 33 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.67 $Y=0.75
+ $X2=1.505 $Y2=0.75
r85 30 33 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=0.895 $Y=0.815
+ $X2=1.505 $Y2=0.815
r86 28 30 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.75
+ $X2=0.895 $Y2=0.75
r87 23 25 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.07 $Y=0.725
+ $X2=4.07 $Y2=0.42
r88 22 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.295 $Y=0.815
+ $X2=3.13 $Y2=0.815
r89 21 23 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=3.905 $Y=0.815
+ $X2=4.07 $Y2=0.725
r90 21 22 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=3.905 $Y=0.815
+ $X2=3.295 $Y2=0.815
r91 17 35 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.13 $Y=0.725 $X2=3.13
+ $Y2=0.815
r92 17 19 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=3.13 $Y=0.725
+ $X2=3.13 $Y2=0.42
r93 15 35 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.965 $Y=0.815
+ $X2=3.13 $Y2=0.815
r94 15 34 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=2.965 $Y=0.815
+ $X2=1.835 $Y2=0.815
r95 4 25 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.42
r96 3 19 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.995
+ $Y=0.235 $X2=3.13 $Y2=0.42
r97 2 32 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.76
r98 1 28 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 48 52 56 60 64 68 72 76 80 84 88 92 96 98 102 104 108 111 112 114 115 117 118
+ 120 121 123 124 126 127 128 130 157 161 166 171 176 181 188 189 192 195 198
+ 201 204 207 210 213 216 220
c300 130 0 1.96891e-19 $X=2.525 $Y=0
c301 126 0 1.96891e-19 $X=10.145 $Y=0
r302 216 217 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.71 $Y=0
+ $X2=17.71 $Y2=0
r303 214 217 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.79 $Y=0
+ $X2=17.71 $Y2=0
r304 213 214 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=16.79 $Y=0
+ $X2=16.79 $Y2=0
r305 211 214 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.79 $Y2=0
r306 210 211 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r307 207 208 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r308 204 205 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r309 201 202 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.11 $Y=0
+ $X2=13.11 $Y2=0
r310 198 199 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r311 195 196 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r312 192 193 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r313 189 217 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=0
+ $X2=17.71 $Y2=0
r314 188 189 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=0
+ $X2=18.17 $Y2=0
r315 186 216 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.935 $Y=0
+ $X2=17.8 $Y2=0
r316 186 188 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=17.935 $Y=0
+ $X2=18.17 $Y2=0
r317 185 211 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=15.87 $Y2=0
r318 185 208 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.41 $Y=0
+ $X2=14.95 $Y2=0
r319 184 185 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.41 $Y=0
+ $X2=15.41 $Y2=0
r320 182 207 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.115 $Y=0
+ $X2=14.98 $Y2=0
r321 182 184 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.115 $Y=0
+ $X2=15.41 $Y2=0
r322 181 210 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=15.785 $Y=0
+ $X2=15.92 $Y2=0
r323 181 184 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=15.785 $Y=0
+ $X2=15.41 $Y2=0
r324 180 208 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r325 180 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.03 $Y2=0
r326 179 180 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r327 177 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.175 $Y=0
+ $X2=14.04 $Y2=0
r328 177 179 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=14.175 $Y=0
+ $X2=14.49 $Y2=0
r329 176 207 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=14.845 $Y=0
+ $X2=14.98 $Y2=0
r330 176 179 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=14.845 $Y=0
+ $X2=14.49 $Y2=0
r331 175 205 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r332 175 202 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=13.11 $Y2=0
r333 174 175 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r334 172 201 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.235 $Y=0
+ $X2=13.1 $Y2=0
r335 172 174 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.235 $Y=0
+ $X2=13.57 $Y2=0
r336 171 204 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=13.905 $Y=0
+ $X2=14.04 $Y2=0
r337 171 174 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=13.905 $Y=0
+ $X2=13.57 $Y2=0
r338 170 202 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r339 170 199 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r340 169 170 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r341 167 198 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.16 $Y2=0
r342 167 169 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=12.295 $Y=0
+ $X2=12.65 $Y2=0
r343 166 201 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=13.1 $Y2=0
r344 166 169 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=12.965 $Y=0
+ $X2=12.65 $Y2=0
r345 165 199 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r346 165 196 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r347 164 165 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r348 162 195 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.22 $Y2=0
r349 162 164 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=11.355 $Y=0
+ $X2=11.73 $Y2=0
r350 161 198 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=12.16 $Y2=0
r351 161 164 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.025 $Y=0
+ $X2=11.73 $Y2=0
r352 160 196 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r353 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r354 157 195 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=11.22 $Y2=0
r355 157 159 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=11.085 $Y=0
+ $X2=10.81 $Y2=0
r356 156 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r357 155 156 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r358 153 156 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.89 $Y2=0
r359 152 155 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=9.89 $Y2=0
r360 152 153 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r361 150 153 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r362 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r363 147 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r364 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r365 144 147 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r366 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r367 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r368 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r369 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r370 138 193 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=2.53 $Y2=0
r371 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r372 135 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=2.66 $Y2=0
r373 135 137 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.795 $Y=0
+ $X2=3.45 $Y2=0
r374 132 220 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r375 130 192 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=2.66 $Y2=0
r376 130 132 149.727 $w=1.68e-07 $l=2.295e-06 $layer=LI1_cond $X=2.525 $Y=0
+ $X2=0.23 $Y2=0
r377 128 193 0.653023 $w=4.8e-07 $l=2.295e-06 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=2.53 $Y2=0
r378 128 220 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r379 126 155 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=9.89 $Y2=0
r380 126 127 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.145 $Y=0
+ $X2=10.28 $Y2=0
r381 125 159 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.81 $Y2=0
r382 125 127 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.415 $Y=0
+ $X2=10.28 $Y2=0
r383 123 149 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.13 $Y2=0
r384 123 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.225 $Y=0
+ $X2=7.36 $Y2=0
r385 122 152 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=7.59 $Y2=0
r386 122 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.495 $Y=0
+ $X2=7.36 $Y2=0
r387 120 146 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.21 $Y2=0
r388 120 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.285 $Y=0
+ $X2=6.42 $Y2=0
r389 119 149 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=7.13 $Y2=0
r390 119 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=6.42 $Y2=0
r391 117 143 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.29 $Y2=0
r392 117 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.345 $Y=0
+ $X2=5.48 $Y2=0
r393 116 146 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=6.21 $Y2=0
r394 116 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=5.48 $Y2=0
r395 114 140 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.37 $Y2=0
r396 114 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.405 $Y=0
+ $X2=4.54 $Y2=0
r397 113 143 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=5.29 $Y2=0
r398 113 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=0
+ $X2=4.54 $Y2=0
r399 111 137 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=0
+ $X2=3.45 $Y2=0
r400 111 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.465 $Y=0
+ $X2=3.6 $Y2=0
r401 110 140 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=4.37 $Y2=0
r402 110 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.735 $Y=0
+ $X2=3.6 $Y2=0
r403 106 216 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.8 $Y=0.085
+ $X2=17.8 $Y2=0
r404 106 108 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.8 $Y=0.085
+ $X2=17.8 $Y2=0.38
r405 105 213 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.995 $Y=0
+ $X2=16.86 $Y2=0
r406 104 216 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.665 $Y=0
+ $X2=17.8 $Y2=0
r407 104 105 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.665 $Y=0
+ $X2=16.995 $Y2=0
r408 100 213 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.86 $Y=0.085
+ $X2=16.86 $Y2=0
r409 100 102 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.86 $Y=0.085
+ $X2=16.86 $Y2=0.38
r410 99 210 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.055 $Y=0
+ $X2=15.92 $Y2=0
r411 98 213 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.725 $Y=0
+ $X2=16.86 $Y2=0
r412 98 99 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.725 $Y=0
+ $X2=16.055 $Y2=0
r413 94 210 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.92 $Y=0.085
+ $X2=15.92 $Y2=0
r414 94 96 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=15.92 $Y=0.085
+ $X2=15.92 $Y2=0.38
r415 90 207 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.98 $Y=0.085
+ $X2=14.98 $Y2=0
r416 90 92 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=14.98 $Y=0.085
+ $X2=14.98 $Y2=0.38
r417 86 204 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=14.04 $Y=0.085
+ $X2=14.04 $Y2=0
r418 86 88 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=14.04 $Y=0.085
+ $X2=14.04 $Y2=0.385
r419 82 201 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.1 $Y=0.085
+ $X2=13.1 $Y2=0
r420 82 84 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.1 $Y=0.085
+ $X2=13.1 $Y2=0.38
r421 78 198 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=12.16 $Y=0.085
+ $X2=12.16 $Y2=0
r422 78 80 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=12.16 $Y=0.085
+ $X2=12.16 $Y2=0.38
r423 74 195 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0
r424 74 76 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.22 $Y=0.085
+ $X2=11.22 $Y2=0.38
r425 70 127 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0
r426 70 72 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.28 $Y=0.085
+ $X2=10.28 $Y2=0.38
r427 66 124 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r428 66 68 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.385
r429 62 121 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r430 62 64 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.38
r431 58 118 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r432 58 60 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.38
r433 54 115 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0
r434 54 56 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.54 $Y=0.085
+ $X2=4.54 $Y2=0.38
r435 50 112 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0
r436 50 52 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.38
r437 46 192 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0
r438 46 48 12.8049 $w=2.68e-07 $l=3e-07 $layer=LI1_cond $X=2.66 $Y=0.085
+ $X2=2.66 $Y2=0.385
r439 15 108 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=17.615
+ $Y=0.235 $X2=17.8 $Y2=0.38
r440 14 102 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=16.675
+ $Y=0.235 $X2=16.86 $Y2=0.38
r441 13 96 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=15.735
+ $Y=0.235 $X2=15.92 $Y2=0.38
r442 12 92 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=14.795
+ $Y=0.235 $X2=14.98 $Y2=0.38
r443 11 88 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=13.855
+ $Y=0.235 $X2=14.04 $Y2=0.385
r444 10 84 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=12.915
+ $Y=0.235 $X2=13.1 $Y2=0.38
r445 9 80 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.975
+ $Y=0.235 $X2=12.16 $Y2=0.38
r446 8 76 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.235 $X2=11.22 $Y2=0.38
r447 7 72 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=10.155
+ $Y=0.235 $X2=10.28 $Y2=0.38
r448 6 68 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=7.175
+ $Y=0.235 $X2=7.36 $Y2=0.385
r449 5 64 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.38
r450 4 60 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.235 $X2=5.48 $Y2=0.38
r451 3 56 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.38
r452 2 52 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.6 $Y2=0.38
r453 1 48 182 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.66 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2_16%A_1163_47# 1 2 3 4 15 17 18 21 27 30 31 33
+ 34
r87 33 34 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=9.29 $Y=0.75
+ $X2=9.125 $Y2=0.75
r88 31 34 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=8.515 $Y=0.815
+ $X2=9.125 $Y2=0.815
r89 29 31 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=0.75
+ $X2=8.515 $Y2=0.75
r90 29 30 8.14364 $w=3.08e-07 $l=1.65e-07 $layer=LI1_cond $X=8.35 $Y=0.75
+ $X2=8.185 $Y2=0.75
r91 24 27 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=6.89 $Y2=0.815
r92 24 30 69.6263 $w=1.78e-07 $l=1.13e-06 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=8.185 $Y2=0.815
r93 19 27 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=6.89 $Y=0.725 $X2=6.89
+ $Y2=0.815
r94 19 21 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.89 $Y=0.725
+ $X2=6.89 $Y2=0.42
r95 17 27 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=0.815
+ $X2=6.89 $Y2=0.815
r96 17 18 37.5859 $w=1.78e-07 $l=6.1e-07 $layer=LI1_cond $X=6.725 $Y=0.815
+ $X2=6.115 $Y2=0.815
r97 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=5.95 $Y=0.725
+ $X2=6.115 $Y2=0.815
r98 13 15 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.95 $Y=0.725
+ $X2=5.95 $Y2=0.42
r99 4 33 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=9.155
+ $Y=0.235 $X2=9.29 $Y2=0.76
r100 3 29 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=8.215
+ $Y=0.235 $X2=8.35 $Y2=0.76
r101 2 21 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=6.755
+ $Y=0.235 $X2=6.89 $Y2=0.42
r102 1 15 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=5.815
+ $Y=0.235 $X2=5.95 $Y2=0.42
.ends

