* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__bufinv_16 A VGND VNB VPB VPWR Y
X0 a_391_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_27_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND a_27_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_391_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VPWR a_27_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_391_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VPWR a_27_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 a_391_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_27_47# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_391_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_391_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 VGND a_27_47# a_391_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 a_27_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X43 VPWR a_391_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 Y a_391_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X45 Y a_391_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X48 VPWR a_27_47# a_391_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X49 VGND a_391_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
