* File: sky130_fd_sc_hdll__a222oi_1.spice
* Created: Wed Sep  2 08:18:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a222oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a222oi_1  VNB VPB C1 C2 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C2	C2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1011 A_119_47# N_C1_M1011_g N_Y_M1011_s VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.1984 PD=0.85 PS=1.9 NRD=9.372 NRS=8.436 M=1 R=4.26667 SA=75000.2
+ SB=75003.3 A=0.096 P=1.58 MULT=1
MM1002 N_VGND_M1002_d N_C2_M1002_g A_119_47# VNB NSHORT L=0.15 W=0.64 AD=0.3648
+ AS=0.0672 PD=1.78 PS=0.85 NRD=8.436 NRS=9.372 M=1 R=4.26667 SA=75000.6
+ SB=75002.9 A=0.096 P=1.58 MULT=1
MM1010 A_449_47# N_B2_M1010_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.64 AD=0.0672
+ AS=0.3648 PD=0.85 PS=1.78 NRD=9.372 NRS=89.052 M=1 R=4.26667 SA=75001.9
+ SB=75001.7 A=0.096 P=1.58 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g A_449_47# VNB NSHORT L=0.15 W=0.64 AD=0.1216
+ AS=0.0672 PD=1.02 PS=0.85 NRD=12.18 NRS=9.372 M=1 R=4.26667 SA=75002.2
+ SB=75001.3 A=0.096 P=1.58 MULT=1
MM1005 A_627_47# N_A1_M1005_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.64 AD=0.1216
+ AS=0.1216 PD=1.02 PS=1.02 NRD=25.308 NRS=6.552 M=1 R=4.26667 SA=75002.8
+ SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g A_627_47# VNB NSHORT L=0.15 W=0.64 AD=0.1984
+ AS=0.1216 PD=1.9 PS=1.02 NRD=0 NRS=25.308 M=1 R=4.26667 SA=75003.3 SB=75000.2
+ A=0.096 P=1.58 MULT=1
MM1006 N_A_117_297#_M1006_d N_C1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_C2_M1001_g N_A_117_297#_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_117_297#_M1004_d N_B2_M1004_g N_A_357_297#_M1004_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1000 N_A_357_297#_M1000_d N_B1_M1000_g N_A_117_297#_M1004_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A1_M1009_g N_A_357_297#_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.145 PD=1.35 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1007 N_A_357_297#_M1007_d N_A2_M1007_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.175 PD=2.54 PS=1.35 NRD=0.9653 NRS=12.7853 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__a222oi_1.pxi.spice"
*
.ends
*
*
