* File: sky130_fd_sc_hdll__and2_6.pxi.spice
* Created: Thu Aug 27 18:57:07 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2_6%B N_B_c_86_n N_B_M1007_g N_B_c_87_n N_B_M1001_g
+ N_B_c_88_n N_B_M1012_g N_B_c_89_n N_B_M1015_g N_B_c_90_n N_B_c_95_n N_B_c_96_n
+ N_B_c_143_p N_B_c_97_n N_B_c_91_n N_B_c_92_n B PM_SKY130_FD_SC_HDLL__AND2_6%B
x_PM_SKY130_FD_SC_HDLL__AND2_6%A N_A_c_171_n N_A_M1002_g N_A_c_167_n N_A_M1008_g
+ N_A_c_168_n N_A_M1009_g N_A_c_172_n N_A_M1018_g A N_A_c_169_n N_A_c_170_n
+ PM_SKY130_FD_SC_HDLL__AND2_6%A
x_PM_SKY130_FD_SC_HDLL__AND2_6%A_117_297# N_A_117_297#_M1008_d
+ N_A_117_297#_M1007_d N_A_117_297#_M1018_s N_A_117_297#_c_225_n
+ N_A_117_297#_M1000_g N_A_117_297#_c_215_n N_A_117_297#_M1004_g
+ N_A_117_297#_c_216_n N_A_117_297#_M1006_g N_A_117_297#_c_226_n
+ N_A_117_297#_M1003_g N_A_117_297#_c_227_n N_A_117_297#_M1005_g
+ N_A_117_297#_c_217_n N_A_117_297#_M1010_g N_A_117_297#_c_218_n
+ N_A_117_297#_M1014_g N_A_117_297#_c_228_n N_A_117_297#_M1011_g
+ N_A_117_297#_c_229_n N_A_117_297#_M1013_g N_A_117_297#_c_219_n
+ N_A_117_297#_M1017_g N_A_117_297#_c_220_n N_A_117_297#_M1019_g
+ N_A_117_297#_c_230_n N_A_117_297#_M1016_g N_A_117_297#_c_237_n
+ N_A_117_297#_c_238_n N_A_117_297#_c_240_n N_A_117_297#_c_244_n
+ N_A_117_297#_c_245_n N_A_117_297#_c_221_n N_A_117_297#_c_222_n
+ N_A_117_297#_c_316_p N_A_117_297#_c_255_n N_A_117_297#_c_258_n
+ N_A_117_297#_c_223_n N_A_117_297#_c_224_n
+ PM_SKY130_FD_SC_HDLL__AND2_6%A_117_297#
x_PM_SKY130_FD_SC_HDLL__AND2_6%VPWR N_VPWR_M1007_s N_VPWR_M1002_d N_VPWR_M1015_s
+ N_VPWR_M1003_d N_VPWR_M1011_d N_VPWR_M1016_d N_VPWR_c_381_n N_VPWR_c_382_n
+ N_VPWR_c_383_n N_VPWR_c_384_n N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n VPWR N_VPWR_c_391_n
+ N_VPWR_c_392_n N_VPWR_c_393_n N_VPWR_c_380_n N_VPWR_c_395_n N_VPWR_c_396_n
+ N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n PM_SKY130_FD_SC_HDLL__AND2_6%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2_6%X N_X_M1004_s N_X_M1010_s N_X_M1017_s N_X_M1000_s
+ N_X_M1005_s N_X_M1013_s N_X_c_537_p N_X_c_522_n N_X_c_482_n N_X_c_472_n
+ N_X_c_476_n N_X_c_477_n N_X_c_541_p N_X_c_526_n N_X_c_498_n N_X_c_478_n
+ N_X_c_545_p N_X_c_530_n N_X_c_473_n N_X_c_479_n N_X_c_474_n N_X_c_480_n X
+ PM_SKY130_FD_SC_HDLL__AND2_6%X
x_PM_SKY130_FD_SC_HDLL__AND2_6%VGND N_VGND_M1001_s N_VGND_M1012_s N_VGND_M1006_d
+ N_VGND_M1014_d N_VGND_M1019_d N_VGND_c_557_n N_VGND_c_558_n N_VGND_c_559_n
+ N_VGND_c_560_n N_VGND_c_561_n N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n
+ N_VGND_c_565_n VGND N_VGND_c_566_n N_VGND_c_567_n N_VGND_c_568_n
+ N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n N_VGND_c_572_n
+ PM_SKY130_FD_SC_HDLL__AND2_6%VGND
cc_1 VNB N_B_c_86_n 0.0298625f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B_c_87_n 0.0219327f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_3 VNB N_B_c_88_n 0.0178693f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_4 VNB N_B_c_89_n 0.022373f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_5 VNB N_B_c_90_n 0.00282996f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.325
cc_6 VNB N_B_c_91_n 0.0154282f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_7 VNB N_B_c_92_n 0.00291745f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_8 VNB N_A_c_167_n 0.0159567f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=0.995
cc_9 VNB N_A_c_168_n 0.0163424f $X=-0.19 $Y=-0.24 $X2=1.82 $Y2=0.995
cc_10 VNB N_A_c_169_n 0.00397755f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_11 VNB N_A_c_170_n 0.0340864f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.16
cc_12 VNB N_A_117_297#_c_215_n 0.0174785f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.325
cc_13 VNB N_A_117_297#_c_216_n 0.0168734f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.55
cc_14 VNB N_A_117_297#_c_217_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_15 VNB N_A_117_297#_c_218_n 0.0168771f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_A_117_297#_c_219_n 0.0168638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_117_297#_c_220_n 0.0194565f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_117_297#_c_221_n 0.00243553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_117_297#_c_222_n 2.27519e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_117_297#_c_223_n 0.00125224f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_117_297#_c_224_n 0.115108f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VPWR_c_380_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_472_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_24 VNB N_X_c_473_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_474_n 6.84655e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB X 0.017142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_557_n 0.0115788f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.55
cc_28 VNB N_VGND_c_558_n 0.0287273f $X=-0.19 $Y=-0.24 $X2=1.795 $Y2=1.465
cc_29 VNB N_VGND_c_559_n 0.00506067f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_30 VNB N_VGND_c_560_n 0.017129f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.16
cc_31 VNB N_VGND_c_561_n 0.00446122f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_32 VNB N_VGND_c_562_n 0.0155206f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_33 VNB N_VGND_c_563_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_564_n 0.0155193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_565_n 0.0174479f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_566_n 0.042283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_567_n 0.014713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_568_n 0.287545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_569_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_570_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_571_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_572_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_B_c_86_n 0.0338412f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_44 VPB N_B_c_89_n 0.0250756f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_45 VPB N_B_c_95_n 0.00142318f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.465
cc_46 VPB N_B_c_96_n 0.0121879f $X=-0.19 $Y=1.305 $X2=1.705 $Y2=1.55
cc_47 VPB N_B_c_97_n 0.00133746f $X=-0.19 $Y=1.305 $X2=1.795 $Y2=1.465
cc_48 VPB N_B_c_91_n 0.00449876f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_49 VPB N_B_c_92_n 2.02246e-19 $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_50 VPB N_A_c_171_n 0.0159868f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_A_c_172_n 0.0160012f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_52 VPB N_A_c_170_n 0.0195372f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.16
cc_53 VPB N_A_117_297#_c_225_n 0.0157647f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_54 VPB N_A_117_297#_c_226_n 0.0157176f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_55 VPB N_A_117_297#_c_227_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_56 VPB N_A_117_297#_c_228_n 0.0157197f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=1.16
cc_57 VPB N_A_117_297#_c_229_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_117_297#_c_230_n 0.0184001f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_117_297#_c_222_n 0.0011823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_117_297#_c_224_n 0.0717921f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_381_n 0.0109725f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_62 VPB N_VPWR_c_382_n 0.0313356f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_63 VPB N_VPWR_c_383_n 3.40287e-19 $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.16
cc_64 VPB N_VPWR_c_384_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_385_n 0.0147329f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=1.16
cc_66 VPB N_VPWR_c_386_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_387_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_388_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_389_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_390_n 0.0300286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_391_n 0.015714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_392_n 0.0135016f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_393_n 0.014713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_380_n 0.0557506f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_395_n 0.00436768f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_396_n 0.0043669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_397_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_398_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_399_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_X_c_476_n 0.00184039f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=1.16
cc_81 VPB N_X_c_477_n 0.00201632f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_82 VPB N_X_c_478_n 0.00185796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_X_c_479_n 0.00165339f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_X_c_480_n 0.00258613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB X 0.00626897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 N_B_c_86_n N_A_c_171_n 0.0224096f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_87 N_B_c_95_n N_A_c_171_n 0.00102484f $X=0.525 $Y=1.465 $X2=-0.19 $Y2=-0.24
cc_88 N_B_c_96_n N_A_c_171_n 0.011867f $X=1.705 $Y=1.55 $X2=-0.19 $Y2=-0.24
cc_89 N_B_c_87_n N_A_c_167_n 0.0469093f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B_c_88_n N_A_c_168_n 0.0404173f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B_c_89_n N_A_c_172_n 0.021892f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B_c_96_n N_A_c_172_n 0.011867f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_93 N_B_c_97_n N_A_c_172_n 0.00112883f $X=1.795 $Y=1.465 $X2=0 $Y2=0
cc_94 N_B_c_86_n N_A_c_169_n 0.00106734f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_89_n N_A_c_169_n 3.41921e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_90_n N_A_c_169_n 0.0181146f $X=0.525 $Y=1.325 $X2=0 $Y2=0
cc_97 N_B_c_96_n N_A_c_169_n 0.0486416f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_98 N_B_c_92_n N_A_c_169_n 0.024537f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_99 N_B_c_86_n N_A_c_170_n 0.024873f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_89_n N_A_c_170_n 0.0252145f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B_c_90_n N_A_c_170_n 5.63263e-19 $X=0.525 $Y=1.325 $X2=0 $Y2=0
cc_102 N_B_c_95_n N_A_c_170_n 0.00160606f $X=0.525 $Y=1.465 $X2=0 $Y2=0
cc_103 N_B_c_96_n N_A_c_170_n 0.0081456f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_104 N_B_c_92_n N_A_c_170_n 0.00340829f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_105 N_B_c_96_n N_A_117_297#_M1007_d 0.00187091f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_106 N_B_c_96_n N_A_117_297#_M1018_s 0.00187127f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_107 N_B_c_89_n N_A_117_297#_c_225_n 0.033347f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B_c_88_n N_A_117_297#_c_215_n 0.0205121f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_c_96_n N_A_117_297#_c_237_n 0.0371166f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_110 N_B_c_87_n N_A_117_297#_c_238_n 0.00119819f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_111 N_B_c_88_n N_A_117_297#_c_238_n 0.0015362f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B_c_88_n N_A_117_297#_c_240_n 0.0124097f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_89_n N_A_117_297#_c_240_n 0.00353141f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_96_n N_A_117_297#_c_240_n 0.0045795f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_115 N_B_c_92_n N_A_117_297#_c_240_n 0.0161726f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B_c_87_n N_A_117_297#_c_244_n 5.07286e-19 $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_117 N_B_c_89_n N_A_117_297#_c_245_n 0.0134453f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B_c_96_n N_A_117_297#_c_245_n 0.0052294f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_119 N_B_c_92_n N_A_117_297#_c_245_n 0.00243107f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_120 N_B_c_88_n N_A_117_297#_c_221_n 0.00343684f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_89_n N_A_117_297#_c_221_n 3.83145e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B_c_92_n N_A_117_297#_c_221_n 0.00439055f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B_c_89_n N_A_117_297#_c_222_n 0.00625836f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_c_96_n N_A_117_297#_c_222_n 0.00994131f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_125 N_B_c_97_n N_A_117_297#_c_222_n 0.00746569f $X=1.795 $Y=1.465 $X2=0 $Y2=0
cc_126 N_B_c_92_n N_A_117_297#_c_222_n 0.00439055f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_127 N_B_c_86_n N_A_117_297#_c_255_n 0.00769618f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B_c_96_n N_A_117_297#_c_255_n 0.0142842f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_129 N_B_c_143_p N_A_117_297#_c_255_n 0.00163947f $X=0.615 $Y=1.55 $X2=0 $Y2=0
cc_130 N_B_c_96_n N_A_117_297#_c_258_n 0.0146933f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_131 N_B_c_89_n N_A_117_297#_c_223_n 0.00156266f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B_c_92_n N_A_117_297#_c_223_n 0.017424f $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_133 N_B_c_89_n N_A_117_297#_c_224_n 0.0218009f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_134 N_B_c_92_n N_A_117_297#_c_224_n 2.86091e-19 $X=1.88 $Y=1.16 $X2=0 $Y2=0
cc_135 N_B_c_96_n N_VPWR_M1002_d 0.00187547f $X=1.705 $Y=1.55 $X2=0 $Y2=0
cc_136 N_B_c_86_n N_VPWR_c_382_n 0.00463531f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_137 N_B_c_91_n N_VPWR_c_382_n 0.0110835f $X=0.435 $Y=1.16 $X2=0 $Y2=0
cc_138 N_B_c_86_n N_VPWR_c_383_n 4.46241e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_139 N_B_c_89_n N_VPWR_c_383_n 5.16374e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_140 N_B_c_89_n N_VPWR_c_384_n 0.00819135f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B_c_86_n N_VPWR_c_391_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B_c_89_n N_VPWR_c_392_n 0.00469105f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B_c_86_n N_VPWR_c_380_n 0.012655f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B_c_89_n N_VPWR_c_380_n 0.00545209f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_145 N_B_c_86_n N_VGND_c_558_n 0.00239208f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_146 N_B_c_87_n N_VGND_c_558_n 0.0207834f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_91_n N_VGND_c_558_n 0.0280967f $X=0.435 $Y=1.16 $X2=0 $Y2=0
cc_148 N_B_c_88_n N_VGND_c_559_n 0.00467817f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_149 N_B_c_87_n N_VGND_c_566_n 0.00585385f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_150 N_B_c_88_n N_VGND_c_566_n 0.00428022f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_87_n N_VGND_c_568_n 0.0117974f $X=0.58 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_88_n N_VGND_c_568_n 0.00622853f $X=1.82 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_171_n N_A_117_297#_c_237_n 0.011717f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_172_n N_A_117_297#_c_237_n 0.011717f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_c_167_n N_A_117_297#_c_238_n 0.00762373f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_168_n N_A_117_297#_c_238_n 0.00771706f $X=1.39 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_168_n N_A_117_297#_c_240_n 0.00826322f $X=1.39 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_169_n N_A_117_297#_c_240_n 0.011531f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_c_170_n N_A_117_297#_c_240_n 0.00169164f $X=1.39 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_c_167_n N_A_117_297#_c_244_n 0.00355778f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_168_n N_A_117_297#_c_244_n 8.67038e-19 $X=1.39 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_169_n N_A_117_297#_c_244_n 0.0214622f $X=1.37 $Y=1.16 $X2=0 $Y2=0
cc_163 N_A_c_170_n N_A_117_297#_c_244_n 0.00208238f $X=1.39 $Y=1.202 $X2=0 $Y2=0
cc_164 N_A_c_171_n N_VPWR_c_383_n 0.00787198f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_172_n N_VPWR_c_383_n 0.00781221f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_172_n N_VPWR_c_384_n 5.12605e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_171_n N_VPWR_c_391_n 0.00469105f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_172_n N_VPWR_c_392_n 0.00469105f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_171_n N_VPWR_c_380_n 0.00545209f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_172_n N_VPWR_c_380_n 0.00545209f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_167_n N_VGND_c_566_n 0.00541359f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_168_n N_VGND_c_566_n 0.00415469f $X=1.39 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_167_n N_VGND_c_568_n 0.00964924f $X=0.97 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_c_168_n N_VGND_c_568_n 0.00579893f $X=1.39 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_117_297#_c_237_n N_VPWR_M1002_d 0.00348603f $X=1.535 $Y=1.89 $X2=0
+ $Y2=0
cc_176 N_A_117_297#_c_245_n N_VPWR_M1015_s 0.00504258f $X=2.135 $Y=1.89 $X2=0
+ $Y2=0
cc_177 N_A_117_297#_c_222_n N_VPWR_M1015_s 0.00336092f $X=2.22 $Y=1.805 $X2=0
+ $Y2=0
cc_178 N_A_117_297#_c_237_n N_VPWR_c_383_n 0.0165599f $X=1.535 $Y=1.89 $X2=0
+ $Y2=0
cc_179 N_A_117_297#_c_225_n N_VPWR_c_384_n 0.00819057f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_117_297#_c_226_n N_VPWR_c_384_n 5.12605e-19 $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_117_297#_c_245_n N_VPWR_c_384_n 0.0161564f $X=2.135 $Y=1.89 $X2=0
+ $Y2=0
cc_182 N_A_117_297#_c_225_n N_VPWR_c_385_n 0.00622633f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_117_297#_c_226_n N_VPWR_c_385_n 0.00622633f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_117_297#_c_225_n N_VPWR_c_386_n 6.06824e-19 $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_117_297#_c_226_n N_VPWR_c_386_n 0.0125911f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_117_297#_c_227_n N_VPWR_c_386_n 0.0125911f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_117_297#_c_228_n N_VPWR_c_386_n 6.06824e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_117_297#_c_227_n N_VPWR_c_387_n 0.00622633f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_117_297#_c_228_n N_VPWR_c_387_n 0.00622633f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_117_297#_c_227_n N_VPWR_c_388_n 6.06824e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_117_297#_c_228_n N_VPWR_c_388_n 0.0125911f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_117_297#_c_229_n N_VPWR_c_388_n 0.0125911f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_117_297#_c_230_n N_VPWR_c_388_n 6.06824e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_117_297#_c_229_n N_VPWR_c_389_n 0.00622633f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_117_297#_c_230_n N_VPWR_c_389_n 0.00622633f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_196 N_A_117_297#_c_229_n N_VPWR_c_390_n 6.06824e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_117_297#_c_230_n N_VPWR_c_390_n 0.0142536f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_117_297#_c_237_n N_VPWR_c_391_n 0.00211388f $X=1.535 $Y=1.89 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_c_255_n N_VPWR_c_391_n 0.017264f $X=0.73 $Y=1.96 $X2=0 $Y2=0
cc_200 N_A_117_297#_c_237_n N_VPWR_c_392_n 0.00211388f $X=1.535 $Y=1.89 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_c_245_n N_VPWR_c_392_n 0.00211388f $X=2.135 $Y=1.89 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_c_258_n N_VPWR_c_392_n 0.0156136f $X=1.67 $Y=1.96 $X2=0
+ $Y2=0
cc_203 N_A_117_297#_M1007_d N_VPWR_c_380_n 0.00235201f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_M1018_s N_VPWR_c_380_n 0.00239141f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_c_225_n N_VPWR_c_380_n 0.0104011f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_c_226_n N_VPWR_c_380_n 0.0104011f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_117_297#_c_227_n N_VPWR_c_380_n 0.0104011f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_117_297#_c_228_n N_VPWR_c_380_n 0.0104011f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_117_297#_c_229_n N_VPWR_c_380_n 0.0104011f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_117_297#_c_230_n N_VPWR_c_380_n 0.0104011f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_117_297#_c_237_n N_VPWR_c_380_n 0.00840516f $X=1.535 $Y=1.89 $X2=0
+ $Y2=0
cc_212 N_A_117_297#_c_245_n N_VPWR_c_380_n 0.00492978f $X=2.135 $Y=1.89 $X2=0
+ $Y2=0
cc_213 N_A_117_297#_c_255_n N_VPWR_c_380_n 0.0113082f $X=0.73 $Y=1.96 $X2=0
+ $Y2=0
cc_214 N_A_117_297#_c_258_n N_VPWR_c_380_n 0.010313f $X=1.67 $Y=1.96 $X2=0 $Y2=0
cc_215 N_A_117_297#_c_216_n N_X_c_482_n 0.0106343f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_117_297#_c_217_n N_X_c_482_n 0.0106343f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_117_297#_c_316_p N_X_c_482_n 0.0428524f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A_117_297#_c_224_n N_X_c_482_n 0.00457246f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A_117_297#_c_215_n N_X_c_472_n 0.00115949f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A_117_297#_c_216_n N_X_c_472_n 0.00145892f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_117_297#_c_316_p N_X_c_472_n 0.01642f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_117_297#_c_224_n N_X_c_472_n 0.00224547f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_223 N_A_117_297#_c_226_n N_X_c_476_n 0.015168f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_117_297#_c_227_n N_X_c_476_n 0.0152439f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_117_297#_c_316_p N_X_c_476_n 0.0451906f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_117_297#_c_224_n N_X_c_476_n 0.00802533f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_227 N_A_117_297#_c_225_n N_X_c_477_n 3.65096e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_117_297#_c_222_n N_X_c_477_n 0.00760681f $X=2.22 $Y=1.805 $X2=0 $Y2=0
cc_229 N_A_117_297#_c_316_p N_X_c_477_n 0.0211577f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_117_297#_c_224_n N_X_c_477_n 0.00748099f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_231 N_A_117_297#_c_218_n N_X_c_498_n 0.0106343f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_117_297#_c_219_n N_X_c_498_n 0.0112061f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_117_297#_c_316_p N_X_c_498_n 0.0394413f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_117_297#_c_224_n N_X_c_498_n 0.00457246f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_235 N_A_117_297#_c_228_n N_X_c_478_n 0.0152439f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_117_297#_c_229_n N_X_c_478_n 0.0156962f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_117_297#_c_316_p N_X_c_478_n 0.0418984f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_117_297#_c_224_n N_X_c_478_n 0.00807f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A_117_297#_c_316_p N_X_c_473_n 0.01642f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_117_297#_c_224_n N_X_c_473_n 0.00224547f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_117_297#_c_316_p N_X_c_479_n 0.0211577f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_117_297#_c_224_n N_X_c_479_n 0.00748099f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_243 N_A_117_297#_c_220_n N_X_c_474_n 0.00924485f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_117_297#_c_224_n N_X_c_474_n 9.29358e-19 $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_245 N_A_117_297#_c_230_n N_X_c_480_n 0.0149179f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_117_297#_c_224_n N_X_c_480_n 0.00407701f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_247 N_A_117_297#_c_219_n X 0.00161795f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_117_297#_c_220_n X 0.0044983f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A_117_297#_c_230_n X 0.00154471f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_117_297#_c_316_p X 0.017118f $X=4.14 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_117_297#_c_224_n X 0.037839f $X=4.7 $Y=1.202 $X2=0 $Y2=0
cc_252 N_A_117_297#_c_240_n N_VGND_M1012_s 0.0094216f $X=2.135 $Y=0.74 $X2=0
+ $Y2=0
cc_253 N_A_117_297#_c_221_n N_VGND_M1012_s 7.20909e-19 $X=2.22 $Y=1.055 $X2=0
+ $Y2=0
cc_254 N_A_117_297#_c_238_n N_VGND_c_558_n 0.0116359f $X=1.18 $Y=0.38 $X2=0
+ $Y2=0
cc_255 N_A_117_297#_c_244_n N_VGND_c_558_n 0.00522624f $X=1.345 $Y=0.74 $X2=0
+ $Y2=0
cc_256 N_A_117_297#_c_215_n N_VGND_c_559_n 0.00323651f $X=2.4 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_117_297#_c_240_n N_VGND_c_559_n 0.0252938f $X=2.135 $Y=0.74 $X2=0
+ $Y2=0
cc_258 N_A_117_297#_c_215_n N_VGND_c_560_n 0.00585385f $X=2.4 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_117_297#_c_216_n N_VGND_c_560_n 0.00436487f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_117_297#_c_216_n N_VGND_c_561_n 0.00185632f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_261 N_A_117_297#_c_217_n N_VGND_c_561_n 0.00181032f $X=3.34 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_117_297#_c_217_n N_VGND_c_562_n 0.00436487f $X=3.34 $Y=0.995 $X2=0
+ $Y2=0
cc_263 N_A_117_297#_c_218_n N_VGND_c_562_n 0.00436487f $X=3.76 $Y=0.995 $X2=0
+ $Y2=0
cc_264 N_A_117_297#_c_218_n N_VGND_c_563_n 0.00181032f $X=3.76 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_117_297#_c_219_n N_VGND_c_563_n 0.00181032f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_266 N_A_117_297#_c_219_n N_VGND_c_564_n 0.00436487f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_267 N_A_117_297#_c_220_n N_VGND_c_564_n 0.00436349f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_268 N_A_117_297#_c_220_n N_VGND_c_565_n 0.00356356f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_269 N_A_117_297#_c_238_n N_VGND_c_566_n 0.018715f $X=1.18 $Y=0.38 $X2=0 $Y2=0
cc_270 N_A_117_297#_c_240_n N_VGND_c_566_n 0.0084616f $X=2.135 $Y=0.74 $X2=0
+ $Y2=0
cc_271 N_A_117_297#_M1008_d N_VGND_c_568_n 0.00215201f $X=1.045 $Y=0.235 $X2=0
+ $Y2=0
cc_272 N_A_117_297#_c_215_n N_VGND_c_568_n 0.011086f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_117_297#_c_216_n N_VGND_c_568_n 0.00612685f $X=2.82 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_117_297#_c_217_n N_VGND_c_568_n 0.00608257f $X=3.34 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_117_297#_c_218_n N_VGND_c_568_n 0.00608257f $X=3.76 $Y=0.995 $X2=0
+ $Y2=0
cc_276 N_A_117_297#_c_219_n N_VGND_c_568_n 0.00608257f $X=4.28 $Y=0.995 $X2=0
+ $Y2=0
cc_277 N_A_117_297#_c_220_n N_VGND_c_568_n 0.00720554f $X=4.7 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_117_297#_c_238_n N_VGND_c_568_n 0.0121647f $X=1.18 $Y=0.38 $X2=0
+ $Y2=0
cc_279 N_A_117_297#_c_240_n N_VGND_c_568_n 0.0177614f $X=2.135 $Y=0.74 $X2=0
+ $Y2=0
cc_280 N_A_117_297#_c_240_n A_131_47# 0.00622249f $X=2.135 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_281 N_VPWR_c_380_n N_X_M1000_s 0.00300692f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_380_n N_X_M1005_s 0.00300692f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_380_n N_X_M1013_s 0.00300692f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_385_n N_X_c_522_n 0.0156407f $X=2.915 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_380_n N_X_c_522_n 0.0103212f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_M1003_d N_X_c_476_n 0.00187091f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_c_386_n N_X_c_476_n 0.0171295f $X=3.08 $Y=1.89 $X2=0 $Y2=0
cc_288 N_VPWR_c_387_n N_X_c_526_n 0.0156407f $X=3.855 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_380_n N_X_c_526_n 0.0103212f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_M1011_d N_X_c_478_n 0.00187091f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_291 N_VPWR_c_388_n N_X_c_478_n 0.0171295f $X=4.02 $Y=1.89 $X2=0 $Y2=0
cc_292 N_VPWR_c_389_n N_X_c_530_n 0.0156407f $X=4.795 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_380_n N_X_c_530_n 0.0103212f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_M1016_d N_X_c_480_n 0.00700419f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_295 N_VPWR_c_390_n N_X_c_480_n 0.0108527f $X=4.96 $Y=1.89 $X2=0 $Y2=0
cc_296 N_X_c_482_n N_VGND_M1006_d 0.00500594f $X=3.415 $Y=0.8 $X2=0 $Y2=0
cc_297 N_X_c_498_n N_VGND_M1014_d 0.00500594f $X=4.355 $Y=0.8 $X2=0 $Y2=0
cc_298 N_X_c_474_n N_VGND_M1019_d 0.00932143f $X=4.665 $Y=0.8 $X2=0 $Y2=0
cc_299 N_X_c_537_p N_VGND_c_560_n 0.0148827f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_300 N_X_c_482_n N_VGND_c_560_n 0.00219745f $X=3.415 $Y=0.8 $X2=0 $Y2=0
cc_301 N_X_c_482_n N_VGND_c_561_n 0.0199861f $X=3.415 $Y=0.8 $X2=0 $Y2=0
cc_302 N_X_c_482_n N_VGND_c_562_n 0.00219745f $X=3.415 $Y=0.8 $X2=0 $Y2=0
cc_303 N_X_c_541_p N_VGND_c_562_n 0.0148827f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_304 N_X_c_498_n N_VGND_c_562_n 0.00219745f $X=4.355 $Y=0.8 $X2=0 $Y2=0
cc_305 N_X_c_498_n N_VGND_c_563_n 0.0199861f $X=4.355 $Y=0.8 $X2=0 $Y2=0
cc_306 N_X_c_498_n N_VGND_c_564_n 0.00219745f $X=4.355 $Y=0.8 $X2=0 $Y2=0
cc_307 N_X_c_545_p N_VGND_c_564_n 0.0149192f $X=4.49 $Y=0.42 $X2=0 $Y2=0
cc_308 N_X_c_474_n N_VGND_c_564_n 0.00240483f $X=4.665 $Y=0.8 $X2=0 $Y2=0
cc_309 N_X_c_474_n N_VGND_c_565_n 0.0123344f $X=4.665 $Y=0.8 $X2=0 $Y2=0
cc_310 N_X_M1004_s N_VGND_c_568_n 0.00215201f $X=2.475 $Y=0.235 $X2=0 $Y2=0
cc_311 N_X_M1010_s N_VGND_c_568_n 0.00215201f $X=3.415 $Y=0.235 $X2=0 $Y2=0
cc_312 N_X_M1017_s N_VGND_c_568_n 0.00215201f $X=4.355 $Y=0.235 $X2=0 $Y2=0
cc_313 N_X_c_537_p N_VGND_c_568_n 0.0103005f $X=2.61 $Y=0.56 $X2=0 $Y2=0
cc_314 N_X_c_482_n N_VGND_c_568_n 0.00879353f $X=3.415 $Y=0.8 $X2=0 $Y2=0
cc_315 N_X_c_541_p N_VGND_c_568_n 0.0103005f $X=3.55 $Y=0.42 $X2=0 $Y2=0
cc_316 N_X_c_498_n N_VGND_c_568_n 0.00877625f $X=4.355 $Y=0.8 $X2=0 $Y2=0
cc_317 N_X_c_545_p N_VGND_c_568_n 0.010312f $X=4.49 $Y=0.42 $X2=0 $Y2=0
cc_318 N_X_c_474_n N_VGND_c_568_n 0.00481487f $X=4.665 $Y=0.8 $X2=0 $Y2=0
cc_319 N_VGND_c_568_n A_293_47# 0.0102589f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
cc_320 N_VGND_c_568_n A_131_47# 0.00335103f $X=5.29 $Y=0 $X2=-0.19 $Y2=-0.24
