* File: sky130_fd_sc_hdll__o221ai_4.pxi.spice
* Created: Wed Sep  2 08:45:07 2020
* 
x_PM_SKY130_FD_SC_HDLL__O221AI_4%C1 N_C1_c_128_n N_C1_M1000_g N_C1_c_122_n
+ N_C1_M1006_g N_C1_c_129_n N_C1_M1008_g N_C1_c_123_n N_C1_M1016_g N_C1_c_130_n
+ N_C1_M1012_g N_C1_c_124_n N_C1_M1020_g N_C1_c_131_n N_C1_M1024_g N_C1_c_125_n
+ N_C1_M1031_g C1 N_C1_c_126_n N_C1_c_127_n C1 PM_SKY130_FD_SC_HDLL__O221AI_4%C1
x_PM_SKY130_FD_SC_HDLL__O221AI_4%B1 N_B1_c_191_n N_B1_M1013_g N_B1_c_183_n
+ N_B1_M1021_g N_B1_c_192_n N_B1_M1018_g N_B1_c_184_n N_B1_M1023_g N_B1_c_193_n
+ N_B1_M1028_g N_B1_c_185_n N_B1_M1033_g N_B1_c_186_n N_B1_M1034_g N_B1_c_187_n
+ N_B1_M1037_g N_B1_c_195_n N_B1_c_196_n N_B1_c_203_p N_B1_c_188_n N_B1_c_189_n
+ B1 N_B1_c_190_n B1 PM_SKY130_FD_SC_HDLL__O221AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O221AI_4%B2 N_B2_c_282_n N_B2_M1007_g N_B2_c_288_n
+ N_B2_M1001_g N_B2_c_283_n N_B2_M1027_g N_B2_c_289_n N_B2_M1010_g N_B2_c_284_n
+ N_B2_M1029_g N_B2_c_290_n N_B2_M1025_g N_B2_c_291_n N_B2_M1030_g N_B2_c_285_n
+ N_B2_M1039_g B2 N_B2_c_286_n N_B2_c_287_n B2 PM_SKY130_FD_SC_HDLL__O221AI_4%B2
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A1 N_A1_c_354_n N_A1_M1003_g N_A1_c_355_n
+ N_A1_M1009_g N_A1_c_356_n N_A1_M1011_g N_A1_c_363_n N_A1_M1022_g N_A1_c_357_n
+ N_A1_M1014_g N_A1_c_364_n N_A1_M1026_g N_A1_c_358_n N_A1_M1032_g N_A1_c_365_n
+ N_A1_M1035_g N_A1_c_366_n N_A1_c_359_n N_A1_c_367_n N_A1_c_360_n A1
+ N_A1_c_425_p N_A1_c_361_n A1 PM_SKY130_FD_SC_HDLL__O221AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A2 N_A2_c_468_n N_A2_M1004_g N_A2_c_474_n
+ N_A2_M1002_g N_A2_c_469_n N_A2_M1017_g N_A2_c_475_n N_A2_M1005_g N_A2_c_470_n
+ N_A2_M1019_g N_A2_c_476_n N_A2_M1015_g N_A2_c_477_n N_A2_M1038_g N_A2_c_471_n
+ N_A2_M1036_g A2 N_A2_c_472_n N_A2_c_473_n A2 PM_SKY130_FD_SC_HDLL__O221AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O221AI_4%VPWR N_VPWR_M1000_s N_VPWR_M1008_s
+ N_VPWR_M1024_s N_VPWR_M1018_d N_VPWR_M1034_d N_VPWR_M1022_s N_VPWR_M1035_s
+ N_VPWR_c_550_n N_VPWR_c_551_n N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n
+ N_VPWR_c_555_n N_VPWR_c_556_n N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n
+ N_VPWR_c_560_n N_VPWR_c_561_n N_VPWR_c_562_n N_VPWR_c_563_n N_VPWR_c_564_n
+ VPWR N_VPWR_c_565_n N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_568_n
+ N_VPWR_c_549_n PM_SKY130_FD_SC_HDLL__O221AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O221AI_4%Y N_Y_M1006_d N_Y_M1020_d N_Y_M1000_d
+ N_Y_M1012_d N_Y_M1001_s N_Y_M1025_s N_Y_M1002_d N_Y_M1015_d N_Y_c_679_n
+ N_Y_c_746_n N_Y_c_681_n N_Y_c_748_n N_Y_c_680_n N_Y_c_683_n N_Y_c_715_n
+ N_Y_c_684_n N_Y_c_685_n Y N_Y_c_717_n PM_SKY130_FD_SC_HDLL__O221AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A_601_297# N_A_601_297#_M1013_s
+ N_A_601_297#_M1028_s N_A_601_297#_M1010_d N_A_601_297#_M1030_d
+ N_A_601_297#_c_808_n N_A_601_297#_c_797_n N_A_601_297#_c_824_n
+ N_A_601_297#_c_825_n N_A_601_297#_c_813_n N_A_601_297#_c_799_n
+ PM_SKY130_FD_SC_HDLL__O221AI_4%A_601_297#
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A_1369_297# N_A_1369_297#_M1003_d
+ N_A_1369_297#_M1005_s N_A_1369_297#_M1038_s N_A_1369_297#_M1026_d
+ N_A_1369_297#_c_836_n N_A_1369_297#_c_871_n N_A_1369_297#_c_838_n
+ N_A_1369_297#_c_843_n N_A_1369_297#_c_831_n N_A_1369_297#_c_864_n
+ PM_SKY130_FD_SC_HDLL__O221AI_4%A_1369_297#
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1016_s
+ N_A_27_47#_M1031_s N_A_27_47#_M1021_d N_A_27_47#_M1033_d N_A_27_47#_M1027_s
+ N_A_27_47#_M1039_s N_A_27_47#_c_873_n N_A_27_47#_c_874_n N_A_27_47#_c_875_n
+ PM_SKY130_FD_SC_HDLL__O221AI_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_4%A_511_47# N_A_511_47#_M1021_s
+ N_A_511_47#_M1023_s N_A_511_47#_M1007_d N_A_511_47#_M1029_d
+ N_A_511_47#_M1037_s N_A_511_47#_M1004_d N_A_511_47#_M1019_d
+ N_A_511_47#_M1011_s N_A_511_47#_M1032_s N_A_511_47#_c_1014_p
+ N_A_511_47#_c_920_n N_A_511_47#_c_950_n N_A_511_47#_c_921_n
+ N_A_511_47#_c_979_n N_A_511_47#_c_922_n N_A_511_47#_c_954_n
+ N_A_511_47#_c_923_n N_A_511_47#_c_924_n N_A_511_47#_c_925_n
+ N_A_511_47#_c_926_n N_A_511_47#_c_927_n N_A_511_47#_c_928_n
+ N_A_511_47#_c_929_n PM_SKY130_FD_SC_HDLL__O221AI_4%A_511_47#
x_PM_SKY130_FD_SC_HDLL__O221AI_4%VGND N_VGND_M1009_d N_VGND_M1017_s
+ N_VGND_M1036_s N_VGND_M1014_d N_VGND_c_1047_n N_VGND_c_1048_n N_VGND_c_1049_n
+ N_VGND_c_1050_n N_VGND_c_1051_n N_VGND_c_1052_n N_VGND_c_1053_n
+ N_VGND_c_1054_n N_VGND_c_1055_n N_VGND_c_1056_n N_VGND_c_1057_n
+ N_VGND_c_1058_n VGND N_VGND_c_1059_n N_VGND_c_1060_n
+ PM_SKY130_FD_SC_HDLL__O221AI_4%VGND
cc_1 VNB N_C1_c_122_n 0.0222098f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB N_C1_c_123_n 0.0169723f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB N_C1_c_124_n 0.0169687f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_4 VNB N_C1_c_125_n 0.0196785f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_C1_c_126_n 0.0153245f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.16
cc_6 VNB N_C1_c_127_n 0.0896685f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_B1_c_183_n 0.0204963f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_8 VNB N_B1_c_184_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_9 VNB N_B1_c_185_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=0.995
cc_10 VNB N_B1_c_186_n 0.0221872f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_11 VNB N_B1_c_187_n 0.0177944f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_12 VNB N_B1_c_188_n 0.0114212f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.16
cc_13 VNB N_B1_c_189_n 0.00353116f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_14 VNB N_B1_c_190_n 0.0621321f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B2_c_282_n 0.0167331f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_16 VNB N_B2_c_283_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_17 VNB N_B2_c_284_n 0.0174163f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_18 VNB N_B2_c_285_n 0.0176273f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_19 VNB N_B2_c_286_n 0.00219191f $X=-0.19 $Y=-0.24 $X2=1.48 $Y2=1.202
cc_20 VNB N_B2_c_287_n 0.0724595f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.202
cc_21 VNB N_A1_c_354_n 0.0222042f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_22 VNB N_A1_c_355_n 0.017338f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_23 VNB N_A1_c_356_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_24 VNB N_A1_c_357_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_25 VNB N_A1_c_358_n 0.0219568f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_26 VNB N_A1_c_359_n 0.00149193f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_27 VNB N_A1_c_360_n 0.00352495f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_28 VNB N_A1_c_361_n 0.0696468f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A2_c_468_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_30 VNB N_A2_c_469_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_31 VNB N_A2_c_470_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.41
cc_32 VNB N_A2_c_471_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_33 VNB N_A2_c_472_n 0.00275279f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.16
cc_34 VNB N_A2_c_473_n 0.0725593f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_35 VNB N_VPWR_c_549_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_679_n 0.00272401f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.105
cc_37 VNB N_Y_c_680_n 0.0106174f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.175
cc_38 VNB N_A_27_47#_c_873_n 0.00926099f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_39 VNB N_A_27_47#_c_874_n 0.0178018f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_40 VNB N_A_27_47#_c_875_n 0.0115835f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.16
cc_41 VNB N_A_511_47#_c_920_n 0.00343671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_511_47#_c_921_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_511_47#_c_922_n 0.00424067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_511_47#_c_923_n 0.0158613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_511_47#_c_924_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_511_47#_c_925_n 0.00253999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_511_47#_c_926_n 0.00878678f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_511_47#_c_927_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_511_47#_c_928_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_511_47#_c_929_n 0.00252071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_1047_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.985
cc_52 VNB N_VGND_c_1048_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_53 VNB N_VGND_c_1049_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_54 VNB N_VGND_c_1050_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_55 VNB N_VGND_c_1051_n 0.158938f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_56 VNB N_VGND_c_1052_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_57 VNB N_VGND_c_1053_n 0.019187f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_58 VNB N_VGND_c_1054_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_59 VNB N_VGND_c_1055_n 0.0193072f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.202
cc_60 VNB N_VGND_c_1056_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.66 $Y2=1.16
cc_61 VNB N_VGND_c_1057_n 0.019187f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_62 VNB N_VGND_c_1058_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_63 VNB N_VGND_c_1059_n 0.0196191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_1060_n 0.490906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VPB N_C1_c_128_n 0.0210739f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_66 VPB N_C1_c_129_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_67 VPB N_C1_c_130_n 0.0158724f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_68 VPB N_C1_c_131_n 0.0191784f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_69 VPB N_C1_c_127_n 0.0523058f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_70 VPB N_B1_c_191_n 0.0194081f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_71 VPB N_B1_c_192_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_72 VPB N_B1_c_193_n 0.0160057f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_73 VPB N_B1_c_186_n 0.0256643f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_74 VPB N_B1_c_195_n 0.00122397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B1_c_196_n 0.0068192f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_76 VPB N_B1_c_189_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.202
cc_77 VPB N_B1_c_190_n 0.034591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_B2_c_288_n 0.015997f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_79 VPB N_B2_c_289_n 0.0158995f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_80 VPB N_B2_c_290_n 0.0158664f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_81 VPB N_B2_c_291_n 0.0159964f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_82 VPB N_B2_c_287_n 0.0456211f $X=-0.19 $Y=1.305 $X2=1.66 $Y2=1.202
cc_83 VPB N_A1_c_354_n 0.0256643f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_84 VPB N_A1_c_363_n 0.0156258f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_85 VPB N_A1_c_364_n 0.01623f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_86 VPB N_A1_c_365_n 0.0200169f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_87 VPB N_A1_c_366_n 0.0123873f $X=-0.19 $Y=1.305 $X2=1.055 $Y2=1.105
cc_88 VPB N_A1_c_367_n 0.00160641f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_89 VPB N_A1_c_360_n 0.00272944f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_90 VPB N_A1_c_361_n 0.0392633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A2_c_474_n 0.0159964f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_92 VPB N_A2_c_475_n 0.0158907f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_93 VPB N_A2_c_476_n 0.0158911f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=0.995
cc_94 VPB N_A2_c_477_n 0.01598f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_95 VPB N_A2_c_473_n 0.0449843f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_96 VPB N_VPWR_c_550_n 0.011928f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_97 VPB N_VPWR_c_551_n 0.00714573f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_98 VPB N_VPWR_c_552_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.16
cc_99 VPB N_VPWR_c_553_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_100 VPB N_VPWR_c_554_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.66 $Y2=1.16
cc_101 VPB N_VPWR_c_555_n 0.00514458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_556_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.66 $Y2=1.175
cc_103 VPB N_VPWR_c_557_n 0.012566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_558_n 0.010808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_559_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_560_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_561_n 0.0611151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_562_n 0.00477752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_563_n 0.0608235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_564_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_565_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_566_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_567_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_568_n 0.0229095f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_549_n 0.0476287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_Y_c_681_n 0.00202374f $X=-0.19 $Y=1.305 $X2=1.66 $Y2=1.16
cc_117 VPB N_Y_c_680_n 0.0043829f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_118 VPB N_Y_c_683_n 0.0170593f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.19
cc_119 VPB N_Y_c_684_n 0.00192677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_Y_c_685_n 0.00378296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_1369_297#_c_831_n 0.00231366f $X=-0.19 $Y=1.305 $X2=0.49
+ $Y2=1.202
cc_122 N_C1_c_128_n N_VPWR_c_551_n 0.00479105f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_123 N_C1_c_126_n N_VPWR_c_551_n 0.0161005f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_124 N_C1_c_127_n N_VPWR_c_551_n 0.00177943f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_125 N_C1_c_128_n N_VPWR_c_552_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_126 N_C1_c_129_n N_VPWR_c_552_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_127 N_C1_c_129_n N_VPWR_c_553_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_128 N_C1_c_130_n N_VPWR_c_553_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_129 N_C1_c_130_n N_VPWR_c_567_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_130 N_C1_c_131_n N_VPWR_c_567_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_131 N_C1_c_131_n N_VPWR_c_568_n 0.00514457f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_132 N_C1_c_128_n N_VPWR_c_549_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_133 N_C1_c_129_n N_VPWR_c_549_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_134 N_C1_c_130_n N_VPWR_c_549_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_135 N_C1_c_131_n N_VPWR_c_549_n 0.00821445f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_136 N_C1_c_122_n N_Y_c_679_n 0.00543615f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_137 N_C1_c_123_n N_Y_c_679_n 0.0103107f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_138 N_C1_c_124_n N_Y_c_679_n 0.0103107f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_139 N_C1_c_125_n N_Y_c_679_n 0.0131153f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_140 N_C1_c_126_n N_Y_c_679_n 0.0719449f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_141 N_C1_c_127_n N_Y_c_679_n 0.0101574f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_142 N_C1_c_128_n N_Y_c_681_n 0.00130685f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_143 N_C1_c_126_n N_Y_c_681_n 0.020385f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_144 N_C1_c_127_n N_Y_c_681_n 0.00664519f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_145 N_C1_c_131_n N_Y_c_680_n 0.00132273f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_146 N_C1_c_125_n N_Y_c_680_n 0.0201428f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_147 N_C1_c_126_n N_Y_c_680_n 0.0131966f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_148 N_C1_c_129_n N_Y_c_684_n 0.015669f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_149 N_C1_c_130_n N_Y_c_684_n 0.0157513f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_150 N_C1_c_126_n N_Y_c_684_n 0.0747653f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_151 N_C1_c_127_n N_Y_c_684_n 0.0156153f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_152 N_C1_c_131_n N_Y_c_685_n 0.0283716f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_153 N_C1_c_127_n N_Y_c_685_n 7.03448e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_154 N_C1_c_122_n N_A_27_47#_c_874_n 0.00489172f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_155 N_C1_c_126_n N_A_27_47#_c_874_n 0.0200862f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_156 N_C1_c_127_n N_A_27_47#_c_874_n 9.92702e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_157 N_C1_c_122_n N_A_27_47#_c_875_n 0.0102623f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_158 N_C1_c_123_n N_A_27_47#_c_875_n 0.00931157f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_159 N_C1_c_124_n N_A_27_47#_c_875_n 0.00931157f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_160 N_C1_c_125_n N_A_27_47#_c_875_n 0.00931157f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_161 N_C1_c_126_n N_A_27_47#_c_875_n 0.00355623f $X=1.66 $Y=1.16 $X2=0 $Y2=0
cc_162 N_C1_c_127_n N_A_27_47#_c_875_n 0.00167844f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_163 N_C1_c_125_n N_A_511_47#_c_925_n 7.32022e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_164 N_C1_c_122_n N_VGND_c_1051_n 0.00357877f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_165 N_C1_c_123_n N_VGND_c_1051_n 0.00357877f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_166 N_C1_c_124_n N_VGND_c_1051_n 0.00357877f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_167 N_C1_c_125_n N_VGND_c_1051_n 0.00357877f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_168 N_C1_c_122_n N_VGND_c_1060_n 0.00637194f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_169 N_C1_c_123_n N_VGND_c_1060_n 0.00548399f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_170 N_C1_c_124_n N_VGND_c_1060_n 0.00548399f $X=1.48 $Y=0.995 $X2=0 $Y2=0
cc_171 N_C1_c_125_n N_VGND_c_1060_n 0.00668309f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_c_185_n N_B2_c_282_n 0.0251408f $X=3.88 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_173 N_B1_c_193_n N_B2_c_288_n 0.0221596f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B1_c_195_n N_B2_c_288_n 2.00551e-19 $X=4.83 $Y=1.445 $X2=0 $Y2=0
cc_175 N_B1_c_195_n N_B2_c_289_n 0.00105606f $X=4.83 $Y=1.445 $X2=0 $Y2=0
cc_176 N_B1_c_203_p N_B2_c_289_n 0.00751689f $X=4.925 $Y=1.53 $X2=0 $Y2=0
cc_177 N_B1_c_195_n N_B2_c_290_n 6.599e-19 $X=4.83 $Y=1.445 $X2=0 $Y2=0
cc_178 N_B1_c_196_n N_B2_c_290_n 0.011867f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_179 N_B1_c_186_n N_B2_c_291_n 0.0406946f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B1_c_196_n N_B2_c_291_n 0.0112841f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_181 N_B1_c_189_n N_B2_c_291_n 0.00101445f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_182 N_B1_c_187_n N_B2_c_285_n 0.0216072f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B1_c_186_n N_B2_c_286_n 7.90451e-19 $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B1_c_196_n N_B2_c_286_n 0.0535758f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_185 N_B1_c_188_n N_B2_c_286_n 0.0168455f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_186 N_B1_c_189_n N_B2_c_286_n 0.0161629f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_187 N_B1_c_186_n N_B2_c_287_n 0.0251091f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B1_c_195_n N_B2_c_287_n 0.0107982f $X=4.83 $Y=1.445 $X2=0 $Y2=0
cc_189 N_B1_c_196_n N_B2_c_287_n 0.0149524f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_190 N_B1_c_188_n N_B2_c_287_n 0.0356609f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_191 N_B1_c_189_n N_B2_c_287_n 0.00395727f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_192 N_B1_c_190_n N_B2_c_287_n 0.0251408f $X=3.855 $Y=1.202 $X2=0 $Y2=0
cc_193 N_B1_c_186_n N_A1_c_354_n 0.0537779f $X=6.205 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_194 N_B1_c_189_n N_A1_c_354_n 0.00168165f $X=6.18 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_195 N_B1_c_187_n N_A1_c_355_n 0.0157982f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_196 N_B1_c_186_n N_A1_c_360_n 0.00168165f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B1_c_189_n N_A1_c_360_n 0.0455154f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B1_c_189_n N_VPWR_M1034_d 0.00156777f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_199 N_B1_c_192_n N_VPWR_c_554_n 0.00300743f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B1_c_193_n N_VPWR_c_554_n 0.00300743f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B1_c_186_n N_VPWR_c_555_n 0.00598445f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B1_c_191_n N_VPWR_c_559_n 0.00702461f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_c_192_n N_VPWR_c_559_n 0.00702461f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B1_c_193_n N_VPWR_c_561_n 0.00702461f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B1_c_186_n N_VPWR_c_561_n 0.00513303f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B1_c_191_n N_VPWR_c_568_n 0.00514457f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B1_c_191_n N_VPWR_c_549_n 0.0136891f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B1_c_192_n N_VPWR_c_549_n 0.00693457f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_193_n N_VPWR_c_549_n 0.00695979f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B1_c_186_n N_VPWR_c_549_n 0.00701287f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B1_c_196_n N_Y_M1025_s 0.00187547f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_212 N_B1_c_191_n N_Y_c_680_n 8.72032e-19 $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B1_c_183_n N_Y_c_680_n 0.00283838f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B1_c_188_n N_Y_c_680_n 0.0134954f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_215 N_B1_c_190_n N_Y_c_680_n 0.00722527f $X=3.855 $Y=1.202 $X2=0 $Y2=0
cc_216 N_B1_c_191_n N_Y_c_683_n 0.0194073f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B1_c_192_n N_Y_c_683_n 0.01191f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B1_c_193_n N_Y_c_683_n 0.011867f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B1_c_203_p N_Y_c_683_n 0.0149286f $X=4.925 $Y=1.53 $X2=0 $Y2=0
cc_220 N_B1_c_188_n N_Y_c_683_n 0.145921f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_221 N_B1_c_190_n N_Y_c_683_n 0.0168148f $X=3.855 $Y=1.202 $X2=0 $Y2=0
cc_222 N_B1_c_193_n N_Y_c_715_n 8.1738e-19 $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B1_c_191_n N_Y_c_685_n 0.0100311f $X=2.915 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B1_c_186_n N_Y_c_717_n 0.0166626f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B1_c_196_n N_Y_c_717_n 0.0607449f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_226 N_B1_c_203_p N_Y_c_717_n 0.0113744f $X=4.925 $Y=1.53 $X2=0 $Y2=0
cc_227 N_B1_c_188_n N_Y_c_717_n 0.00418222f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_228 N_B1_c_189_n N_Y_c_717_n 0.0205262f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_229 N_B1_c_196_n N_A_601_297#_M1010_d 0.00187547f $X=6.015 $Y=1.53 $X2=0
+ $Y2=0
cc_230 N_B1_c_196_n N_A_601_297#_M1030_d 0.00172342f $X=6.015 $Y=1.53 $X2=0
+ $Y2=0
cc_231 N_B1_c_189_n N_A_601_297#_M1030_d 7.76441e-19 $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_232 N_B1_c_192_n N_A_601_297#_c_797_n 0.011229f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B1_c_193_n N_A_601_297#_c_797_n 0.011272f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_234 N_B1_c_186_n N_A_601_297#_c_799_n 0.0028452f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_235 N_B1_c_183_n N_A_27_47#_c_875_n 0.0116561f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B1_c_184_n N_A_27_47#_c_875_n 0.00931157f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B1_c_185_n N_A_27_47#_c_875_n 0.00931157f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B1_c_183_n N_A_511_47#_c_925_n 0.00929111f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B1_c_184_n N_A_511_47#_c_925_n 0.00929111f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B1_c_185_n N_A_511_47#_c_925_n 0.00894065f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B1_c_196_n N_A_511_47#_c_925_n 0.00926609f $X=6.015 $Y=1.53 $X2=0 $Y2=0
cc_242 N_B1_c_188_n N_A_511_47#_c_925_n 0.10875f $X=4.735 $Y=1.175 $X2=0 $Y2=0
cc_243 N_B1_c_190_n N_A_511_47#_c_925_n 0.00871767f $X=3.855 $Y=1.202 $X2=0
+ $Y2=0
cc_244 N_B1_c_186_n N_A_511_47#_c_926_n 0.0044163f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B1_c_187_n N_A_511_47#_c_926_n 0.0159827f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B1_c_189_n N_A_511_47#_c_926_n 0.0302712f $X=6.18 $Y=1.16 $X2=0 $Y2=0
cc_247 N_B1_c_183_n N_VGND_c_1051_n 0.00357877f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_c_184_n N_VGND_c_1051_n 0.00357877f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B1_c_185_n N_VGND_c_1051_n 0.00357877f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_187_n N_VGND_c_1051_n 0.00426565f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_183_n N_VGND_c_1060_n 0.00672921f $X=2.94 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_184_n N_VGND_c_1060_n 0.00548399f $X=3.41 $Y=0.995 $X2=0 $Y2=0
cc_253 N_B1_c_185_n N_VGND_c_1060_n 0.00538422f $X=3.88 $Y=0.995 $X2=0 $Y2=0
cc_254 N_B1_c_187_n N_VGND_c_1060_n 0.00632911f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_255 N_B2_c_288_n N_VPWR_c_561_n 0.00429453f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B2_c_289_n N_VPWR_c_561_n 0.00429453f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B2_c_290_n N_VPWR_c_561_n 0.00429453f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B2_c_291_n N_VPWR_c_561_n 0.00429453f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B2_c_288_n N_VPWR_c_549_n 0.00609021f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B2_c_289_n N_VPWR_c_549_n 0.00606499f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B2_c_290_n N_VPWR_c_549_n 0.00606499f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B2_c_291_n N_VPWR_c_549_n 0.00609021f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B2_c_288_n N_Y_c_683_n 0.0117685f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B2_c_289_n N_Y_c_683_n 0.00119625f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B2_c_287_n N_Y_c_683_n 0.00423254f $X=5.735 $Y=1.202 $X2=0 $Y2=0
cc_266 N_B2_c_288_n N_Y_c_715_n 0.00877192f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B2_c_289_n N_Y_c_715_n 0.00361268f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B2_c_289_n N_Y_c_717_n 0.012227f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B2_c_290_n N_Y_c_717_n 0.011914f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B2_c_291_n N_Y_c_717_n 0.0118581f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B2_c_287_n N_Y_c_717_n 0.00275505f $X=5.735 $Y=1.202 $X2=0 $Y2=0
cc_272 N_B2_c_288_n N_A_601_297#_c_799_n 0.0116484f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B2_c_289_n N_A_601_297#_c_799_n 0.0103969f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B2_c_290_n N_A_601_297#_c_799_n 0.0104142f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B2_c_291_n N_A_601_297#_c_799_n 0.0104142f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B2_c_282_n N_A_27_47#_c_875_n 0.00931157f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_277 N_B2_c_283_n N_A_27_47#_c_875_n 0.00931157f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_278 N_B2_c_284_n N_A_27_47#_c_875_n 0.00964761f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_279 N_B2_c_285_n N_A_27_47#_c_875_n 0.00964761f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_280 N_B2_c_282_n N_A_511_47#_c_925_n 0.00894065f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B2_c_283_n N_A_511_47#_c_925_n 0.00928704f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B2_c_284_n N_A_511_47#_c_925_n 0.00882716f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B2_c_285_n N_A_511_47#_c_925_n 0.00877034f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B2_c_286_n N_A_511_47#_c_925_n 0.0459672f $X=5.65 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B2_c_287_n N_A_511_47#_c_925_n 0.0112676f $X=5.735 $Y=1.202 $X2=0 $Y2=0
cc_286 N_B2_c_285_n N_A_511_47#_c_926_n 0.00232072f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_287 N_B2_c_282_n N_VGND_c_1051_n 0.00357877f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_288 N_B2_c_283_n N_VGND_c_1051_n 0.00357877f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_289 N_B2_c_284_n N_VGND_c_1051_n 0.00357877f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_290 N_B2_c_285_n N_VGND_c_1051_n 0.00357877f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_291 N_B2_c_282_n N_VGND_c_1060_n 0.00538422f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_292 N_B2_c_283_n N_VGND_c_1060_n 0.00548399f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_293 N_B2_c_284_n N_VGND_c_1060_n 0.00560377f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_294 N_B2_c_285_n N_VGND_c_1060_n 0.00562222f $X=5.76 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A1_c_355_n N_A2_c_468_n 0.0258949f $X=6.78 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_296 N_A1_c_354_n N_A2_c_474_n 0.0406946f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A1_c_366_n N_A2_c_474_n 0.0112841f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_298 N_A1_c_360_n N_A2_c_474_n 0.00101445f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A1_c_366_n N_A2_c_475_n 0.011867f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_300 N_A1_c_366_n N_A2_c_476_n 0.01191f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_301 N_A1_c_363_n N_A2_c_477_n 0.0226278f $X=9.105 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A1_c_366_n N_A2_c_477_n 0.0142273f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_303 N_A1_c_367_n N_A2_c_477_n 7.03078e-19 $X=9.162 $Y=1.445 $X2=0 $Y2=0
cc_304 N_A1_c_356_n N_A2_c_471_n 0.0239161f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A1_c_354_n N_A2_c_472_n 2.32333e-19 $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_306 N_A1_c_366_n N_A2_c_472_n 0.113835f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_307 N_A1_c_359_n N_A2_c_472_n 0.0115402f $X=9.162 $Y=1.275 $X2=0 $Y2=0
cc_308 N_A1_c_360_n N_A2_c_472_n 0.0160817f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_309 N_A1_c_361_n N_A2_c_472_n 2.49913e-19 $X=10.02 $Y=1.202 $X2=0 $Y2=0
cc_310 N_A1_c_354_n N_A2_c_473_n 0.0263635f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A1_c_366_n N_A2_c_473_n 0.0231495f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_312 N_A1_c_359_n N_A2_c_473_n 2.49913e-19 $X=9.162 $Y=1.275 $X2=0 $Y2=0
cc_313 N_A1_c_367_n N_A2_c_473_n 9.22604e-19 $X=9.162 $Y=1.445 $X2=0 $Y2=0
cc_314 N_A1_c_360_n N_A2_c_473_n 0.00395386f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_315 N_A1_c_361_n N_A2_c_473_n 0.0239161f $X=10.02 $Y=1.202 $X2=0 $Y2=0
cc_316 N_A1_c_360_n N_VPWR_M1034_d 0.00156777f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A1_c_366_n N_VPWR_M1022_s 0.00230525f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_318 N_A1_c_354_n N_VPWR_c_555_n 0.00582761f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A1_c_363_n N_VPWR_c_556_n 0.00300743f $X=9.105 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A1_c_364_n N_VPWR_c_556_n 0.00300743f $X=9.575 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A1_c_365_n N_VPWR_c_558_n 0.00578236f $X=10.045 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A1_c_361_n N_VPWR_c_558_n 0.00103985f $X=10.02 $Y=1.202 $X2=0 $Y2=0
cc_323 N_A1_c_354_n N_VPWR_c_563_n 0.004871f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A1_c_363_n N_VPWR_c_563_n 0.00702461f $X=9.105 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A1_c_364_n N_VPWR_c_565_n 0.00702461f $X=9.575 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A1_c_365_n N_VPWR_c_565_n 0.00702461f $X=10.045 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A1_c_354_n N_VPWR_c_549_n 0.00674306f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A1_c_363_n N_VPWR_c_549_n 0.00695979f $X=9.105 $Y=1.41 $X2=0 $Y2=0
cc_329 N_A1_c_364_n N_VPWR_c_549_n 0.00693457f $X=9.575 $Y=1.41 $X2=0 $Y2=0
cc_330 N_A1_c_365_n N_VPWR_c_549_n 0.0133558f $X=10.045 $Y=1.41 $X2=0 $Y2=0
cc_331 N_A1_c_366_n N_Y_M1002_d 0.00187547f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_332 N_A1_c_366_n N_Y_M1015_d 0.00187547f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_333 N_A1_c_354_n N_Y_c_717_n 0.0162681f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_334 N_A1_c_366_n N_Y_c_717_n 0.0875398f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_335 N_A1_c_360_n N_Y_c_717_n 0.0205262f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A1_c_366_n N_A_1369_297#_M1003_d 0.00172342f $X=9.005 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_337 N_A1_c_360_n N_A_1369_297#_M1003_d 7.76441e-19 $X=6.73 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_338 N_A1_c_366_n N_A_1369_297#_M1005_s 0.00187547f $X=9.005 $Y=1.53 $X2=0
+ $Y2=0
cc_339 N_A1_c_366_n N_A_1369_297#_M1038_s 0.00183902f $X=9.005 $Y=1.53 $X2=0
+ $Y2=0
cc_340 N_A1_c_354_n N_A_1369_297#_c_836_n 0.00458775f $X=6.755 $Y=1.41 $X2=0
+ $Y2=0
cc_341 N_A1_c_366_n N_A_1369_297#_c_836_n 0.00362004f $X=9.005 $Y=1.53 $X2=0
+ $Y2=0
cc_342 N_A1_c_363_n N_A_1369_297#_c_838_n 0.0112647f $X=9.105 $Y=1.41 $X2=0
+ $Y2=0
cc_343 N_A1_c_364_n N_A_1369_297#_c_838_n 0.0132594f $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_344 N_A1_c_366_n N_A_1369_297#_c_838_n 0.0188459f $X=9.005 $Y=1.53 $X2=0
+ $Y2=0
cc_345 N_A1_c_425_p N_A_1369_297#_c_838_n 0.00936841f $X=9.95 $Y=1.16 $X2=0
+ $Y2=0
cc_346 N_A1_c_361_n N_A_1369_297#_c_838_n 0.00332181f $X=10.02 $Y=1.202 $X2=0
+ $Y2=0
cc_347 N_A1_c_366_n N_A_1369_297#_c_843_n 0.014075f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_348 N_A1_c_364_n N_A_1369_297#_c_831_n 4.44016e-19 $X=9.575 $Y=1.41 $X2=0
+ $Y2=0
cc_349 N_A1_c_365_n N_A_1369_297#_c_831_n 3.55815e-19 $X=10.045 $Y=1.41 $X2=0
+ $Y2=0
cc_350 N_A1_c_366_n N_A_1369_297#_c_831_n 0.00532569f $X=9.005 $Y=1.53 $X2=0
+ $Y2=0
cc_351 N_A1_c_425_p N_A_1369_297#_c_831_n 0.0202219f $X=9.95 $Y=1.16 $X2=0 $Y2=0
cc_352 N_A1_c_361_n N_A_1369_297#_c_831_n 0.00658737f $X=10.02 $Y=1.202 $X2=0
+ $Y2=0
cc_353 N_A1_c_354_n N_A_511_47#_c_920_n 0.001478f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A1_c_355_n N_A_511_47#_c_920_n 0.0103956f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_355 N_A1_c_366_n N_A_511_47#_c_920_n 0.00608471f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_356 N_A1_c_355_n N_A_511_47#_c_950_n 5.34052e-19 $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_357 N_A1_c_356_n N_A_511_47#_c_922_n 0.00845282f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_358 N_A1_c_366_n N_A_511_47#_c_922_n 0.00911016f $X=9.005 $Y=1.53 $X2=0 $Y2=0
cc_359 N_A1_c_359_n N_A_511_47#_c_922_n 0.00893273f $X=9.162 $Y=1.275 $X2=0
+ $Y2=0
cc_360 N_A1_c_356_n N_A_511_47#_c_954_n 0.00644736f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A1_c_357_n N_A_511_47#_c_954_n 0.00686626f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A1_c_358_n N_A_511_47#_c_954_n 5.45498e-19 $X=10.02 $Y=0.995 $X2=0
+ $Y2=0
cc_363 N_A1_c_357_n N_A_511_47#_c_923_n 0.00901745f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A1_c_358_n N_A_511_47#_c_923_n 0.0103267f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A1_c_425_p N_A_511_47#_c_923_n 0.0452977f $X=9.95 $Y=1.16 $X2=0 $Y2=0
cc_366 N_A1_c_361_n N_A_511_47#_c_923_n 0.00674339f $X=10.02 $Y=1.202 $X2=0
+ $Y2=0
cc_367 N_A1_c_357_n N_A_511_47#_c_924_n 5.24597e-19 $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A1_c_358_n N_A_511_47#_c_924_n 0.00651696f $X=10.02 $Y=0.995 $X2=0
+ $Y2=0
cc_369 N_A1_c_354_n N_A_511_47#_c_926_n 0.00291462f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_370 N_A1_c_360_n N_A_511_47#_c_926_n 0.0296144f $X=6.73 $Y=1.16 $X2=0 $Y2=0
cc_371 N_A1_c_356_n N_A_511_47#_c_929_n 0.00132031f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_372 N_A1_c_357_n N_A_511_47#_c_929_n 0.00116636f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A1_c_359_n N_A_511_47#_c_929_n 0.0169059f $X=9.162 $Y=1.275 $X2=0 $Y2=0
cc_374 N_A1_c_425_p N_A_511_47#_c_929_n 0.0148598f $X=9.95 $Y=1.16 $X2=0 $Y2=0
cc_375 N_A1_c_361_n N_A_511_47#_c_929_n 0.00358162f $X=10.02 $Y=1.202 $X2=0
+ $Y2=0
cc_376 N_A1_c_355_n N_VGND_c_1047_n 0.00268723f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_377 N_A1_c_356_n N_VGND_c_1049_n 0.00268723f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_378 N_A1_c_357_n N_VGND_c_1050_n 0.00379224f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_379 N_A1_c_358_n N_VGND_c_1050_n 0.00276126f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_380 N_A1_c_355_n N_VGND_c_1051_n 0.00439206f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_381 N_A1_c_356_n N_VGND_c_1057_n 0.00424416f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_382 N_A1_c_357_n N_VGND_c_1057_n 0.00423334f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_383 N_A1_c_358_n N_VGND_c_1059_n 0.00423334f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_384 N_A1_c_355_n N_VGND_c_1060_n 0.00625209f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_385 N_A1_c_356_n N_VGND_c_1060_n 0.00589024f $X=9.08 $Y=0.995 $X2=0 $Y2=0
cc_386 N_A1_c_357_n N_VGND_c_1060_n 0.006093f $X=9.55 $Y=0.995 $X2=0 $Y2=0
cc_387 N_A1_c_358_n N_VGND_c_1060_n 0.0068733f $X=10.02 $Y=0.995 $X2=0 $Y2=0
cc_388 N_A2_c_474_n N_VPWR_c_563_n 0.00429453f $X=7.225 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A2_c_475_n N_VPWR_c_563_n 0.00429453f $X=7.695 $Y=1.41 $X2=0 $Y2=0
cc_390 N_A2_c_476_n N_VPWR_c_563_n 0.00429453f $X=8.165 $Y=1.41 $X2=0 $Y2=0
cc_391 N_A2_c_477_n N_VPWR_c_563_n 0.00429453f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_392 N_A2_c_474_n N_VPWR_c_549_n 0.00609021f $X=7.225 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A2_c_475_n N_VPWR_c_549_n 0.00606499f $X=7.695 $Y=1.41 $X2=0 $Y2=0
cc_394 N_A2_c_476_n N_VPWR_c_549_n 0.00606499f $X=8.165 $Y=1.41 $X2=0 $Y2=0
cc_395 N_A2_c_477_n N_VPWR_c_549_n 0.00609021f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_396 N_A2_c_474_n N_Y_c_717_n 0.0118581f $X=7.225 $Y=1.41 $X2=0 $Y2=0
cc_397 N_A2_c_475_n N_Y_c_717_n 0.011914f $X=7.695 $Y=1.41 $X2=0 $Y2=0
cc_398 N_A2_c_476_n N_Y_c_717_n 0.011914f $X=8.165 $Y=1.41 $X2=0 $Y2=0
cc_399 N_A2_c_477_n N_Y_c_717_n 0.00313253f $X=8.635 $Y=1.41 $X2=0 $Y2=0
cc_400 N_A2_c_474_n N_A_1369_297#_c_836_n 0.0104142f $X=7.225 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A2_c_475_n N_A_1369_297#_c_836_n 0.0104142f $X=7.695 $Y=1.41 $X2=0
+ $Y2=0
cc_402 N_A2_c_476_n N_A_1369_297#_c_836_n 0.0104142f $X=8.165 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_A2_c_477_n N_A_1369_297#_c_836_n 0.0122183f $X=8.635 $Y=1.41 $X2=0
+ $Y2=0
cc_404 N_A2_c_468_n N_A_511_47#_c_920_n 0.00845772f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A2_c_472_n N_A_511_47#_c_920_n 0.00820272f $X=8.46 $Y=1.16 $X2=0 $Y2=0
cc_406 N_A2_c_468_n N_A_511_47#_c_950_n 0.00643055f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A2_c_469_n N_A_511_47#_c_950_n 0.00686626f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A2_c_470_n N_A_511_47#_c_950_n 5.45498e-19 $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A2_c_469_n N_A_511_47#_c_921_n 0.00901745f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A2_c_470_n N_A_511_47#_c_921_n 0.00901745f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A2_c_472_n N_A_511_47#_c_921_n 0.0397461f $X=8.46 $Y=1.16 $X2=0 $Y2=0
cc_412 N_A2_c_473_n N_A_511_47#_c_921_n 0.00345541f $X=8.635 $Y=1.202 $X2=0
+ $Y2=0
cc_413 N_A2_c_469_n N_A_511_47#_c_979_n 5.24597e-19 $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_414 N_A2_c_470_n N_A_511_47#_c_979_n 0.00651696f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_415 N_A2_c_471_n N_A_511_47#_c_922_n 0.0103942f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_416 N_A2_c_472_n N_A_511_47#_c_922_n 0.0117061f $X=8.46 $Y=1.16 $X2=0 $Y2=0
cc_417 N_A2_c_471_n N_A_511_47#_c_954_n 5.32212e-19 $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_418 N_A2_c_468_n N_A_511_47#_c_927_n 0.00132158f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_419 N_A2_c_469_n N_A_511_47#_c_927_n 0.00116636f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_420 N_A2_c_472_n N_A_511_47#_c_927_n 0.0306016f $X=8.46 $Y=1.16 $X2=0 $Y2=0
cc_421 N_A2_c_473_n N_A_511_47#_c_927_n 0.00358305f $X=8.635 $Y=1.202 $X2=0
+ $Y2=0
cc_422 N_A2_c_470_n N_A_511_47#_c_928_n 0.00119564f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_423 N_A2_c_472_n N_A_511_47#_c_928_n 0.0307352f $X=8.46 $Y=1.16 $X2=0 $Y2=0
cc_424 N_A2_c_473_n N_A_511_47#_c_928_n 0.00486271f $X=8.635 $Y=1.202 $X2=0
+ $Y2=0
cc_425 N_A2_c_468_n N_VGND_c_1047_n 0.00268723f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A2_c_469_n N_VGND_c_1048_n 0.00379224f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A2_c_470_n N_VGND_c_1048_n 0.00276126f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A2_c_471_n N_VGND_c_1049_n 0.00268723f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A2_c_468_n N_VGND_c_1053_n 0.00424416f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_430 N_A2_c_469_n N_VGND_c_1053_n 0.00423334f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A2_c_470_n N_VGND_c_1055_n 0.00423334f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_432 N_A2_c_471_n N_VGND_c_1055_n 0.00439206f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A2_c_468_n N_VGND_c_1060_n 0.00589024f $X=7.2 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A2_c_469_n N_VGND_c_1060_n 0.006093f $X=7.67 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A2_c_470_n N_VGND_c_1060_n 0.00608558f $X=8.14 $Y=0.995 $X2=0 $Y2=0
cc_436 N_A2_c_471_n N_VGND_c_1060_n 0.00618081f $X=8.66 $Y=0.995 $X2=0 $Y2=0
cc_437 N_VPWR_c_549_n N_Y_M1000_d 0.00370124f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_438 N_VPWR_c_549_n N_Y_M1012_d 0.00307556f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_439 N_VPWR_c_549_n N_Y_M1001_s 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_440 N_VPWR_c_549_n N_Y_M1025_s 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_441 N_VPWR_c_549_n N_Y_M1002_d 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_442 N_VPWR_c_549_n N_Y_M1015_d 0.00232895f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_443 N_VPWR_c_552_n N_Y_c_746_n 0.0149311f $X=1.095 $Y=2.72 $X2=0 $Y2=0
cc_444 N_VPWR_c_549_n N_Y_c_746_n 0.00955092f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_c_567_n N_Y_c_748_n 0.014675f $X=2.035 $Y=2.465 $X2=0 $Y2=0
cc_446 N_VPWR_c_549_n N_Y_c_748_n 0.00948039f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_447 N_VPWR_M1024_s N_Y_c_683_n 0.0103462f $X=2.015 $Y=1.485 $X2=0 $Y2=0
cc_448 N_VPWR_M1018_d N_Y_c_683_n 0.00187547f $X=3.475 $Y=1.485 $X2=0 $Y2=0
cc_449 N_VPWR_c_568_n N_Y_c_683_n 0.0158748f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_450 N_VPWR_M1008_s N_Y_c_684_n 0.00205023f $X=1.075 $Y=1.485 $X2=0 $Y2=0
cc_451 N_VPWR_c_553_n N_Y_c_684_n 0.0122355f $X=1.22 $Y=1.99 $X2=0 $Y2=0
cc_452 N_VPWR_M1024_s N_Y_c_685_n 0.0122767f $X=2.015 $Y=1.485 $X2=0 $Y2=0
cc_453 N_VPWR_c_568_n N_Y_c_685_n 0.0214276f $X=2.805 $Y=2.465 $X2=0 $Y2=0
cc_454 N_VPWR_c_549_n N_Y_c_685_n 0.00865749f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_455 N_VPWR_M1034_d N_Y_c_717_n 0.0103467f $X=6.295 $Y=1.485 $X2=0 $Y2=0
cc_456 N_VPWR_c_555_n N_Y_c_717_n 0.0196908f $X=6.48 $Y=2.35 $X2=0 $Y2=0
cc_457 N_VPWR_c_561_n N_Y_c_717_n 0.0027165f $X=6.355 $Y=2.72 $X2=0 $Y2=0
cc_458 N_VPWR_c_563_n N_Y_c_717_n 0.00202091f $X=9.215 $Y=2.72 $X2=0 $Y2=0
cc_459 N_VPWR_c_549_n N_Y_c_717_n 0.0184019f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_549_n N_A_601_297#_M1013_s 0.0031047f $X=10.35 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_461 N_VPWR_c_549_n N_A_601_297#_M1028_s 0.00241848f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_549_n N_A_601_297#_M1010_d 0.00231289f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_549_n N_A_601_297#_M1030_d 0.00231289f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_559_n N_A_601_297#_c_808_n 0.0149311f $X=3.495 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_549_n N_A_601_297#_c_808_n 0.00955092f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_466 N_VPWR_M1018_d N_A_601_297#_c_797_n 0.00347905f $X=3.475 $Y=1.485 $X2=0
+ $Y2=0
cc_467 N_VPWR_c_554_n N_A_601_297#_c_797_n 0.0139109f $X=3.62 $Y=2.3 $X2=0 $Y2=0
cc_468 N_VPWR_c_549_n N_A_601_297#_c_797_n 0.0141598f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_561_n N_A_601_297#_c_813_n 0.0134783f $X=6.355 $Y=2.72 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_549_n N_A_601_297#_c_813_n 0.00808747f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_555_n N_A_601_297#_c_799_n 0.0130957f $X=6.48 $Y=2.35 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_561_n N_A_601_297#_c_799_n 0.109166f $X=6.355 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_c_549_n N_A_601_297#_c_799_n 0.0695192f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_549_n N_A_1369_297#_M1003_d 0.00231289f $X=10.35 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_475 N_VPWR_c_549_n N_A_1369_297#_M1005_s 0.00231289f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_549_n N_A_1369_297#_M1038_s 0.00241848f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_549_n N_A_1369_297#_M1026_d 0.0031047f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_478 N_VPWR_c_555_n N_A_1369_297#_c_836_n 0.0159918f $X=6.48 $Y=2.35 $X2=0
+ $Y2=0
cc_479 N_VPWR_c_563_n N_A_1369_297#_c_836_n 0.125753f $X=9.215 $Y=2.72 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_549_n N_A_1369_297#_c_836_n 0.0792478f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_481 N_VPWR_M1022_s N_A_1369_297#_c_838_n 0.00409206f $X=9.195 $Y=1.485 $X2=0
+ $Y2=0
cc_482 N_VPWR_c_556_n N_A_1369_297#_c_838_n 0.0139109f $X=9.34 $Y=2.3 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_549_n N_A_1369_297#_c_838_n 0.0141598f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_484 N_VPWR_c_558_n N_A_1369_297#_c_831_n 0.00259649f $X=10.28 $Y=1.62 $X2=0
+ $Y2=0
cc_485 N_VPWR_c_565_n N_A_1369_297#_c_864_n 0.0149311f $X=10.155 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_549_n N_A_1369_297#_c_864_n 0.00955092f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_558_n N_A_511_47#_c_923_n 0.0103208f $X=10.28 $Y=1.62 $X2=0
+ $Y2=0
cc_488 N_Y_c_683_n N_A_601_297#_M1013_s 0.00187091f $X=4.345 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_489 N_Y_c_683_n N_A_601_297#_M1028_s 0.00183902f $X=4.345 $Y=1.53 $X2=0 $Y2=0
cc_490 N_Y_c_717_n N_A_601_297#_M1010_d 0.00387132f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_491 N_Y_c_717_n N_A_601_297#_M1030_d 0.00406208f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_492 N_Y_c_683_n N_A_601_297#_c_797_n 0.0511916f $X=4.345 $Y=1.53 $X2=0 $Y2=0
cc_493 N_Y_c_715_n N_A_601_297#_c_797_n 0.0148585f $X=4.455 $Y=1.785 $X2=0 $Y2=0
cc_494 N_Y_c_683_n N_A_601_297#_c_824_n 0.0143191f $X=4.345 $Y=1.53 $X2=0 $Y2=0
cc_495 N_Y_c_715_n N_A_601_297#_c_825_n 0.00395094f $X=4.455 $Y=1.785 $X2=0
+ $Y2=0
cc_496 N_Y_M1001_s N_A_601_297#_c_799_n 0.00394064f $X=4.415 $Y=1.485 $X2=0
+ $Y2=0
cc_497 N_Y_M1025_s N_A_601_297#_c_799_n 0.00394288f $X=5.355 $Y=1.485 $X2=0
+ $Y2=0
cc_498 N_Y_c_683_n N_A_601_297#_c_799_n 0.00248657f $X=4.345 $Y=1.53 $X2=0 $Y2=0
cc_499 N_Y_c_715_n N_A_601_297#_c_799_n 0.0083207f $X=4.455 $Y=1.785 $X2=0 $Y2=0
cc_500 N_Y_c_717_n N_A_601_297#_c_799_n 0.0554154f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_501 N_Y_c_717_n N_A_1369_297#_M1003_d 0.00406208f $X=8.4 $Y=1.92 $X2=-0.19
+ $Y2=-0.24
cc_502 N_Y_c_717_n N_A_1369_297#_M1005_s 0.00387132f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_503 N_Y_M1002_d N_A_1369_297#_c_836_n 0.00394288f $X=7.315 $Y=1.485 $X2=0
+ $Y2=0
cc_504 N_Y_M1015_d N_A_1369_297#_c_836_n 0.00394288f $X=8.255 $Y=1.485 $X2=0
+ $Y2=0
cc_505 N_Y_c_717_n N_A_1369_297#_c_836_n 0.0631991f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_506 N_Y_c_717_n N_A_1369_297#_c_871_n 0.00316953f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_507 N_Y_c_717_n N_A_1369_297#_c_843_n 0.0120899f $X=8.4 $Y=1.92 $X2=0 $Y2=0
cc_508 N_Y_c_679_n N_A_27_47#_M1016_s 0.00417498f $X=2.12 $Y=0.755 $X2=0 $Y2=0
cc_509 N_Y_c_679_n N_A_27_47#_M1031_s 0.00379863f $X=2.12 $Y=0.755 $X2=0 $Y2=0
cc_510 N_Y_c_680_n N_A_27_47#_M1031_s 3.00511e-19 $X=2.222 $Y=1.445 $X2=0 $Y2=0
cc_511 N_Y_c_679_n N_A_27_47#_c_874_n 0.0176073f $X=2.12 $Y=0.755 $X2=0 $Y2=0
cc_512 N_Y_M1006_d N_A_27_47#_c_875_n 0.00400389f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_513 N_Y_M1020_d N_A_27_47#_c_875_n 0.00400389f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_514 N_Y_c_679_n N_A_27_47#_c_875_n 0.0985423f $X=2.12 $Y=0.755 $X2=0 $Y2=0
cc_515 N_Y_c_679_n N_A_511_47#_c_925_n 0.0149754f $X=2.12 $Y=0.755 $X2=0 $Y2=0
cc_516 N_Y_c_683_n N_A_511_47#_c_925_n 0.00136402f $X=4.345 $Y=1.53 $X2=0 $Y2=0
cc_517 N_Y_M1006_d N_VGND_c_1060_n 0.00256987f $X=0.615 $Y=0.235 $X2=0 $Y2=0
cc_518 N_Y_M1020_d N_VGND_c_1060_n 0.00256987f $X=1.555 $Y=0.235 $X2=0 $Y2=0
cc_519 N_A_27_47#_c_875_n N_A_511_47#_M1021_s 0.00663816f $X=5.97 $Y=0.39
+ $X2=-0.19 $Y2=-0.24
cc_520 N_A_27_47#_c_875_n N_A_511_47#_M1023_s 0.00400389f $X=5.97 $Y=0.39 $X2=0
+ $Y2=0
cc_521 N_A_27_47#_c_875_n N_A_511_47#_M1007_d 0.00400389f $X=5.97 $Y=0.39 $X2=0
+ $Y2=0
cc_522 N_A_27_47#_c_875_n N_A_511_47#_M1029_d 0.00507817f $X=5.97 $Y=0.39 $X2=0
+ $Y2=0
cc_523 N_A_27_47#_M1021_d N_A_511_47#_c_925_n 0.00434237f $X=3.015 $Y=0.235
+ $X2=0 $Y2=0
cc_524 N_A_27_47#_M1033_d N_A_511_47#_c_925_n 0.0035985f $X=3.955 $Y=0.235 $X2=0
+ $Y2=0
cc_525 N_A_27_47#_M1027_s N_A_511_47#_c_925_n 0.00518226f $X=4.845 $Y=0.235
+ $X2=0 $Y2=0
cc_526 N_A_27_47#_M1039_s N_A_511_47#_c_925_n 0.00373854f $X=5.835 $Y=0.235
+ $X2=0 $Y2=0
cc_527 N_A_27_47#_c_875_n N_A_511_47#_c_925_n 0.191551f $X=5.97 $Y=0.39 $X2=0
+ $Y2=0
cc_528 N_A_27_47#_M1039_s N_A_511_47#_c_926_n 0.00176035f $X=5.835 $Y=0.235
+ $X2=0 $Y2=0
cc_529 N_A_27_47#_c_873_n N_VGND_c_1051_n 0.01753f $X=0.24 $Y=0.475 $X2=0 $Y2=0
cc_530 N_A_27_47#_c_875_n N_VGND_c_1051_n 0.331222f $X=5.97 $Y=0.39 $X2=0 $Y2=0
cc_531 N_A_27_47#_M1006_s N_VGND_c_1060_n 0.00266714f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_532 N_A_27_47#_M1016_s N_VGND_c_1060_n 0.00255381f $X=1.085 $Y=0.235 $X2=0
+ $Y2=0
cc_533 N_A_27_47#_M1031_s N_VGND_c_1060_n 0.00209344f $X=2.025 $Y=0.235 $X2=0
+ $Y2=0
cc_534 N_A_27_47#_M1021_d N_VGND_c_1060_n 0.00255381f $X=3.015 $Y=0.235 $X2=0
+ $Y2=0
cc_535 N_A_27_47#_M1033_d N_VGND_c_1060_n 0.00215227f $X=3.955 $Y=0.235 $X2=0
+ $Y2=0
cc_536 N_A_27_47#_M1027_s N_VGND_c_1060_n 0.00255381f $X=4.845 $Y=0.235 $X2=0
+ $Y2=0
cc_537 N_A_27_47#_M1039_s N_VGND_c_1060_n 0.00262586f $X=5.835 $Y=0.235 $X2=0
+ $Y2=0
cc_538 N_A_27_47#_c_873_n N_VGND_c_1060_n 0.00961275f $X=0.24 $Y=0.475 $X2=0
+ $Y2=0
cc_539 N_A_27_47#_c_875_n N_VGND_c_1060_n 0.207811f $X=5.97 $Y=0.39 $X2=0 $Y2=0
cc_540 N_A_511_47#_c_920_n N_VGND_M1009_d 0.00165819f $X=7.245 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_541 N_A_511_47#_c_921_n N_VGND_M1017_s 0.00251047f $X=8.185 $Y=0.815 $X2=0
+ $Y2=0
cc_542 N_A_511_47#_c_922_n N_VGND_M1036_s 0.00165819f $X=9.125 $Y=0.82 $X2=0
+ $Y2=0
cc_543 N_A_511_47#_c_923_n N_VGND_M1014_d 0.00251047f $X=10.065 $Y=0.815 $X2=0
+ $Y2=0
cc_544 N_A_511_47#_c_920_n N_VGND_c_1047_n 0.0116528f $X=7.245 $Y=0.82 $X2=0
+ $Y2=0
cc_545 N_A_511_47#_c_950_n N_VGND_c_1048_n 0.0183628f $X=7.46 $Y=0.39 $X2=0
+ $Y2=0
cc_546 N_A_511_47#_c_921_n N_VGND_c_1048_n 0.0127273f $X=8.185 $Y=0.815 $X2=0
+ $Y2=0
cc_547 N_A_511_47#_c_922_n N_VGND_c_1049_n 0.0116529f $X=9.125 $Y=0.82 $X2=0
+ $Y2=0
cc_548 N_A_511_47#_c_954_n N_VGND_c_1050_n 0.0183628f $X=9.34 $Y=0.39 $X2=0
+ $Y2=0
cc_549 N_A_511_47#_c_923_n N_VGND_c_1050_n 0.0127273f $X=10.065 $Y=0.815 $X2=0
+ $Y2=0
cc_550 N_A_511_47#_c_1014_p N_VGND_c_1051_n 0.0208133f $X=6.52 $Y=0.39 $X2=0
+ $Y2=0
cc_551 N_A_511_47#_c_920_n N_VGND_c_1051_n 0.00248202f $X=7.245 $Y=0.82 $X2=0
+ $Y2=0
cc_552 N_A_511_47#_c_926_n N_VGND_c_1051_n 0.00315004f $X=6.685 $Y=0.775 $X2=0
+ $Y2=0
cc_553 N_A_511_47#_c_920_n N_VGND_c_1053_n 0.00193763f $X=7.245 $Y=0.82 $X2=0
+ $Y2=0
cc_554 N_A_511_47#_c_950_n N_VGND_c_1053_n 0.0223596f $X=7.46 $Y=0.39 $X2=0
+ $Y2=0
cc_555 N_A_511_47#_c_921_n N_VGND_c_1053_n 0.00266636f $X=8.185 $Y=0.815 $X2=0
+ $Y2=0
cc_556 N_A_511_47#_c_921_n N_VGND_c_1055_n 0.00198695f $X=8.185 $Y=0.815 $X2=0
+ $Y2=0
cc_557 N_A_511_47#_c_979_n N_VGND_c_1055_n 0.0231806f $X=8.4 $Y=0.39 $X2=0 $Y2=0
cc_558 N_A_511_47#_c_922_n N_VGND_c_1055_n 0.00248202f $X=9.125 $Y=0.82 $X2=0
+ $Y2=0
cc_559 N_A_511_47#_c_922_n N_VGND_c_1057_n 0.00193763f $X=9.125 $Y=0.82 $X2=0
+ $Y2=0
cc_560 N_A_511_47#_c_954_n N_VGND_c_1057_n 0.0223596f $X=9.34 $Y=0.39 $X2=0
+ $Y2=0
cc_561 N_A_511_47#_c_923_n N_VGND_c_1057_n 0.00266636f $X=10.065 $Y=0.815 $X2=0
+ $Y2=0
cc_562 N_A_511_47#_c_923_n N_VGND_c_1059_n 0.00198695f $X=10.065 $Y=0.815 $X2=0
+ $Y2=0
cc_563 N_A_511_47#_c_924_n N_VGND_c_1059_n 0.0244796f $X=10.28 $Y=0.39 $X2=0
+ $Y2=0
cc_564 N_A_511_47#_M1021_s N_VGND_c_1060_n 0.00251142f $X=2.555 $Y=0.235 $X2=0
+ $Y2=0
cc_565 N_A_511_47#_M1023_s N_VGND_c_1060_n 0.00256987f $X=3.485 $Y=0.235 $X2=0
+ $Y2=0
cc_566 N_A_511_47#_M1007_d N_VGND_c_1060_n 0.00256987f $X=4.375 $Y=0.235 $X2=0
+ $Y2=0
cc_567 N_A_511_47#_M1029_d N_VGND_c_1060_n 0.00297142f $X=5.315 $Y=0.235 $X2=0
+ $Y2=0
cc_568 N_A_511_47#_M1037_s N_VGND_c_1060_n 0.00348662f $X=6.305 $Y=0.235 $X2=0
+ $Y2=0
cc_569 N_A_511_47#_M1004_d N_VGND_c_1060_n 0.0025535f $X=7.275 $Y=0.235 $X2=0
+ $Y2=0
cc_570 N_A_511_47#_M1019_d N_VGND_c_1060_n 0.00304426f $X=8.215 $Y=0.235 $X2=0
+ $Y2=0
cc_571 N_A_511_47#_M1011_s N_VGND_c_1060_n 0.0025535f $X=9.155 $Y=0.235 $X2=0
+ $Y2=0
cc_572 N_A_511_47#_M1032_s N_VGND_c_1060_n 0.00250309f $X=10.095 $Y=0.235 $X2=0
+ $Y2=0
cc_573 N_A_511_47#_c_1014_p N_VGND_c_1060_n 0.0124562f $X=6.52 $Y=0.39 $X2=0
+ $Y2=0
cc_574 N_A_511_47#_c_920_n N_VGND_c_1060_n 0.00938601f $X=7.245 $Y=0.82 $X2=0
+ $Y2=0
cc_575 N_A_511_47#_c_950_n N_VGND_c_1060_n 0.0141302f $X=7.46 $Y=0.39 $X2=0
+ $Y2=0
cc_576 N_A_511_47#_c_921_n N_VGND_c_1060_n 0.00972452f $X=8.185 $Y=0.815 $X2=0
+ $Y2=0
cc_577 N_A_511_47#_c_979_n N_VGND_c_1060_n 0.0143352f $X=8.4 $Y=0.39 $X2=0 $Y2=0
cc_578 N_A_511_47#_c_922_n N_VGND_c_1060_n 0.00938601f $X=9.125 $Y=0.82 $X2=0
+ $Y2=0
cc_579 N_A_511_47#_c_954_n N_VGND_c_1060_n 0.0141302f $X=9.34 $Y=0.39 $X2=0
+ $Y2=0
cc_580 N_A_511_47#_c_923_n N_VGND_c_1060_n 0.00972452f $X=10.065 $Y=0.815 $X2=0
+ $Y2=0
cc_581 N_A_511_47#_c_924_n N_VGND_c_1060_n 0.0143352f $X=10.28 $Y=0.39 $X2=0
+ $Y2=0
cc_582 N_A_511_47#_c_925_n N_VGND_c_1060_n 0.0121332f $X=6.015 $Y=0.775 $X2=0
+ $Y2=0
