* NGSPICE file created from sky130_fd_sc_hdll__o21ba_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 VPWR a_186_21# X VPB phighvt w=1e+06u l=180000u
+  ad=1.3807e+12p pd=8.86e+06u as=3.15e+11p ps=2.63e+06u
M1001 a_186_21# a_27_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.45e+11p pd=2.69e+06u as=0p ps=0u
M1002 VGND a_186_21# X VNB nshort w=650000u l=150000u
+  ad=5.66e+11p pd=5.73e+06u as=2.5675e+11p ps=2.09e+06u
M1003 X a_186_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_518_47# a_27_93# a_186_21# VNB nshort w=650000u l=150000u
+  ad=4.4525e+11p pd=3.97e+06u as=1.69e+11p ps=1.82e+06u
M1005 VPWR B1_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1006 VGND A2 a_518_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_518_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_186_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR A1 a_621_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.35e+11p ps=2.47e+06u
M1010 a_621_297# A2 a_186_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B1_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends

