* File: sky130_fd_sc_hdll__einvn_8.pxi.spice
* Created: Wed Sep  2 08:31:26 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVN_8%TE_B N_TE_B_c_146_n N_TE_B_M1014_g
+ N_TE_B_c_141_n N_TE_B_M1024_g N_TE_B_c_142_n N_TE_B_c_143_n N_TE_B_c_149_n
+ N_TE_B_M1000_g N_TE_B_c_150_n N_TE_B_c_151_n N_TE_B_M1002_g N_TE_B_c_152_n
+ N_TE_B_c_153_n N_TE_B_M1005_g N_TE_B_c_154_n N_TE_B_c_155_n N_TE_B_M1011_g
+ N_TE_B_c_156_n N_TE_B_c_157_n N_TE_B_M1012_g N_TE_B_c_158_n N_TE_B_c_159_n
+ N_TE_B_M1016_g N_TE_B_c_160_n N_TE_B_c_161_n N_TE_B_M1026_g N_TE_B_c_162_n
+ N_TE_B_c_163_n N_TE_B_M1031_g N_TE_B_c_144_n N_TE_B_c_165_n N_TE_B_c_166_n
+ N_TE_B_c_167_n N_TE_B_c_168_n N_TE_B_c_169_n N_TE_B_c_170_n TE_B
+ PM_SKY130_FD_SC_HDLL__EINVN_8%TE_B
x_PM_SKY130_FD_SC_HDLL__EINVN_8%A_27_47# N_A_27_47#_M1024_s N_A_27_47#_M1014_s
+ N_A_27_47#_c_278_n N_A_27_47#_M1004_g N_A_27_47#_c_279_n N_A_27_47#_c_280_n
+ N_A_27_47#_c_281_n N_A_27_47#_M1007_g N_A_27_47#_c_282_n N_A_27_47#_c_283_n
+ N_A_27_47#_M1008_g N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_M1015_g
+ N_A_27_47#_c_286_n N_A_27_47#_c_287_n N_A_27_47#_M1018_g N_A_27_47#_c_288_n
+ N_A_27_47#_c_289_n N_A_27_47#_M1025_g N_A_27_47#_c_290_n N_A_27_47#_c_291_n
+ N_A_27_47#_M1028_g N_A_27_47#_c_292_n N_A_27_47#_M1029_g N_A_27_47#_c_293_n
+ N_A_27_47#_c_294_n N_A_27_47#_c_295_n N_A_27_47#_c_296_n N_A_27_47#_c_297_n
+ N_A_27_47#_c_298_n N_A_27_47#_c_299_n N_A_27_47#_c_300_n N_A_27_47#_c_305_n
+ N_A_27_47#_c_301_n N_A_27_47#_c_302_n PM_SKY130_FD_SC_HDLL__EINVN_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVN_8%A N_A_c_435_n N_A_M1009_g N_A_c_445_n
+ N_A_M1001_g N_A_c_436_n N_A_M1010_g N_A_c_446_n N_A_M1003_g N_A_c_437_n
+ N_A_M1019_g N_A_c_447_n N_A_M1006_g N_A_c_438_n N_A_M1020_g N_A_c_448_n
+ N_A_M1013_g N_A_c_439_n N_A_M1021_g N_A_c_449_n N_A_M1017_g N_A_c_440_n
+ N_A_M1022_g N_A_c_450_n N_A_M1023_g N_A_c_441_n N_A_M1030_g N_A_c_451_n
+ N_A_M1027_g N_A_c_452_n N_A_M1032_g N_A_c_442_n N_A_M1033_g A A A A A A A A
+ N_A_c_443_n A A A A A A A A PM_SKY130_FD_SC_HDLL__EINVN_8%A
x_PM_SKY130_FD_SC_HDLL__EINVN_8%VPWR N_VPWR_M1014_d N_VPWR_M1002_d
+ N_VPWR_M1011_d N_VPWR_M1016_d N_VPWR_M1031_d N_VPWR_c_571_n N_VPWR_c_572_n
+ N_VPWR_c_573_n N_VPWR_c_574_n N_VPWR_c_575_n N_VPWR_c_576_n N_VPWR_c_577_n
+ N_VPWR_c_578_n VPWR N_VPWR_c_579_n N_VPWR_c_580_n N_VPWR_c_581_n
+ N_VPWR_c_570_n N_VPWR_c_583_n N_VPWR_c_584_n N_VPWR_c_585_n N_VPWR_c_586_n
+ N_VPWR_c_587_n PM_SKY130_FD_SC_HDLL__EINVN_8%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVN_8%A_222_309# N_A_222_309#_M1000_s
+ N_A_222_309#_M1005_s N_A_222_309#_M1012_s N_A_222_309#_M1026_s
+ N_A_222_309#_M1001_s N_A_222_309#_M1003_s N_A_222_309#_M1013_s
+ N_A_222_309#_M1023_s N_A_222_309#_M1032_s N_A_222_309#_c_712_n
+ N_A_222_309#_c_700_n N_A_222_309#_c_701_n N_A_222_309#_c_720_n
+ N_A_222_309#_c_702_n N_A_222_309#_c_725_n N_A_222_309#_c_703_n
+ N_A_222_309#_c_730_n N_A_222_309#_c_704_n N_A_222_309#_c_705_n
+ N_A_222_309#_c_757_n N_A_222_309#_c_706_n N_A_222_309#_c_822_p
+ N_A_222_309#_c_759_n N_A_222_309#_c_830_p N_A_222_309#_c_761_n
+ N_A_222_309#_c_837_p N_A_222_309#_c_707_n N_A_222_309#_c_708_n
+ N_A_222_309#_c_709_n N_A_222_309#_c_710_n N_A_222_309#_c_711_n
+ N_A_222_309#_c_809_n N_A_222_309#_c_811_n N_A_222_309#_c_813_n
+ PM_SKY130_FD_SC_HDLL__EINVN_8%A_222_309#
x_PM_SKY130_FD_SC_HDLL__EINVN_8%Z N_Z_M1009_d N_Z_M1019_d N_Z_M1021_d
+ N_Z_M1030_d N_Z_M1001_d N_Z_M1006_d N_Z_M1017_d N_Z_M1027_d N_Z_c_860_n
+ N_Z_c_851_n N_Z_c_852_n N_Z_c_871_n N_Z_c_853_n N_Z_c_854_n N_Z_c_855_n
+ N_Z_c_856_n N_Z_c_857_n N_Z_c_858_n Z Z Z Z N_Z_c_908_n N_Z_c_912_n
+ N_Z_c_849_n Z PM_SKY130_FD_SC_HDLL__EINVN_8%Z
x_PM_SKY130_FD_SC_HDLL__EINVN_8%VGND N_VGND_M1024_d N_VGND_M1004_s
+ N_VGND_M1008_s N_VGND_M1018_s N_VGND_M1028_s N_VGND_c_971_n N_VGND_c_972_n
+ N_VGND_c_973_n N_VGND_c_974_n N_VGND_c_975_n N_VGND_c_976_n N_VGND_c_977_n
+ N_VGND_c_978_n N_VGND_c_979_n N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n
+ VGND N_VGND_c_983_n N_VGND_c_984_n N_VGND_c_985_n N_VGND_c_986_n
+ N_VGND_c_987_n PM_SKY130_FD_SC_HDLL__EINVN_8%VGND
x_PM_SKY130_FD_SC_HDLL__EINVN_8%A_235_47# N_A_235_47#_M1004_d
+ N_A_235_47#_M1007_d N_A_235_47#_M1015_d N_A_235_47#_M1025_d
+ N_A_235_47#_M1029_d N_A_235_47#_M1010_s N_A_235_47#_M1020_s
+ N_A_235_47#_M1022_s N_A_235_47#_M1033_s N_A_235_47#_c_1093_n
+ N_A_235_47#_c_1100_n N_A_235_47#_c_1094_n N_A_235_47#_c_1106_n
+ N_A_235_47#_c_1107_n N_A_235_47#_c_1111_n N_A_235_47#_c_1112_n
+ N_A_235_47#_c_1116_n N_A_235_47#_c_1117_n N_A_235_47#_c_1191_n
+ N_A_235_47#_c_1095_n N_A_235_47#_c_1121_n N_A_235_47#_c_1123_n
+ N_A_235_47#_c_1125_n PM_SKY130_FD_SC_HDLL__EINVN_8%A_235_47#
cc_1 VNB N_TE_B_c_141_n 0.0247359f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_TE_B_c_142_n 0.0136496f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_3 VNB N_TE_B_c_143_n 0.0391648f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.25
cc_4 VNB N_TE_B_c_144_n 0.0121778f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.25
cc_5 VNB TE_B 0.0135358f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_27_47#_c_278_n 0.0186317f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_7 VNB N_A_27_47#_c_279_n 0.0137618f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=2.015
cc_8 VNB N_A_27_47#_c_280_n 0.00835566f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=2.015
cc_9 VNB N_A_27_47#_c_281_n 0.0154576f $X=-0.19 $Y=-0.24 $X2=1.4 $Y2=1.395
cc_10 VNB N_A_27_47#_c_282_n 0.0113195f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_11 VNB N_A_27_47#_c_283_n 0.01485f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.395
cc_12 VNB N_A_27_47#_c_284_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=2.015
cc_13 VNB N_A_27_47#_c_285_n 0.0150799f $X=-0.19 $Y=-0.24 $X2=2.34 $Y2=1.395
cc_14 VNB N_A_27_47#_c_286_n 0.0113195f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_15 VNB N_A_27_47#_c_287_n 0.01485f $X=-0.19 $Y=-0.24 $X2=2.81 $Y2=1.395
cc_16 VNB N_A_27_47#_c_288_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=2.9 $Y2=2.015
cc_17 VNB N_A_27_47#_c_289_n 0.0150799f $X=-0.19 $Y=-0.24 $X2=3.28 $Y2=1.395
cc_18 VNB N_A_27_47#_c_290_n 0.0113195f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=2.015
cc_19 VNB N_A_27_47#_c_291_n 0.0149644f $X=-0.19 $Y=-0.24 $X2=3.75 $Y2=1.395
cc_20 VNB N_A_27_47#_c_292_n 0.0397388f $X=-0.19 $Y=-0.24 $X2=4.22 $Y2=1.395
cc_21 VNB N_A_27_47#_c_293_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=2.015
cc_22 VNB N_A_27_47#_c_294_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=2.015
cc_23 VNB N_A_27_47#_c_295_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.25
cc_24 VNB N_A_27_47#_c_296_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_297_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.395
cc_26 VNB N_A_27_47#_c_298_n 0.00473803f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=1.395
cc_27 VNB N_A_27_47#_c_299_n 0.0153763f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.395
cc_28 VNB N_A_27_47#_c_300_n 0.012479f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=1.395
cc_29 VNB N_A_27_47#_c_301_n 0.012178f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_30 VNB N_A_27_47#_c_302_n 0.00887388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_c_435_n 0.0171013f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_32 VNB N_A_c_436_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_33 VNB N_A_c_437_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=1.395
cc_34 VNB N_A_c_438_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.47
cc_35 VNB N_A_c_439_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_36 VNB N_A_c_440_n 0.0169727f $X=-0.19 $Y=-0.24 $X2=2.9 $Y2=2.015
cc_37 VNB N_A_c_441_n 0.0174134f $X=-0.19 $Y=-0.24 $X2=3.75 $Y2=1.395
cc_38 VNB N_A_c_442_n 0.0201569f $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=2.015
cc_39 VNB N_A_c_443_n 0.152272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB A 0.00545171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_570_n 0.383598f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_42 VNB N_Z_c_849_n 0.00954692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB Z 0.0235222f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_971_n 0.00547736f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.395
cc_45 VNB N_VGND_c_972_n 0.0185905f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=2.015
cc_46 VNB N_VGND_c_973_n 0.00501792f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=1.47
cc_47 VNB N_VGND_c_974_n 0.00213025f $X=-0.19 $Y=-0.24 $X2=2.52 $Y2=1.395
cc_48 VNB N_VGND_c_975_n 0.00213025f $X=-0.19 $Y=-0.24 $X2=3.28 $Y2=1.395
cc_49 VNB N_VGND_c_976_n 0.00278323f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=2.015
cc_50 VNB N_VGND_c_977_n 0.0148248f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=1.47
cc_51 VNB N_VGND_c_978_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=3.84 $Y2=2.015
cc_52 VNB N_VGND_c_979_n 0.0148248f $X=-0.19 $Y=-0.24 $X2=4.22 $Y2=1.395
cc_53 VNB N_VGND_c_980_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=3.93 $Y2=1.395
cc_54 VNB N_VGND_c_981_n 0.0148248f $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=2.015
cc_55 VNB N_VGND_c_982_n 0.00526505f $X=-0.19 $Y=-0.24 $X2=4.31 $Y2=2.015
cc_56 VNB N_VGND_c_983_n 0.0143689f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.395
cc_57 VNB N_VGND_c_984_n 0.102609f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_985_n 0.437475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_986_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_987_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_235_47#_c_1093_n 0.00632144f $X=-0.19 $Y=-0.24 $X2=2.52 $Y2=1.395
cc_62 VNB N_A_235_47#_c_1094_n 0.0026801f $X=-0.19 $Y=-0.24 $X2=3.28 $Y2=1.395
cc_63 VNB N_A_235_47#_c_1095_n 0.00962047f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_64 VPB N_TE_B_c_146_n 0.0207069f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB N_TE_B_c_142_n 0.0103502f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.25
cc_66 VPB N_TE_B_c_143_n 0.0172515f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.25
cc_67 VPB N_TE_B_c_149_n 0.0164357f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.47
cc_68 VPB N_TE_B_c_150_n 0.0146992f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_69 VPB N_TE_B_c_151_n 0.0153558f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.47
cc_70 VPB N_TE_B_c_152_n 0.00980191f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.395
cc_71 VPB N_TE_B_c_153_n 0.0156362f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.47
cc_72 VPB N_TE_B_c_154_n 0.00984228f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_73 VPB N_TE_B_c_155_n 0.0153569f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.47
cc_74 VPB N_TE_B_c_156_n 0.00984251f $X=-0.19 $Y=1.305 $X2=2.81 $Y2=1.395
cc_75 VPB N_TE_B_c_157_n 0.0156362f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=1.47
cc_76 VPB N_TE_B_c_158_n 0.00984228f $X=-0.19 $Y=1.305 $X2=3.28 $Y2=1.395
cc_77 VPB N_TE_B_c_159_n 0.0153569f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.47
cc_78 VPB N_TE_B_c_160_n 0.00984251f $X=-0.19 $Y=1.305 $X2=3.75 $Y2=1.395
cc_79 VPB N_TE_B_c_161_n 0.0156362f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=1.47
cc_80 VPB N_TE_B_c_162_n 0.0230223f $X=-0.19 $Y=1.305 $X2=4.22 $Y2=1.395
cc_81 VPB N_TE_B_c_163_n 0.0187512f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.47
cc_82 VPB N_TE_B_c_144_n 0.00718766f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.25
cc_83 VPB N_TE_B_c_165_n 0.00533627f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.395
cc_84 VPB N_TE_B_c_166_n 0.0046927f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.395
cc_85 VPB N_TE_B_c_167_n 0.0046927f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.395
cc_86 VPB N_TE_B_c_168_n 0.0046927f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=1.395
cc_87 VPB N_TE_B_c_169_n 0.0046927f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.395
cc_88 VPB N_TE_B_c_170_n 0.0046927f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=1.395
cc_89 VPB TE_B 0.00306416f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_90 VPB N_A_27_47#_c_292_n 0.00961856f $X=-0.19 $Y=1.305 $X2=4.22 $Y2=1.395
cc_91 VPB N_A_27_47#_c_300_n 0.00959511f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.395
cc_92 VPB N_A_27_47#_c_305_n 0.0304719f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_93 VPB N_A_27_47#_c_301_n 0.00251088f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_94 VPB N_A_c_445_n 0.0209413f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_95 VPB N_A_c_446_n 0.0159705f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=2.015
cc_96 VPB N_A_c_447_n 0.0159705f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_97 VPB N_A_c_448_n 0.0159705f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_98 VPB N_A_c_449_n 0.0159705f $X=-0.19 $Y=1.305 $X2=2.52 $Y2=1.395
cc_99 VPB N_A_c_450_n 0.0159705f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.47
cc_100 VPB N_A_c_451_n 0.0159697f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=2.015
cc_101 VPB N_A_c_452_n 0.019165f $X=-0.19 $Y=1.305 $X2=3.93 $Y2=1.395
cc_102 VPB N_A_c_443_n 0.0997785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_571_n 0.00222504f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=1.395
cc_104 VPB N_VPWR_c_572_n 3.28479e-19 $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_105 VPB N_VPWR_c_573_n 0.0140826f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.47
cc_106 VPB N_VPWR_c_574_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=2.52 $Y2=1.395
cc_107 VPB N_VPWR_c_575_n 0.0140826f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=2.015
cc_108 VPB N_VPWR_c_576_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=3.37 $Y2=1.47
cc_109 VPB N_VPWR_c_577_n 0.0140826f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=2.015
cc_110 VPB N_VPWR_c_578_n 0.0100775f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=2.015
cc_111 VPB N_VPWR_c_579_n 0.0151047f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.47
cc_112 VPB N_VPWR_c_580_n 0.0157606f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.395
cc_113 VPB N_VPWR_c_581_n 0.104313f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_114 VPB N_VPWR_c_570_n 0.0552226f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_115 VPB N_VPWR_c_583_n 0.00580052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_584_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_585_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_586_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_VPWR_c_587_n 0.00618855f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_222_309#_c_700_n 0.00278842f $X=-0.19 $Y=1.305 $X2=3.28 $Y2=1.395
cc_121 VPB N_A_222_309#_c_701_n 0.00177529f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.395
cc_122 VPB N_A_222_309#_c_702_n 0.0026444f $X=-0.19 $Y=1.305 $X2=3.46 $Y2=1.395
cc_123 VPB N_A_222_309#_c_703_n 0.0026444f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=1.47
cc_124 VPB N_A_222_309#_c_704_n 0.0144968f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.395
cc_125 VPB N_A_222_309#_c_705_n 0.00697069f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=1.395
cc_126 VPB N_A_222_309#_c_706_n 0.00193066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_222_309#_c_707_n 0.00820528f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_222_309#_c_708_n 0.021034f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_222_309#_c_709_n 0.00106199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_222_309#_c_710_n 0.00106199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_222_309#_c_711_n 0.00106199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_Z_c_851_n 0.00171122f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=1.47
cc_133 VPB N_Z_c_852_n 0.00174853f $X=-0.19 $Y=1.305 $X2=2.9 $Y2=2.015
cc_134 VPB N_Z_c_853_n 0.00171122f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=2.015
cc_135 VPB N_Z_c_854_n 0.00171122f $X=-0.19 $Y=1.305 $X2=3.75 $Y2=1.395
cc_136 VPB N_Z_c_855_n 0.0104709f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=1.47
cc_137 VPB N_Z_c_856_n 0.00174853f $X=-0.19 $Y=1.305 $X2=3.84 $Y2=2.015
cc_138 VPB N_Z_c_857_n 0.00174853f $X=-0.19 $Y=1.305 $X2=3.93 $Y2=1.395
cc_139 VPB N_Z_c_858_n 0.00174853f $X=-0.19 $Y=1.305 $X2=4.31 $Y2=2.015
cc_140 VPB Z 0.00775893f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 N_TE_B_c_152_n N_A_27_47#_c_279_n 0.0160826f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_142 N_TE_B_c_165_n N_A_27_47#_c_280_n 0.0160826f $X=1.49 $Y=1.395 $X2=0 $Y2=0
cc_143 N_TE_B_c_154_n N_A_27_47#_c_282_n 0.0160826f $X=2.34 $Y=1.395 $X2=0 $Y2=0
cc_144 N_TE_B_c_156_n N_A_27_47#_c_284_n 0.0160826f $X=2.81 $Y=1.395 $X2=0 $Y2=0
cc_145 N_TE_B_c_158_n N_A_27_47#_c_286_n 0.0160826f $X=3.28 $Y=1.395 $X2=0 $Y2=0
cc_146 N_TE_B_c_160_n N_A_27_47#_c_288_n 0.0160826f $X=3.75 $Y=1.395 $X2=0 $Y2=0
cc_147 N_TE_B_c_162_n N_A_27_47#_c_290_n 0.0160826f $X=4.22 $Y=1.395 $X2=0 $Y2=0
cc_148 N_TE_B_c_162_n N_A_27_47#_c_292_n 3.39336e-19 $X=4.22 $Y=1.395 $X2=0
+ $Y2=0
cc_149 N_TE_B_c_166_n N_A_27_47#_c_293_n 0.0160826f $X=1.96 $Y=1.395 $X2=0 $Y2=0
cc_150 N_TE_B_c_167_n N_A_27_47#_c_294_n 0.0160826f $X=2.43 $Y=1.395 $X2=0 $Y2=0
cc_151 N_TE_B_c_168_n N_A_27_47#_c_295_n 0.0160826f $X=2.9 $Y=1.395 $X2=0 $Y2=0
cc_152 N_TE_B_c_169_n N_A_27_47#_c_296_n 0.0160826f $X=3.37 $Y=1.395 $X2=0 $Y2=0
cc_153 N_TE_B_c_170_n N_A_27_47#_c_297_n 0.0160826f $X=3.84 $Y=1.395 $X2=0 $Y2=0
cc_154 N_TE_B_c_141_n N_A_27_47#_c_299_n 0.00611572f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_155 N_TE_B_c_146_n N_A_27_47#_c_300_n 0.0192728f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_156 N_TE_B_c_141_n N_A_27_47#_c_300_n 0.0215796f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_157 N_TE_B_c_142_n N_A_27_47#_c_300_n 0.0171587f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_158 N_TE_B_c_143_n N_A_27_47#_c_300_n 0.0243661f $X=0.595 $Y=1.25 $X2=0 $Y2=0
cc_159 N_TE_B_c_149_n N_A_27_47#_c_300_n 0.00196252f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_160 N_TE_B_c_144_n N_A_27_47#_c_300_n 0.00472039f $X=1.02 $Y=1.25 $X2=0 $Y2=0
cc_161 TE_B N_A_27_47#_c_300_n 0.0678691f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_162 N_TE_B_c_146_n N_A_27_47#_c_305_n 0.00781263f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_163 N_TE_B_c_142_n N_A_27_47#_c_301_n 0.00164242f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_164 N_TE_B_c_150_n N_A_27_47#_c_301_n 0.00914812f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_165 N_TE_B_c_152_n N_A_27_47#_c_301_n 0.00618718f $X=1.87 $Y=1.395 $X2=0
+ $Y2=0
cc_166 N_TE_B_c_154_n N_A_27_47#_c_301_n 0.00621851f $X=2.34 $Y=1.395 $X2=0
+ $Y2=0
cc_167 N_TE_B_c_156_n N_A_27_47#_c_301_n 0.00622389f $X=2.81 $Y=1.395 $X2=0
+ $Y2=0
cc_168 N_TE_B_c_158_n N_A_27_47#_c_301_n 0.00621851f $X=3.28 $Y=1.395 $X2=0
+ $Y2=0
cc_169 N_TE_B_c_160_n N_A_27_47#_c_301_n 0.00622389f $X=3.75 $Y=1.395 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_162_n N_A_27_47#_c_301_n 0.0106577f $X=4.22 $Y=1.395 $X2=0 $Y2=0
cc_171 N_TE_B_c_144_n N_A_27_47#_c_301_n 0.0176781f $X=1.02 $Y=1.25 $X2=0 $Y2=0
cc_172 N_TE_B_c_165_n N_A_27_47#_c_301_n 0.00465183f $X=1.49 $Y=1.395 $X2=0
+ $Y2=0
cc_173 N_TE_B_c_166_n N_A_27_47#_c_301_n 0.00425603f $X=1.96 $Y=1.395 $X2=0
+ $Y2=0
cc_174 N_TE_B_c_167_n N_A_27_47#_c_301_n 0.00425603f $X=2.43 $Y=1.395 $X2=0
+ $Y2=0
cc_175 N_TE_B_c_168_n N_A_27_47#_c_301_n 0.00425603f $X=2.9 $Y=1.395 $X2=0 $Y2=0
cc_176 N_TE_B_c_169_n N_A_27_47#_c_301_n 0.00425603f $X=3.37 $Y=1.395 $X2=0
+ $Y2=0
cc_177 N_TE_B_c_170_n N_A_27_47#_c_301_n 0.00425603f $X=3.84 $Y=1.395 $X2=0
+ $Y2=0
cc_178 N_TE_B_c_146_n N_VPWR_c_571_n 0.0170835f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_179 N_TE_B_c_142_n N_VPWR_c_571_n 0.00105584f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_180 N_TE_B_c_149_n N_VPWR_c_571_n 0.00524796f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_181 N_TE_B_c_149_n N_VPWR_c_572_n 7.75802e-19 $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_182 N_TE_B_c_151_n N_VPWR_c_572_n 0.0154334f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_183 N_TE_B_c_153_n N_VPWR_c_572_n 0.0117009f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_184 N_TE_B_c_155_n N_VPWR_c_572_n 6.61031e-19 $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_185 N_TE_B_c_153_n N_VPWR_c_573_n 0.00622633f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_186 N_TE_B_c_155_n N_VPWR_c_573_n 0.00427505f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_187 N_TE_B_c_153_n N_VPWR_c_574_n 6.99539e-19 $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_188 N_TE_B_c_155_n N_VPWR_c_574_n 0.0153088f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_189 N_TE_B_c_157_n N_VPWR_c_574_n 0.0117009f $X=2.9 $Y=1.47 $X2=0 $Y2=0
cc_190 N_TE_B_c_159_n N_VPWR_c_574_n 6.61031e-19 $X=3.37 $Y=1.47 $X2=0 $Y2=0
cc_191 N_TE_B_c_157_n N_VPWR_c_575_n 0.00622633f $X=2.9 $Y=1.47 $X2=0 $Y2=0
cc_192 N_TE_B_c_159_n N_VPWR_c_575_n 0.00427505f $X=3.37 $Y=1.47 $X2=0 $Y2=0
cc_193 N_TE_B_c_157_n N_VPWR_c_576_n 6.99539e-19 $X=2.9 $Y=1.47 $X2=0 $Y2=0
cc_194 N_TE_B_c_159_n N_VPWR_c_576_n 0.0153088f $X=3.37 $Y=1.47 $X2=0 $Y2=0
cc_195 N_TE_B_c_161_n N_VPWR_c_576_n 0.0117009f $X=3.84 $Y=1.47 $X2=0 $Y2=0
cc_196 N_TE_B_c_163_n N_VPWR_c_576_n 6.61031e-19 $X=4.31 $Y=1.47 $X2=0 $Y2=0
cc_197 N_TE_B_c_161_n N_VPWR_c_577_n 0.00622633f $X=3.84 $Y=1.47 $X2=0 $Y2=0
cc_198 N_TE_B_c_163_n N_VPWR_c_577_n 0.00427505f $X=4.31 $Y=1.47 $X2=0 $Y2=0
cc_199 N_TE_B_c_161_n N_VPWR_c_578_n 7.00525e-19 $X=3.84 $Y=1.47 $X2=0 $Y2=0
cc_200 N_TE_B_c_163_n N_VPWR_c_578_n 0.0163735f $X=4.31 $Y=1.47 $X2=0 $Y2=0
cc_201 N_TE_B_c_146_n N_VPWR_c_579_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_202 N_TE_B_c_149_n N_VPWR_c_580_n 0.00635665f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_203 N_TE_B_c_151_n N_VPWR_c_580_n 0.00427505f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_204 N_TE_B_c_146_n N_VPWR_c_570_n 0.00835414f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_205 N_TE_B_c_149_n N_VPWR_c_570_n 0.0111139f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_206 N_TE_B_c_151_n N_VPWR_c_570_n 0.00740765f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_207 N_TE_B_c_153_n N_VPWR_c_570_n 0.010479f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_208 N_TE_B_c_155_n N_VPWR_c_570_n 0.00740765f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_209 N_TE_B_c_157_n N_VPWR_c_570_n 0.010479f $X=2.9 $Y=1.47 $X2=0 $Y2=0
cc_210 N_TE_B_c_159_n N_VPWR_c_570_n 0.00740765f $X=3.37 $Y=1.47 $X2=0 $Y2=0
cc_211 N_TE_B_c_161_n N_VPWR_c_570_n 0.010479f $X=3.84 $Y=1.47 $X2=0 $Y2=0
cc_212 N_TE_B_c_163_n N_VPWR_c_570_n 0.00740765f $X=4.31 $Y=1.47 $X2=0 $Y2=0
cc_213 N_TE_B_c_146_n N_A_222_309#_c_712_n 7.83445e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_TE_B_c_149_n N_A_222_309#_c_712_n 0.0127872f $X=1.02 $Y=1.47 $X2=0
+ $Y2=0
cc_215 N_TE_B_c_151_n N_A_222_309#_c_712_n 0.00614066f $X=1.49 $Y=1.47 $X2=0
+ $Y2=0
cc_216 N_TE_B_c_151_n N_A_222_309#_c_700_n 0.014571f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_217 N_TE_B_c_152_n N_A_222_309#_c_700_n 0.00250384f $X=1.87 $Y=1.395 $X2=0
+ $Y2=0
cc_218 N_TE_B_c_153_n N_A_222_309#_c_700_n 0.0160672f $X=1.96 $Y=1.47 $X2=0
+ $Y2=0
cc_219 N_TE_B_c_149_n N_A_222_309#_c_701_n 0.00430535f $X=1.02 $Y=1.47 $X2=0
+ $Y2=0
cc_220 N_TE_B_c_150_n N_A_222_309#_c_701_n 0.0026331f $X=1.4 $Y=1.395 $X2=0
+ $Y2=0
cc_221 N_TE_B_c_153_n N_A_222_309#_c_720_n 0.00600706f $X=1.96 $Y=1.47 $X2=0
+ $Y2=0
cc_222 N_TE_B_c_155_n N_A_222_309#_c_720_n 0.00555086f $X=2.43 $Y=1.47 $X2=0
+ $Y2=0
cc_223 N_TE_B_c_155_n N_A_222_309#_c_702_n 0.0145381f $X=2.43 $Y=1.47 $X2=0
+ $Y2=0
cc_224 N_TE_B_c_156_n N_A_222_309#_c_702_n 0.00250384f $X=2.81 $Y=1.395 $X2=0
+ $Y2=0
cc_225 N_TE_B_c_157_n N_A_222_309#_c_702_n 0.0160672f $X=2.9 $Y=1.47 $X2=0 $Y2=0
cc_226 N_TE_B_c_157_n N_A_222_309#_c_725_n 0.00600706f $X=2.9 $Y=1.47 $X2=0
+ $Y2=0
cc_227 N_TE_B_c_159_n N_A_222_309#_c_725_n 0.00555086f $X=3.37 $Y=1.47 $X2=0
+ $Y2=0
cc_228 N_TE_B_c_159_n N_A_222_309#_c_703_n 0.0145381f $X=3.37 $Y=1.47 $X2=0
+ $Y2=0
cc_229 N_TE_B_c_160_n N_A_222_309#_c_703_n 0.00250384f $X=3.75 $Y=1.395 $X2=0
+ $Y2=0
cc_230 N_TE_B_c_161_n N_A_222_309#_c_703_n 0.0160672f $X=3.84 $Y=1.47 $X2=0
+ $Y2=0
cc_231 N_TE_B_c_161_n N_A_222_309#_c_730_n 0.00600706f $X=3.84 $Y=1.47 $X2=0
+ $Y2=0
cc_232 N_TE_B_c_163_n N_A_222_309#_c_730_n 0.00555086f $X=4.31 $Y=1.47 $X2=0
+ $Y2=0
cc_233 N_TE_B_c_162_n N_A_222_309#_c_704_n 2.27622e-19 $X=4.22 $Y=1.395 $X2=0
+ $Y2=0
cc_234 N_TE_B_c_163_n N_A_222_309#_c_704_n 0.0165379f $X=4.31 $Y=1.47 $X2=0
+ $Y2=0
cc_235 N_TE_B_c_163_n N_A_222_309#_c_705_n 0.00381329f $X=4.31 $Y=1.47 $X2=0
+ $Y2=0
cc_236 N_TE_B_c_154_n N_A_222_309#_c_709_n 0.0026331f $X=2.34 $Y=1.395 $X2=0
+ $Y2=0
cc_237 N_TE_B_c_158_n N_A_222_309#_c_710_n 0.0026331f $X=3.28 $Y=1.395 $X2=0
+ $Y2=0
cc_238 N_TE_B_c_162_n N_A_222_309#_c_711_n 0.0026331f $X=4.22 $Y=1.395 $X2=0
+ $Y2=0
cc_239 N_TE_B_c_141_n N_VGND_c_971_n 0.0126377f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_240 N_TE_B_c_142_n N_VGND_c_971_n 7.86225e-19 $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_241 N_TE_B_c_141_n N_VGND_c_983_n 0.00198948f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_242 N_TE_B_c_141_n N_VGND_c_985_n 0.00369246f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_243 N_TE_B_c_141_n N_A_235_47#_c_1093_n 0.00345847f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_TE_B_c_141_n N_A_235_47#_c_1094_n 7.1239e-19 $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_TE_B_c_150_n N_A_235_47#_c_1094_n 0.00101478f $X=1.4 $Y=1.395 $X2=0
+ $Y2=0
cc_246 N_TE_B_c_144_n N_A_235_47#_c_1094_n 2.76908e-19 $X=1.02 $Y=1.25 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_292_n N_A_c_435_n 0.017141f $X=4.865 $Y=0.96 $X2=-0.19
+ $Y2=-0.24
cc_248 N_A_27_47#_c_292_n N_A_c_443_n 0.017141f $X=4.865 $Y=0.96 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_301_n N_A_c_443_n 0.00195057f $X=4.755 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_292_n A 0.00107674f $X=4.865 $Y=0.96 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_301_n A 0.0269779f $X=4.755 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_300_n N_VPWR_M1014_d 0.00340372f $X=0.217 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_253 N_A_27_47#_c_300_n N_VPWR_c_571_n 0.0266259f $X=0.217 $Y=1.665 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_305_n N_VPWR_c_571_n 0.048465f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_305_n N_VPWR_c_579_n 0.0178516f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_256 N_A_27_47#_M1014_s N_VPWR_c_570_n 0.00430086f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_305_n N_VPWR_c_570_n 0.00974347f $X=0.26 $Y=1.815 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_280_n N_A_222_309#_c_700_n 4.62969e-19 $X=1.585 $Y=1.035
+ $X2=0 $Y2=0
cc_259 N_A_27_47#_c_301_n N_A_222_309#_c_700_n 0.0563004f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_c_300_n N_A_222_309#_c_701_n 0.00948929f $X=0.217 $Y=1.665
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_301_n N_A_222_309#_c_701_n 0.0229519f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_282_n N_A_222_309#_c_702_n 2.26097e-19 $X=2.425 $Y=1.035
+ $X2=0 $Y2=0
cc_263 N_A_27_47#_c_294_n N_A_222_309#_c_702_n 3.6695e-19 $X=2.5 $Y=1.035 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_301_n N_A_222_309#_c_702_n 0.0563002f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_286_n N_A_222_309#_c_703_n 2.26097e-19 $X=3.365 $Y=1.035
+ $X2=0 $Y2=0
cc_266 N_A_27_47#_c_296_n N_A_222_309#_c_703_n 3.6695e-19 $X=3.44 $Y=1.035 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_301_n N_A_222_309#_c_703_n 0.0563002f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_290_n N_A_222_309#_c_704_n 2.26097e-19 $X=4.305 $Y=1.035
+ $X2=0 $Y2=0
cc_269 N_A_27_47#_c_292_n N_A_222_309#_c_704_n 0.0081578f $X=4.865 $Y=0.96 $X2=0
+ $Y2=0
cc_270 N_A_27_47#_c_298_n N_A_222_309#_c_704_n 8.94605e-19 $X=4.38 $Y=1.035
+ $X2=0 $Y2=0
cc_271 N_A_27_47#_c_301_n N_A_222_309#_c_704_n 0.0617071f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_272 N_A_27_47#_c_301_n N_A_222_309#_c_709_n 0.0143361f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_301_n N_A_222_309#_c_710_n 0.0143361f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_301_n N_A_222_309#_c_711_n 0.0143361f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_300_n N_VGND_M1024_d 0.0031873f $X=0.217 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_276 N_A_27_47#_c_278_n N_VGND_c_971_n 0.00270009f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_299_n N_VGND_c_971_n 0.0176937f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_300_n N_VGND_c_971_n 0.026897f $X=0.217 $Y=1.665 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_278_n N_VGND_c_972_n 0.00428022f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_278_n N_VGND_c_973_n 0.00320532f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_281_n N_VGND_c_973_n 0.00175624f $X=2.03 $Y=0.96 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_281_n N_VGND_c_974_n 5.76807e-19 $X=2.03 $Y=0.96 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_283_n N_VGND_c_974_n 0.00733819f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_285_n N_VGND_c_974_n 0.00167984f $X=2.97 $Y=0.96 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_285_n N_VGND_c_975_n 5.76807e-19 $X=2.97 $Y=0.96 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_287_n N_VGND_c_975_n 0.00733819f $X=3.44 $Y=0.96 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_289_n N_VGND_c_975_n 0.00167984f $X=3.91 $Y=0.96 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_289_n N_VGND_c_976_n 5.77428e-19 $X=3.91 $Y=0.96 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_291_n N_VGND_c_976_n 0.0073999f $X=4.38 $Y=0.96 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_292_n N_VGND_c_976_n 0.00443615f $X=4.865 $Y=0.96 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_281_n N_VGND_c_977_n 0.00428022f $X=2.03 $Y=0.96 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_283_n N_VGND_c_977_n 0.00341689f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_285_n N_VGND_c_979_n 0.00428022f $X=2.97 $Y=0.96 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_287_n N_VGND_c_979_n 0.00341689f $X=3.44 $Y=0.96 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_289_n N_VGND_c_981_n 0.00428022f $X=3.91 $Y=0.96 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_291_n N_VGND_c_981_n 0.00341689f $X=4.38 $Y=0.96 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_299_n N_VGND_c_983_n 0.0176218f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_298 N_A_27_47#_c_300_n N_VGND_c_983_n 0.00233482f $X=0.217 $Y=1.665 $X2=0
+ $Y2=0
cc_299 N_A_27_47#_c_292_n N_VGND_c_984_n 0.00428022f $X=4.865 $Y=0.96 $X2=0
+ $Y2=0
cc_300 N_A_27_47#_M1024_s N_VGND_c_985_n 0.00292082f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_c_278_n N_VGND_c_985_n 0.00730356f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_281_n N_VGND_c_985_n 0.00605834f $X=2.03 $Y=0.96 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_283_n N_VGND_c_985_n 0.00415805f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_285_n N_VGND_c_985_n 0.005943f $X=2.97 $Y=0.96 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_287_n N_VGND_c_985_n 0.00415805f $X=3.44 $Y=0.96 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_289_n N_VGND_c_985_n 0.005943f $X=3.91 $Y=0.96 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_291_n N_VGND_c_985_n 0.00415805f $X=4.38 $Y=0.96 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_292_n N_VGND_c_985_n 0.00603614f $X=4.865 $Y=0.96 $X2=0
+ $Y2=0
cc_309 N_A_27_47#_c_299_n N_VGND_c_985_n 0.00969887f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_310 N_A_27_47#_c_300_n N_VGND_c_985_n 0.00623299f $X=0.217 $Y=1.665 $X2=0
+ $Y2=0
cc_311 N_A_27_47#_c_278_n N_A_235_47#_c_1100_n 0.0117709f $X=1.51 $Y=0.96 $X2=0
+ $Y2=0
cc_312 N_A_27_47#_c_279_n N_A_235_47#_c_1100_n 0.00378178f $X=1.955 $Y=1.035
+ $X2=0 $Y2=0
cc_313 N_A_27_47#_c_281_n N_A_235_47#_c_1100_n 0.0112338f $X=2.03 $Y=0.96 $X2=0
+ $Y2=0
cc_314 N_A_27_47#_c_301_n N_A_235_47#_c_1100_n 0.048449f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_315 N_A_27_47#_c_300_n N_A_235_47#_c_1094_n 0.0159283f $X=0.217 $Y=1.665
+ $X2=0 $Y2=0
cc_316 N_A_27_47#_c_301_n N_A_235_47#_c_1094_n 0.0272529f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_317 N_A_27_47#_c_283_n N_A_235_47#_c_1106_n 0.00437226f $X=2.5 $Y=0.96 $X2=0
+ $Y2=0
cc_318 N_A_27_47#_c_283_n N_A_235_47#_c_1107_n 0.0106628f $X=2.5 $Y=0.96 $X2=0
+ $Y2=0
cc_319 N_A_27_47#_c_284_n N_A_235_47#_c_1107_n 0.00278658f $X=2.895 $Y=1.035
+ $X2=0 $Y2=0
cc_320 N_A_27_47#_c_285_n N_A_235_47#_c_1107_n 0.0109748f $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_321 N_A_27_47#_c_301_n N_A_235_47#_c_1107_n 0.0479154f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_322 N_A_27_47#_c_287_n N_A_235_47#_c_1111_n 0.00437226f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_287_n N_A_235_47#_c_1112_n 0.0106628f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_288_n N_A_235_47#_c_1112_n 0.00278658f $X=3.835 $Y=1.035
+ $X2=0 $Y2=0
cc_325 N_A_27_47#_c_289_n N_A_235_47#_c_1112_n 0.0109748f $X=3.91 $Y=0.96 $X2=0
+ $Y2=0
cc_326 N_A_27_47#_c_301_n N_A_235_47#_c_1112_n 0.0479154f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_291_n N_A_235_47#_c_1116_n 0.00437226f $X=4.38 $Y=0.96 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_291_n N_A_235_47#_c_1117_n 0.0107736f $X=4.38 $Y=0.96 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_292_n N_A_235_47#_c_1117_n 0.0109528f $X=4.865 $Y=0.96 $X2=0
+ $Y2=0
cc_330 N_A_27_47#_c_301_n N_A_235_47#_c_1117_n 0.0486416f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_302_n N_A_235_47#_c_1117_n 0.00338335f $X=4.62 $Y=1.142
+ $X2=0 $Y2=0
cc_332 N_A_27_47#_c_282_n N_A_235_47#_c_1121_n 0.00268716f $X=2.425 $Y=1.035
+ $X2=0 $Y2=0
cc_333 N_A_27_47#_c_301_n N_A_235_47#_c_1121_n 0.0135367f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_286_n N_A_235_47#_c_1123_n 0.00268716f $X=3.365 $Y=1.035
+ $X2=0 $Y2=0
cc_335 N_A_27_47#_c_301_n N_A_235_47#_c_1123_n 0.0135367f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_336 N_A_27_47#_c_290_n N_A_235_47#_c_1125_n 0.00268716f $X=4.305 $Y=1.035
+ $X2=0 $Y2=0
cc_337 N_A_27_47#_c_301_n N_A_235_47#_c_1125_n 0.0135367f $X=4.755 $Y=1.16 $X2=0
+ $Y2=0
cc_338 N_A_c_445_n N_VPWR_c_578_n 0.00302791f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_339 N_A_c_445_n N_VPWR_c_581_n 0.00429453f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A_c_446_n N_VPWR_c_581_n 0.00429453f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_c_447_n N_VPWR_c_581_n 0.00429453f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A_c_448_n N_VPWR_c_581_n 0.00429453f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_c_449_n N_VPWR_c_581_n 0.00429453f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_c_450_n N_VPWR_c_581_n 0.00429453f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_345 N_A_c_451_n N_VPWR_c_581_n 0.00429453f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_346 N_A_c_452_n N_VPWR_c_581_n 0.00429453f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_c_445_n N_VPWR_c_570_n 0.00743756f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_348 N_A_c_446_n N_VPWR_c_570_n 0.00606499f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_349 N_A_c_447_n N_VPWR_c_570_n 0.00606499f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A_c_448_n N_VPWR_c_570_n 0.00606499f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A_c_449_n N_VPWR_c_570_n 0.00606499f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A_c_450_n N_VPWR_c_570_n 0.00606499f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A_c_451_n N_VPWR_c_570_n 0.00606499f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A_c_452_n N_VPWR_c_570_n 0.00703152f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A_c_445_n N_A_222_309#_c_704_n 0.00313169f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_356 A N_A_222_309#_c_704_n 0.00405228f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_357 N_A_c_445_n N_A_222_309#_c_757_n 0.0145788f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_358 N_A_c_446_n N_A_222_309#_c_757_n 0.0112917f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_359 N_A_c_447_n N_A_222_309#_c_759_n 0.0105301f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_360 N_A_c_448_n N_A_222_309#_c_759_n 0.0112917f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_361 N_A_c_449_n N_A_222_309#_c_761_n 0.0105301f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_362 N_A_c_450_n N_A_222_309#_c_761_n 0.0112917f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_363 N_A_c_451_n N_A_222_309#_c_707_n 0.0105301f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_364 N_A_c_452_n N_A_222_309#_c_707_n 0.0112917f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_365 N_A_c_445_n N_Z_c_860_n 0.00820493f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_366 N_A_c_446_n N_Z_c_860_n 0.00722372f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_367 N_A_c_447_n N_Z_c_860_n 5.29188e-19 $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_368 N_A_c_446_n N_Z_c_851_n 0.0113508f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_369 N_A_c_447_n N_Z_c_851_n 0.00843151f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_370 N_A_c_443_n N_Z_c_851_n 0.00749091f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_371 A N_Z_c_851_n 0.040596f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_372 N_A_c_445_n N_Z_c_852_n 0.00555082f $X=5.35 $Y=1.41 $X2=0 $Y2=0
cc_373 N_A_c_446_n N_Z_c_852_n 0.0011994f $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_374 N_A_c_443_n N_Z_c_852_n 0.00775434f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_375 A N_Z_c_852_n 0.0313201f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_376 N_A_c_446_n N_Z_c_871_n 5.6266e-19 $X=5.82 $Y=1.41 $X2=0 $Y2=0
cc_377 N_A_c_447_n N_Z_c_871_n 0.00926808f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_378 N_A_c_448_n N_Z_c_871_n 0.00722372f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_379 N_A_c_449_n N_Z_c_871_n 5.29188e-19 $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_380 N_A_c_448_n N_Z_c_853_n 0.0113508f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_381 N_A_c_449_n N_Z_c_853_n 0.00843151f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_382 N_A_c_443_n N_Z_c_853_n 0.00749091f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_383 A N_Z_c_853_n 0.040596f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_384 N_A_c_450_n N_Z_c_854_n 0.0113508f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_385 N_A_c_451_n N_Z_c_854_n 0.00843151f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_386 N_A_c_443_n N_Z_c_854_n 0.00749091f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_387 A N_Z_c_854_n 0.040596f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_388 N_A_c_452_n N_Z_c_855_n 0.0139227f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_389 N_A_c_443_n N_Z_c_855_n 3.62918e-19 $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_390 A N_Z_c_855_n 0.00562029f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_391 N_A_c_447_n N_Z_c_856_n 0.00272414f $X=6.29 $Y=1.41 $X2=0 $Y2=0
cc_392 N_A_c_448_n N_Z_c_856_n 0.0011994f $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_393 N_A_c_443_n N_Z_c_856_n 0.00775434f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_394 A N_Z_c_856_n 0.0313201f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_395 N_A_c_449_n N_Z_c_857_n 0.00272414f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_396 N_A_c_450_n N_Z_c_857_n 0.0011994f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_397 N_A_c_443_n N_Z_c_857_n 0.00775434f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_398 A N_Z_c_857_n 0.0313201f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_399 N_A_c_451_n N_Z_c_858_n 0.00272414f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_400 N_A_c_452_n N_Z_c_858_n 0.0011994f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_401 N_A_c_443_n N_Z_c_858_n 0.00754839f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_402 A N_Z_c_858_n 0.0313201f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_403 N_A_c_435_n Z 0.00292377f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_404 N_A_c_436_n Z 0.0096418f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_405 N_A_c_437_n Z 0.0096418f $X=6.265 $Y=0.995 $X2=0 $Y2=0
cc_406 N_A_c_438_n Z 0.0096418f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_407 N_A_c_439_n Z 0.0096418f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_408 N_A_c_440_n Z 0.0096418f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_409 N_A_c_441_n Z 0.0096418f $X=8.145 $Y=0.995 $X2=0 $Y2=0
cc_410 N_A_c_442_n Z 0.0123957f $X=8.665 $Y=0.995 $X2=0 $Y2=0
cc_411 N_A_c_443_n Z 0.0231929f $X=8.64 $Y=1.202 $X2=0 $Y2=0
cc_412 A Z 0.210639f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_413 N_A_c_448_n N_Z_c_908_n 5.6266e-19 $X=6.76 $Y=1.41 $X2=0 $Y2=0
cc_414 N_A_c_449_n N_Z_c_908_n 0.00926808f $X=7.23 $Y=1.41 $X2=0 $Y2=0
cc_415 N_A_c_450_n N_Z_c_908_n 0.00722372f $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_416 N_A_c_451_n N_Z_c_908_n 5.29188e-19 $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_417 N_A_c_450_n N_Z_c_912_n 5.6266e-19 $X=7.7 $Y=1.41 $X2=0 $Y2=0
cc_418 N_A_c_451_n N_Z_c_912_n 0.00926808f $X=8.17 $Y=1.41 $X2=0 $Y2=0
cc_419 N_A_c_452_n N_Z_c_912_n 0.0117662f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_420 N_A_c_452_n Z 0.00164139f $X=8.64 $Y=1.41 $X2=0 $Y2=0
cc_421 N_A_c_442_n Z 0.0195504f $X=8.665 $Y=0.995 $X2=0 $Y2=0
cc_422 A Z 0.0193293f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_423 N_A_c_435_n N_VGND_c_984_n 0.00357877f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_424 N_A_c_436_n N_VGND_c_984_n 0.00357877f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_425 N_A_c_437_n N_VGND_c_984_n 0.00357877f $X=6.265 $Y=0.995 $X2=0 $Y2=0
cc_426 N_A_c_438_n N_VGND_c_984_n 0.00357877f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_427 N_A_c_439_n N_VGND_c_984_n 0.00357877f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_428 N_A_c_440_n N_VGND_c_984_n 0.00357877f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_429 N_A_c_441_n N_VGND_c_984_n 0.00357877f $X=8.145 $Y=0.995 $X2=0 $Y2=0
cc_430 N_A_c_442_n N_VGND_c_984_n 0.00357877f $X=8.665 $Y=0.995 $X2=0 $Y2=0
cc_431 N_A_c_435_n N_VGND_c_985_n 0.00552325f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_432 N_A_c_436_n N_VGND_c_985_n 0.00548399f $X=5.795 $Y=0.995 $X2=0 $Y2=0
cc_433 N_A_c_437_n N_VGND_c_985_n 0.00548399f $X=6.265 $Y=0.995 $X2=0 $Y2=0
cc_434 N_A_c_438_n N_VGND_c_985_n 0.00548399f $X=6.735 $Y=0.995 $X2=0 $Y2=0
cc_435 N_A_c_439_n N_VGND_c_985_n 0.00548399f $X=7.205 $Y=0.995 $X2=0 $Y2=0
cc_436 N_A_c_440_n N_VGND_c_985_n 0.00548399f $X=7.675 $Y=0.995 $X2=0 $Y2=0
cc_437 N_A_c_441_n N_VGND_c_985_n 0.00560377f $X=8.145 $Y=0.995 $X2=0 $Y2=0
cc_438 N_A_c_442_n N_VGND_c_985_n 0.00648779f $X=8.665 $Y=0.995 $X2=0 $Y2=0
cc_439 A N_A_235_47#_c_1117_n 0.00435364f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_440 N_A_c_435_n N_A_235_47#_c_1095_n 0.0112485f $X=5.325 $Y=0.995 $X2=0 $Y2=0
cc_441 N_A_c_436_n N_A_235_47#_c_1095_n 0.00861661f $X=5.795 $Y=0.995 $X2=0
+ $Y2=0
cc_442 N_A_c_437_n N_A_235_47#_c_1095_n 0.00861661f $X=6.265 $Y=0.995 $X2=0
+ $Y2=0
cc_443 N_A_c_438_n N_A_235_47#_c_1095_n 0.00861661f $X=6.735 $Y=0.995 $X2=0
+ $Y2=0
cc_444 N_A_c_439_n N_A_235_47#_c_1095_n 0.00861661f $X=7.205 $Y=0.995 $X2=0
+ $Y2=0
cc_445 N_A_c_440_n N_A_235_47#_c_1095_n 0.00861661f $X=7.675 $Y=0.995 $X2=0
+ $Y2=0
cc_446 N_A_c_441_n N_A_235_47#_c_1095_n 0.00891411f $X=8.145 $Y=0.995 $X2=0
+ $Y2=0
cc_447 N_A_c_442_n N_A_235_47#_c_1095_n 0.00891411f $X=8.665 $Y=0.995 $X2=0
+ $Y2=0
cc_448 A N_A_235_47#_c_1095_n 0.00419156f $X=8.525 $Y=1.19 $X2=0 $Y2=0
cc_449 N_VPWR_c_570_n N_A_222_309#_M1000_s 0.00444633f $X=8.97 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_450 N_VPWR_c_570_n N_A_222_309#_M1005_s 0.00656398f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_451 N_VPWR_c_570_n N_A_222_309#_M1012_s 0.00656398f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_452 N_VPWR_c_570_n N_A_222_309#_M1026_s 0.00656398f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_453 N_VPWR_c_570_n N_A_222_309#_M1001_s 0.00218326f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_454 N_VPWR_c_570_n N_A_222_309#_M1003_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_455 N_VPWR_c_570_n N_A_222_309#_M1013_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_456 N_VPWR_c_570_n N_A_222_309#_M1023_s 0.00231272f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_457 N_VPWR_c_570_n N_A_222_309#_M1032_s 0.00217523f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_458 N_VPWR_c_572_n N_A_222_309#_c_712_n 0.0487409f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_459 N_VPWR_c_580_n N_A_222_309#_c_712_n 0.0171175f $X=1.51 $Y=2.72 $X2=0
+ $Y2=0
cc_460 N_VPWR_c_570_n N_A_222_309#_c_712_n 0.0103125f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_461 N_VPWR_M1002_d N_A_222_309#_c_700_n 0.00187091f $X=1.58 $Y=1.545 $X2=0
+ $Y2=0
cc_462 N_VPWR_c_572_n N_A_222_309#_c_700_n 0.0209383f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_463 N_VPWR_c_572_n N_A_222_309#_c_720_n 0.0385613f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_464 N_VPWR_c_573_n N_A_222_309#_c_720_n 0.0118139f $X=2.45 $Y=2.72 $X2=0
+ $Y2=0
cc_465 N_VPWR_c_574_n N_A_222_309#_c_720_n 0.0470327f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_466 N_VPWR_c_570_n N_A_222_309#_c_720_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_467 N_VPWR_M1011_d N_A_222_309#_c_702_n 0.00187091f $X=2.52 $Y=1.545 $X2=0
+ $Y2=0
cc_468 N_VPWR_c_574_n N_A_222_309#_c_702_n 0.0209383f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_469 N_VPWR_c_574_n N_A_222_309#_c_725_n 0.0385613f $X=2.665 $Y=2.02 $X2=0
+ $Y2=0
cc_470 N_VPWR_c_575_n N_A_222_309#_c_725_n 0.0118139f $X=3.39 $Y=2.72 $X2=0
+ $Y2=0
cc_471 N_VPWR_c_576_n N_A_222_309#_c_725_n 0.0470327f $X=3.605 $Y=2.02 $X2=0
+ $Y2=0
cc_472 N_VPWR_c_570_n N_A_222_309#_c_725_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_473 N_VPWR_M1016_d N_A_222_309#_c_703_n 0.00187091f $X=3.46 $Y=1.545 $X2=0
+ $Y2=0
cc_474 N_VPWR_c_576_n N_A_222_309#_c_703_n 0.0209383f $X=3.605 $Y=2.02 $X2=0
+ $Y2=0
cc_475 N_VPWR_c_576_n N_A_222_309#_c_730_n 0.0385613f $X=3.605 $Y=2.02 $X2=0
+ $Y2=0
cc_476 N_VPWR_c_577_n N_A_222_309#_c_730_n 0.0118139f $X=4.33 $Y=2.72 $X2=0
+ $Y2=0
cc_477 N_VPWR_c_578_n N_A_222_309#_c_730_n 0.047223f $X=4.545 $Y=2 $X2=0 $Y2=0
cc_478 N_VPWR_c_570_n N_A_222_309#_c_730_n 0.00646998f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_479 N_VPWR_M1031_d N_A_222_309#_c_704_n 0.00285703f $X=4.4 $Y=1.545 $X2=0
+ $Y2=0
cc_480 N_VPWR_c_578_n N_A_222_309#_c_704_n 0.0275265f $X=4.545 $Y=2 $X2=0 $Y2=0
cc_481 N_VPWR_c_578_n N_A_222_309#_c_705_n 0.0317623f $X=4.545 $Y=2 $X2=0 $Y2=0
cc_482 N_VPWR_c_581_n N_A_222_309#_c_757_n 0.0415295f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_570_n N_A_222_309#_c_757_n 0.026948f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_484 N_VPWR_c_578_n N_A_222_309#_c_706_n 0.0127186f $X=4.545 $Y=2 $X2=0 $Y2=0
cc_485 N_VPWR_c_581_n N_A_222_309#_c_706_n 0.0176351f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_486 N_VPWR_c_570_n N_A_222_309#_c_706_n 0.00962794f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_487 N_VPWR_c_581_n N_A_222_309#_c_759_n 0.0415032f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_488 N_VPWR_c_570_n N_A_222_309#_c_759_n 0.0268781f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_489 N_VPWR_c_581_n N_A_222_309#_c_761_n 0.0415032f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_490 N_VPWR_c_570_n N_A_222_309#_c_761_n 0.0268781f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_491 N_VPWR_c_581_n N_A_222_309#_c_707_n 0.0630218f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_492 N_VPWR_c_570_n N_A_222_309#_c_707_n 0.0386144f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_493 N_VPWR_c_581_n N_A_222_309#_c_809_n 0.0119417f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_494 N_VPWR_c_570_n N_A_222_309#_c_809_n 0.00654447f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_495 N_VPWR_c_581_n N_A_222_309#_c_811_n 0.0119417f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_496 N_VPWR_c_570_n N_A_222_309#_c_811_n 0.00654447f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_497 N_VPWR_c_581_n N_A_222_309#_c_813_n 0.0119417f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_498 N_VPWR_c_570_n N_A_222_309#_c_813_n 0.00654447f $X=8.97 $Y=2.72 $X2=0
+ $Y2=0
cc_499 N_VPWR_c_570_n N_Z_M1001_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_c_570_n N_Z_M1006_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_501 N_VPWR_c_570_n N_Z_M1017_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_502 N_VPWR_c_570_n N_Z_M1027_d 0.00232895f $X=8.97 $Y=2.72 $X2=0 $Y2=0
cc_503 N_A_222_309#_c_757_n N_Z_M1001_d 0.00352392f $X=5.97 $Y=2.38 $X2=0 $Y2=0
cc_504 N_A_222_309#_c_759_n N_Z_M1006_d 0.00352392f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_505 N_A_222_309#_c_761_n N_Z_M1017_d 0.00352392f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_506 N_A_222_309#_c_707_n N_Z_M1027_d 0.00352392f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_507 N_A_222_309#_c_704_n N_Z_c_860_n 0.00329755f $X=4.95 $Y=1.58 $X2=0 $Y2=0
cc_508 N_A_222_309#_c_705_n N_Z_c_860_n 0.0352962f $X=5.115 $Y=1.815 $X2=0 $Y2=0
cc_509 N_A_222_309#_c_757_n N_Z_c_860_n 0.0195903f $X=5.97 $Y=2.38 $X2=0 $Y2=0
cc_510 N_A_222_309#_c_822_p N_Z_c_860_n 0.0201988f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_511 N_A_222_309#_M1003_s N_Z_c_851_n 0.00178587f $X=5.91 $Y=1.485 $X2=0 $Y2=0
cc_512 N_A_222_309#_c_757_n N_Z_c_851_n 0.00346334f $X=5.97 $Y=2.38 $X2=0 $Y2=0
cc_513 N_A_222_309#_c_822_p N_Z_c_851_n 0.0136517f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_514 N_A_222_309#_c_759_n N_Z_c_851_n 0.00238643f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_515 N_A_222_309#_c_704_n N_Z_c_852_n 0.0113624f $X=4.95 $Y=1.58 $X2=0 $Y2=0
cc_516 N_A_222_309#_c_822_p N_Z_c_871_n 0.0246362f $X=6.055 $Y=1.96 $X2=0 $Y2=0
cc_517 N_A_222_309#_c_759_n N_Z_c_871_n 0.0195903f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_518 N_A_222_309#_c_830_p N_Z_c_871_n 0.0201988f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_519 N_A_222_309#_M1013_s N_Z_c_853_n 0.00178587f $X=6.85 $Y=1.485 $X2=0 $Y2=0
cc_520 N_A_222_309#_c_759_n N_Z_c_853_n 0.00346334f $X=6.91 $Y=2.38 $X2=0 $Y2=0
cc_521 N_A_222_309#_c_830_p N_Z_c_853_n 0.0136517f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_522 N_A_222_309#_c_761_n N_Z_c_853_n 0.00238643f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_523 N_A_222_309#_M1023_s N_Z_c_854_n 0.00178587f $X=7.79 $Y=1.485 $X2=0 $Y2=0
cc_524 N_A_222_309#_c_761_n N_Z_c_854_n 0.00346334f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_525 N_A_222_309#_c_837_p N_Z_c_854_n 0.0136517f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_526 N_A_222_309#_c_707_n N_Z_c_854_n 0.00238643f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_527 N_A_222_309#_M1032_s N_Z_c_855_n 0.00296518f $X=8.73 $Y=1.485 $X2=0 $Y2=0
cc_528 N_A_222_309#_c_707_n N_Z_c_855_n 0.00346334f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_529 N_A_222_309#_c_708_n N_Z_c_855_n 0.026889f $X=8.875 $Y=1.96 $X2=0 $Y2=0
cc_530 N_A_222_309#_c_830_p N_Z_c_908_n 0.0246362f $X=6.995 $Y=1.96 $X2=0 $Y2=0
cc_531 N_A_222_309#_c_761_n N_Z_c_908_n 0.0195903f $X=7.85 $Y=2.38 $X2=0 $Y2=0
cc_532 N_A_222_309#_c_837_p N_Z_c_908_n 0.0201988f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_533 N_A_222_309#_c_837_p N_Z_c_912_n 0.0246362f $X=7.935 $Y=1.96 $X2=0 $Y2=0
cc_534 N_A_222_309#_c_707_n N_Z_c_912_n 0.0195903f $X=8.79 $Y=2.38 $X2=0 $Y2=0
cc_535 N_A_222_309#_c_708_n N_Z_c_912_n 0.021104f $X=8.875 $Y=1.96 $X2=0 $Y2=0
cc_536 N_A_222_309#_c_704_n N_A_235_47#_c_1117_n 0.00485941f $X=4.95 $Y=1.58
+ $X2=0 $Y2=0
cc_537 N_Z_M1009_d N_VGND_c_985_n 0.00256987f $X=5.4 $Y=0.235 $X2=0 $Y2=0
cc_538 N_Z_M1019_d N_VGND_c_985_n 0.00256987f $X=6.34 $Y=0.235 $X2=0 $Y2=0
cc_539 N_Z_M1021_d N_VGND_c_985_n 0.00256987f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_540 N_Z_M1030_d N_VGND_c_985_n 0.00297142f $X=8.22 $Y=0.235 $X2=0 $Y2=0
cc_541 Z N_A_235_47#_M1010_s 0.00400356f $X=8.87 $Y=0.765 $X2=0 $Y2=0
cc_542 Z N_A_235_47#_M1020_s 0.00400356f $X=8.87 $Y=0.765 $X2=0 $Y2=0
cc_543 Z N_A_235_47#_M1022_s 0.00400356f $X=8.87 $Y=0.765 $X2=0 $Y2=0
cc_544 Z N_A_235_47#_M1033_s 0.00212897f $X=8.87 $Y=0.765 $X2=0 $Y2=0
cc_545 N_Z_c_849_n N_A_235_47#_M1033_s 0.00273062f $X=8.982 $Y=0.825 $X2=0 $Y2=0
cc_546 Z N_A_235_47#_M1033_s 0.00101757f $X=8.955 $Y=0.85 $X2=0 $Y2=0
cc_547 N_Z_M1009_d N_A_235_47#_c_1095_n 0.00399896f $X=5.4 $Y=0.235 $X2=0 $Y2=0
cc_548 N_Z_M1019_d N_A_235_47#_c_1095_n 0.00399896f $X=6.34 $Y=0.235 $X2=0 $Y2=0
cc_549 N_Z_M1021_d N_A_235_47#_c_1095_n 0.00399896f $X=7.28 $Y=0.235 $X2=0 $Y2=0
cc_550 N_Z_M1030_d N_A_235_47#_c_1095_n 0.00505942f $X=8.22 $Y=0.235 $X2=0 $Y2=0
cc_551 Z N_A_235_47#_c_1095_n 0.180698f $X=8.87 $Y=0.765 $X2=0 $Y2=0
cc_552 N_Z_c_849_n N_A_235_47#_c_1095_n 0.0176261f $X=8.982 $Y=0.825 $X2=0 $Y2=0
cc_553 N_VGND_c_985_n N_A_235_47#_M1004_d 0.00229009f $X=8.97 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_554 N_VGND_c_985_n N_A_235_47#_M1007_d 0.00314422f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_985_n N_A_235_47#_M1015_d 0.00314422f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_985_n N_A_235_47#_M1025_d 0.00314422f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_985_n N_A_235_47#_M1029_d 0.00266653f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_985_n N_A_235_47#_M1010_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_985_n N_A_235_47#_M1020_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_985_n N_A_235_47#_M1022_s 0.00255381f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_985_n N_A_235_47#_M1033_s 0.00225742f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_971_n N_A_235_47#_c_1093_n 0.0193138f $X=0.73 $Y=0.38 $X2=0
+ $Y2=0
cc_563 N_VGND_c_972_n N_A_235_47#_c_1093_n 0.0220167f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_c_985_n N_A_235_47#_c_1093_n 0.0121907f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_M1004_s N_A_235_47#_c_1100_n 0.00491295f $X=1.585 $Y=0.235 $X2=0
+ $Y2=0
cc_566 N_VGND_c_972_n N_A_235_47#_c_1100_n 0.0029785f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_973_n N_A_235_47#_c_1100_n 0.0196524f $X=1.77 $Y=0.36 $X2=0
+ $Y2=0
cc_568 N_VGND_c_977_n N_A_235_47#_c_1100_n 0.0029785f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_569 N_VGND_c_985_n N_A_235_47#_c_1100_n 0.0120605f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_974_n N_A_235_47#_c_1106_n 0.0139248f $X=2.71 $Y=0.36 $X2=0
+ $Y2=0
cc_571 N_VGND_c_977_n N_A_235_47#_c_1106_n 0.011459f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_985_n N_A_235_47#_c_1106_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_M1008_s N_A_235_47#_c_1107_n 0.0038973f $X=2.575 $Y=0.235 $X2=0
+ $Y2=0
cc_574 N_VGND_c_974_n N_A_235_47#_c_1107_n 0.0178569f $X=2.71 $Y=0.36 $X2=0
+ $Y2=0
cc_575 N_VGND_c_977_n N_A_235_47#_c_1107_n 0.00310196f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_576 N_VGND_c_979_n N_A_235_47#_c_1107_n 0.0029785f $X=3.485 $Y=0 $X2=0 $Y2=0
cc_577 N_VGND_c_985_n N_A_235_47#_c_1107_n 0.0122777f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_578 N_VGND_c_975_n N_A_235_47#_c_1111_n 0.0139248f $X=3.65 $Y=0.36 $X2=0
+ $Y2=0
cc_579 N_VGND_c_979_n N_A_235_47#_c_1111_n 0.011459f $X=3.485 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_985_n N_A_235_47#_c_1111_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_581 N_VGND_M1018_s N_A_235_47#_c_1112_n 0.0038973f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_582 N_VGND_c_975_n N_A_235_47#_c_1112_n 0.0178569f $X=3.65 $Y=0.36 $X2=0
+ $Y2=0
cc_583 N_VGND_c_979_n N_A_235_47#_c_1112_n 0.00310196f $X=3.485 $Y=0 $X2=0 $Y2=0
cc_584 N_VGND_c_981_n N_A_235_47#_c_1112_n 0.0029785f $X=4.425 $Y=0 $X2=0 $Y2=0
cc_585 N_VGND_c_985_n N_A_235_47#_c_1112_n 0.0122777f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_586 N_VGND_c_976_n N_A_235_47#_c_1116_n 0.013957f $X=4.59 $Y=0.36 $X2=0 $Y2=0
cc_587 N_VGND_c_981_n N_A_235_47#_c_1116_n 0.011459f $X=4.425 $Y=0 $X2=0 $Y2=0
cc_588 N_VGND_c_985_n N_A_235_47#_c_1116_n 0.00644035f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_589 N_VGND_M1028_s N_A_235_47#_c_1117_n 0.00425468f $X=4.455 $Y=0.235 $X2=0
+ $Y2=0
cc_590 N_VGND_c_976_n N_A_235_47#_c_1117_n 0.0190084f $X=4.59 $Y=0.36 $X2=0
+ $Y2=0
cc_591 N_VGND_c_981_n N_A_235_47#_c_1117_n 0.00310196f $X=4.425 $Y=0 $X2=0 $Y2=0
cc_592 N_VGND_c_984_n N_A_235_47#_c_1117_n 0.0029785f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_593 N_VGND_c_985_n N_A_235_47#_c_1117_n 0.0123613f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_594 N_VGND_c_984_n N_A_235_47#_c_1191_n 0.0142806f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_595 N_VGND_c_985_n N_A_235_47#_c_1191_n 0.00824212f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_596 N_VGND_c_984_n N_A_235_47#_c_1095_n 0.220821f $X=8.97 $Y=0 $X2=0 $Y2=0
cc_597 N_VGND_c_985_n N_A_235_47#_c_1095_n 0.13954f $X=8.97 $Y=0 $X2=0 $Y2=0
