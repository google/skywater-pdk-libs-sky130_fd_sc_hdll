* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb4to1_2 D[3] D[2] D[1] D[0] S[3] S[2] S[1] S[0] VGND
+ VNB VPB VPWR Z
X0 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_2112_333# a_1989_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X2 Z a_278_265# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X3 Z S[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 a_845_69# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X5 VPWR D[3] a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_27_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND D[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 VGND D[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_1566_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 Z a_701_47# a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_845_69# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_2133_69# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR S[1] a_701_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_824_333# a_701_47# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X15 a_27_297# a_278_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X17 a_27_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 VGND S[1] a_701_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X19 a_278_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_2112_333# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR D[1] a_824_333# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VPWR D[2] a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 VGND D[0] a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_27_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X26 Z S[3] a_2133_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X27 a_824_333# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_1315_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_2133_69# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X31 VPWR D[0] a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 Z S[1] a_845_69# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X33 VGND S[3] a_1989_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_278_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 Z a_1566_265# a_1315_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X36 VPWR S[3] a_1989_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 a_1315_297# a_1566_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 a_1566_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X39 Z a_1989_47# a_2112_333# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
.ends
