* File: sky130_fd_sc_hdll__clkbuf_2.pxi.spice
* Created: Thu Aug 27 19:01:42 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_2%A N_A_c_40_n N_A_M1002_g N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__CLKBUF_2%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_2%A_27_47# N_A_27_47#_M1000_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_69_n N_A_27_47#_M1001_g N_A_27_47#_c_74_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_75_n N_A_27_47#_M1005_g N_A_27_47#_c_70_n N_A_27_47#_M1003_g
+ N_A_27_47#_c_71_n N_A_27_47#_c_77_n N_A_27_47#_c_86_n N_A_27_47#_c_78_n
+ N_A_27_47#_c_72_n N_A_27_47#_c_79_n N_A_27_47#_c_73_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_2%VPWR N_VPWR_M1002_d N_VPWR_M1005_d
+ N_VPWR_c_133_n N_VPWR_c_134_n VPWR N_VPWR_c_135_n N_VPWR_c_136_n
+ N_VPWR_c_137_n N_VPWR_c_132_n N_VPWR_c_139_n N_VPWR_c_140_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_2%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_2%X N_X_M1001_s N_X_M1004_s N_X_c_165_n
+ N_X_c_176_n X X X X X X PM_SKY130_FD_SC_HDLL__CLKBUF_2%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_2%VGND N_VGND_M1000_d N_VGND_M1003_d
+ N_VGND_c_205_n N_VGND_c_206_n VGND N_VGND_c_207_n N_VGND_c_208_n
+ N_VGND_c_209_n N_VGND_c_210_n N_VGND_c_211_n N_VGND_c_212_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_2%VGND
cc_1 VNB N_A_c_40_n 0.0323065f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_A_M1000_g 0.0325693f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.445
cc_3 VNB A 0.00879335f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.765
cc_4 VNB N_A_27_47#_c_69_n 0.016451f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_27_47#_c_70_n 0.0179824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_71_n 0.0330785f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_c_72_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_73_n 0.0716888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VPWR_c_132_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_X_c_165_n 4.05749e-19 $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_11 VNB X 0.0134156f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=0.85
cc_12 VNB X 0.020783f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_205_n 0.00474165f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_14 VNB N_VGND_c_206_n 0.013686f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_15 VNB N_VGND_c_207_n 0.0182778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_208_n 0.0164481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_209_n 0.0148721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_210_n 0.154942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_211_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_212_n 0.0058339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_A_c_40_n 0.0318843f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_22 VPB A 0.00123495f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.765
cc_23 VPB N_A_27_47#_c_74_n 0.0165244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_24 VPB N_A_27_47#_c_75_n 0.0184706f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_25 VPB N_A_27_47#_c_71_n 0.0090886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_47#_c_77_n 0.0297332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_A_27_47#_c_78_n 5.29992e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_27_47#_c_79_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_A_27_47#_c_73_n 0.0213144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_133_n 0.00229023f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.105
cc_31 VPB N_VPWR_c_134_n 0.0147361f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_32 VPB N_VPWR_c_135_n 0.0154253f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_136_n 0.0159877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_137_n 0.0148721f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_VPWR_c_132_n 0.0557756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_139_n 0.00583344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_140_n 0.00589477f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB X 0.00743383f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_39 VPB X 0.0218946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 N_A_M1000_g N_A_27_47#_c_69_n 0.00975348f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_41 N_A_c_40_n N_A_27_47#_c_74_n 0.0169499f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_42 N_A_c_40_n N_A_27_47#_c_71_n 0.0152606f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_43 N_A_M1000_g N_A_27_47#_c_71_n 0.00636688f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_44 A N_A_27_47#_c_71_n 0.0452976f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_45 N_A_c_40_n N_A_27_47#_c_86_n 0.0180013f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_46 A N_A_27_47#_c_86_n 0.0297086f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_47 N_A_c_40_n N_A_27_47#_c_78_n 0.00121365f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_78_n 0.0252837f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_49 N_A_c_40_n N_A_27_47#_c_79_n 4.39692e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A_c_40_n N_A_27_47#_c_73_n 0.0377942f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_51 A N_A_27_47#_c_73_n 0.00616608f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_52 N_A_c_40_n N_VPWR_c_133_n 0.0175719f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A_c_40_n N_VPWR_c_135_n 0.00447018f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_54 N_A_c_40_n N_VPWR_c_132_n 0.00866609f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_55 A X 0.00434654f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_56 A X 0.00495573f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_57 N_A_c_40_n N_VGND_c_205_n 4.03454e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_M1000_g N_VGND_c_205_n 0.00317144f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_59 A N_VGND_c_205_n 0.0168184f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_60 N_A_M1000_g N_VGND_c_207_n 0.00440413f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_61 A N_VGND_c_207_n 0.00256127f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_62 N_A_M1000_g N_VGND_c_210_n 0.00698017f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_63 A N_VGND_c_210_n 0.00504947f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_64 N_A_27_47#_c_86_n N_VPWR_M1002_d 0.00607473f $X=1.015 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_27_47#_c_74_n N_VPWR_c_133_n 0.00175741f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_27_47#_c_86_n N_VPWR_c_133_n 0.021715f $X=1.015 $Y=1.58 $X2=0 $Y2=0
cc_67 N_A_27_47#_c_74_n N_VPWR_c_134_n 6.30662e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A_27_47#_c_75_n N_VPWR_c_134_n 0.0115029f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A_27_47#_c_77_n N_VPWR_c_135_n 0.0158305f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_70 N_A_27_47#_c_74_n N_VPWR_c_136_n 0.00702461f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_71 N_A_27_47#_c_75_n N_VPWR_c_136_n 0.00316784f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_27_47#_M1002_s N_VPWR_c_132_n 0.0041805f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_73 N_A_27_47#_c_74_n N_VPWR_c_132_n 0.0127459f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_27_47#_c_75_n N_VPWR_c_132_n 0.00385556f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_77_n N_VPWR_c_132_n 0.0101646f $X=0.26 $Y=1.745 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_86_n N_X_M1004_s 0.00314634f $X=1.015 $Y=1.58 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_69_n N_X_c_165_n 0.00332787f $X=1 $Y=0.745 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_70_n N_X_c_165_n 0.00412399f $X=1.52 $Y=0.745 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_73_n N_X_c_165_n 0.00122054f $X=1.495 $Y=1.077 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_75_n N_X_c_176_n 0.00442044f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_69_n X 0.00287689f $X=1 $Y=0.745 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_70_n X 0.00678842f $X=1.52 $Y=0.745 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_78_n X 0.013238f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_73_n X 0.0191794f $X=1.495 $Y=1.077 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_75_n X 0.0156204f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_86_n X 0.0106739f $X=1.015 $Y=1.58 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_73_n X 0.00242395f $X=1.495 $Y=1.077 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_74_n X 0.00123218f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_75_n X 0.0179872f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_86_n X 0.0142044f $X=1.015 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_78_n X 0.0380469f $X=1.1 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_73_n X 0.0283687f $X=1.495 $Y=1.077 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_69_n N_VGND_c_205_n 0.00158701f $X=1 $Y=0.745 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_69_n N_VGND_c_206_n 5.58224e-19 $X=1 $Y=0.745 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_70_n N_VGND_c_206_n 0.0112285f $X=1.52 $Y=0.745 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_72_n N_VGND_c_207_n 0.0173041f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_69_n N_VGND_c_208_n 0.00585385f $X=1 $Y=0.745 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_70_n N_VGND_c_208_n 0.00199015f $X=1.52 $Y=0.745 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1000_s N_VGND_c_210_n 0.00547712f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_69_n N_VGND_c_210_n 0.0109235f $X=1 $Y=0.745 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_70_n N_VGND_c_210_n 0.00285558f $X=1.52 $Y=0.745 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_72_n N_VGND_c_210_n 0.00982816f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_103 N_VPWR_c_132_n N_X_M1004_s 0.00416463f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_104 N_VPWR_c_134_n N_X_c_176_n 0.016919f $X=1.73 $Y=2.295 $X2=0 $Y2=0
cc_105 N_VPWR_c_136_n N_X_c_176_n 0.0101029f $X=1.515 $Y=2.72 $X2=0 $Y2=0
cc_106 N_VPWR_c_132_n N_X_c_176_n 0.00684471f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_107 N_VPWR_M1005_d X 0.00374364f $X=1.585 $Y=1.485 $X2=0 $Y2=0
cc_108 N_VPWR_c_134_n X 0.0219654f $X=1.73 $Y=2.295 $X2=0 $Y2=0
cc_109 N_VPWR_c_136_n X 0.00213799f $X=1.515 $Y=2.72 $X2=0 $Y2=0
cc_110 N_VPWR_c_132_n X 0.00561876f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_M1005_d X 0.00241487f $X=1.585 $Y=1.485 $X2=0 $Y2=0
cc_112 N_X_c_165_n N_VGND_c_206_n 0.0174262f $X=1.26 $Y=0.42 $X2=0 $Y2=0
cc_113 X N_VGND_c_206_n 0.0250101f $X=1.675 $Y=0.765 $X2=0 $Y2=0
cc_114 N_X_c_165_n N_VGND_c_208_n 0.0137398f $X=1.26 $Y=0.42 $X2=0 $Y2=0
cc_115 X N_VGND_c_208_n 0.00287214f $X=1.675 $Y=0.765 $X2=0 $Y2=0
cc_116 N_X_M1001_s N_VGND_c_210_n 0.00558965f $X=1.075 $Y=0.235 $X2=0 $Y2=0
cc_117 N_X_c_165_n N_VGND_c_210_n 0.00771386f $X=1.26 $Y=0.42 $X2=0 $Y2=0
cc_118 X N_VGND_c_210_n 0.00595232f $X=1.675 $Y=0.765 $X2=0 $Y2=0
