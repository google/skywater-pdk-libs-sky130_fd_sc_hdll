* File: sky130_fd_sc_hdll__inv_12.pxi.spice
* Created: Thu Aug 27 19:08:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_12%A N_A_c_88_n N_A_M1000_g N_A_c_101_n N_A_M1002_g
+ N_A_c_89_n N_A_M1001_g N_A_c_102_n N_A_M1003_g N_A_c_90_n N_A_M1005_g
+ N_A_c_103_n N_A_M1004_g N_A_c_91_n N_A_M1007_g N_A_c_104_n N_A_M1006_g
+ N_A_c_92_n N_A_M1011_g N_A_c_105_n N_A_M1008_g N_A_c_93_n N_A_M1012_g
+ N_A_c_106_n N_A_M1009_g N_A_c_94_n N_A_M1013_g N_A_c_107_n N_A_M1010_g
+ N_A_c_95_n N_A_M1014_g N_A_c_108_n N_A_M1015_g N_A_c_96_n N_A_M1016_g
+ N_A_c_109_n N_A_M1017_g N_A_c_97_n N_A_M1020_g N_A_c_110_n N_A_M1018_g
+ N_A_c_98_n N_A_M1022_g N_A_c_111_n N_A_M1019_g N_A_c_112_n N_A_M1021_g
+ N_A_c_99_n N_A_M1023_g A A A A A A A A A N_A_c_161_p N_A_c_100_n A A A A A A A
+ A PM_SKY130_FD_SC_HDLL__INV_12%A
x_PM_SKY130_FD_SC_HDLL__INV_12%VPWR N_VPWR_M1002_s N_VPWR_M1003_s N_VPWR_M1006_s
+ N_VPWR_M1009_s N_VPWR_M1015_s N_VPWR_M1018_s N_VPWR_M1021_s N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ N_VPWR_c_331_n N_VPWR_c_332_n N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n
+ N_VPWR_c_336_n N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n N_VPWR_c_340_n
+ N_VPWR_c_341_n N_VPWR_c_342_n N_VPWR_c_343_n VPWR N_VPWR_c_344_n
+ N_VPWR_c_324_n PM_SKY130_FD_SC_HDLL__INV_12%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_12%Y N_Y_M1000_d N_Y_M1005_d N_Y_M1011_d N_Y_M1013_d
+ N_Y_M1016_d N_Y_M1022_d N_Y_M1002_d N_Y_M1004_d N_Y_M1008_d N_Y_M1010_d
+ N_Y_M1017_d N_Y_M1019_d N_Y_c_444_n N_Y_c_447_n N_Y_c_426_n N_Y_c_427_n
+ N_Y_c_457_n N_Y_c_440_n N_Y_c_464_n N_Y_c_468_n N_Y_c_428_n N_Y_c_476_n
+ N_Y_c_480_n N_Y_c_484_n N_Y_c_429_n N_Y_c_492_n N_Y_c_496_n N_Y_c_500_n
+ N_Y_c_430_n N_Y_c_508_n N_Y_c_512_n N_Y_c_516_n N_Y_c_431_n N_Y_c_524_n
+ N_Y_c_528_n N_Y_c_530_n N_Y_c_432_n N_Y_c_441_n N_Y_c_433_n N_Y_c_541_n
+ N_Y_c_434_n N_Y_c_549_n N_Y_c_435_n N_Y_c_557_n N_Y_c_436_n N_Y_c_565_n
+ N_Y_c_437_n N_Y_c_572_n Y Y PM_SKY130_FD_SC_HDLL__INV_12%Y
x_PM_SKY130_FD_SC_HDLL__INV_12%VGND N_VGND_M1000_s N_VGND_M1001_s N_VGND_M1007_s
+ N_VGND_M1012_s N_VGND_M1014_s N_VGND_M1020_s N_VGND_M1023_s N_VGND_c_683_n
+ N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n N_VGND_c_698_n
+ N_VGND_c_699_n N_VGND_c_700_n N_VGND_c_701_n VGND N_VGND_c_702_n
+ N_VGND_c_703_n PM_SKY130_FD_SC_HDLL__INV_12%VGND
cc_1 VNB N_A_c_88_n 0.0196289f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=0.995
cc_2 VNB N_A_c_89_n 0.0167438f $X=-0.19 $Y=-0.24 $X2=1.105 $Y2=0.995
cc_3 VNB N_A_c_90_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.575 $Y2=0.995
cc_4 VNB N_A_c_91_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.045 $Y2=0.995
cc_5 VNB N_A_c_92_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.515 $Y2=0.995
cc_6 VNB N_A_c_93_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=2.985 $Y2=0.995
cc_7 VNB N_A_c_94_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=3.455 $Y2=0.995
cc_8 VNB N_A_c_95_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.995
cc_9 VNB N_A_c_96_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=0.995
cc_10 VNB N_A_c_97_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=4.865 $Y2=0.995
cc_11 VNB N_A_c_98_n 0.0171975f $X=-0.19 $Y=-0.24 $X2=5.335 $Y2=0.995
cc_12 VNB N_A_c_99_n 0.0200652f $X=-0.19 $Y=-0.24 $X2=5.855 $Y2=0.995
cc_13 VNB N_A_c_100_n 0.229146f $X=-0.19 $Y=-0.24 $X2=5.83 $Y2=1.202
cc_14 VNB N_VPWR_c_324_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.202
cc_15 VNB N_Y_c_426_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.56
cc_16 VNB N_Y_c_427_n 0.0163883f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.41
cc_17 VNB N_Y_c_428_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=4.865 $Y2=0.56
cc_18 VNB N_Y_c_429_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=5.83 $Y2=1.985
cc_19 VNB N_Y_c_430_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=5.085 $Y2=1.105
cc_20 VNB N_Y_c_431_n 0.00247508f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.202
cc_21 VNB N_Y_c_432_n 0.0109332f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.202
cc_22 VNB N_Y_c_433_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=5.595 $Y2=1.16
cc_23 VNB N_Y_c_434_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0.895 $Y2=1.2
cc_24 VNB N_Y_c_435_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.19
cc_25 VNB N_Y_c_436_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=1.19
cc_26 VNB N_Y_c_437_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB Y 0.0249933f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.19
cc_28 VNB Y 0.0221428f $X=-0.19 $Y=-0.24 $X2=3.005 $Y2=1.2
cc_29 VNB N_VGND_c_683_n 0.0145634f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=1.41
cc_30 VNB N_VGND_c_684_n 0.0171601f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=1.985
cc_31 VNB N_VGND_c_685_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.54 $Y2=1.41
cc_32 VNB N_VGND_c_686_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.985 $Y2=0.56
cc_33 VNB N_VGND_c_687_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.01 $Y2=1.985
cc_34 VNB N_VGND_c_688_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=1.41
cc_35 VNB N_VGND_c_689_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=3.925 $Y2=0.56
cc_36 VNB N_VGND_c_690_n 0.0137227f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.41
cc_37 VNB N_VGND_c_691_n 0.0170519f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=1.985
cc_38 VNB N_VGND_c_692_n 0.0191635f $X=-0.19 $Y=-0.24 $X2=4.395 $Y2=0.56
cc_39 VNB N_VGND_c_693_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=1.41
cc_40 VNB N_VGND_c_694_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=4.42 $Y2=1.985
cc_41 VNB N_VGND_c_695_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=4.865 $Y2=0.995
cc_42 VNB N_VGND_c_696_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=4.865 $Y2=0.56
cc_43 VNB N_VGND_c_697_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=4.89 $Y2=1.41
cc_44 VNB N_VGND_c_698_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=4.89 $Y2=1.985
cc_45 VNB N_VGND_c_699_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=5.335 $Y2=0.995
cc_46 VNB N_VGND_c_700_n 0.0191455f $X=-0.19 $Y=-0.24 $X2=5.335 $Y2=0.56
cc_47 VNB N_VGND_c_701_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=5.36 $Y2=1.41
cc_48 VNB N_VGND_c_702_n 0.0187013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_703_n 0.31707f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.202
cc_50 VPB N_A_c_101_n 0.0191437f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.41
cc_51 VPB N_A_c_102_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.13 $Y2=1.41
cc_52 VPB N_A_c_103_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.6 $Y2=1.41
cc_53 VPB N_A_c_104_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=1.41
cc_54 VPB N_A_c_105_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.41
cc_55 VPB N_A_c_106_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.41
cc_56 VPB N_A_c_107_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.41
cc_57 VPB N_A_c_108_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.41
cc_58 VPB N_A_c_109_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.42 $Y2=1.41
cc_59 VPB N_A_c_110_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.89 $Y2=1.41
cc_60 VPB N_A_c_111_n 0.0162608f $X=-0.19 $Y=1.305 $X2=5.36 $Y2=1.41
cc_61 VPB N_A_c_112_n 0.0191402f $X=-0.19 $Y=1.305 $X2=5.83 $Y2=1.41
cc_62 VPB N_A_c_100_n 0.15021f $X=-0.19 $Y=1.305 $X2=5.83 $Y2=1.202
cc_63 VPB N_VPWR_c_325_n 0.0152107f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=1.41
cc_64 VPB N_VPWR_c_326_n 0.0300039f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=1.985
cc_65 VPB N_VPWR_c_327_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.54 $Y2=1.41
cc_66 VPB N_VPWR_c_328_n 0.00469739f $X=-0.19 $Y=1.305 $X2=2.985 $Y2=0.56
cc_67 VPB N_VPWR_c_329_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.01 $Y2=1.985
cc_68 VPB N_VPWR_c_330_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.41
cc_69 VPB N_VPWR_c_331_n 0.00469739f $X=-0.19 $Y=1.305 $X2=3.925 $Y2=0.56
cc_70 VPB N_VPWR_c_332_n 0.0137786f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.41
cc_71 VPB N_VPWR_c_333_n 0.0295331f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.985
cc_72 VPB N_VPWR_c_334_n 0.0206409f $X=-0.19 $Y=1.305 $X2=4.395 $Y2=0.56
cc_73 VPB N_VPWR_c_335_n 0.00324069f $X=-0.19 $Y=1.305 $X2=4.42 $Y2=1.41
cc_74 VPB N_VPWR_c_336_n 0.0206409f $X=-0.19 $Y=1.305 $X2=4.42 $Y2=1.985
cc_75 VPB N_VPWR_c_337_n 0.00324069f $X=-0.19 $Y=1.305 $X2=4.865 $Y2=0.995
cc_76 VPB N_VPWR_c_338_n 0.0206409f $X=-0.19 $Y=1.305 $X2=4.865 $Y2=0.56
cc_77 VPB N_VPWR_c_339_n 0.00324069f $X=-0.19 $Y=1.305 $X2=4.89 $Y2=1.41
cc_78 VPB N_VPWR_c_340_n 0.0206409f $X=-0.19 $Y=1.305 $X2=4.89 $Y2=1.985
cc_79 VPB N_VPWR_c_341_n 0.00324069f $X=-0.19 $Y=1.305 $X2=5.335 $Y2=0.995
cc_80 VPB N_VPWR_c_342_n 0.0206409f $X=-0.19 $Y=1.305 $X2=5.335 $Y2=0.56
cc_81 VPB N_VPWR_c_343_n 0.00324069f $X=-0.19 $Y=1.305 $X2=5.36 $Y2=1.41
cc_82 VPB N_VPWR_c_344_n 0.0204049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_324_n 0.0548481f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.202
cc_84 VPB N_Y_c_440_n 0.0150327f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=1.985
cc_85 VPB N_Y_c_441_n 0.0116155f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.202
cc_86 VPB Y 0.0117999f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.19
cc_87 VPB Y 0.0103262f $X=-0.19 $Y=1.305 $X2=3.005 $Y2=1.2
cc_88 N_A_c_101_n N_VPWR_c_326_n 0.00674649f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_c_102_n N_VPWR_c_327_n 0.0052072f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_103_n N_VPWR_c_327_n 0.004751f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_104_n N_VPWR_c_328_n 0.0052072f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_105_n N_VPWR_c_328_n 0.004751f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_c_106_n N_VPWR_c_329_n 0.0052072f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_107_n N_VPWR_c_329_n 0.004751f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_c_108_n N_VPWR_c_330_n 0.0052072f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_c_109_n N_VPWR_c_330_n 0.004751f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_110_n N_VPWR_c_331_n 0.0052072f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_111_n N_VPWR_c_331_n 0.004751f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_c_112_n N_VPWR_c_333_n 0.0045102f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_101_n N_VPWR_c_334_n 0.00597712f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_102_n N_VPWR_c_334_n 0.00673617f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_103_n N_VPWR_c_336_n 0.00597712f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_104_n N_VPWR_c_336_n 0.00673617f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_105_n N_VPWR_c_338_n 0.00597712f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_106_n N_VPWR_c_338_n 0.00673617f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_c_107_n N_VPWR_c_340_n 0.00597712f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_c_108_n N_VPWR_c_340_n 0.00673617f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_c_109_n N_VPWR_c_342_n 0.00597712f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_c_110_n N_VPWR_c_342_n 0.00673617f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_111_n N_VPWR_c_344_n 0.00597712f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_112_n N_VPWR_c_344_n 0.00673617f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_101_n N_VPWR_c_324_n 0.0110272f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_102_n N_VPWR_c_324_n 0.0118438f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_103_n N_VPWR_c_324_n 0.00999457f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_104_n N_VPWR_c_324_n 0.0118438f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_c_105_n N_VPWR_c_324_n 0.00999457f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_106_n N_VPWR_c_324_n 0.0118438f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_107_n N_VPWR_c_324_n 0.00999457f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_c_108_n N_VPWR_c_324_n 0.0118438f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_109_n N_VPWR_c_324_n 0.00999457f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_110_n N_VPWR_c_324_n 0.0118438f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A_c_111_n N_VPWR_c_324_n 0.00999457f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_112_n N_VPWR_c_324_n 0.0128334f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_88_n N_Y_c_444_n 0.0110698f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_c_89_n N_Y_c_444_n 0.00685623f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_90_n N_Y_c_444_n 5.4298e-19 $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_101_n N_Y_c_447_n 0.0181026f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_c_102_n N_Y_c_447_n 0.0107003f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_103_n N_Y_c_447_n 6.25403e-19 $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_89_n N_Y_c_426_n 0.00923615f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_131 N_A_c_90_n N_Y_c_426_n 0.00923615f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_c_100_n N_Y_c_426_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_133 N_A_c_88_n N_Y_c_427_n 0.0138364f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_89_n N_Y_c_427_n 0.00133134f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A_c_161_p N_Y_c_427_n 0.068576f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A_c_100_n N_Y_c_427_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_c_102_n N_Y_c_457_n 0.0137916f $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_103_n N_Y_c_457_n 0.0101048f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_100_n N_Y_c_457_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_140 N_A_c_101_n N_Y_c_440_n 0.01557f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_102_n N_Y_c_440_n 6.17393e-19 $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_161_p N_Y_c_440_n 0.0586497f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_c_100_n N_Y_c_440_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_144 N_A_c_89_n N_Y_c_464_n 5.22028e-19 $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_90_n N_Y_c_464_n 0.00641183f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_91_n N_Y_c_464_n 0.00674948f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_c_92_n N_Y_c_464_n 5.42233e-19 $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_c_102_n N_Y_c_468_n 6.48386e-19 $X=1.13 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_103_n N_Y_c_468_n 0.0130707f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_104_n N_Y_c_468_n 0.0106251f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_105_n N_Y_c_468_n 6.24674e-19 $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_91_n N_Y_c_428_n 0.00923615f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_92_n N_Y_c_428_n 0.00923615f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_161_p N_Y_c_428_n 0.0405926f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_c_100_n N_Y_c_428_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_c_104_n N_Y_c_476_n 0.0137916f $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_c_105_n N_Y_c_476_n 0.0101048f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_161_p N_Y_c_476_n 0.0356113f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_c_100_n N_Y_c_476_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_160 N_A_c_91_n N_Y_c_480_n 5.22028e-19 $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_92_n N_Y_c_480_n 0.00641183f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_93_n N_Y_c_480_n 0.00674948f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_94_n N_Y_c_480_n 5.42233e-19 $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_104_n N_Y_c_484_n 6.48386e-19 $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_c_105_n N_Y_c_484_n 0.0130707f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_c_106_n N_Y_c_484_n 0.0106251f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_c_107_n N_Y_c_484_n 6.24674e-19 $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_93_n N_Y_c_429_n 0.00923615f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_169 N_A_c_94_n N_Y_c_429_n 0.00923615f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_161_p N_Y_c_429_n 0.0405926f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_100_n N_Y_c_429_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_c_106_n N_Y_c_492_n 0.0137916f $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_c_107_n N_Y_c_492_n 0.0101048f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_161_p N_Y_c_492_n 0.0356113f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_c_100_n N_Y_c_492_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_176 N_A_c_93_n N_Y_c_496_n 5.22028e-19 $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_94_n N_Y_c_496_n 0.00641183f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_95_n N_Y_c_496_n 0.00674948f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_96_n N_Y_c_496_n 5.42233e-19 $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_106_n N_Y_c_500_n 6.48386e-19 $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_c_107_n N_Y_c_500_n 0.0130707f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_c_108_n N_Y_c_500_n 0.0106251f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_c_109_n N_Y_c_500_n 6.24674e-19 $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_c_95_n N_Y_c_430_n 0.00923615f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A_c_96_n N_Y_c_430_n 0.00923615f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_c_161_p N_Y_c_430_n 0.0405926f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_c_100_n N_Y_c_430_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_188 N_A_c_108_n N_Y_c_508_n 0.0137916f $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_109_n N_Y_c_508_n 0.0101048f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_161_p N_Y_c_508_n 0.0356113f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A_c_100_n N_Y_c_508_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_192 N_A_c_95_n N_Y_c_512_n 5.22028e-19 $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_96_n N_Y_c_512_n 0.00641183f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_97_n N_Y_c_512_n 0.00674948f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_98_n N_Y_c_512_n 5.42233e-19 $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_108_n N_Y_c_516_n 6.48386e-19 $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_109_n N_Y_c_516_n 0.0130707f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_110_n N_Y_c_516_n 0.0106251f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_111_n N_Y_c_516_n 6.24674e-19 $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_97_n N_Y_c_431_n 0.00923615f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_98_n N_Y_c_431_n 0.00923615f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_161_p N_Y_c_431_n 0.0405926f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_c_100_n N_Y_c_431_n 0.00346f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_204 N_A_c_110_n N_Y_c_524_n 0.0137916f $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_111_n N_Y_c_524_n 0.0101048f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_161_p N_Y_c_524_n 0.0356113f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_c_100_n N_Y_c_524_n 0.00635951f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_208 N_A_c_97_n N_Y_c_528_n 5.22028e-19 $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_c_98_n N_Y_c_528_n 0.00641183f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_110_n N_Y_c_530_n 6.48386e-19 $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_111_n N_Y_c_530_n 0.0130707f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_112_n N_Y_c_530_n 0.0152835f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_c_99_n N_Y_c_432_n 0.0143569f $X=5.855 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_161_p N_Y_c_432_n 0.00285544f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_c_112_n N_Y_c_441_n 0.0168658f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_161_p N_Y_c_441_n 0.00276009f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_217 N_A_c_90_n N_Y_c_433_n 0.00119366f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_c_91_n N_Y_c_433_n 0.00119366f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_161_p N_Y_c_433_n 0.031064f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_c_100_n N_Y_c_433_n 0.00358305f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_221 N_A_c_103_n N_Y_c_541_n 0.00210477f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_104_n N_Y_c_541_n 5.79575e-19 $X=2.07 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_161_p N_Y_c_541_n 0.0253353f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_c_100_n N_Y_c_541_n 0.00651614f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_225 N_A_c_92_n N_Y_c_434_n 0.00119366f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_c_93_n N_Y_c_434_n 0.00119366f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_227 N_A_c_161_p N_Y_c_434_n 0.031064f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A_c_100_n N_Y_c_434_n 0.00358305f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_229 N_A_c_105_n N_Y_c_549_n 0.00210477f $X=2.54 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_c_106_n N_Y_c_549_n 5.79575e-19 $X=3.01 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_c_161_p N_Y_c_549_n 0.0253353f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_232 N_A_c_100_n N_Y_c_549_n 0.00651614f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_233 N_A_c_94_n N_Y_c_435_n 0.00119366f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_c_95_n N_Y_c_435_n 0.00119366f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_c_161_p N_Y_c_435_n 0.031064f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_c_100_n N_Y_c_435_n 0.00358305f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_237 N_A_c_107_n N_Y_c_557_n 0.00210477f $X=3.48 $Y=1.41 $X2=0 $Y2=0
cc_238 N_A_c_108_n N_Y_c_557_n 5.79575e-19 $X=3.95 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_161_p N_Y_c_557_n 0.0253353f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_c_100_n N_Y_c_557_n 0.00651614f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_c_96_n N_Y_c_436_n 0.00119366f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_97_n N_Y_c_436_n 0.00119366f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_161_p N_Y_c_436_n 0.031064f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_c_100_n N_Y_c_436_n 0.00358305f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_245 N_A_c_109_n N_Y_c_565_n 0.00210477f $X=4.42 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_110_n N_Y_c_565_n 5.79575e-19 $X=4.89 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_161_p N_Y_c_565_n 0.0253353f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_100_n N_Y_c_565_n 0.00651614f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_249 N_A_c_98_n N_Y_c_437_n 0.00122295f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_161_p N_Y_c_437_n 0.0311977f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_251 N_A_c_100_n N_Y_c_437_n 0.00486271f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_252 N_A_c_111_n N_Y_c_572_n 0.00210477f $X=5.36 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_112_n N_Y_c_572_n 5.79575e-19 $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_161_p N_Y_c_572_n 0.0253353f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_c_100_n N_Y_c_572_n 0.00631893f $X=5.83 $Y=1.202 $X2=0 $Y2=0
cc_256 N_A_c_88_n Y 0.0196788f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_c_101_n Y 0.00371943f $X=0.66 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_161_p Y 0.0212121f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_c_112_n Y 0.00341357f $X=5.83 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_99_n Y 0.0195682f $X=5.855 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_c_161_p Y 0.0209006f $X=5.595 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_c_88_n N_VGND_c_684_n 0.00450113f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_c_89_n N_VGND_c_685_n 0.00376026f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_c_90_n N_VGND_c_685_n 0.00276126f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_c_91_n N_VGND_c_686_n 0.00376026f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_c_92_n N_VGND_c_686_n 0.00276126f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_93_n N_VGND_c_687_n 0.00376026f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_c_94_n N_VGND_c_687_n 0.00276126f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_c_95_n N_VGND_c_688_n 0.00376026f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_c_96_n N_VGND_c_688_n 0.00276126f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_c_97_n N_VGND_c_689_n 0.00376026f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_c_98_n N_VGND_c_689_n 0.00276126f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_c_99_n N_VGND_c_691_n 0.0046798f $X=5.855 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_c_88_n N_VGND_c_692_n 0.00421248f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_275 N_A_c_89_n N_VGND_c_692_n 0.00421248f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_276 N_A_c_90_n N_VGND_c_694_n 0.00422241f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A_c_91_n N_VGND_c_694_n 0.00422241f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_c_92_n N_VGND_c_696_n 0.00422241f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_93_n N_VGND_c_696_n 0.00422241f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A_c_94_n N_VGND_c_698_n 0.00422241f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A_c_95_n N_VGND_c_698_n 0.00422241f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_c_96_n N_VGND_c_700_n 0.00422241f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_283 N_A_c_97_n N_VGND_c_700_n 0.00422241f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_284 N_A_c_98_n N_VGND_c_702_n 0.00422241f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A_c_99_n N_VGND_c_702_n 0.00436487f $X=5.855 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_c_88_n N_VGND_c_703_n 0.00691717f $X=0.635 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_c_89_n N_VGND_c_703_n 0.00608774f $X=1.105 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_c_90_n N_VGND_c_703_n 0.0059505f $X=1.575 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_c_91_n N_VGND_c_703_n 0.00607326f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_c_92_n N_VGND_c_703_n 0.0059505f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_291 N_A_c_93_n N_VGND_c_703_n 0.00607326f $X=2.985 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A_c_94_n N_VGND_c_703_n 0.0059505f $X=3.455 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_c_95_n N_VGND_c_703_n 0.00607326f $X=3.925 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_c_96_n N_VGND_c_703_n 0.0059505f $X=4.395 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_c_97_n N_VGND_c_703_n 0.00607326f $X=4.865 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_c_98_n N_VGND_c_703_n 0.00606584f $X=5.335 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_c_99_n N_VGND_c_703_n 0.00710196f $X=5.855 $Y=0.995 $X2=0 $Y2=0
cc_298 N_VPWR_c_324_n N_Y_M1002_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_299 N_VPWR_c_324_n N_Y_M1004_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_300 N_VPWR_c_324_n N_Y_M1008_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_324_n N_Y_M1010_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_324_n N_Y_M1017_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_303 N_VPWR_c_324_n N_Y_M1019_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_304 N_VPWR_c_326_n N_Y_c_447_n 0.048465f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_305 N_VPWR_c_327_n N_Y_c_447_n 0.0385613f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_306 N_VPWR_c_334_n N_Y_c_447_n 0.0223557f $X=1.28 $Y=2.72 $X2=0 $Y2=0
cc_307 N_VPWR_c_324_n N_Y_c_447_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_308 N_VPWR_M1003_s N_Y_c_457_n 0.00325884f $X=1.22 $Y=1.485 $X2=0 $Y2=0
cc_309 N_VPWR_c_327_n N_Y_c_457_n 0.0136682f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_310 N_VPWR_M1002_s N_Y_c_440_n 0.0036766f $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_311 N_VPWR_c_326_n N_Y_c_440_n 0.0207202f $X=0.425 $Y=2 $X2=0 $Y2=0
cc_312 N_VPWR_c_327_n N_Y_c_468_n 0.0470327f $X=1.365 $Y=2 $X2=0 $Y2=0
cc_313 N_VPWR_c_328_n N_Y_c_468_n 0.0385613f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_314 N_VPWR_c_336_n N_Y_c_468_n 0.0223557f $X=2.22 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_324_n N_Y_c_468_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_M1006_s N_Y_c_476_n 0.00325884f $X=2.16 $Y=1.485 $X2=0 $Y2=0
cc_317 N_VPWR_c_328_n N_Y_c_476_n 0.0136682f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_318 N_VPWR_c_328_n N_Y_c_484_n 0.0470327f $X=2.305 $Y=2 $X2=0 $Y2=0
cc_319 N_VPWR_c_329_n N_Y_c_484_n 0.0385613f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_320 N_VPWR_c_338_n N_Y_c_484_n 0.0223557f $X=3.16 $Y=2.72 $X2=0 $Y2=0
cc_321 N_VPWR_c_324_n N_Y_c_484_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_M1009_s N_Y_c_492_n 0.00325884f $X=3.1 $Y=1.485 $X2=0 $Y2=0
cc_323 N_VPWR_c_329_n N_Y_c_492_n 0.0136682f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_324 N_VPWR_c_329_n N_Y_c_500_n 0.0470327f $X=3.245 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_c_330_n N_Y_c_500_n 0.0385613f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_326 N_VPWR_c_340_n N_Y_c_500_n 0.0223557f $X=4.1 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_324_n N_Y_c_500_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_M1015_s N_Y_c_508_n 0.00325884f $X=4.04 $Y=1.485 $X2=0 $Y2=0
cc_329 N_VPWR_c_330_n N_Y_c_508_n 0.0136682f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_330 N_VPWR_c_330_n N_Y_c_516_n 0.0470327f $X=4.185 $Y=2 $X2=0 $Y2=0
cc_331 N_VPWR_c_331_n N_Y_c_516_n 0.0385613f $X=5.125 $Y=2 $X2=0 $Y2=0
cc_332 N_VPWR_c_342_n N_Y_c_516_n 0.0223557f $X=5.04 $Y=2.72 $X2=0 $Y2=0
cc_333 N_VPWR_c_324_n N_Y_c_516_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_334 N_VPWR_M1018_s N_Y_c_524_n 0.00325884f $X=4.98 $Y=1.485 $X2=0 $Y2=0
cc_335 N_VPWR_c_331_n N_Y_c_524_n 0.0136682f $X=5.125 $Y=2 $X2=0 $Y2=0
cc_336 N_VPWR_c_331_n N_Y_c_530_n 0.0470327f $X=5.125 $Y=2 $X2=0 $Y2=0
cc_337 N_VPWR_c_344_n N_Y_c_530_n 0.0223557f $X=5.975 $Y=2.72 $X2=0 $Y2=0
cc_338 N_VPWR_c_324_n N_Y_c_530_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_339 N_VPWR_M1021_s N_Y_c_441_n 0.00340873f $X=5.92 $Y=1.485 $X2=0 $Y2=0
cc_340 N_VPWR_c_333_n N_Y_c_441_n 0.0228233f $X=6.065 $Y=2 $X2=0 $Y2=0
cc_341 N_VPWR_M1002_s Y 7.90669e-19 $X=0.3 $Y=1.485 $X2=0 $Y2=0
cc_342 N_Y_c_427_n N_VGND_M1000_s 0.00285834f $X=1.06 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_343 N_Y_c_426_n N_VGND_M1001_s 0.0025045f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_344 N_Y_c_428_n N_VGND_M1007_s 0.0025045f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_345 N_Y_c_429_n N_VGND_M1012_s 0.0025045f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_346 N_Y_c_430_n N_VGND_M1014_s 0.0025045f $X=4.44 $Y=0.81 $X2=0 $Y2=0
cc_347 N_Y_c_431_n N_VGND_M1020_s 0.0025045f $X=5.38 $Y=0.81 $X2=0 $Y2=0
cc_348 N_Y_c_432_n N_VGND_M1023_s 0.00314359f $X=5.97 $Y=0.81 $X2=0 $Y2=0
cc_349 N_Y_c_427_n N_VGND_c_683_n 0.00267039f $X=1.06 $Y=0.81 $X2=0 $Y2=0
cc_350 N_Y_c_427_n N_VGND_c_684_n 0.0195556f $X=1.06 $Y=0.81 $X2=0 $Y2=0
cc_351 N_Y_c_444_n N_VGND_c_685_n 0.0177507f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_352 N_Y_c_426_n N_VGND_c_685_n 0.0127393f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_353 N_Y_c_464_n N_VGND_c_686_n 0.0177507f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_354 N_Y_c_428_n N_VGND_c_686_n 0.0127393f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_355 N_Y_c_480_n N_VGND_c_687_n 0.0177507f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_356 N_Y_c_429_n N_VGND_c_687_n 0.0127393f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_357 N_Y_c_496_n N_VGND_c_688_n 0.0177507f $X=3.715 $Y=0.38 $X2=0 $Y2=0
cc_358 N_Y_c_430_n N_VGND_c_688_n 0.0127393f $X=4.44 $Y=0.81 $X2=0 $Y2=0
cc_359 N_Y_c_512_n N_VGND_c_689_n 0.0177507f $X=4.655 $Y=0.38 $X2=0 $Y2=0
cc_360 N_Y_c_431_n N_VGND_c_689_n 0.0127393f $X=5.38 $Y=0.81 $X2=0 $Y2=0
cc_361 N_Y_c_432_n N_VGND_c_690_n 0.00156502f $X=5.97 $Y=0.81 $X2=0 $Y2=0
cc_362 N_Y_c_432_n N_VGND_c_691_n 0.0209716f $X=5.97 $Y=0.81 $X2=0 $Y2=0
cc_363 N_Y_c_444_n N_VGND_c_692_n 0.02191f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_364 N_Y_c_427_n N_VGND_c_692_n 0.00480429f $X=1.06 $Y=0.81 $X2=0 $Y2=0
cc_365 N_Y_c_426_n N_VGND_c_694_n 0.00203746f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_366 N_Y_c_464_n N_VGND_c_694_n 0.0223596f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_367 N_Y_c_428_n N_VGND_c_694_n 0.00273345f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_368 N_Y_c_428_n N_VGND_c_696_n 0.00203746f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_369 N_Y_c_480_n N_VGND_c_696_n 0.0223596f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_370 N_Y_c_429_n N_VGND_c_696_n 0.00273345f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_371 N_Y_c_429_n N_VGND_c_698_n 0.00203746f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_372 N_Y_c_496_n N_VGND_c_698_n 0.0223596f $X=3.715 $Y=0.38 $X2=0 $Y2=0
cc_373 N_Y_c_430_n N_VGND_c_698_n 0.00273345f $X=4.44 $Y=0.81 $X2=0 $Y2=0
cc_374 N_Y_c_430_n N_VGND_c_700_n 0.00203746f $X=4.44 $Y=0.81 $X2=0 $Y2=0
cc_375 N_Y_c_512_n N_VGND_c_700_n 0.0223596f $X=4.655 $Y=0.38 $X2=0 $Y2=0
cc_376 N_Y_c_431_n N_VGND_c_700_n 0.00273345f $X=5.38 $Y=0.81 $X2=0 $Y2=0
cc_377 N_Y_c_431_n N_VGND_c_702_n 0.00203746f $X=5.38 $Y=0.81 $X2=0 $Y2=0
cc_378 N_Y_c_528_n N_VGND_c_702_n 0.0231806f $X=5.595 $Y=0.38 $X2=0 $Y2=0
cc_379 N_Y_c_432_n N_VGND_c_702_n 0.00245083f $X=5.97 $Y=0.81 $X2=0 $Y2=0
cc_380 N_Y_M1000_d N_VGND_c_703_n 0.0025535f $X=0.71 $Y=0.235 $X2=0 $Y2=0
cc_381 N_Y_M1005_d N_VGND_c_703_n 0.0025535f $X=1.65 $Y=0.235 $X2=0 $Y2=0
cc_382 N_Y_M1011_d N_VGND_c_703_n 0.0025535f $X=2.59 $Y=0.235 $X2=0 $Y2=0
cc_383 N_Y_M1013_d N_VGND_c_703_n 0.0025535f $X=3.53 $Y=0.235 $X2=0 $Y2=0
cc_384 N_Y_M1016_d N_VGND_c_703_n 0.0025535f $X=4.47 $Y=0.235 $X2=0 $Y2=0
cc_385 N_Y_M1022_d N_VGND_c_703_n 0.0030386f $X=5.41 $Y=0.235 $X2=0 $Y2=0
cc_386 N_Y_c_444_n N_VGND_c_703_n 0.0140045f $X=0.895 $Y=0.38 $X2=0 $Y2=0
cc_387 N_Y_c_426_n N_VGND_c_703_n 0.00455756f $X=1.62 $Y=0.81 $X2=0 $Y2=0
cc_388 N_Y_c_427_n N_VGND_c_703_n 0.0148078f $X=1.06 $Y=0.81 $X2=0 $Y2=0
cc_389 N_Y_c_464_n N_VGND_c_703_n 0.0141302f $X=1.835 $Y=0.38 $X2=0 $Y2=0
cc_390 N_Y_c_428_n N_VGND_c_703_n 0.00983903f $X=2.56 $Y=0.81 $X2=0 $Y2=0
cc_391 N_Y_c_480_n N_VGND_c_703_n 0.0141302f $X=2.775 $Y=0.38 $X2=0 $Y2=0
cc_392 N_Y_c_429_n N_VGND_c_703_n 0.00983903f $X=3.5 $Y=0.81 $X2=0 $Y2=0
cc_393 N_Y_c_496_n N_VGND_c_703_n 0.0141302f $X=3.715 $Y=0.38 $X2=0 $Y2=0
cc_394 N_Y_c_430_n N_VGND_c_703_n 0.00983903f $X=4.44 $Y=0.81 $X2=0 $Y2=0
cc_395 N_Y_c_512_n N_VGND_c_703_n 0.0141302f $X=4.655 $Y=0.38 $X2=0 $Y2=0
cc_396 N_Y_c_431_n N_VGND_c_703_n 0.00983903f $X=5.38 $Y=0.81 $X2=0 $Y2=0
cc_397 N_Y_c_528_n N_VGND_c_703_n 0.0143352f $X=5.595 $Y=0.38 $X2=0 $Y2=0
cc_398 N_Y_c_432_n N_VGND_c_703_n 0.00827125f $X=5.97 $Y=0.81 $X2=0 $Y2=0
