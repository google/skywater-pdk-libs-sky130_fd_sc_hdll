* File: sky130_fd_sc_hdll__dfstp_2.pex.spice
* Created: Thu Aug 27 19:04:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%CLK 4 5 7 8 10 13 19 20 24 26
c41 13 0 2.71124e-20 $X=0.52 $Y=0.805
r42 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r43 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r44 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r45 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r46 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r47 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r48 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r49 5 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r51 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r52 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r53 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r54 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_27_47# 1 2 8 9 11 14 16 18 19 21 22 24
+ 25 27 30 34 35 36 39 41 45 46 49 50 51 53 54 68 72 73 75 76 77 82 90 96
c262 73 0 3.46126e-20 $X=2.875 $Y=1.825
c263 50 0 1.75333e-19 $X=6.37 $Y=0.81
c264 46 0 9.81997e-20 $X=2.585 $Y=0.87
c265 36 0 1.76957e-19 $X=0.66 $Y=1.88
c266 22 0 1.37207e-19 $X=5.54 $Y=1.99
c267 19 0 2.53929e-20 $X=2.96 $Y=1.99
r268 93 104 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.605 $Y=1.81
+ $X2=5.415 $Y2=1.81
r269 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.605
+ $Y=1.74 $X2=5.605 $Y2=1.74
r270 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.74 $X2=2.965 $Y2=1.74
r271 81 82 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r272 76 93 6.87748 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=5.79 $Y=1.81
+ $X2=5.605 $Y2=1.81
r273 75 77 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.79 $Y=1.825
+ $X2=5.645 $Y2=1.825
r274 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.79 $Y=1.825
+ $X2=5.79 $Y2=1.825
r275 73 77 3.42821 $w=1.4e-07 $l=2.77e-06 $layer=MET1_cond $X=2.875 $Y=1.87
+ $X2=5.645 $Y2=1.87
r276 71 90 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.73 $Y=1.765
+ $X2=2.965 $Y2=1.765
r277 71 99 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.73 $Y=1.765
+ $X2=2.635 $Y2=1.765
r278 70 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.73 $Y=1.825
+ $X2=2.875 $Y2=1.825
r279 70 72 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.73 $Y=1.825
+ $X2=2.585 $Y2=1.825
r280 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.73 $Y=1.825
+ $X2=2.73 $Y2=1.825
r281 68 72 2.09158 $w=1.4e-07 $l=1.69e-06 $layer=MET1_cond $X=0.895 $Y=1.87
+ $X2=2.585 $Y2=1.87
r282 65 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.75 $Y=1.825
+ $X2=0.895 $Y2=1.825
r283 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.75 $Y=1.825
+ $X2=0.75 $Y2=1.825
r284 58 96 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.535 $Y=0.93
+ $X2=6.645 $Y2=0.93
r285 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.535
+ $Y=0.93 $X2=6.535 $Y2=0.93
r286 54 57 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.56 $Y=0.81
+ $X2=6.56 $Y2=0.93
r287 50 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.37 $Y=0.81
+ $X2=6.56 $Y2=0.81
r288 50 51 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.37 $Y=0.81
+ $X2=5.5 $Y2=0.81
r289 49 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.415 $Y=1.655
+ $X2=5.415 $Y2=1.81
r290 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=0.895
+ $X2=5.5 $Y2=0.81
r291 48 49 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.415 $Y=0.895
+ $X2=5.415 $Y2=1.655
r292 46 84 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.585 $Y=0.87
+ $X2=2.455 $Y2=0.87
r293 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.87 $X2=2.585 $Y2=0.87
r294 43 99 2.7393 $w=2.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.635 $Y=1.575
+ $X2=2.635 $Y2=1.765
r295 43 45 30.0916 $w=2.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.635 $Y=1.575
+ $X2=2.635 $Y2=0.87
r296 42 81 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r297 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r298 39 66 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.88
r299 39 41 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.235
r300 38 41 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=1.235
r301 37 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r302 36 66 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.775 $Y2=1.88
r303 36 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r304 34 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.775 $Y2=0.805
r305 34 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r306 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r307 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r308 25 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=0.765
+ $X2=6.645 $Y2=0.93
r309 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.645 $Y=0.765
+ $X2=6.645 $Y2=0.445
r310 22 92 46.5577 $w=3.26e-07 $l=2.91548e-07 $layer=POLY_cond $X=5.54 $Y=1.99
+ $X2=5.63 $Y2=1.74
r311 22 24 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.54 $Y=1.99
+ $X2=5.54 $Y2=2.275
r312 19 89 46.5577 $w=3.26e-07 $l=2.64575e-07 $layer=POLY_cond $X=2.96 $Y=1.99
+ $X2=2.99 $Y2=1.74
r313 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.96 $Y=1.99
+ $X2=2.96 $Y2=2.275
r314 16 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=0.705
+ $X2=2.455 $Y2=0.87
r315 16 18 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.455 $Y=0.705
+ $X2=2.455 $Y2=0.415
r316 12 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r317 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r318 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r319 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r320 7 81 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r321 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r322 2 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r323 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%D 1 3 6 8 9 14
c38 1 0 1.46624e-19 $X=1.955 $Y=1.57
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.17 $X2=1.955 $Y2=1.17
r40 8 9 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.1 $Y=1.19 $X2=2.1
+ $Y2=1.53
r41 8 14 0.520034 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=2.1 $Y=1.19 $X2=2.1
+ $Y2=1.17
r42 4 13 38.9026 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.005
+ $X2=1.98 $Y2=1.17
r43 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.98 $Y=1.005 $X2=1.98
+ $Y2=0.555
r44 1 13 76.7755 $w=2.7e-07 $l=4.12311e-07 $layer=POLY_cond $X=1.955 $Y=1.57
+ $X2=1.98 $Y2=1.17
r45 1 3 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=1.955 $Y=1.57
+ $X2=1.955 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_211_363# 1 2 8 9 11 12 13 16 19 21 24 26
+ 28 29 30 31 34 36 41 43 44 49 50 51 58 63
c199 51 0 1.51904e-19 $X=5.665 $Y=1.195
c200 50 0 4.09811e-20 $X=5.81 $Y=1.195
c201 49 0 2.54518e-19 $X=5.81 $Y=1.195
c202 36 0 2.53929e-20 $X=3.385 $Y=1.19
c203 34 0 9.81997e-20 $X=3.277 $Y=1.12
c204 30 0 1.75333e-19 $X=5.97 $Y=1.125
c205 21 0 1.7977e-19 $X=6.13 $Y=1.89
c206 8 0 4.36039e-20 $X=2.49 $Y=1.89
r207 58 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=0.93
+ $X2=3.165 $Y2=1.095
r208 58 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=0.93
+ $X2=3.165 $Y2=0.765
r209 50 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.815
+ $Y=1.26 $X2=5.815 $Y2=1.26
r210 49 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.81 $Y=1.195
+ $X2=5.665 $Y2=1.195
r211 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.81 $Y=1.195
+ $X2=5.81 $Y2=1.195
r212 46 47 0.0440827 $w=2.9e-07 $l=7e-08 $layer=MET1_cond $X=3.24 $Y=0.85
+ $X2=3.24 $Y2=0.92
r213 44 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=0.93 $X2=3.165 $Y2=0.93
r214 43 46 0.0220415 $w=2.9e-07 $l=4.5e-08 $layer=MET1_cond $X=3.24 $Y=0.805
+ $X2=3.24 $Y2=0.85
r215 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.24 $Y=0.805
+ $X2=3.24 $Y2=0.805
r216 39 67 59.1587 $w=2.23e-07 $l=1.155e-06 $layer=LI1_cond $X=1.227 $Y=0.805
+ $X2=1.227 $Y2=1.96
r217 39 63 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.227 $Y=0.805
+ $X2=1.227 $Y2=0.51
r218 38 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.25 $Y=0.805
+ $X2=1.395 $Y2=0.805
r219 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.25 $Y=0.805
+ $X2=1.25 $Y2=0.805
r220 36 51 2.82178 $w=1.4e-07 $l=2.28e-06 $layer=MET1_cond $X=3.385 $Y=1.19
+ $X2=5.665 $Y2=1.19
r221 34 36 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.277 $Y=1.12
+ $X2=3.385 $Y2=1.19
r222 34 47 0.142799 $w=2.15e-07 $l=2e-07 $layer=MET1_cond $X=3.277 $Y=1.12
+ $X2=3.277 $Y2=0.92
r223 31 46 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=3.095 $Y=0.85
+ $X2=3.24 $Y2=0.85
r224 31 41 2.10396 $w=1.4e-07 $l=1.7e-06 $layer=MET1_cond $X=3.095 $Y=0.85
+ $X2=1.395 $Y2=0.85
r225 29 54 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.97 $Y=1.26
+ $X2=5.815 $Y2=1.26
r226 29 30 0.63749 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.97 $Y=1.26
+ $X2=5.97 $Y2=1.125
r227 26 28 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.13 $Y=1.99
+ $X2=6.13 $Y2=2.275
r228 22 30 28.793 $w=1.75e-07 $l=1.45e-07 $layer=POLY_cond $X=6.115 $Y=1.125
+ $X2=5.97 $Y2=1.125
r229 22 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.115 $Y=1.125
+ $X2=6.115 $Y2=0.445
r230 21 26 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.13 $Y=1.89 $X2=6.13
+ $Y2=1.99
r231 20 30 28.793 $w=1.75e-07 $l=4.02119e-07 $layer=POLY_cond $X=6.13 $Y=1.455
+ $X2=5.97 $Y2=1.125
r232 20 21 144.236 $w=2e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=1.455
+ $X2=6.13 $Y2=1.89
r233 19 61 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.105 $Y=1.245
+ $X2=3.105 $Y2=1.095
r234 16 60 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.105 $Y=0.415
+ $X2=3.105 $Y2=0.765
r235 12 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.03 $Y=1.32
+ $X2=3.105 $Y2=1.245
r236 12 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.03 $Y=1.32
+ $X2=2.59 $Y2=1.32
r237 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.49 $Y=1.99
+ $X2=2.49 $Y2=2.275
r238 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.49 $Y=1.89 $X2=2.49
+ $Y2=1.99
r239 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=2.49 $Y=1.395
+ $X2=2.59 $Y2=1.32
r240 7 8 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=2.49 $Y=1.395 $X2=2.49
+ $Y2=1.89
r241 2 67 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r242 1 63 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_702_21# 1 2 9 11 13 14 18 20 24 27 29 34
+ 36
c108 36 0 2.23858e-19 $X=4.95 $Y=1.065
c109 34 0 2.11834e-19 $X=4.425 $Y=1.96
c110 29 0 1.15651e-19 $X=3.695 $Y=1.74
r111 35 36 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=0.725
+ $X2=4.95 $Y2=1.065
r112 29 32 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=3.76 $Y=1.74
+ $X2=3.76 $Y2=1.96
r113 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.74 $X2=3.695 $Y2=1.74
r114 27 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.025 $Y=1.835
+ $X2=5.025 $Y2=1.065
r115 24 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.875 $Y=0.46
+ $X2=4.875 $Y2=0.725
r116 21 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=1.96
+ $X2=4.425 $Y2=1.96
r117 20 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.94 $Y=1.96
+ $X2=5.025 $Y2=1.835
r118 20 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.94 $Y=1.96
+ $X2=4.51 $Y2=1.96
r119 16 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.085
+ $X2=4.425 $Y2=1.96
r120 16 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.085
+ $X2=4.425 $Y2=2.21
r121 15 32 1.80669 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.91 $Y=1.96
+ $X2=3.76 $Y2=1.96
r122 14 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=1.96
+ $X2=4.425 $Y2=1.96
r123 14 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.34 $Y=1.96
+ $X2=3.91 $Y2=1.96
r124 11 30 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=3.61 $Y=1.99
+ $X2=3.695 $Y2=1.74
r125 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.61 $Y=1.99
+ $X2=3.61 $Y2=2.275
r126 7 30 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=3.585 $Y=1.575
+ $X2=3.695 $Y2=1.74
r127 7 9 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.585 $Y=1.575
+ $X2=3.585 $Y2=0.445
r128 2 18 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=2.065 $X2=4.425 $Y2=2.21
r129 1 24 182 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=1 $X=4.69
+ $Y=0.235 $X2=4.875 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%SET_B 2 3 5 8 12 17 18 20 21 22 23 24 26
+ 29 34 37 38 44
c129 44 0 7.40925e-20 $X=4.365 $Y=0.85
c130 26 0 1.71107e-19 $X=7.59 $Y=0.85
c131 24 0 3.91725e-20 $X=4.51 $Y=0.85
c132 23 0 1.86694e-20 $X=7.445 $Y=0.85
c133 8 0 1.90694e-19 $X=4.255 $Y=0.445
c134 3 0 1.15651e-19 $X=4.19 $Y=1.99
r135 37 40 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=0.98
+ $X2=7.45 $Y2=1.145
r136 37 39 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=0.98
+ $X2=7.45 $Y2=0.815
r137 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.425
+ $Y=0.98 $X2=7.425 $Y2=0.98
r138 34 35 10.074 $w=3.11e-07 $l=6.5e-08 $layer=POLY_cond $X=4.19 $Y=0.98
+ $X2=4.255 $Y2=0.98
r139 33 44 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.075 $Y=0.9
+ $X2=4.365 $Y2=0.9
r140 32 34 17.8232 $w=3.11e-07 $l=1.15e-07 $layer=POLY_cond $X=4.075 $Y=0.98
+ $X2=4.19 $Y2=0.98
r141 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=0.98 $X2=4.075 $Y2=0.98
r142 29 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.365 $Y=0.85
+ $X2=4.365 $Y2=0.85
r143 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0.85
+ $X2=7.59 $Y2=0.85
r144 24 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.51 $Y=0.85
+ $X2=4.365 $Y2=0.85
r145 23 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=0.85
+ $X2=7.59 $Y2=0.85
r146 23 24 3.63242 $w=1.4e-07 $l=2.935e-06 $layer=MET1_cond $X=7.445 $Y=0.85
+ $X2=4.51 $Y2=0.85
r147 21 22 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.52 $Y=1.535
+ $X2=7.52 $Y2=1.685
r148 21 40 129.315 $w=2e-07 $l=3.9e-07 $layer=POLY_cond $X=7.51 $Y=1.535
+ $X2=7.51 $Y2=1.145
r149 18 20 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.53 $Y=1.99
+ $X2=7.53 $Y2=2.275
r150 17 18 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.53 $Y=1.89 $X2=7.53
+ $Y2=1.99
r151 17 22 67.9733 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=7.53 $Y=1.89
+ $X2=7.53 $Y2=1.685
r152 12 39 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.365 $Y=0.445
+ $X2=7.365 $Y2=0.815
r153 6 35 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=0.815
+ $X2=4.255 $Y2=0.98
r154 6 8 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.255 $Y=0.815
+ $X2=4.255 $Y2=0.445
r155 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.19 $Y=1.99
+ $X2=4.19 $Y2=2.275
r156 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.19 $Y=1.89 $X2=4.19
+ $Y2=1.99
r157 1 34 13.1188 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.145
+ $X2=4.19 $Y2=0.98
r158 1 2 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=4.19 $Y=1.145 $X2=4.19
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_506_47# 1 2 7 9 11 13 14 16 17 20 21 23
+ 24 26 27 28 32 37 39 40 45 46 56
c160 56 0 1.34022e-19 $X=5.13 $Y=1.4
c161 46 0 3.91725e-20 $X=4.62 $Y=1.32
c162 45 0 4.36039e-20 $X=3.74 $Y=1.317
c163 24 0 3.31643e-20 $X=5.705 $Y=0.735
c164 17 0 1.50733e-19 $X=5.63 $Y=0.825
r165 55 56 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=4.66 $Y=1.4
+ $X2=5.13 $Y2=1.4
r166 54 55 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.64 $Y=1.4 $X2=4.66
+ $Y2=1.4
r167 50 54 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.635 $Y=1.4
+ $X2=4.64 $Y2=1.4
r168 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.4 $X2=4.635 $Y2=1.4
r169 46 49 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=4.62 $Y=1.32 $X2=4.62
+ $Y2=1.4
r170 40 46 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.47 $Y=1.32 $X2=4.62
+ $Y2=1.32
r171 40 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.47 $Y=1.32
+ $X2=3.74 $Y2=1.32
r172 39 45 6.97143 $w=1.73e-07 $l=1.1e-07 $layer=LI1_cond $X=3.63 $Y=1.317
+ $X2=3.74 $Y2=1.317
r173 39 42 17.4286 $w=1.73e-07 $l=2.75e-07 $layer=LI1_cond $X=3.63 $Y=1.317
+ $X2=3.355 $Y2=1.317
r174 38 39 40.0736 $w=2.18e-07 $l=7.65e-07 $layer=LI1_cond $X=3.63 $Y=0.465
+ $X2=3.63 $Y2=1.23
r175 36 42 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=3.355 $Y=1.405
+ $X2=3.355 $Y2=1.317
r176 36 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.355 $Y=1.405
+ $X2=3.355 $Y2=2.25
r177 32 38 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=3.63 $Y2=0.465
r178 32 34 40.4818 $w=1.98e-07 $l=7.3e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=2.79 $Y2=0.365
r179 28 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.335
+ $X2=3.355 $Y2=2.25
r180 28 30 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.27 $Y=2.335
+ $X2=2.725 $Y2=2.335
r181 24 26 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.705 $Y=0.735
+ $X2=5.705 $Y2=0.445
r182 21 23 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.13 $Y=1.99
+ $X2=5.13 $Y2=2.275
r183 20 21 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.13 $Y=1.89 $X2=5.13
+ $Y2=1.99
r184 19 56 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.565
+ $X2=5.13 $Y2=1.4
r185 19 20 107.763 $w=2e-07 $l=3.25e-07 $layer=POLY_cond $X=5.13 $Y=1.565
+ $X2=5.13 $Y2=1.89
r186 18 27 4.90422 $w=1.8e-07 $l=1e-07 $layer=POLY_cond $X=4.74 $Y=0.825
+ $X2=4.64 $Y2=0.825
r187 17 24 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.63 $Y=0.825
+ $X2=5.705 $Y2=0.735
r188 17 18 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=5.63 $Y=0.825
+ $X2=4.74 $Y2=0.825
r189 14 16 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.66 $Y=1.99
+ $X2=4.66 $Y2=2.275
r190 13 14 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.66 $Y=1.89 $X2=4.66
+ $Y2=1.99
r191 12 55 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.565
+ $X2=4.66 $Y2=1.4
r192 12 13 107.763 $w=2e-07 $l=3.25e-07 $layer=POLY_cond $X=4.66 $Y=1.565
+ $X2=4.66 $Y2=1.89
r193 11 54 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=1.235
+ $X2=4.64 $Y2=1.4
r194 10 27 20.8929 $w=1.75e-07 $l=9e-08 $layer=POLY_cond $X=4.64 $Y=0.915
+ $X2=4.64 $Y2=0.825
r195 10 11 106.105 $w=2e-07 $l=3.2e-07 $layer=POLY_cond $X=4.64 $Y=0.915
+ $X2=4.64 $Y2=1.235
r196 7 27 20.8929 $w=1.75e-07 $l=1.01735e-07 $layer=POLY_cond $X=4.615 $Y=0.735
+ $X2=4.64 $Y2=0.825
r197 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.615 $Y=0.735
+ $X2=4.615 $Y2=0.445
r198 2 30 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.065 $X2=2.725 $Y2=2.335
r199 1 34 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.79 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_1288_261# 1 2 7 9 12 21 24 28 31 32
c69 31 0 1.7977e-19 $X=8.21 $Y=1.67
c70 7 0 5.96505e-20 $X=6.54 $Y=1.99
r71 30 32 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=8.295 $Y=1.67
+ $X2=8.445 $Y2=1.67
r72 30 31 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=1.67
+ $X2=8.21 $Y2=1.67
r73 26 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.295 $Y=0.515
+ $X2=8.445 $Y2=0.515
r74 24 32 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=8.445 $Y=1.575
+ $X2=8.445 $Y2=1.67
r75 23 28 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=8.445 $Y=0.68
+ $X2=8.445 $Y2=0.515
r76 23 24 47.2684 $w=2.08e-07 $l=8.95e-07 $layer=LI1_cond $X=8.445 $Y=0.68
+ $X2=8.445 $Y2=1.575
r77 19 30 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.295 $Y=1.765
+ $X2=8.295 $Y2=1.67
r78 19 21 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.295 $Y=1.765
+ $X2=8.295 $Y2=1.87
r79 16 31 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=6.625 $Y=1.66
+ $X2=8.21 $Y2=1.66
r80 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.625
+ $Y=1.66 $X2=6.625 $Y2=1.66
r81 10 17 62.9618 $w=3.88e-07 $l=4.61519e-07 $layer=POLY_cond $X=7.005 $Y=1.305
+ $X2=6.76 $Y2=1.66
r82 10 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.005 $Y=1.305
+ $X2=7.005 $Y2=0.445
r83 7 17 54.9609 $w=3.88e-07 $l=4.26028e-07 $layer=POLY_cond $X=6.54 $Y=1.99
+ $X2=6.76 $Y2=1.66
r84 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.54 $Y=1.99 $X2=6.54
+ $Y2=2.275
r85 2 21 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=8.15
+ $Y=1.645 $X2=8.295 $Y2=1.87
r86 1 26 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=8.16
+ $Y=0.235 $X2=8.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_1126_413# 1 2 3 10 12 15 17 19 21 24 26
+ 27 32 33 37 38 39 42 47 49 52 54 56
c156 52 0 9.39049e-20 $X=7.005 $Y=1.32
c157 24 0 1.24715e-19 $X=9.075 $Y=0.56
r158 55 58 1.29832 $w=2.97e-07 $l=8e-09 $layer=POLY_cond $X=7.99 $Y=1.26
+ $X2=7.99 $Y2=1.252
r159 54 56 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=1.29
+ $X2=7.79 $Y2=1.29
r160 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=1.26 $X2=7.955 $Y2=1.26
r161 45 47 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=7.26 $Y=2.085
+ $X2=7.26 $Y2=2.21
r162 44 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.32
+ $X2=7.005 $Y2=1.32
r163 44 56 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.09 $Y=1.32 $X2=7.79
+ $Y2=1.32
r164 42 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=1.235
+ $X2=7.005 $Y2=1.32
r165 41 42 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.005 $Y=0.475
+ $X2=7.005 $Y2=1.235
r166 40 49 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.29 $Y=2 $X2=6.18
+ $Y2=2
r167 39 45 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.14 $Y=2
+ $X2=7.26 $Y2=2.085
r168 39 40 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.14 $Y=2 $X2=6.29
+ $Y2=2
r169 37 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=1.32
+ $X2=7.005 $Y2=1.32
r170 37 38 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.92 $Y=1.32
+ $X2=6.29 $Y2=1.32
r171 33 41 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.92 $Y=0.39
+ $X2=7.005 $Y2=0.475
r172 33 35 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.92 $Y=0.39
+ $X2=6.355 $Y2=0.39
r173 32 49 4.45262 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=1.915
+ $X2=6.18 $Y2=2
r174 31 38 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.18 $Y=1.405
+ $X2=6.29 $Y2=1.32
r175 31 32 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=6.18 $Y=1.405
+ $X2=6.18 $Y2=1.915
r176 27 49 15.1913 $w=2.18e-07 $l=2.9e-07 $layer=LI1_cond $X=6.18 $Y=2.29
+ $X2=6.18 $Y2=2
r177 27 29 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.07 $Y=2.29
+ $X2=5.775 $Y2=2.29
r178 22 26 33.6231 $w=1.65e-07 $l=1.667e-07 $layer=POLY_cond $X=9.075 $Y=1.095
+ $X2=9.055 $Y2=1.252
r179 22 24 274.33 $w=1.5e-07 $l=5.35e-07 $layer=POLY_cond $X=9.075 $Y=1.095
+ $X2=9.075 $Y2=0.56
r180 19 26 33.6231 $w=1.65e-07 $l=1.60481e-07 $layer=POLY_cond $X=9.05 $Y=1.41
+ $X2=9.055 $Y2=1.252
r181 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.05 $Y=1.41
+ $X2=9.05 $Y2=1.985
r182 18 58 1.48158 $w=3.15e-07 $l=1.7e-07 $layer=POLY_cond $X=8.16 $Y=1.252
+ $X2=7.99 $Y2=1.252
r183 17 26 3.33671 $w=3.15e-07 $l=9.5e-08 $layer=POLY_cond $X=8.96 $Y=1.252
+ $X2=9.055 $Y2=1.252
r184 17 18 146.55 $w=3.15e-07 $l=8e-07 $layer=POLY_cond $X=8.96 $Y=1.252
+ $X2=8.16 $Y2=1.252
r185 13 58 37.2679 $w=2.97e-07 $l=1.98907e-07 $layer=POLY_cond $X=8.085 $Y=1.095
+ $X2=7.99 $Y2=1.252
r186 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.085 $Y=1.095
+ $X2=8.085 $Y2=0.505
r187 10 55 57.7348 $w=2.97e-07 $l=3.4322e-07 $layer=POLY_cond $X=8.06 $Y=1.57
+ $X2=7.99 $Y2=1.26
r188 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.06 $Y=1.57
+ $X2=8.06 $Y2=2.065
r189 3 47 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.17
+ $Y=2.065 $X2=7.295 $Y2=2.21
r190 2 29 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=2.065 $X2=5.775 $Y2=2.33
r191 1 35 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.235 $X2=6.355 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_1738_47# 1 2 7 9 10 12 13 15 16 18 23 28
+ 31 35 37 40
r77 40 41 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=9.99 $Y=1.202
+ $X2=10.015 $Y2=1.202
r78 39 40 60.25 $w=3.76e-07 $l=4.7e-07 $layer=POLY_cond $X=9.52 $Y=1.202
+ $X2=9.99 $Y2=1.202
r79 35 36 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=2 $X2=8.815
+ $Y2=1.915
r80 32 39 3.20479 $w=3.76e-07 $l=2.5e-08 $layer=POLY_cond $X=9.495 $Y=1.202
+ $X2=9.52 $Y2=1.202
r81 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.495
+ $Y=1.16 $X2=9.495 $Y2=1.16
r82 29 37 0.221902 $w=3.3e-07 $l=1.25e-07 $layer=LI1_cond $X=8.98 $Y=1.16
+ $X2=8.855 $Y2=1.16
r83 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=8.98 $Y=1.16
+ $X2=9.495 $Y2=1.16
r84 28 36 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.855 $Y=1.66
+ $X2=8.855 $Y2=1.915
r85 25 37 7.38875 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=8.855 $Y=1.325
+ $X2=8.855 $Y2=1.16
r86 25 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.855 $Y=1.325
+ $X2=8.855 $Y2=1.66
r87 21 37 7.38875 $w=2.1e-07 $l=1.83916e-07 $layer=LI1_cond $X=8.815 $Y=0.995
+ $X2=8.855 $Y2=1.16
r88 21 23 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.815 $Y=0.995
+ $X2=8.815 $Y2=0.51
r89 16 41 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.015 $Y=0.995
+ $X2=10.015 $Y2=1.202
r90 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.015 $Y=0.995
+ $X2=10.015 $Y2=0.56
r91 13 40 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.99 $Y=1.41
+ $X2=9.99 $Y2=1.202
r92 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.99 $Y=1.41
+ $X2=9.99 $Y2=1.985
r93 10 39 19.9938 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.52 $Y=1.41
+ $X2=9.52 $Y2=1.202
r94 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.52 $Y=1.41
+ $X2=9.52 $Y2=1.985
r95 7 32 24.356 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.495 $Y=0.995
+ $X2=9.495 $Y2=1.202
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.495 $Y=0.995
+ $X2=9.495 $Y2=0.56
r97 2 35 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=8.69
+ $Y=1.485 $X2=8.815 $Y2=2
r98 2 28 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=8.69
+ $Y=1.485 $X2=8.815 $Y2=1.66
r99 1 23 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.69
+ $Y=0.235 $X2=8.815 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%VPWR 1 2 3 4 5 6 7 8 27 29 33 37 41 45 47
+ 50 51 53 54 55 57 59 65 73 78 96 101 104 107 114 121 129
c173 8 0 6.22691e-20 $X=10.08 $Y=1.485
c174 1 0 1.76957e-19 $X=0.585 $Y=1.815
r175 128 129 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r176 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r177 121 124 9.67042 $w=4.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.705 $Y=2.34
+ $X2=6.705 $Y2=2.72
r178 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r179 114 117 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.87 $Y=2.34
+ $X2=4.87 $Y2=2.72
r180 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r181 107 110 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.92 $Y=2.34
+ $X2=3.92 $Y2=2.72
r182 104 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r183 102 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r184 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r185 99 129 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r186 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r187 96 128 4.11489 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=10.185 $Y=2.72
+ $X2=10.382 $Y2=2.72
r188 96 98 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.185 $Y=2.72
+ $X2=9.89 $Y2=2.72
r189 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r190 94 95 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r191 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r192 91 94 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r193 91 92 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r194 89 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r195 89 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r196 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r197 86 124 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.705 $Y2=2.72
r198 86 88 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.59 $Y2=2.72
r199 85 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r200 84 85 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r201 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r202 82 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r203 81 84 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r204 81 82 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r205 79 117 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=4.87 $Y2=2.72
r206 79 81 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=5.29 $Y2=2.72
r207 78 124 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=6.47 $Y=2.72
+ $X2=6.705 $Y2=2.72
r208 78 84 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.47 $Y=2.72
+ $X2=6.21 $Y2=2.72
r209 77 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r210 77 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r211 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r212 74 110 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=3.92 $Y2=2.72
r213 74 76 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=4.37 $Y2=2.72
r214 73 117 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.68 $Y=2.72
+ $X2=4.87 $Y2=2.72
r215 73 76 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.68 $Y=2.72
+ $X2=4.37 $Y2=2.72
r216 72 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r217 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r218 69 72 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r219 69 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r220 68 71 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r221 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r222 66 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=1.72 $Y2=2.72
r223 66 68 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=2.07 $Y2=2.72
r224 65 110 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.92 $Y2=2.72
r225 65 71 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r226 59 101 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r227 57 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r228 55 59 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r229 55 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r230 53 94 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=9.2 $Y=2.72
+ $X2=8.97 $Y2=2.72
r231 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.2 $Y=2.72
+ $X2=9.285 $Y2=2.72
r232 52 98 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=9.37 $Y=2.72
+ $X2=9.89 $Y2=2.72
r233 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.37 $Y=2.72
+ $X2=9.285 $Y2=2.72
r234 50 88 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r235 50 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.875 $Y2=2.72
r236 49 91 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=8.05 $Y2=2.72
r237 49 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=7.875 $Y2=2.72
r238 45 128 3.13317 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=10.317
+ $Y=2.635 $X2=10.382 $Y2=2.72
r239 45 47 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=10.317 $Y=2.635
+ $X2=10.317 $Y2=1.955
r240 41 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=9.285 $Y=1.66
+ $X2=9.285 $Y2=2.34
r241 39 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.285 $Y=2.635
+ $X2=9.285 $Y2=2.72
r242 39 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.285 $Y=2.635
+ $X2=9.285 $Y2=2.34
r243 35 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.72
r244 35 37 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.21
r245 31 104 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r246 31 33 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.22
r247 30 101 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r248 29 104 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.72 $Y2=2.72
r249 29 30 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.895 $Y2=2.72
r250 25 101 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r251 25 27 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r252 8 47 300 $w=1.7e-07 $l=5.56956e-07 $layer=licon1_PDIFF $count=2 $X=10.08
+ $Y=1.485 $X2=10.27 $Y2=1.955
r253 7 44 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.485 $X2=9.285 $Y2=2.34
r254 7 41 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.14
+ $Y=1.485 $X2=9.285 $Y2=1.66
r255 6 37 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=7.62
+ $Y=2.065 $X2=7.825 $Y2=2.21
r256 5 121 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=6.63
+ $Y=2.065 $X2=6.775 $Y2=2.34
r257 4 114 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=2.065 $X2=4.895 $Y2=2.34
r258 3 107 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.065 $X2=3.895 $Y2=2.34
r259 2 33 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.645 $X2=1.72 $Y2=2.22
r260 1 27 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%A_409_329# 1 2 8 9 10 11 12 15 20
c59 20 0 1.81236e-19 $X=2.19 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0.635
+ $X2=2.19 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=1.88
+ $X2=2.19 $Y2=1.88
r62 11 12 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.105 $Y=1.88
+ $X2=1.7 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.105 $Y=0.73
+ $X2=2.19 $Y2=0.635
r64 9 10 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=2.105 $Y=0.73
+ $X2=1.7 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=1.795
+ $X2=1.7 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.7 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.615 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.645 $X2=2.19 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%Q 1 2 7 8 9 10 11 12 23 40 49
c38 40 0 1.86984e-19 $X=10.25 $Y=0.85
r39 49 50 1.08688 $w=9.43e-07 $l=3.5e-08 $layer=LI1_cond $X=10.012 $Y=1.53
+ $X2=10.012 $Y2=1.495
r40 40 47 0.406829 $w=7.33e-07 $l=2.5e-08 $layer=LI1_cond $X=10.117 $Y=0.85
+ $X2=10.117 $Y2=0.825
r41 36 46 4.01609 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=9.85 $Y=0.63
+ $X2=9.85 $Y2=0.745
r42 23 52 1.13313 $w=4.73e-07 $l=4.5e-08 $layer=LI1_cond $X=9.777 $Y=1.66
+ $X2=9.777 $Y2=1.615
r43 12 52 3.78883 $w=9.43e-07 $l=6e-08 $layer=LI1_cond $X=10.012 $Y=1.555
+ $X2=10.012 $Y2=1.615
r44 12 49 0.322751 $w=9.43e-07 $l=2.5e-08 $layer=LI1_cond $X=10.012 $Y=1.555
+ $X2=10.012 $Y2=1.53
r45 12 50 0.406829 $w=7.33e-07 $l=2.5e-08 $layer=LI1_cond $X=10.117 $Y=1.47
+ $X2=10.117 $Y2=1.495
r46 11 12 4.55649 $w=7.33e-07 $l=2.8e-07 $layer=LI1_cond $X=10.117 $Y=1.19
+ $X2=10.117 $Y2=1.47
r47 10 47 0.548694 $w=7.98e-07 $l=3e-08 $layer=LI1_cond $X=10.085 $Y=0.795
+ $X2=10.085 $Y2=0.825
r48 10 46 4.9885 $w=7.98e-07 $l=5e-08 $layer=LI1_cond $X=10.085 $Y=0.795
+ $X2=10.085 $Y2=0.745
r49 10 11 5.04468 $w=7.33e-07 $l=3.1e-07 $layer=LI1_cond $X=10.117 $Y=0.88
+ $X2=10.117 $Y2=1.19
r50 10 40 0.488195 $w=7.33e-07 $l=3e-08 $layer=LI1_cond $X=10.117 $Y=0.88
+ $X2=10.117 $Y2=0.85
r51 9 36 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=9.85 $Y=0.51 $X2=9.85
+ $Y2=0.63
r52 8 29 3.27348 $w=4.73e-07 $l=1.3e-07 $layer=LI1_cond $X=9.777 $Y=2.21
+ $X2=9.777 $Y2=2.34
r53 7 8 8.5614 $w=4.73e-07 $l=3.4e-07 $layer=LI1_cond $X=9.777 $Y=1.87 $X2=9.777
+ $Y2=2.21
r54 7 23 5.28793 $w=4.73e-07 $l=2.1e-07 $layer=LI1_cond $X=9.777 $Y=1.87
+ $X2=9.777 $Y2=1.66
r55 2 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.61
+ $Y=1.485 $X2=9.755 $Y2=2.34
r56 2 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.61
+ $Y=1.485 $X2=9.755 $Y2=1.66
r57 1 36 182 $w=1.7e-07 $l=4.96865e-07 $layer=licon1_NDIFF $count=1 $X=9.57
+ $Y=0.235 $X2=9.8 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_2%VGND 1 2 3 4 5 6 7 22 26 30 34 36 38 41 42
+ 43 45 47 53 58 78 84 90 93 100 105 108 111
c170 111 0 2.71124e-20 $X=10.35 $Y=0
c171 105 0 3.3422e-20 $X=7.32 $Y=0.24
c172 5 0 1.71107e-19 $X=7.44 $Y=0.235
r173 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r174 107 108 13.0581 $w=6.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.725 $Y=0.24
+ $X2=8.03 $Y2=0.24
r175 103 107 2.48416 $w=6.48e-07 $l=1.35e-07 $layer=LI1_cond $X=7.59 $Y=0.24
+ $X2=7.725 $Y2=0.24
r176 103 105 12.4141 $w=6.48e-07 $l=2.7e-07 $layer=LI1_cond $X=7.59 $Y=0.24
+ $X2=7.32 $Y2=0.24
r177 103 104 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r178 100 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r179 93 97 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=4.14 $Y=0 $X2=4.14
+ $Y2=0.36
r180 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r181 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r182 85 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r183 84 87 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r184 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r185 81 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r186 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r187 78 110 4.11489 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=10.382 $Y2=0
r188 78 80 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=10.185 $Y=0
+ $X2=9.89 $Y2=0
r189 77 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r190 76 77 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r191 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r192 74 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r193 73 76 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r194 73 108 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.03
+ $Y2=0
r195 73 74 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r196 70 104 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r197 69 105 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=7.32
+ $Y2=0
r198 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r199 67 70 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r200 67 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r201 66 69 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=7.13
+ $Y2=0
r202 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r203 64 100 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.335
+ $Y2=0
r204 64 66 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.75
+ $Y2=0
r205 62 101 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r206 62 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r207 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r208 59 93 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.14
+ $Y2=0
r209 59 61 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r210 58 100 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.335
+ $Y2=0
r211 58 61 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=4.83
+ $Y2=0
r212 57 94 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.91 $Y2=0
r213 57 91 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r214 56 57 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r215 54 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.72
+ $Y2=0
r216 54 56 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=2.07 $Y2=0
r217 53 93 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.14
+ $Y2=0
r218 53 56 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=2.07
+ $Y2=0
r219 47 84 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r220 45 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r221 43 47 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r222 43 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r223 41 76 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=9.07 $Y=0 $X2=8.97
+ $Y2=0
r224 41 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.07 $Y=0 $X2=9.26
+ $Y2=0
r225 40 80 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=9.45 $Y=0 $X2=9.89
+ $Y2=0
r226 40 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.45 $Y=0 $X2=9.26
+ $Y2=0
r227 36 110 3.13317 $w=2.65e-07 $l=1.12916e-07 $layer=LI1_cond $X=10.317
+ $Y=0.085 $X2=10.382 $Y2=0
r228 36 38 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=10.317 $Y=0.085
+ $X2=10.317 $Y2=0.38
r229 32 42 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0
r230 32 34 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=9.26 $Y=0.085
+ $X2=9.26 $Y2=0.38
r231 28 100 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.335 $Y=0.085
+ $X2=5.335 $Y2=0
r232 28 30 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0.085
+ $X2=5.335 $Y2=0.38
r233 24 90 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r234 24 26 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.38
r235 23 84 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r236 22 90 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=0 $X2=1.72
+ $Y2=0
r237 22 23 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=0.895 $Y2=0
r238 7 38 182 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=1 $X=10.09
+ $Y=0.235 $X2=10.27 $Y2=0.38
r239 6 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=9.15
+ $Y=0.235 $X2=9.285 $Y2=0.38
r240 5 107 182 $w=1.7e-07 $l=3.88652e-07 $layer=licon1_NDIFF $count=1 $X=7.44
+ $Y=0.235 $X2=7.725 $Y2=0.48
r241 4 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.235 $X2=5.445 $Y2=0.38
r242 3 97 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.235 $X2=3.995 $Y2=0.36
r243 2 26 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.38
r244 1 87 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

