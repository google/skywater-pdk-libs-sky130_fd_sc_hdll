* File: sky130_fd_sc_hdll__clkinv_4.pex.spice
* Created: Wed Sep  2 08:26:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_4%A 1 3 6 8 10 11 15 17 19 20 24 26 28 29
+ 33 35 37 38 40 41 42 43 44 45 47 48 49 50 51 52 53 67 70 74 78 82
c108 48 0 1.9478e-19 $X=2.84 $Y=1.16
c109 42 0 1.9478e-19 $X=0.92 $Y=1.16
r110 63 82 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.56
+ $Y=1.16 $X2=2.56 $Y2=1.16
r111 60 67 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.66
+ $Y=1.16 $X2=0.66 $Y2=1.16
r112 53 82 12.8049 $w=2.23e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=1.177
+ $X2=2.53 $Y2=1.177
r113 52 82 13.3171 $w=2.23e-07 $l=2.6e-07 $layer=LI1_cond $X=2.27 $Y=1.177
+ $X2=2.53 $Y2=1.177
r114 52 78 10.2439 $w=2.23e-07 $l=2e-07 $layer=LI1_cond $X=2.27 $Y=1.177
+ $X2=2.07 $Y2=1.177
r115 51 78 15.8781 $w=2.23e-07 $l=3.1e-07 $layer=LI1_cond $X=1.76 $Y=1.177
+ $X2=2.07 $Y2=1.177
r116 51 74 7.68295 $w=2.23e-07 $l=1.5e-07 $layer=LI1_cond $X=1.76 $Y=1.177
+ $X2=1.61 $Y2=1.177
r117 50 74 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=1.25 $Y=1.177
+ $X2=1.61 $Y2=1.177
r118 50 70 5.12197 $w=2.23e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=1.177
+ $X2=1.15 $Y2=1.177
r119 49 70 21.0001 $w=2.23e-07 $l=4.1e-07 $layer=LI1_cond $X=0.74 $Y=1.177
+ $X2=1.15 $Y2=1.177
r120 49 67 4.09758 $w=2.23e-07 $l=8e-08 $layer=LI1_cond $X=0.74 $Y=1.177
+ $X2=0.66 $Y2=1.177
r121 48 63 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.84 $Y=1.16
+ $X2=2.56 $Y2=1.16
r122 47 63 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=2.46 $Y=1.217
+ $X2=2.56 $Y2=1.16
r123 42 60 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=0.66 $Y2=1.16
r124 42 43 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=0.92 $Y=1.16
+ $X2=1.02 $Y2=1.217
r125 41 60 4.44347 $w=2.7e-07 $l=2e-08 $layer=POLY_cond $X=0.64 $Y=1.16 $X2=0.66
+ $Y2=1.16
r126 38 48 28.3559 $w=2.7e-07 $l=2.95804e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.84 $Y2=1.16
r127 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.94 $Y=1.41
+ $X2=2.94 $Y2=1.985
r128 35 47 18.4447 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.46 $Y2=1.217
r129 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.46 $Y=1.41
+ $X2=2.46 $Y2=1.985
r130 31 47 18.4447 $w=1.5e-07 $l=2.04118e-07 $layer=POLY_cond $X=2.435 $Y=1.025
+ $X2=2.46 $Y2=1.217
r131 31 33 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=2.435 $Y=1.025
+ $X2=2.435 $Y2=0.445
r132 30 45 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=2.08 $Y=1.16
+ $X2=1.98 $Y2=1.217
r133 29 47 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=2.36 $Y=1.16
+ $X2=2.46 $Y2=1.217
r134 29 30 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=2.36 $Y=1.16
+ $X2=2.08 $Y2=1.16
r135 26 45 18.4447 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.98 $Y=1.41
+ $X2=1.98 $Y2=1.217
r136 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.98 $Y=1.41
+ $X2=1.98 $Y2=1.985
r137 22 45 18.4447 $w=1.5e-07 $l=2.04118e-07 $layer=POLY_cond $X=1.955 $Y=1.025
+ $X2=1.98 $Y2=1.217
r138 22 24 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.955 $Y=1.025
+ $X2=1.955 $Y2=0.445
r139 21 44 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=1.6 $Y=1.16
+ $X2=1.5 $Y2=1.217
r140 20 45 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.98 $Y2=1.217
r141 20 21 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.88 $Y=1.16
+ $X2=1.6 $Y2=1.16
r142 17 44 18.4447 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.217
r143 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.5 $Y2=1.985
r144 13 44 18.4447 $w=1.5e-07 $l=2.04118e-07 $layer=POLY_cond $X=1.475 $Y=1.025
+ $X2=1.5 $Y2=1.217
r145 13 15 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=1.475 $Y=1.025
+ $X2=1.475 $Y2=0.445
r146 12 43 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=1.12 $Y=1.16
+ $X2=1.02 $Y2=1.217
r147 11 44 6.70161 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=1.4 $Y=1.16
+ $X2=1.5 $Y2=1.217
r148 11 12 62.2086 $w=2.7e-07 $l=2.8e-07 $layer=POLY_cond $X=1.4 $Y=1.16
+ $X2=1.12 $Y2=1.16
r149 8 43 18.4447 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.217
r150 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r151 4 43 18.4447 $w=1.5e-07 $l=2.04118e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=1.02 $Y2=1.217
r152 4 6 297.404 $w=1.5e-07 $l=5.8e-07 $layer=POLY_cond $X=0.995 $Y=1.025
+ $X2=0.995 $Y2=0.445
r153 1 41 28.3559 $w=2.7e-07 $l=2.95804e-07 $layer=POLY_cond $X=0.54 $Y=1.41
+ $X2=0.64 $Y2=1.16
r154 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.54 $Y=1.41
+ $X2=0.54 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_4%VPWR 1 2 3 4 13 15 17 21 25 27 29 32 33
+ 34 40 48 52
r52 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r53 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r54 43 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 42 43 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r56 40 51 4.96304 $w=1.7e-07 $l=3.15e-07 $layer=LI1_cond $X=3.05 $Y=2.72
+ $X2=3.365 $Y2=2.72
r57 40 42 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.05 $Y=2.72 $X2=2.99
+ $Y2=2.72
r58 39 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 39 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r60 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r61 36 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.39 $Y=2.72 $X2=1.26
+ $Y2=2.72
r62 36 38 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.39 $Y=2.72
+ $X2=2.07 $Y2=2.72
r63 34 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 34 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 32 38 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=2.09 $Y=2.72 $X2=2.07
+ $Y2=2.72
r66 32 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.09 $Y=2.72 $X2=2.22
+ $Y2=2.72
r67 31 42 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=2.35 $Y=2.72 $X2=2.99
+ $Y2=2.72
r68 31 33 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.35 $Y=2.72 $X2=2.22
+ $Y2=2.72
r69 27 51 3.27718 $w=3.85e-07 $l=1.5995e-07 $layer=LI1_cond $X=3.242 $Y=2.635
+ $X2=3.365 $Y2=2.72
r70 27 29 20.0555 $w=3.83e-07 $l=6.7e-07 $layer=LI1_cond $X=3.242 $Y=2.635
+ $X2=3.242 $Y2=1.965
r71 23 33 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.635
+ $X2=2.22 $Y2=2.72
r72 23 25 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=2.22 $Y=2.635
+ $X2=2.22 $Y2=1.965
r73 19 48 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=2.635
+ $X2=1.26 $Y2=2.72
r74 19 21 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.26 $Y=2.635
+ $X2=1.26 $Y2=1.965
r75 18 45 4.96256 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=0.43 $Y=2.72
+ $X2=0.215 $Y2=2.72
r76 17 48 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.13 $Y=2.72 $X2=1.26
+ $Y2=2.72
r77 17 18 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.13 $Y=2.72 $X2=0.43
+ $Y2=2.72
r78 13 45 2.93137 $w=3.45e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.215 $Y2=2.72
r79 13 15 22.3808 $w=3.43e-07 $l=6.7e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=1.965
r80 4 29 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=3.03
+ $Y=1.485 $X2=3.18 $Y2=1.965
r81 3 25 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=2.07
+ $Y=1.485 $X2=2.22 $Y2=1.965
r82 2 21 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.485 $X2=1.26 $Y2=1.965
r83 1 15 300 $w=1.7e-07 $l=5.56417e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.3 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_4%Y 1 2 3 4 5 17 18 19 20 21 24 26 30 32 36
+ 38 42 44 48 50 52 53 54 55 56 57 58 59 65 66
c117 38 0 1.9478e-19 $X=2.57 $Y=1.545
c118 26 0 1.9478e-19 $X=1.615 $Y=1.545
r119 59 66 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=1.545 $X2=3.42
+ $Y2=1.46
r120 59 66 0.307318 $w=2.98e-07 $l=8e-09 $layer=LI1_cond $X=3.42 $Y=1.452
+ $X2=3.42 $Y2=1.46
r121 58 59 10.0647 $w=2.98e-07 $l=2.62e-07 $layer=LI1_cond $X=3.42 $Y=1.19
+ $X2=3.42 $Y2=1.452
r122 57 65 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.42 $Y=0.81 $X2=3.42
+ $Y2=0.895
r123 57 58 10.5641 $w=2.98e-07 $l=2.75e-07 $layer=LI1_cond $X=3.42 $Y=0.915
+ $X2=3.42 $Y2=1.19
r124 57 65 0.768295 $w=2.98e-07 $l=2e-08 $layer=LI1_cond $X=3.42 $Y=0.915
+ $X2=3.42 $Y2=0.895
r125 51 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.83 $Y=1.545
+ $X2=2.7 $Y2=1.545
r126 50 59 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.27 $Y=1.545
+ $X2=3.42 $Y2=1.545
r127 50 51 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=3.27 $Y=1.545
+ $X2=2.83 $Y2=1.545
r128 46 56 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=1.63 $X2=2.7
+ $Y2=1.545
r129 46 48 8.86495 $w=2.58e-07 $l=2e-07 $layer=LI1_cond $X=2.7 $Y=1.63 $X2=2.7
+ $Y2=1.83
r130 45 55 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.345 $Y=0.81
+ $X2=2.217 $Y2=0.81
r131 44 57 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=3.27 $Y=0.81
+ $X2=3.42 $Y2=0.81
r132 44 45 60.3476 $w=1.68e-07 $l=9.25e-07 $layer=LI1_cond $X=3.27 $Y=0.81
+ $X2=2.345 $Y2=0.81
r133 40 55 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.217 $Y=0.725
+ $X2=2.217 $Y2=0.81
r134 40 42 12.6543 $w=2.53e-07 $l=2.8e-07 $layer=LI1_cond $X=2.217 $Y=0.725
+ $X2=2.217 $Y2=0.445
r135 39 54 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=1.87 $Y=1.545
+ $X2=1.742 $Y2=1.545
r136 38 56 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.57 $Y=1.545
+ $X2=2.7 $Y2=1.545
r137 38 39 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.57 $Y=1.545
+ $X2=1.87 $Y2=1.545
r138 34 54 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.742 $Y=1.63
+ $X2=1.742 $Y2=1.545
r139 34 36 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=1.742 $Y=1.63
+ $X2=1.742 $Y2=1.83
r140 33 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.39 $Y=0.81
+ $X2=1.26 $Y2=0.81
r141 32 55 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.09 $Y=0.81
+ $X2=2.217 $Y2=0.81
r142 32 33 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.09 $Y=0.81 $X2=1.39
+ $Y2=0.81
r143 28 53 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=0.725
+ $X2=1.26 $Y2=0.81
r144 28 30 12.4109 $w=2.58e-07 $l=2.8e-07 $layer=LI1_cond $X=1.26 $Y=0.725
+ $X2=1.26 $Y2=0.445
r145 27 52 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.91 $Y=1.545
+ $X2=0.782 $Y2=1.545
r146 26 54 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=1.615 $Y=1.545
+ $X2=1.742 $Y2=1.545
r147 26 27 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=1.615 $Y=1.545
+ $X2=0.91 $Y2=1.545
r148 22 52 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.782 $Y=1.63
+ $X2=0.782 $Y2=1.545
r149 22 24 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=0.782 $Y=1.63
+ $X2=0.782 $Y2=1.83
r150 20 52 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.655 $Y=1.545
+ $X2=0.782 $Y2=1.545
r151 20 21 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.655 $Y=1.545
+ $X2=0.275 $Y2=1.545
r152 18 53 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.13 $Y=0.81
+ $X2=1.26 $Y2=0.81
r153 18 19 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.13 $Y=0.81
+ $X2=0.275 $Y2=0.81
r154 17 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=1.46
+ $X2=0.275 $Y2=1.545
r155 16 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.275 $Y2=0.81
r156 16 17 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=0.19 $Y=0.895
+ $X2=0.19 $Y2=1.46
r157 5 48 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=2.55
+ $Y=1.485 $X2=2.7 $Y2=1.83
r158 4 36 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=1.59
+ $Y=1.485 $X2=1.74 $Y2=1.83
r159 3 24 300 $w=1.7e-07 $l=4.13249e-07 $layer=licon1_PDIFF $count=2 $X=0.63
+ $Y=1.485 $X2=0.78 $Y2=1.83
r160 2 42 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.03
+ $Y=0.235 $X2=2.22 $Y2=0.445
r161 1 30 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_4%VGND 1 2 3 12 14 18 22 25 26 27 29 39 40
+ 43 46
r45 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r46 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r47 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r50 37 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r51 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 34 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=1.74
+ $Y2=0
r53 34 36 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.87 $Y=0 $X2=2.53
+ $Y2=0
r54 29 43 8.88104 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.737
+ $Y2=0
r55 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.23
+ $Y2=0
r56 27 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r57 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 25 36 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.53
+ $Y2=0
r59 25 26 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.565 $Y=0 $X2=2.715
+ $Y2=0
r60 24 39 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=3.45
+ $Y2=0
r61 24 26 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.715
+ $Y2=0
r62 20 26 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0
r63 20 22 11.7165 $w=2.98e-07 $l=3.05e-07 $layer=LI1_cond $X=2.715 $Y=0.085
+ $X2=2.715 $Y2=0.39
r64 16 46 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0
r65 16 18 13.519 $w=2.58e-07 $l=3.05e-07 $layer=LI1_cond $X=1.74 $Y=0.085
+ $X2=1.74 $Y2=0.39
r66 15 43 8.88104 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.91 $Y=0 $X2=0.737
+ $Y2=0
r67 14 46 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.74
+ $Y2=0
r68 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=0.91
+ $Y2=0
r69 10 43 1.03204 $w=3.45e-07 $l=8.5e-08 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0
r70 10 12 10.1883 $w=3.43e-07 $l=3.05e-07 $layer=LI1_cond $X=0.737 $Y=0.085
+ $X2=0.737 $Y2=0.39
r71 3 22 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=2.51
+ $Y=0.235 $X2=2.7 $Y2=0.39
r72 2 18 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=1.55
+ $Y=0.235 $X2=1.74 $Y2=0.39
r73 1 12 182 $w=1.7e-07 $l=3.07896e-07 $layer=licon1_NDIFF $count=1 $X=0.54
+ $Y=0.235 $X2=0.78 $Y2=0.39
.ends

