* File: sky130_fd_sc_hdll__buf_2.pxi.spice
* Created: Wed Sep  2 08:24:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_2%A N_A_c_47_n N_A_c_48_n N_A_M1002_g N_A_M1000_g A
+ N_A_c_46_n PM_SKY130_FD_SC_HDLL__BUF_2%A
x_PM_SKY130_FD_SC_HDLL__BUF_2%A_27_47# N_A_27_47#_M1000_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_79_n N_A_27_47#_M1001_g N_A_27_47#_c_88_n N_A_27_47#_M1003_g
+ N_A_27_47#_c_80_n N_A_27_47#_c_81_n N_A_27_47#_c_91_n N_A_27_47#_M1004_g
+ N_A_27_47#_c_82_n N_A_27_47#_M1005_g N_A_27_47#_c_83_n N_A_27_47#_c_153_p
+ N_A_27_47#_c_93_n N_A_27_47#_c_84_n N_A_27_47#_c_85_n N_A_27_47#_c_94_n
+ N_A_27_47#_c_95_n N_A_27_47#_c_96_n N_A_27_47#_c_86_n N_A_27_47#_c_87_n
+ PM_SKY130_FD_SC_HDLL__BUF_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUF_2%VPWR N_VPWR_M1002_d N_VPWR_M1004_s N_VPWR_c_161_n
+ N_VPWR_c_162_n N_VPWR_c_163_n VPWR VPWR N_VPWR_c_164_n N_VPWR_c_165_n
+ N_VPWR_c_166_n N_VPWR_c_160_n PM_SKY130_FD_SC_HDLL__BUF_2%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_2%X N_X_M1001_d N_X_M1003_d X X X X X X
+ PM_SKY130_FD_SC_HDLL__BUF_2%X
x_PM_SKY130_FD_SC_HDLL__BUF_2%VGND N_VGND_M1000_d N_VGND_M1005_s N_VGND_c_211_n
+ N_VGND_c_212_n N_VGND_c_213_n VGND VGND N_VGND_c_214_n N_VGND_c_215_n
+ N_VGND_c_216_n N_VGND_c_217_n PM_SKY130_FD_SC_HDLL__BUF_2%VGND
cc_1 VNB N_A_M1000_g 0.0380428f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A 0.01798f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_A_c_46_n 0.0380199f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_47#_c_79_n 0.0175635f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_47#_c_80_n 0.0231971f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_6 VNB N_A_27_47#_c_81_n 0.0167981f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_7 VNB N_A_27_47#_c_82_n 0.0221394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_83_n 0.0237142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_84_n 0.00320505f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_85_n 0.0076639f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_86_n 0.00219346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_87_n 0.00102979f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VPWR_c_160_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB X 8.55205e-19 $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_15 VNB N_VGND_c_211_n 0.00285908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_212_n 0.0127809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_213_n 0.0358086f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_18 VNB N_VGND_c_214_n 0.0241666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_215_n 0.0187885f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_216_n 0.00513086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_217_n 0.147212f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A_c_47_n 0.0245065f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.63
cc_23 VPB N_A_c_48_n 0.0302378f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.73
cc_24 VPB A 0.00733067f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_25 VPB N_A_c_46_n 0.00931503f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_26 VPB N_A_27_47#_c_88_n 0.0175385f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_27 VPB N_A_27_47#_c_80_n 0.0149858f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_28 VPB N_A_27_47#_c_81_n 0.0102818f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_29 VPB N_A_27_47#_c_91_n 0.0200594f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A_27_47#_c_83_n 0.009426f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_A_27_47#_c_93_n 0.00661021f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_47#_c_94_n 0.00540387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_47#_c_95_n 0.00830608f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_47#_c_96_n 0.00261949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_47#_c_86_n 5.32814e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_161_n 0.00606664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_162_n 0.0127584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_163_n 0.0470309f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_39 VPB N_VPWR_c_164_n 0.019656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_165_n 0.0255311f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_166_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_160_n 0.0540136f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB X 0.00412346f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_44 N_A_M1000_g N_A_27_47#_c_79_n 0.0199163f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_45 N_A_c_47_n N_A_27_47#_c_88_n 0.00977992f $X=0.495 $Y=1.63 $X2=0 $Y2=0
cc_46 N_A_c_48_n N_A_27_47#_c_88_n 0.00769771f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_47 N_A_c_47_n N_A_27_47#_c_81_n 0.00250317f $X=0.495 $Y=1.63 $X2=0 $Y2=0
cc_48 A N_A_27_47#_c_81_n 2.91038e-19 $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_c_46_n N_A_27_47#_c_81_n 0.0211074f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_50 N_A_c_48_n N_A_27_47#_c_93_n 0.00802728f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_51 N_A_M1000_g N_A_27_47#_c_84_n 0.0178499f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_52 A N_A_27_47#_c_84_n 0.00726338f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_53 N_A_c_46_n N_A_27_47#_c_84_n 8.41031e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_54 A N_A_27_47#_c_85_n 0.0143207f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_55 N_A_c_46_n N_A_27_47#_c_85_n 0.00127129f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_c_47_n N_A_27_47#_c_94_n 0.0120572f $X=0.495 $Y=1.63 $X2=0 $Y2=0
cc_57 N_A_c_48_n N_A_27_47#_c_94_n 0.0123398f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_58 A N_A_27_47#_c_94_n 0.00690389f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_59 N_A_c_46_n N_A_27_47#_c_94_n 3.19113e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_60 A N_A_27_47#_c_95_n 0.0145573f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_61 N_A_c_46_n N_A_27_47#_c_95_n 0.00123585f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_c_47_n N_A_27_47#_c_96_n 0.00372007f $X=0.495 $Y=1.63 $X2=0 $Y2=0
cc_63 N_A_c_46_n N_A_27_47#_c_86_n 0.00372007f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_64 N_A_M1000_g N_A_27_47#_c_87_n 0.00372007f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_65 A N_A_27_47#_c_87_n 0.0197071f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_A_c_48_n N_VPWR_c_161_n 0.00395131f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_67 N_A_c_48_n N_VPWR_c_164_n 0.00702461f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_68 N_A_c_48_n N_VPWR_c_160_n 0.0136548f $X=0.495 $Y=1.73 $X2=0 $Y2=0
cc_69 N_A_M1000_g N_VGND_c_211_n 0.00316741f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_70 N_A_M1000_g N_VGND_c_215_n 0.00425094f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_71 N_A_M1000_g N_VGND_c_217_n 0.00681735f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_72 N_A_27_47#_c_94_n N_VPWR_M1002_d 0.0051833f $X=0.725 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_27_47#_c_96_n N_VPWR_M1002_d 7.12055e-19 $X=0.81 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_27_47#_c_88_n N_VPWR_c_161_n 0.0032688f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_27_47#_c_81_n N_VPWR_c_161_n 2.89388e-19 $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_27_47#_c_93_n N_VPWR_c_161_n 0.0165113f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_77 N_A_27_47#_c_94_n N_VPWR_c_161_n 0.0216025f $X=0.725 $Y=1.62 $X2=0 $Y2=0
cc_78 N_A_27_47#_c_91_n N_VPWR_c_163_n 0.0112858f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_27_47#_c_93_n N_VPWR_c_164_n 0.0120448f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_80 N_A_27_47#_c_88_n N_VPWR_c_165_n 0.00700684f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_47#_c_91_n N_VPWR_c_165_n 0.00429201f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_27_47#_c_88_n N_VPWR_c_160_n 0.0128328f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_27_47#_c_91_n N_VPWR_c_160_n 0.00745584f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_27_47#_c_93_n N_VPWR_c_160_n 0.00646998f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_85 N_A_27_47#_c_79_n X 0.00984749f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_27_47#_c_88_n X 0.0134185f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_80_n X 0.0225098f $X=1.495 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_81_n X 8.92342e-19 $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_89 N_A_27_47#_c_91_n X 0.0372272f $X=1.595 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_82_n X 0.0223942f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_83_n X 0.0260495f $X=1.595 $Y=1.202 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_84_n X 0.00855591f $X=0.725 $Y=0.72 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_96_n X 0.00858054f $X=0.81 $Y=1.535 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_86_n X 0.0187248f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_87_n X 0.00892895f $X=0.875 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_84_n N_VGND_M1000_d 0.00426581f $X=0.725 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_27_47#_c_87_n N_VGND_M1000_d 9.20178e-19 $X=0.875 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_27_47#_c_79_n N_VGND_c_211_n 0.00817114f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_27_47#_c_81_n N_VGND_c_211_n 3.34628e-19 $X=1.12 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_47#_c_82_n N_VGND_c_211_n 9.57539e-19 $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_84_n N_VGND_c_211_n 0.01863f $X=0.725 $Y=0.72 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_82_n N_VGND_c_213_n 0.0172406f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_79_n N_VGND_c_214_n 0.00505556f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_82_n N_VGND_c_214_n 0.00359186f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_153_p N_VGND_c_215_n 0.0116326f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_84_n N_VGND_c_215_n 0.00388761f $X=0.725 $Y=0.72 $X2=0 $Y2=0
cc_107 N_A_27_47#_M1000_s N_VGND_c_217_n 0.00429125f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_108 N_A_27_47#_c_79_n N_VGND_c_217_n 0.0090506f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_82_n N_VGND_c_217_n 0.00686961f $X=1.62 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_27_47#_c_153_p N_VGND_c_217_n 0.00643448f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_84_n N_VGND_c_217_n 0.00827273f $X=0.725 $Y=0.72 $X2=0 $Y2=0
cc_112 N_VPWR_c_160_n N_X_M1003_d 0.00876103f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_113 N_VPWR_c_161_n X 0.0298999f $X=0.765 $Y=1.96 $X2=0 $Y2=0
cc_114 N_VPWR_c_165_n X 0.0270609f $X=1.865 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_c_160_n X 0.0154673f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_116 N_VPWR_c_163_n N_VGND_c_213_n 0.0101002f $X=1.95 $Y=1.66 $X2=0 $Y2=0
cc_117 X N_VGND_c_211_n 0.0100008f $X=1.52 $Y=0.425 $X2=0 $Y2=0
cc_118 X N_VGND_c_213_n 0.0521193f $X=1.52 $Y=0.425 $X2=0 $Y2=0
cc_119 X N_VGND_c_214_n 0.0274408f $X=1.52 $Y=0.425 $X2=0 $Y2=0
cc_120 N_X_M1001_d N_VGND_c_217_n 0.0108114f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_121 X N_VGND_c_217_n 0.0156091f $X=1.52 $Y=0.425 $X2=0 $Y2=0
