* File: sky130_fd_sc_hdll__nand4_4.pxi.spice
* Created: Thu Aug 27 19:14:33 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4_4%D N_D_c_122_n N_D_M1001_g N_D_M1002_g
+ N_D_c_123_n N_D_M1014_g N_D_M1022_g N_D_c_124_n N_D_M1020_g N_D_M1023_g
+ N_D_c_125_n N_D_M1028_g N_D_M1031_g D D D D N_D_c_119_n N_D_c_120_n D D D
+ PM_SKY130_FD_SC_HDLL__NAND4_4%D
x_PM_SKY130_FD_SC_HDLL__NAND4_4%C N_C_M1012_g N_C_c_202_n N_C_M1000_g
+ N_C_M1018_g N_C_c_203_n N_C_M1006_g N_C_M1025_g N_C_c_204_n N_C_M1011_g
+ N_C_c_205_n N_C_M1017_g N_C_M1027_g C C C C N_C_c_201_n C C C C
+ PM_SKY130_FD_SC_HDLL__NAND4_4%C
x_PM_SKY130_FD_SC_HDLL__NAND4_4%B N_B_c_281_n N_B_M1003_g N_B_M1005_g
+ N_B_c_282_n N_B_M1009_g N_B_M1007_g N_B_c_283_n N_B_M1019_g N_B_M1015_g
+ N_B_c_284_n N_B_M1029_g N_B_M1021_g B B B B N_B_c_278_n N_B_c_279_n
+ N_B_c_280_n B B B B PM_SKY130_FD_SC_HDLL__NAND4_4%B
x_PM_SKY130_FD_SC_HDLL__NAND4_4%A N_A_M1008_g N_A_c_360_n N_A_M1004_g
+ N_A_M1010_g N_A_c_361_n N_A_M1013_g N_A_M1024_g N_A_c_362_n N_A_M1016_g
+ N_A_M1026_g N_A_c_363_n N_A_M1030_g A A A N_A_c_358_n N_A_c_359_n A A A
+ PM_SKY130_FD_SC_HDLL__NAND4_4%A
x_PM_SKY130_FD_SC_HDLL__NAND4_4%VPWR N_VPWR_M1001_d N_VPWR_M1014_d
+ N_VPWR_M1028_d N_VPWR_M1006_d N_VPWR_M1017_d N_VPWR_M1009_s N_VPWR_M1029_s
+ N_VPWR_M1013_s N_VPWR_M1030_s N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_436_n N_VPWR_c_437_n N_VPWR_c_438_n
+ N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_441_n N_VPWR_c_442_n N_VPWR_c_443_n
+ N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n N_VPWR_c_447_n N_VPWR_c_448_n
+ N_VPWR_c_449_n N_VPWR_c_450_n N_VPWR_c_451_n VPWR N_VPWR_c_452_n
+ N_VPWR_c_453_n N_VPWR_c_454_n N_VPWR_c_455_n N_VPWR_c_456_n N_VPWR_c_430_n
+ PM_SKY130_FD_SC_HDLL__NAND4_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4_4%Y N_Y_M1008_s N_Y_M1024_s N_Y_M1001_s
+ N_Y_M1020_s N_Y_M1000_s N_Y_M1011_s N_Y_M1003_d N_Y_M1019_d N_Y_M1004_d
+ N_Y_M1016_d N_Y_c_571_n N_Y_c_591_n N_Y_c_572_n N_Y_c_598_n N_Y_c_573_n
+ N_Y_c_603_n N_Y_c_574_n N_Y_c_619_n N_Y_c_575_n N_Y_c_637_n N_Y_c_576_n
+ N_Y_c_644_n N_Y_c_577_n N_Y_c_649_n N_Y_c_650_n N_Y_c_569_n N_Y_c_578_n
+ N_Y_c_579_n N_Y_c_680_n N_Y_c_580_n N_Y_c_581_n N_Y_c_582_n N_Y_c_583_n
+ N_Y_c_584_n N_Y_c_585_n Y PM_SKY130_FD_SC_HDLL__NAND4_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND4_4%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1022_d
+ N_A_27_47#_M1031_d N_A_27_47#_M1018_d N_A_27_47#_M1027_d N_A_27_47#_c_761_n
+ N_A_27_47#_c_762_n N_A_27_47#_c_763_n N_A_27_47#_c_775_n N_A_27_47#_c_764_n
+ N_A_27_47#_c_803_p N_A_27_47#_c_765_n N_A_27_47#_c_766_n
+ PM_SKY130_FD_SC_HDLL__NAND4_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4_4%VGND N_VGND_M1002_s N_VGND_M1023_s
+ N_VGND_c_823_n N_VGND_c_824_n VGND N_VGND_c_825_n N_VGND_c_826_n
+ N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n
+ PM_SKY130_FD_SC_HDLL__NAND4_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4_4%A_485_47# N_A_485_47#_M1012_s
+ N_A_485_47#_M1025_s N_A_485_47#_M1005_s N_A_485_47#_M1015_s
+ N_A_485_47#_c_910_n PM_SKY130_FD_SC_HDLL__NAND4_4%A_485_47#
x_PM_SKY130_FD_SC_HDLL__NAND4_4%A_883_47# N_A_883_47#_M1005_d
+ N_A_883_47#_M1007_d N_A_883_47#_M1021_d N_A_883_47#_M1010_d
+ N_A_883_47#_M1026_d N_A_883_47#_c_943_n N_A_883_47#_c_944_n
+ N_A_883_47#_c_945_n PM_SKY130_FD_SC_HDLL__NAND4_4%A_883_47#
cc_1 VNB N_D_M1002_g 0.0239286f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_D_M1022_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_D_M1023_g 0.0178804f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB N_D_M1031_g 0.018112f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_5 VNB N_D_c_119_n 0.0254432f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.165
cc_6 VNB N_D_c_120_n 0.0843311f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.217
cc_7 VNB D 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.615 $Y2=1.19
cc_8 VNB N_C_M1012_g 0.018242f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_9 VNB N_C_M1018_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_10 VNB N_C_M1025_g 0.0188863f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_11 VNB N_C_M1027_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_12 VNB C 0.00749491f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.105
cc_13 VNB N_C_c_201_n 0.0890066f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_14 VNB N_B_M1005_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_B_M1007_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_16 VNB N_B_M1015_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_17 VNB N_B_M1021_g 0.0189127f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_18 VNB N_B_c_278_n 0.0304355f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.165
cc_19 VNB N_B_c_279_n 0.00322659f $X=-0.19 $Y=-0.24 $X2=1.67 $Y2=1.16
cc_20 VNB N_B_c_280_n 0.0854483f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.217
cc_21 VNB N_A_M1008_g 0.0174843f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_22 VNB N_A_M1010_g 0.0183438f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_23 VNB N_A_M1024_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_24 VNB N_A_M1026_g 0.0243191f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_25 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.17 $Y2=1.105
cc_26 VNB N_A_c_358_n 0.0835269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_c_359_n 0.0255357f $X=-0.19 $Y=-0.24 $X2=0.395 $Y2=1.165
cc_28 VNB N_VPWR_c_430_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_569_n 0.00765946f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB Y 0.00536016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_761_n 0.015377f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_32 VNB N_A_27_47#_c_762_n 0.00353458f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_33 VNB N_A_27_47#_c_763_n 0.01229f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_34 VNB N_A_27_47#_c_764_n 0.00678264f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_35 VNB N_A_27_47#_c_765_n 0.00275309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_27_47#_c_766_n 0.00114174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_823_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_38 VNB N_VGND_c_824_n 0.00272154f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_39 VNB N_VGND_c_825_n 0.0143703f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_40 VNB N_VGND_c_826_n 0.0134472f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.41
cc_41 VNB N_VGND_c_827_n 0.159402f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=1.105
cc_42 VNB N_VGND_c_828_n 0.417956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_829_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_830_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_45 VNB N_A_485_47#_c_910_n 0.0288293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_883_47#_c_943_n 0.00263528f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_47 VNB N_A_883_47#_c_944_n 0.0100703f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_48 VNB N_A_883_47#_c_945_n 0.0177047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VPB N_D_c_122_n 0.0198486f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_50 VPB N_D_c_123_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_51 VPB N_D_c_124_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_52 VPB N_D_c_125_n 0.0160015f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_53 VPB N_D_c_119_n 0.0080961f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.165
cc_54 VPB N_D_c_120_n 0.028998f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_55 VPB N_C_c_202_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_56 VPB N_C_c_203_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_57 VPB N_C_c_204_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_58 VPB N_C_c_205_n 0.0201049f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_59 VPB N_C_c_201_n 0.0287283f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.16
cc_60 VPB N_B_c_281_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_61 VPB N_B_c_282_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_62 VPB N_B_c_283_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_63 VPB N_B_c_284_n 0.0164193f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_64 VPB N_B_c_280_n 0.0289224f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.217
cc_65 VPB N_A_c_360_n 0.0160739f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_66 VPB N_A_c_361_n 0.0158811f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_67 VPB N_A_c_362_n 0.0158869f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_68 VPB N_A_c_363_n 0.0198539f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_69 VPB N_A_c_358_n 0.0282303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_c_359_n 0.00797922f $X=-0.19 $Y=1.305 $X2=0.395 $Y2=1.165
cc_71 VPB N_VPWR_c_431_n 0.00994749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_432_n 0.0464216f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_73 VPB N_VPWR_c_433_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_434_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.165
cc_75 VPB N_VPWR_c_435_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_76 VPB N_VPWR_c_436_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.217
cc_77 VPB N_VPWR_c_437_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.67 $Y2=1.217
cc_78 VPB N_VPWR_c_438_n 0.00760606f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=1.217
cc_79 VPB N_VPWR_c_439_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.175
cc_80 VPB N_VPWR_c_440_n 0.00474148f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.19
cc_81 VPB N_VPWR_c_441_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.175
cc_82 VPB N_VPWR_c_442_n 0.0137153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_443_n 0.0470546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_444_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_445_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_446_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_447_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_448_n 0.0217546f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_449_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_450_n 0.0214331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_451_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_452_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_453_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_454_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_455_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_456_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_430_n 0.0481532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_571_n 0.00176159f $X=-0.19 $Y=1.305 $X2=1.17 $Y2=1.105
cc_99 VPB N_Y_c_572_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_Y_c_573_n 0.00373025f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_Y_c_574_n 0.00173134f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.217
cc_102 VPB N_Y_c_575_n 0.00821225f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_103 VPB N_Y_c_576_n 0.00173134f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.175
cc_104 VPB N_Y_c_577_n 0.00927763f $X=-0.19 $Y=1.305 $X2=1.615 $Y2=1.19
cc_105 VPB N_Y_c_578_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_Y_c_579_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_Y_c_580_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_Y_c_581_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_582_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_583_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_584_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_Y_c_585_n 0.00213755f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB Y 0.00304907f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 N_D_M1031_g N_C_M1012_g 0.0227918f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_115 N_D_c_125_n N_C_c_202_n 0.0231619f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_116 N_D_c_120_n C 0.00202552f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_117 D C 0.0101544f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_118 N_D_c_120_n N_C_c_201_n 0.0227918f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_119 N_D_c_122_n N_VPWR_c_432_n 0.00871449f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_D_c_119_n N_VPWR_c_432_n 0.00558889f $X=0.395 $Y=1.165 $X2=0 $Y2=0
cc_121 D N_VPWR_c_432_n 0.0194886f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_122 N_D_c_122_n N_VPWR_c_433_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_123 N_D_c_123_n N_VPWR_c_433_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_124 N_D_c_123_n N_VPWR_c_434_n 0.0052072f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_125 N_D_c_124_n N_VPWR_c_434_n 0.004751f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_126 N_D_c_124_n N_VPWR_c_435_n 0.00597712f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_127 N_D_c_125_n N_VPWR_c_435_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_128 N_D_c_125_n N_VPWR_c_436_n 0.0052072f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_129 N_D_c_122_n N_VPWR_c_430_n 0.010906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_130 N_D_c_123_n N_VPWR_c_430_n 0.0118438f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_131 N_D_c_124_n N_VPWR_c_430_n 0.00999457f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_132 N_D_c_125_n N_VPWR_c_430_n 0.011869f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_133 N_D_c_122_n N_Y_c_571_n 0.0046976f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_134 N_D_c_123_n N_Y_c_571_n 0.00116723f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_135 N_D_c_120_n N_Y_c_571_n 0.0074788f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_136 D N_Y_c_571_n 0.0305808f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_137 N_D_c_122_n N_Y_c_591_n 0.0121679f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_D_c_123_n N_Y_c_591_n 0.0106251f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_D_c_124_n N_Y_c_591_n 6.24674e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_140 N_D_c_123_n N_Y_c_572_n 0.0153933f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_D_c_124_n N_Y_c_572_n 0.0113962f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_D_c_120_n N_Y_c_572_n 0.00725062f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_143 D N_Y_c_572_n 0.040258f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_144 N_D_c_123_n N_Y_c_598_n 6.48386e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_D_c_124_n N_Y_c_598_n 0.0130707f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_D_c_125_n N_Y_c_598_n 0.0106251f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_147 N_D_c_125_n N_Y_c_573_n 0.0172899f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_148 N_D_c_120_n N_Y_c_573_n 3.62813e-19 $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_149 N_D_c_125_n N_Y_c_603_n 6.48386e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_150 N_D_c_124_n N_Y_c_580_n 0.00292783f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_151 N_D_c_125_n N_Y_c_580_n 0.00116723f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_152 N_D_c_120_n N_Y_c_580_n 0.0074788f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_153 D N_Y_c_580_n 0.0305808f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_154 N_D_M1002_g N_A_27_47#_c_761_n 0.00730084f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_155 N_D_M1002_g N_A_27_47#_c_762_n 0.0133303f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_156 N_D_M1022_g N_A_27_47#_c_762_n 0.0134984f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_157 N_D_c_119_n N_A_27_47#_c_762_n 0.00251219f $X=0.395 $Y=1.165 $X2=0 $Y2=0
cc_158 N_D_c_120_n N_A_27_47#_c_762_n 0.00322716f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_159 D N_A_27_47#_c_762_n 0.0561869f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_160 N_D_c_119_n N_A_27_47#_c_763_n 0.00573234f $X=0.395 $Y=1.165 $X2=0 $Y2=0
cc_161 D N_A_27_47#_c_763_n 0.0194942f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_162 N_D_M1023_g N_A_27_47#_c_775_n 0.004499f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_163 N_D_M1023_g N_A_27_47#_c_764_n 0.0126116f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_164 N_D_M1031_g N_A_27_47#_c_764_n 0.0149379f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_165 N_D_c_120_n N_A_27_47#_c_764_n 0.00345502f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_166 D N_A_27_47#_c_764_n 0.0404306f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_167 N_D_c_120_n N_A_27_47#_c_766_n 0.00308294f $X=1.905 $Y=1.217 $X2=0 $Y2=0
cc_168 D N_A_27_47#_c_766_n 0.0138098f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_169 N_D_M1002_g N_VGND_c_823_n 0.0115037f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_170 N_D_M1022_g N_VGND_c_823_n 0.00162962f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_171 N_D_M1022_g N_VGND_c_824_n 6.16486e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_172 N_D_M1023_g N_VGND_c_824_n 0.00988033f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_173 N_D_M1031_g N_VGND_c_824_n 0.00317372f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_174 N_D_M1002_g N_VGND_c_825_n 0.00199015f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_175 N_D_M1022_g N_VGND_c_826_n 0.00428022f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_176 N_D_M1023_g N_VGND_c_826_n 0.00199015f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_177 N_D_M1031_g N_VGND_c_827_n 0.00428022f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_178 N_D_M1002_g N_VGND_c_828_n 0.00369362f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_179 N_D_M1022_g N_VGND_c_828_n 0.005943f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_180 N_D_M1023_g N_VGND_c_828_n 0.00278819f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_181 N_D_M1031_g N_VGND_c_828_n 0.00583939f $X=1.93 $Y=0.56 $X2=0 $Y2=0
cc_182 C N_B_c_278_n 7.55054e-19 $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_183 N_C_c_201_n N_B_c_278_n 0.00741568f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_184 C N_B_c_279_n 0.0152145f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_185 N_C_c_201_n N_B_c_279_n 6.88356e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_186 N_C_c_202_n N_VPWR_c_436_n 0.004751f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_187 N_C_c_203_n N_VPWR_c_437_n 0.0052072f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_188 N_C_c_204_n N_VPWR_c_437_n 0.004751f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_189 N_C_c_205_n N_VPWR_c_438_n 0.00825342f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_190 N_C_c_202_n N_VPWR_c_444_n 0.00597712f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_191 N_C_c_203_n N_VPWR_c_444_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_192 N_C_c_204_n N_VPWR_c_452_n 0.00597712f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_193 N_C_c_205_n N_VPWR_c_452_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_194 N_C_c_202_n N_VPWR_c_430_n 0.0100198f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_195 N_C_c_203_n N_VPWR_c_430_n 0.0118438f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_196 N_C_c_204_n N_VPWR_c_430_n 0.00999457f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_197 N_C_c_205_n N_VPWR_c_430_n 0.0131262f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_198 N_C_c_202_n N_Y_c_598_n 6.24674e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_199 N_C_c_202_n N_Y_c_573_n 0.0113403f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_200 C N_Y_c_573_n 0.0150129f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_201 N_C_c_201_n N_Y_c_573_n 3.10838e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_202 N_C_c_202_n N_Y_c_603_n 0.0130707f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_203 N_C_c_203_n N_Y_c_603_n 0.0106251f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_204 N_C_c_204_n N_Y_c_603_n 6.24674e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_205 N_C_c_203_n N_Y_c_574_n 0.0153933f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_206 N_C_c_204_n N_Y_c_574_n 0.0113962f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_207 C N_Y_c_574_n 0.040258f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_208 N_C_c_201_n N_Y_c_574_n 0.00725062f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_209 N_C_c_203_n N_Y_c_619_n 6.48386e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_210 N_C_c_204_n N_Y_c_619_n 0.0130707f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_211 N_C_c_205_n N_Y_c_619_n 0.0153658f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_212 N_C_c_205_n N_Y_c_575_n 0.0179883f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_213 C N_Y_c_575_n 0.0227895f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_214 N_C_c_201_n N_Y_c_575_n 3.10838e-19 $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_215 N_C_c_202_n N_Y_c_581_n 0.00292783f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_216 N_C_c_203_n N_Y_c_581_n 0.00116723f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_217 C N_Y_c_581_n 0.0305808f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_218 N_C_c_201_n N_Y_c_581_n 0.0074788f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_219 N_C_c_204_n N_Y_c_582_n 0.00292783f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_220 N_C_c_205_n N_Y_c_582_n 0.00116723f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_221 C N_Y_c_582_n 0.0305808f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_222 N_C_c_201_n N_Y_c_582_n 0.00723098f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_223 N_C_M1012_g N_A_27_47#_c_764_n 4.48192e-19 $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_224 C N_A_27_47#_c_764_n 0.00297817f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_225 N_C_M1012_g N_A_27_47#_c_765_n 0.0127488f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_226 N_C_M1018_g N_A_27_47#_c_765_n 0.00951434f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_227 N_C_M1025_g N_A_27_47#_c_765_n 0.00994068f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_228 N_C_M1027_g N_A_27_47#_c_765_n 0.00994068f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_229 C N_A_27_47#_c_765_n 0.00381697f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_230 N_C_M1012_g N_VGND_c_827_n 0.00357877f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_231 N_C_M1018_g N_VGND_c_827_n 0.00357877f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_232 N_C_M1025_g N_VGND_c_827_n 0.00357877f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_233 N_C_M1027_g N_VGND_c_827_n 0.00357877f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_234 N_C_M1012_g N_VGND_c_828_n 0.00542415f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_235 N_C_M1018_g N_VGND_c_828_n 0.00548399f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_236 N_C_M1025_g N_VGND_c_828_n 0.00560377f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_237 N_C_M1027_g N_VGND_c_828_n 0.00680287f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_238 N_C_M1012_g N_A_485_47#_c_910_n 0.00365114f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_239 N_C_M1018_g N_A_485_47#_c_910_n 0.0111698f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_240 N_C_M1025_g N_A_485_47#_c_910_n 0.0111976f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_241 N_C_M1027_g N_A_485_47#_c_910_n 0.0138648f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_242 C N_A_485_47#_c_910_n 0.120337f $X=3.72 $Y=1.105 $X2=0 $Y2=0
cc_243 N_C_c_201_n N_A_485_47#_c_910_n 0.010834f $X=3.785 $Y=1.217 $X2=0 $Y2=0
cc_244 N_B_M1021_g N_A_M1008_g 0.0171433f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B_c_284_n N_A_c_360_n 0.0180767f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_280_n N_A_c_358_n 0.0171433f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_247 N_B_c_281_n N_VPWR_c_438_n 0.00762417f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_282_n N_VPWR_c_439_n 0.0052072f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_283_n N_VPWR_c_439_n 0.004751f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_284_n N_VPWR_c_440_n 0.00523168f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_251 N_B_c_281_n N_VPWR_c_446_n 0.00597712f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_252 N_B_c_282_n N_VPWR_c_446_n 0.00673617f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_283_n N_VPWR_c_448_n 0.00597712f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_284_n N_VPWR_c_448_n 0.00673617f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_281_n N_VPWR_c_430_n 0.0112769f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_282_n N_VPWR_c_430_n 0.0118438f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_283_n N_VPWR_c_430_n 0.00999457f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_284_n N_VPWR_c_430_n 0.0120928f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B_c_281_n N_Y_c_575_n 0.0139912f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B_c_278_n N_Y_c_575_n 0.00729564f $X=4.675 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B_c_279_n N_Y_c_575_n 0.0401373f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_262 N_B_c_280_n N_Y_c_575_n 2.73568e-19 $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_263 N_B_c_281_n N_Y_c_637_n 0.0178402f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B_c_282_n N_Y_c_637_n 0.0106251f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B_c_283_n N_Y_c_637_n 6.24674e-19 $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_282_n N_Y_c_576_n 0.0153933f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B_c_283_n N_Y_c_576_n 0.0113962f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B_c_279_n N_Y_c_576_n 0.040258f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B_c_280_n N_Y_c_576_n 0.00725062f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_270 N_B_c_282_n N_Y_c_644_n 6.48386e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B_c_283_n N_Y_c_644_n 0.0130707f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B_c_284_n N_Y_c_644_n 0.0114282f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B_c_284_n N_Y_c_577_n 0.0207993f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_280_n N_Y_c_577_n 4.93319e-19 $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_275 N_B_c_284_n N_Y_c_649_n 6.5624e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B_M1021_g N_Y_c_650_n 0.00231614f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_277 N_B_c_281_n N_Y_c_583_n 0.00292783f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B_c_282_n N_Y_c_583_n 0.00116723f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_279_n N_Y_c_583_n 0.0305808f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B_c_280_n N_Y_c_583_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_281 N_B_c_283_n N_Y_c_584_n 0.00292783f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B_c_284_n N_Y_c_584_n 0.00116723f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B_c_279_n N_Y_c_584_n 0.0305808f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_284 N_B_c_280_n N_Y_c_584_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_285 N_B_c_284_n Y 7.1348e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B_M1021_g Y 0.00838538f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_287 N_B_c_279_n Y 0.00815753f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_288 N_B_M1005_g N_VGND_c_827_n 0.00357877f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_289 N_B_M1007_g N_VGND_c_827_n 0.00357877f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_290 N_B_M1015_g N_VGND_c_827_n 0.00357877f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_291 N_B_M1021_g N_VGND_c_827_n 0.00357877f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_292 N_B_M1005_g N_VGND_c_828_n 0.00668309f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_293 N_B_M1007_g N_VGND_c_828_n 0.00548399f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_294 N_B_M1015_g N_VGND_c_828_n 0.00548399f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_295 N_B_M1021_g N_VGND_c_828_n 0.00552482f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_296 N_B_M1005_g N_A_485_47#_c_910_n 0.013837f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_297 N_B_M1007_g N_A_485_47#_c_910_n 0.0111698f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_298 N_B_M1015_g N_A_485_47#_c_910_n 0.0111333f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_299 N_B_M1021_g N_A_485_47#_c_910_n 2.64848e-19 $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_300 N_B_c_278_n N_A_485_47#_c_910_n 0.00896085f $X=4.675 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B_c_279_n N_A_485_47#_c_910_n 0.137788f $X=5.95 $Y=1.16 $X2=0 $Y2=0
cc_302 N_B_c_280_n N_A_485_47#_c_910_n 0.00968149f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_303 N_B_M1005_g N_A_883_47#_c_943_n 0.00958923f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_304 N_B_M1007_g N_A_883_47#_c_943_n 0.00958923f $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_305 N_B_M1015_g N_A_883_47#_c_943_n 0.00958923f $X=5.74 $Y=0.56 $X2=0 $Y2=0
cc_306 N_B_M1021_g N_A_883_47#_c_943_n 0.0143475f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_c_360_n N_VPWR_c_440_n 0.00482668f $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A_c_361_n N_VPWR_c_441_n 0.0052072f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_c_362_n N_VPWR_c_441_n 0.004751f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_c_363_n N_VPWR_c_443_n 0.00955005f $X=8.125 $Y=1.41 $X2=0 $Y2=0
cc_311 A N_VPWR_c_443_n 0.0190809f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_312 N_A_c_359_n N_VPWR_c_443_n 0.00547197f $X=8.345 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_c_360_n N_VPWR_c_450_n 0.00597712f $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_c_361_n N_VPWR_c_450_n 0.00673617f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_315 N_A_c_362_n N_VPWR_c_453_n 0.00597712f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_c_363_n N_VPWR_c_453_n 0.00673617f $X=8.125 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_c_360_n N_VPWR_c_430_n 0.0102184f $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_c_361_n N_VPWR_c_430_n 0.0118438f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_c_362_n N_VPWR_c_430_n 0.00999457f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A_c_363_n N_VPWR_c_430_n 0.0128492f $X=8.125 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A_c_360_n N_Y_c_644_n 6.36264e-19 $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_c_360_n N_Y_c_649_n 0.0137121f $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_c_361_n N_Y_c_649_n 0.0106251f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A_c_362_n N_Y_c_649_n 6.24674e-19 $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A_M1008_g N_Y_c_650_n 0.00746826f $X=6.69 $Y=0.56 $X2=0 $Y2=0
cc_326 N_A_M1010_g N_Y_c_569_n 0.0114825f $X=7.16 $Y=0.56 $X2=0 $Y2=0
cc_327 N_A_M1024_g N_Y_c_569_n 0.0111698f $X=7.63 $Y=0.56 $X2=0 $Y2=0
cc_328 N_A_M1026_g N_Y_c_569_n 0.00411914f $X=8.1 $Y=0.56 $X2=0 $Y2=0
cc_329 A N_Y_c_569_n 0.0689943f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_330 N_A_c_358_n N_Y_c_569_n 0.0103204f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_331 N_A_c_361_n N_Y_c_578_n 0.0153933f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A_c_362_n N_Y_c_578_n 0.0113962f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_333 A N_Y_c_578_n 0.040258f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_334 N_A_c_358_n N_Y_c_578_n 0.00725062f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_335 N_A_c_362_n N_Y_c_579_n 0.00292783f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_336 N_A_c_363_n N_Y_c_579_n 0.00349846f $X=8.125 $Y=1.41 $X2=0 $Y2=0
cc_337 A N_Y_c_579_n 0.0305808f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_338 N_A_c_358_n N_Y_c_579_n 0.0074788f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_339 N_A_c_361_n N_Y_c_680_n 6.48386e-19 $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_340 N_A_c_362_n N_Y_c_680_n 0.0130707f $X=7.655 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_c_363_n N_Y_c_680_n 0.0100147f $X=8.125 $Y=1.41 $X2=0 $Y2=0
cc_342 N_A_c_360_n N_Y_c_585_n 0.0129747f $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_c_361_n N_Y_c_585_n 0.00137869f $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_c_358_n N_Y_c_585_n 0.00838779f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_345 N_A_M1008_g Y 0.00308843f $X=6.69 $Y=0.56 $X2=0 $Y2=0
cc_346 N_A_c_360_n Y 9.13911e-19 $X=6.715 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_M1010_g Y 0.00247878f $X=7.16 $Y=0.56 $X2=0 $Y2=0
cc_348 N_A_c_361_n Y 6.95088e-19 $X=7.185 $Y=1.41 $X2=0 $Y2=0
cc_349 A Y 0.010172f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_350 N_A_c_358_n Y 0.0203356f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_351 N_A_M1008_g N_VGND_c_827_n 0.00357877f $X=6.69 $Y=0.56 $X2=0 $Y2=0
cc_352 N_A_M1010_g N_VGND_c_827_n 0.00357877f $X=7.16 $Y=0.56 $X2=0 $Y2=0
cc_353 N_A_M1024_g N_VGND_c_827_n 0.00357877f $X=7.63 $Y=0.56 $X2=0 $Y2=0
cc_354 N_A_M1026_g N_VGND_c_827_n 0.00357877f $X=8.1 $Y=0.56 $X2=0 $Y2=0
cc_355 N_A_M1008_g N_VGND_c_828_n 0.00552482f $X=6.69 $Y=0.56 $X2=0 $Y2=0
cc_356 N_A_M1010_g N_VGND_c_828_n 0.00548399f $X=7.16 $Y=0.56 $X2=0 $Y2=0
cc_357 N_A_M1024_g N_VGND_c_828_n 0.00548399f $X=7.63 $Y=0.56 $X2=0 $Y2=0
cc_358 N_A_M1026_g N_VGND_c_828_n 0.00643908f $X=8.1 $Y=0.56 $X2=0 $Y2=0
cc_359 N_A_M1008_g N_A_883_47#_c_943_n 0.00958301f $X=6.69 $Y=0.56 $X2=0 $Y2=0
cc_360 N_A_M1010_g N_A_883_47#_c_943_n 0.00958923f $X=7.16 $Y=0.56 $X2=0 $Y2=0
cc_361 N_A_M1024_g N_A_883_47#_c_943_n 0.00958923f $X=7.63 $Y=0.56 $X2=0 $Y2=0
cc_362 N_A_M1026_g N_A_883_47#_c_943_n 0.0112037f $X=8.1 $Y=0.56 $X2=0 $Y2=0
cc_363 A N_A_883_47#_c_943_n 0.00486515f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_364 N_A_c_358_n N_A_883_47#_c_943_n 0.00160151f $X=8.225 $Y=1.165 $X2=0 $Y2=0
cc_365 N_A_M1026_g N_A_883_47#_c_945_n 0.00474438f $X=8.1 $Y=0.56 $X2=0 $Y2=0
cc_366 A N_A_883_47#_c_945_n 0.0190066f $X=8.3 $Y=1.105 $X2=0 $Y2=0
cc_367 N_A_c_359_n N_A_883_47#_c_945_n 0.00558895f $X=8.345 $Y=1.16 $X2=0 $Y2=0
cc_368 N_VPWR_c_430_n N_Y_M1001_s 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_369 N_VPWR_c_430_n N_Y_M1020_s 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_370 N_VPWR_c_430_n N_Y_M1000_s 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_371 N_VPWR_c_430_n N_Y_M1011_s 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_372 N_VPWR_c_430_n N_Y_M1003_d 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_373 N_VPWR_c_430_n N_Y_M1019_d 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_374 N_VPWR_c_430_n N_Y_M1004_d 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_375 N_VPWR_c_430_n N_Y_M1016_d 0.00231261f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_432_n N_Y_c_571_n 0.0178509f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_377 N_VPWR_c_432_n N_Y_c_591_n 0.0615045f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_378 N_VPWR_c_433_n N_Y_c_591_n 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_379 N_VPWR_c_434_n N_Y_c_591_n 0.0385613f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_380 N_VPWR_c_430_n N_Y_c_591_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_M1014_d N_Y_c_572_n 0.00180012f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_382 N_VPWR_c_434_n N_Y_c_572_n 0.0139097f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_383 N_VPWR_c_434_n N_Y_c_598_n 0.0470327f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_384 N_VPWR_c_435_n N_Y_c_598_n 0.0223557f $X=2.055 $Y=2.72 $X2=0 $Y2=0
cc_385 N_VPWR_c_436_n N_Y_c_598_n 0.0385613f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_386 N_VPWR_c_430_n N_Y_c_598_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_M1028_d N_Y_c_573_n 0.00180012f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_388 N_VPWR_c_436_n N_Y_c_573_n 0.0139097f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_389 N_VPWR_c_436_n N_Y_c_603_n 0.0470327f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_390 N_VPWR_c_437_n N_Y_c_603_n 0.0385613f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_391 N_VPWR_c_444_n N_Y_c_603_n 0.0223557f $X=2.995 $Y=2.72 $X2=0 $Y2=0
cc_392 N_VPWR_c_430_n N_Y_c_603_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_M1006_d N_Y_c_574_n 0.00180012f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_394 N_VPWR_c_437_n N_Y_c_574_n 0.0139097f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_395 N_VPWR_c_437_n N_Y_c_619_n 0.0470327f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_438_n N_Y_c_619_n 0.0429581f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_397 N_VPWR_c_452_n N_Y_c_619_n 0.0223557f $X=3.935 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_430_n N_Y_c_619_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_M1017_d N_Y_c_575_n 0.0118304f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_400 N_VPWR_c_438_n N_Y_c_575_n 0.0569634f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_401 N_VPWR_c_438_n N_Y_c_637_n 0.0523533f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_402 N_VPWR_c_439_n N_Y_c_637_n 0.0385613f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_446_n N_Y_c_637_n 0.0223557f $X=5.395 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_430_n N_Y_c_637_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1009_s N_Y_c_576_n 0.00180012f $X=5.335 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_c_439_n N_Y_c_576_n 0.0139097f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_407 N_VPWR_c_439_n N_Y_c_644_n 0.0470327f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_c_440_n N_Y_c_644_n 0.0344369f $X=6.455 $Y=2 $X2=0 $Y2=0
cc_409 N_VPWR_c_448_n N_Y_c_644_n 0.0223557f $X=6.37 $Y=2.72 $X2=0 $Y2=0
cc_410 N_VPWR_c_430_n N_Y_c_644_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_411 N_VPWR_M1029_s N_Y_c_577_n 0.00353218f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_412 N_VPWR_c_440_n N_Y_c_577_n 0.0139097f $X=6.455 $Y=2 $X2=0 $Y2=0
cc_413 N_VPWR_c_440_n N_Y_c_649_n 0.0423054f $X=6.455 $Y=2 $X2=0 $Y2=0
cc_414 N_VPWR_c_441_n N_Y_c_649_n 0.0385613f $X=7.42 $Y=2 $X2=0 $Y2=0
cc_415 N_VPWR_c_450_n N_Y_c_649_n 0.0223557f $X=7.335 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_430_n N_Y_c_649_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_M1013_s N_Y_c_578_n 0.00180012f $X=7.275 $Y=1.485 $X2=0 $Y2=0
cc_418 N_VPWR_c_441_n N_Y_c_578_n 0.0139097f $X=7.42 $Y=2 $X2=0 $Y2=0
cc_419 N_VPWR_c_443_n N_Y_c_579_n 0.0146524f $X=8.36 $Y=1.66 $X2=0 $Y2=0
cc_420 N_VPWR_c_441_n N_Y_c_680_n 0.0470327f $X=7.42 $Y=2 $X2=0 $Y2=0
cc_421 N_VPWR_c_443_n N_Y_c_680_n 0.0505127f $X=8.36 $Y=1.66 $X2=0 $Y2=0
cc_422 N_VPWR_c_453_n N_Y_c_680_n 0.0223557f $X=8.275 $Y=2.72 $X2=0 $Y2=0
cc_423 N_VPWR_c_430_n N_Y_c_680_n 0.0140101f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_M1029_s N_Y_c_585_n 0.00103754f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_425 N_VPWR_c_432_n N_A_27_47#_c_763_n 5.83538e-19 $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_426 N_VPWR_c_443_n N_A_883_47#_c_945_n 7.91944e-19 $X=8.36 $Y=1.66 $X2=0
+ $Y2=0
cc_427 N_Y_c_573_n N_A_27_47#_c_764_n 0.0117299f $X=2.395 $Y=1.555 $X2=0 $Y2=0
cc_428 N_Y_M1008_s N_VGND_c_828_n 0.00256987f $X=6.765 $Y=0.235 $X2=0 $Y2=0
cc_429 N_Y_M1024_s N_VGND_c_828_n 0.00256987f $X=7.705 $Y=0.235 $X2=0 $Y2=0
cc_430 N_Y_c_575_n N_A_485_47#_c_910_n 0.00798715f $X=4.795 $Y=1.555 $X2=0 $Y2=0
cc_431 N_Y_c_650_n N_A_485_47#_c_910_n 0.00607984f $X=6.825 $Y=0.78 $X2=0 $Y2=0
cc_432 N_Y_c_650_n N_A_883_47#_M1021_d 0.00320255f $X=6.825 $Y=0.78 $X2=0 $Y2=0
cc_433 N_Y_c_569_n N_A_883_47#_M1010_d 0.00214463f $X=7.89 $Y=0.74 $X2=0 $Y2=0
cc_434 N_Y_M1008_s N_A_883_47#_c_943_n 0.00398513f $X=6.765 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1024_s N_A_883_47#_c_943_n 0.00401739f $X=7.705 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_c_650_n N_A_883_47#_c_943_n 0.0122599f $X=6.825 $Y=0.78 $X2=0 $Y2=0
cc_437 N_Y_c_569_n N_A_883_47#_c_943_n 0.0670225f $X=7.89 $Y=0.74 $X2=0 $Y2=0
cc_438 N_Y_c_569_n N_A_883_47#_c_945_n 0.016455f $X=7.89 $Y=0.74 $X2=0 $Y2=0
cc_439 N_A_27_47#_c_762_n N_VGND_M1002_s 0.00213962f $X=1.115 $Y=0.78 $X2=-0.19
+ $Y2=-0.24
cc_440 N_A_27_47#_c_764_n N_VGND_M1023_s 0.00213962f $X=2.055 $Y=0.78 $X2=0
+ $Y2=0
cc_441 N_A_27_47#_c_761_n N_VGND_c_823_n 0.0176937f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_442 N_A_27_47#_c_762_n N_VGND_c_823_n 0.0220033f $X=1.115 $Y=0.78 $X2=0 $Y2=0
cc_443 N_A_27_47#_c_775_n N_VGND_c_824_n 0.0171708f $X=1.2 $Y=0.655 $X2=0 $Y2=0
cc_444 N_A_27_47#_c_764_n N_VGND_c_824_n 0.0220033f $X=2.055 $Y=0.78 $X2=0 $Y2=0
cc_445 N_A_27_47#_c_761_n N_VGND_c_825_n 0.0177923f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_446 N_A_27_47#_c_762_n N_VGND_c_825_n 0.00236597f $X=1.115 $Y=0.78 $X2=0
+ $Y2=0
cc_447 N_A_27_47#_c_762_n N_VGND_c_826_n 0.00303619f $X=1.115 $Y=0.78 $X2=0
+ $Y2=0
cc_448 N_A_27_47#_c_775_n N_VGND_c_826_n 0.0115672f $X=1.2 $Y=0.655 $X2=0 $Y2=0
cc_449 N_A_27_47#_c_764_n N_VGND_c_826_n 0.00236597f $X=2.055 $Y=0.78 $X2=0
+ $Y2=0
cc_450 N_A_27_47#_c_764_n N_VGND_c_827_n 0.00303619f $X=2.055 $Y=0.78 $X2=0
+ $Y2=0
cc_451 N_A_27_47#_c_803_p N_VGND_c_827_n 0.0114305f $X=2.225 $Y=0.37 $X2=0 $Y2=0
cc_452 N_A_27_47#_c_765_n N_VGND_c_827_n 0.112394f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_453 N_A_27_47#_M1002_d N_VGND_c_828_n 0.00292228f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_454 N_A_27_47#_M1022_d N_VGND_c_828_n 0.00316288f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_455 N_A_27_47#_M1031_d N_VGND_c_828_n 0.00236502f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_456 N_A_27_47#_M1018_d N_VGND_c_828_n 0.00255381f $X=2.895 $Y=0.235 $X2=0
+ $Y2=0
cc_457 N_A_27_47#_M1027_d N_VGND_c_828_n 0.00209344f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_458 N_A_27_47#_c_761_n N_VGND_c_828_n 0.00973192f $X=0.217 $Y=0.655 $X2=0
+ $Y2=0
cc_459 N_A_27_47#_c_762_n N_VGND_c_828_n 0.0115443f $X=1.115 $Y=0.78 $X2=0 $Y2=0
cc_460 N_A_27_47#_c_775_n N_VGND_c_828_n 0.0064623f $X=1.2 $Y=0.655 $X2=0 $Y2=0
cc_461 N_A_27_47#_c_764_n N_VGND_c_828_n 0.0115443f $X=2.055 $Y=0.78 $X2=0 $Y2=0
cc_462 N_A_27_47#_c_803_p N_VGND_c_828_n 0.00653924f $X=2.225 $Y=0.37 $X2=0
+ $Y2=0
cc_463 N_A_27_47#_c_765_n N_VGND_c_828_n 0.070531f $X=4.02 $Y=0.4 $X2=0 $Y2=0
cc_464 N_A_27_47#_c_765_n N_A_485_47#_M1012_s 0.00401739f $X=4.02 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_465 N_A_27_47#_c_765_n N_A_485_47#_M1025_s 0.00510139f $X=4.02 $Y=0.4 $X2=0
+ $Y2=0
cc_466 N_A_27_47#_M1018_d N_A_485_47#_c_910_n 0.00214463f $X=2.895 $Y=0.235
+ $X2=0 $Y2=0
cc_467 N_A_27_47#_M1027_d N_A_485_47#_c_910_n 0.00312742f $X=3.885 $Y=0.235
+ $X2=0 $Y2=0
cc_468 N_A_27_47#_c_764_n N_A_485_47#_c_910_n 0.0113394f $X=2.055 $Y=0.78 $X2=0
+ $Y2=0
cc_469 N_A_27_47#_c_765_n N_A_485_47#_c_910_n 0.0988536f $X=4.02 $Y=0.4 $X2=0
+ $Y2=0
cc_470 N_A_27_47#_c_765_n N_A_883_47#_c_943_n 0.0197364f $X=4.02 $Y=0.4 $X2=0
+ $Y2=0
cc_471 N_VGND_c_828_n N_A_485_47#_M1012_s 0.00256987f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_472 N_VGND_c_828_n N_A_485_47#_M1025_s 0.00297142f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_473 N_VGND_c_828_n N_A_485_47#_M1005_s 0.00256987f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_474 N_VGND_c_828_n N_A_485_47#_M1015_s 0.00256987f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_475 N_VGND_c_827_n N_A_485_47#_c_910_n 0.00342407f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_476 N_VGND_c_828_n N_A_485_47#_c_910_n 0.0121765f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_477 N_VGND_c_828_n N_A_883_47#_M1005_d 0.00250339f $X=8.51 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_478 N_VGND_c_828_n N_A_883_47#_M1007_d 0.00255381f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_479 N_VGND_c_828_n N_A_883_47#_M1021_d 0.00263412f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_480 N_VGND_c_828_n N_A_883_47#_M1010_d 0.00255381f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_481 N_VGND_c_828_n N_A_883_47#_M1026_d 0.00250318f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_482 N_VGND_c_827_n N_A_883_47#_c_943_n 0.222953f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_483 N_VGND_c_828_n N_A_883_47#_c_943_n 0.140176f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_484 N_VGND_c_827_n N_A_883_47#_c_944_n 0.0179343f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_485 N_VGND_c_828_n N_A_883_47#_c_944_n 0.00980895f $X=8.51 $Y=0 $X2=0 $Y2=0
cc_486 N_A_485_47#_c_910_n N_A_883_47#_M1005_d 0.00428172f $X=5.95 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_487 N_A_485_47#_c_910_n N_A_883_47#_M1007_d 0.00214463f $X=5.95 $Y=0.74 $X2=0
+ $Y2=0
cc_488 N_A_485_47#_M1005_s N_A_883_47#_c_943_n 0.00401739f $X=4.875 $Y=0.235
+ $X2=0 $Y2=0
cc_489 N_A_485_47#_M1015_s N_A_883_47#_c_943_n 0.00401739f $X=5.815 $Y=0.235
+ $X2=0 $Y2=0
cc_490 N_A_485_47#_c_910_n N_A_883_47#_c_943_n 0.0968451f $X=5.95 $Y=0.74 $X2=0
+ $Y2=0
