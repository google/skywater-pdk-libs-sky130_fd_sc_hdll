* File: sky130_fd_sc_hdll__and2b_1.pex.spice
* Created: Thu Aug 27 18:57:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%A_N 2 3 5 8 10 11 12 17
c35 17 0 1.89169e-19 $X=0.36 $Y=1.16
r36 17 20 36.8359 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=1.325
r37 17 19 45.6753 $w=4e-07 $l=1.65e-07 $layer=POLY_cond $X=0.395 $Y=1.16
+ $X2=0.395 $Y2=0.995
r38 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.36
+ $Y=1.16 $X2=0.36 $Y2=1.16
r39 11 12 13.061 $w=2.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.53
r40 11 18 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=0.295 $Y=1.19
+ $X2=0.295 $Y2=1.16
r41 10 18 11.9086 $w=2.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.295 $Y=0.85
+ $X2=0.295 $Y2=1.16
r42 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.445
+ $X2=0.52 $Y2=0.995
r43 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r44 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r45 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%A_27_413# 1 2 8 9 11 12 16 20 22 23 25 27
+ 29 36 42
c71 36 0 1.14278e-19 $X=1.115 $Y=0.97
c72 22 0 2.5987e-19 $X=0.665 $Y=1.9
c73 12 0 1.56867e-21 $X=1.485 $Y=0.88
c74 8 0 1.63204e-19 $X=1.035 $Y=1.89
r75 37 42 54.9546 $w=3.3e-07 $l=2.15e-07 $layer=POLY_cond $X=1.115 $Y=0.97
+ $X2=1.33 $Y2=0.97
r76 37 39 13.9889 $w=3.3e-07 $l=8e-08 $layer=POLY_cond $X=1.115 $Y=0.97
+ $X2=1.035 $Y2=0.97
r77 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.115
+ $Y=0.97 $X2=1.115 $Y2=0.97
r78 34 36 11.6292 $w=3.28e-07 $l=3.33e-07 $layer=LI1_cond $X=0.782 $Y=0.97
+ $X2=1.115 $Y2=0.97
r79 32 34 0.244458 $w=3.28e-07 $l=7e-09 $layer=LI1_cond $X=0.775 $Y=0.97
+ $X2=0.782 $Y2=0.97
r80 29 31 10.1849 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.765 $Y=0.445
+ $X2=0.765 $Y2=0.655
r81 26 34 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.782 $Y=1.135
+ $X2=0.782 $Y2=0.97
r82 26 27 31.8761 $w=2.33e-07 $l=6.5e-07 $layer=LI1_cond $X=0.782 $Y=1.135
+ $X2=0.782 $Y2=1.785
r83 25 32 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=0.97
r84 25 31 7.85757 $w=2.18e-07 $l=1.5e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=0.655
r85 22 27 6.81752 $w=2.3e-07 $l=1.64754e-07 $layer=LI1_cond $X=0.665 $Y=1.9
+ $X2=0.782 $Y2=1.785
r86 22 23 16.034 $w=2.28e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=1.9
+ $X2=0.345 $Y2=1.9
r87 18 23 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.345 $Y2=1.9
r88 18 20 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=2.225
r89 14 16 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.56 $Y=0.805
+ $X2=1.56 $Y2=0.445
r90 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.485 $Y=0.88
+ $X2=1.56 $Y2=0.805
r91 12 42 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=1.485 $Y=0.88
+ $X2=1.33 $Y2=0.88
r92 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.035 $Y=1.99
+ $X2=1.035 $Y2=2.275
r93 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.035 $Y=1.89 $X2=1.035
+ $Y2=1.99
r94 7 39 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.035 $Y=1.135
+ $X2=1.035 $Y2=0.97
r95 7 8 250.341 $w=2e-07 $l=7.55e-07 $layer=POLY_cond $X=1.035 $Y=1.135
+ $X2=1.035 $Y2=1.89
r96 2 20 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.225
r97 1 29 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%B 1 3 6 8
c31 8 0 1.64772e-19 $X=2.07 $Y=1.87
c32 6 0 1.14278e-19 $X=2 $Y=0.445
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.795
+ $Y=1.73 $X2=1.795 $Y2=1.73
r34 8 12 10.2233 $w=3.08e-07 $l=2.75e-07 $layer=LI1_cond $X=2.07 $Y=1.8
+ $X2=1.795 $Y2=1.8
r35 4 11 81.5239 $w=4.81e-07 $l=6.78583e-07 $layer=POLY_cond $X=2 $Y=1.165
+ $X2=1.75 $Y2=1.73
r36 4 6 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2 $Y=1.165 $X2=2
+ $Y2=0.445
r37 1 11 45.8146 $w=4.81e-07 $l=3.55106e-07 $layer=POLY_cond $X=1.525 $Y=1.99
+ $X2=1.75 $Y2=1.73
r38 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.525 $Y=1.99
+ $X2=1.525 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%A_225_413# 1 2 7 9 10 12 15 18 19 21 27
r61 27 28 11.0909 $w=2.53e-07 $l=2.3e-07 $layer=LI1_cond $X=1.3 $Y=0.44 $X2=1.53
+ $Y2=0.44
r62 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.42
+ $Y=1.16 $X2=2.42 $Y2=1.16
r63 19 25 16.6301 $w=4.05e-07 $l=5.86302e-07 $layer=LI1_cond $X=2.08 $Y=1.135
+ $X2=1.53 $Y2=1.21
r64 19 21 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=2.08 $Y=1.135
+ $X2=2.42 $Y2=1.135
r65 18 25 4.30998 $w=2.2e-07 $l=2.65e-07 $layer=LI1_cond $X=1.53 $Y=0.945
+ $X2=1.53 $Y2=1.21
r66 17 28 1.55539 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=1.53 $Y=0.61 $X2=1.53
+ $Y2=0.44
r67 17 18 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.53 $Y=0.61
+ $X2=1.53 $Y2=0.945
r68 13 25 8.82617 $w=4.05e-07 $l=4.04344e-07 $layer=LI1_cond $X=1.237 $Y=1.475
+ $X2=1.53 $Y2=1.21
r69 13 15 25.801 $w=3.33e-07 $l=7.5e-07 $layer=LI1_cond $X=1.237 $Y=1.475
+ $X2=1.237 $Y2=2.225
r70 10 22 40.1245 $w=3.04e-07 $l=2.15349e-07 $layer=POLY_cond $X=2.54 $Y=0.985
+ $X2=2.45 $Y2=1.16
r71 10 12 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.54 $Y=0.985
+ $X2=2.54 $Y2=0.56
r72 7 22 47.5924 $w=3.04e-07 $l=2.80624e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.45 $Y2=1.16
r73 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.515 $Y=1.41
+ $X2=2.515 $Y2=1.985
r74 2 15 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=2.065 $X2=1.28 $Y2=2.225
r75 1 27 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%VPWR 1 2 9 11 13 25 26 29 34 37
c37 34 0 7.07005e-20 $X=1.635 $Y=2.485
r38 36 37 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.485
+ $X2=2.275 $Y2=2.485
r39 32 36 2.24265 $w=6.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=2.19 $Y2=2.485
r40 32 34 15.4628 $w=6.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=1.635 $Y2=2.485
r41 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 26 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 25 37 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.275 $Y2=2.72
r45 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 22 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 21 34 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.635 $Y2=2.72
r49 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 19 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r51 19 21 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 13 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r53 13 15 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 11 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 7 29 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r57 7 9 11.0695 $w=3.78e-07 $l=3.65e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.27
r58 2 36 300 $w=1.7e-07 $l=6.94982e-07 $layer=licon1_PDIFF $count=2 $X=1.615
+ $Y=2.065 $X2=2.19 $Y2=2.33
r59 1 9 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%X 1 2 9 10 11 16 17
r19 28 29 7.295 $w=3.73e-07 $l=2.25e-07 $layer=LI1_cond $X=2.892 $Y=0.55
+ $X2=2.892 $Y2=0.775
r20 17 29 29.9263 $w=3.08e-07 $l=8.05e-07 $layer=LI1_cond $X=2.925 $Y=1.58
+ $X2=2.925 $Y2=0.775
r21 16 17 7.94212 $w=6.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.762 $Y=1.835
+ $X2=2.762 $Y2=1.58
r22 11 28 1.22927 $w=3.73e-07 $l=4e-08 $layer=LI1_cond $X=2.892 $Y=0.51
+ $X2=2.892 $Y2=0.55
r23 10 16 0.659256 $w=6.33e-07 $l=3.5e-08 $layer=LI1_cond $X=2.762 $Y=1.87
+ $X2=2.762 $Y2=1.835
r24 9 10 6.4042 $w=6.33e-07 $l=3.4e-07 $layer=LI1_cond $X=2.762 $Y=2.21
+ $X2=2.762 $Y2=1.87
r25 2 16 300 $w=1.7e-07 $l=4.32724e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.485 $X2=2.79 $Y2=1.835
r26 1 28 182 $w=1.7e-07 $l=3.92874e-07 $layer=licon1_NDIFF $count=1 $X=2.615
+ $Y=0.235 $X2=2.79 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_1%VGND 1 2 7 9 13 15 17 24 25 31
r38 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r39 25 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r40 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r41 22 31 10.508 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.222
+ $Y2=0
r42 22 24 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.99
+ $Y2=0
r43 21 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r44 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 18 28 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r46 18 20 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r47 17 31 10.508 $w=1.7e-07 $l=2.22e-07 $layer=LI1_cond $X=2 $Y=0 $X2=2.222
+ $Y2=0
r48 17 20 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=2 $Y=0 $X2=0.69
+ $Y2=0
r49 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r50 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r51 11 31 1.76584 $w=4.45e-07 $l=8.5e-08 $layer=LI1_cond $X=2.222 $Y=0.085
+ $X2=2.222 $Y2=0
r52 11 13 9.97057 $w=4.43e-07 $l=3.85e-07 $layer=LI1_cond $X=2.222 $Y=0.085
+ $X2=2.222 $Y2=0.47
r53 7 28 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r54 7 9 12.3845 $w=3.33e-07 $l=3.6e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.445
r55 2 13 182 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_NDIFF $count=1 $X=2.075
+ $Y=0.235 $X2=2.28 $Y2=0.47
r56 1 9 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

