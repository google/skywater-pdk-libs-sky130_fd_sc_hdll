* File: sky130_fd_sc_hdll__a22oi_1.pxi.spice
* Created: Thu Aug 27 18:54:23 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22OI_1%B2 N_B2_c_46_n N_B2_M1002_g N_B2_c_47_n
+ N_B2_M1007_g B2 B2 PM_SKY130_FD_SC_HDLL__A22OI_1%B2
x_PM_SKY130_FD_SC_HDLL__A22OI_1%B1 N_B1_c_74_n N_B1_M1001_g N_B1_c_75_n
+ N_B1_M1000_g B1 B1 B1 PM_SKY130_FD_SC_HDLL__A22OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A22OI_1%A1 N_A1_c_109_n N_A1_M1005_g N_A1_c_110_n
+ N_A1_M1003_g A1 A1 N_A1_c_112_n N_A1_c_113_n PM_SKY130_FD_SC_HDLL__A22OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A22OI_1%A2 N_A2_c_141_n N_A2_M1006_g N_A2_c_142_n
+ N_A2_M1004_g A2 PM_SKY130_FD_SC_HDLL__A22OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A22OI_1%Y N_Y_M1001_d N_Y_M1003_s N_Y_M1002_s
+ N_Y_M1000_d N_Y_c_168_n N_Y_c_169_n N_Y_c_207_n N_Y_c_170_n N_Y_c_172_n
+ N_Y_c_173_n N_Y_c_180_n N_Y_c_174_n Y Y Y N_Y_c_176_n
+ PM_SKY130_FD_SC_HDLL__A22OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A22OI_1%A_117_297# N_A_117_297#_M1002_d
+ N_A_117_297#_M1005_d N_A_117_297#_c_246_n N_A_117_297#_c_257_n
+ PM_SKY130_FD_SC_HDLL__A22OI_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A22OI_1%VPWR N_VPWR_M1005_s N_VPWR_M1004_d
+ N_VPWR_c_268_n N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n VPWR
+ N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_267_n N_VPWR_c_275_n
+ PM_SKY130_FD_SC_HDLL__A22OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A22OI_1%VGND N_VGND_M1007_s N_VGND_M1006_d
+ N_VGND_c_305_n N_VGND_c_306_n N_VGND_c_307_n VGND N_VGND_c_308_n
+ N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n
+ PM_SKY130_FD_SC_HDLL__A22OI_1%VGND
cc_1 VNB N_B2_c_46_n 0.0290841f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B2_c_47_n 0.0179427f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB B2 0.0247369f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_4 VNB N_B1_c_74_n 0.0193893f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B1_c_75_n 0.0245333f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B1 0.00497176f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_7 VNB B1 0.00718303f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A1_c_109_n 0.0249024f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_A1_c_110_n 0.0195233f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB A1 0.00612079f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_11 VNB N_A1_c_112_n 0.00334202f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=0.85
cc_12 VNB N_A1_c_113_n 0.00419735f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A2_c_141_n 0.0197842f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_A2_c_142_n 0.0252086f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_15 VNB A2 0.00728035f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_16 VNB N_Y_c_168_n 0.0135712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_169_n 0.0130311f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_170_n 0.0271896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_267_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_305_n 0.0128699f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_21 VNB N_VGND_c_306_n 0.0189114f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_307_n 0.0149922f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_23 VNB N_VGND_c_308_n 0.0452217f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=1.19
cc_24 VNB N_VGND_c_309_n 0.0131156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_310_n 0.185944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_311_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VPB N_B2_c_46_n 0.0331309f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_28 VPB N_B1_c_75_n 0.0314673f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_29 VPB N_A1_c_109_n 0.0304842f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_A2_c_142_n 0.0284447f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_31 VPB N_Y_c_170_n 0.00849929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_Y_c_172_n 0.00746643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_Y_c_173_n 0.00372117f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_Y_c_174_n 0.05251f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB Y 0.0106991f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_Y_c_176_n 0.0262461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_117_297#_c_246_n 0.00789503f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_38 VPB N_VPWR_c_268_n 0.00540402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_VPWR_c_269_n 0.00471756f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_40 VPB N_VPWR_c_270_n 0.0179855f $X=-0.19 $Y=1.305 $X2=0.375 $Y2=1.16
cc_41 VPB N_VPWR_c_271_n 0.00507132f $X=-0.19 $Y=1.305 $X2=0.375 $Y2=1.19
cc_42 VPB N_VPWR_c_272_n 0.0386414f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_273_n 0.014713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_267_n 0.058714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_275_n 0.00546324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 N_B2_c_47_n N_B1_c_74_n 0.0304806f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_47 B2 N_B1_c_74_n 0.00201099f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_48 N_B2_c_46_n N_B1_c_75_n 0.0669432f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_49 B2 N_B1_c_75_n 6.76553e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_50 B2 B1 0.00789857f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_51 N_B2_c_46_n B1 7.09664e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 B2 B1 0.0162938f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_53 N_B2_c_47_n N_Y_c_168_n 8.14295e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 N_B2_c_46_n N_Y_c_172_n 4.66918e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_B2_c_46_n N_Y_c_173_n 2.90944e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 N_B2_c_46_n N_Y_c_180_n 0.0129415f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_B2_c_46_n N_Y_c_174_n 0.0140509f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_58 B2 N_Y_c_174_n 0.0150384f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_59 N_B2_c_46_n Y 0.00464281f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 B2 Y 0.0266757f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_61 N_B2_c_46_n N_Y_c_176_n 0.0103831f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_B2_c_46_n N_VPWR_c_272_n 0.00429425f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B2_c_46_n N_VPWR_c_267_n 0.00700259f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 B2 N_VGND_M1007_s 0.00308023f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_65 N_B2_c_46_n N_VGND_c_306_n 6.83682e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_B2_c_47_n N_VGND_c_306_n 0.0214982f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_67 B2 N_VGND_c_306_n 0.0343697f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_68 N_B2_c_47_n N_VGND_c_310_n 8.26999e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_69 B2 N_VGND_c_310_n 0.00294983f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_70 N_B1_c_75_n N_A1_c_109_n 0.00447051f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_71 B1 N_A1_c_109_n 5.42314e-19 $X=1.145 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_72 B1 A1 0.0257888f $X=1.145 $Y=0.765 $X2=0 $Y2=0
cc_73 N_B1_c_75_n N_A1_c_113_n 7.13069e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 B1 N_A1_c_113_n 0.0014727f $X=1.145 $Y=0.765 $X2=0 $Y2=0
cc_75 B1 N_A1_c_113_n 0.0153799f $X=1.145 $Y=1.105 $X2=0 $Y2=0
cc_76 B1 N_Y_M1001_d 0.00384172f $X=1.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_77 N_B1_c_74_n N_Y_c_168_n 0.0101792f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_78 N_B1_c_75_n N_Y_c_168_n 2.43125e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_79 B1 N_Y_c_168_n 0.0185907f $X=1.145 $Y=0.765 $X2=0 $Y2=0
cc_80 B1 N_Y_c_168_n 0.00446124f $X=1.145 $Y=1.105 $X2=0 $Y2=0
cc_81 N_B1_c_75_n N_Y_c_173_n 0.0026712f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B1_c_75_n N_Y_c_180_n 0.00895143f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B1_c_75_n N_Y_c_174_n 0.0161165f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 B1 N_Y_c_174_n 0.0364046f $X=1.145 $Y=1.105 $X2=0 $Y2=0
cc_85 N_B1_c_75_n N_Y_c_176_n 0.00136747f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B1_c_75_n N_A_117_297#_c_246_n 0.0137257f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B1_c_75_n N_VPWR_c_268_n 0.00236094f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B1_c_75_n N_VPWR_c_272_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B1_c_75_n N_VPWR_c_267_n 0.00737353f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B1_c_74_n N_VGND_c_306_n 0.00288877f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_91 N_B1_c_74_n N_VGND_c_308_n 0.00365461f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_92 N_B1_c_74_n N_VGND_c_310_n 0.0067644f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A1_c_110_n N_A2_c_141_n 0.0299352f $X=1.98 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_94 N_A1_c_109_n N_A2_c_142_n 0.0669249f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A1_c_112_n N_A2_c_142_n 7.32912e-19 $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A1_c_109_n A2 0.00134543f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_97 A1 A2 0.00217377f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A1_c_112_n A2 0.0183474f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_99 A1 N_Y_M1003_s 0.00545883f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A1_c_109_n N_Y_c_168_n 0.00209545f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A1_c_110_n N_Y_c_168_n 0.0108835f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_102 A1 N_Y_c_168_n 0.0166025f $X=1.565 $Y=0.765 $X2=0 $Y2=0
cc_103 N_A1_c_112_n N_Y_c_168_n 0.00885963f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A1_c_109_n N_Y_c_174_n 0.0161165f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A1_c_112_n N_Y_c_174_n 0.0251124f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A1_c_113_n N_Y_c_174_n 0.0175558f $X=1.63 $Y=1.055 $X2=0 $Y2=0
cc_107 N_A1_c_109_n N_A_117_297#_c_246_n 0.0147263f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_109_n N_VPWR_c_268_n 0.0113334f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_109_n N_VPWR_c_270_n 0.00395083f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A1_c_109_n N_VPWR_c_267_n 0.00473008f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A1_c_110_n N_VGND_c_308_n 0.00357877f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_110_n N_VGND_c_310_n 0.00657948f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_141_n N_Y_c_169_n 0.013406f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A2_c_142_n N_Y_c_169_n 7.17521e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_115 A2 N_Y_c_169_n 0.0216257f $X=2.4 $Y=1.105 $X2=0 $Y2=0
cc_116 A2 N_Y_c_207_n 4.56812e-19 $X=2.4 $Y=1.105 $X2=0 $Y2=0
cc_117 N_A2_c_141_n N_Y_c_170_n 0.00536237f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A2_c_142_n N_Y_c_170_n 0.00792014f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_119 A2 N_Y_c_170_n 0.0235186f $X=2.4 $Y=1.105 $X2=0 $Y2=0
cc_120 N_A2_c_142_n N_Y_c_174_n 0.0214678f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_121 A2 N_Y_c_174_n 0.0263866f $X=2.4 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A2_c_142_n N_A_117_297#_c_246_n 0.00281218f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A2_c_142_n N_VPWR_c_268_n 0.00117667f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A2_c_142_n N_VPWR_c_269_n 0.00327906f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_142_n N_VPWR_c_270_n 0.00702461f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A2_c_142_n N_VPWR_c_267_n 0.0136712f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A2_c_141_n N_VGND_c_307_n 0.00474118f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A2_c_141_n N_VGND_c_308_n 0.00428022f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_141_n N_VGND_c_310_n 0.00706358f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_130 N_Y_c_180_n N_A_117_297#_M1002_d 0.00348224f $X=1.035 $Y=2.33 $X2=-0.19
+ $Y2=-0.24
cc_131 N_Y_c_174_n N_A_117_297#_M1002_d 0.00178587f $X=2.795 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_132 N_Y_c_174_n N_A_117_297#_M1005_d 0.00178587f $X=2.795 $Y=1.53 $X2=0 $Y2=0
cc_133 N_Y_M1000_d N_A_117_297#_c_246_n 0.00566948f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_Y_c_173_n N_A_117_297#_c_246_n 0.0170129f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_135 N_Y_c_180_n N_A_117_297#_c_246_n 0.00597357f $X=1.035 $Y=2.33 $X2=0 $Y2=0
cc_136 N_Y_c_174_n N_A_117_297#_c_246_n 0.0899206f $X=2.795 $Y=1.53 $X2=0 $Y2=0
cc_137 N_Y_c_180_n N_A_117_297#_c_257_n 0.0115453f $X=1.035 $Y=2.33 $X2=0 $Y2=0
cc_138 N_Y_c_174_n N_A_117_297#_c_257_n 0.0129015f $X=2.795 $Y=1.53 $X2=0 $Y2=0
cc_139 N_Y_c_176_n N_A_117_297#_c_257_n 0.0199789f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_140 N_Y_c_174_n N_VPWR_M1005_s 0.00291237f $X=2.795 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_141 N_Y_c_174_n N_VPWR_M1004_d 0.00404786f $X=2.795 $Y=1.53 $X2=0 $Y2=0
cc_142 N_Y_c_173_n N_VPWR_c_268_n 0.0176695f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_143 N_Y_c_174_n N_VPWR_c_269_n 0.0160432f $X=2.795 $Y=1.53 $X2=0 $Y2=0
cc_144 N_Y_c_172_n N_VPWR_c_272_n 0.0211994f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_145 N_Y_c_180_n N_VPWR_c_272_n 0.0553209f $X=1.035 $Y=2.33 $X2=0 $Y2=0
cc_146 N_Y_M1002_s N_VPWR_c_267_n 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_147 N_Y_M1000_d N_VPWR_c_267_n 0.00217543f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_148 N_Y_c_172_n N_VPWR_c_267_n 0.012545f $X=0.26 $Y=2.295 $X2=0 $Y2=0
cc_149 N_Y_c_180_n N_VPWR_c_267_n 0.0338884f $X=1.035 $Y=2.33 $X2=0 $Y2=0
cc_150 N_Y_c_169_n N_VGND_M1006_d 0.00860556f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_151 N_Y_c_170_n N_VGND_M1006_d 9.34528e-19 $X=2.965 $Y=1.445 $X2=0 $Y2=0
cc_152 N_Y_c_168_n N_VGND_c_306_n 0.0138717f $X=2.095 $Y=0.38 $X2=0 $Y2=0
cc_153 N_Y_c_169_n N_VGND_c_307_n 0.0234938f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_154 N_Y_c_168_n N_VGND_c_308_n 0.0865139f $X=2.095 $Y=0.38 $X2=0 $Y2=0
cc_155 N_Y_c_169_n N_VGND_c_308_n 0.0030777f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_156 N_Y_c_169_n N_VGND_c_309_n 0.00583805f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_157 N_Y_M1001_d N_VGND_c_310_n 0.00217543f $X=1.015 $Y=0.235 $X2=0 $Y2=0
cc_158 N_Y_M1003_s N_VGND_c_310_n 0.00250339f $X=1.595 $Y=0.235 $X2=0 $Y2=0
cc_159 N_Y_c_168_n N_VGND_c_310_n 0.051421f $X=2.095 $Y=0.38 $X2=0 $Y2=0
cc_160 N_Y_c_169_n N_VGND_c_310_n 0.0159836f $X=2.795 $Y=0.74 $X2=0 $Y2=0
cc_161 N_Y_c_168_n A_411_47# 0.00192108f $X=2.095 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_162 N_Y_c_207_n A_411_47# 0.00319553f $X=2.275 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_163 N_A_117_297#_c_246_n N_VPWR_M1005_s 0.00595501f $X=2.105 $Y=1.882
+ $X2=-0.19 $Y2=1.305
cc_164 N_A_117_297#_c_246_n N_VPWR_c_268_n 0.0151429f $X=2.105 $Y=1.882 $X2=0
+ $Y2=0
cc_165 N_A_117_297#_c_246_n N_VPWR_c_270_n 0.00596559f $X=2.105 $Y=1.882 $X2=0
+ $Y2=0
cc_166 N_A_117_297#_c_246_n N_VPWR_c_272_n 0.0026864f $X=2.105 $Y=1.882 $X2=0
+ $Y2=0
cc_167 N_A_117_297#_M1002_d N_VPWR_c_267_n 0.00232092f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_168 N_A_117_297#_M1005_d N_VPWR_c_267_n 0.00517304f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_169 N_A_117_297#_c_246_n N_VPWR_c_267_n 0.0173552f $X=2.105 $Y=1.882 $X2=0
+ $Y2=0
cc_170 N_VGND_c_310_n A_119_47# 0.010682f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_171 N_VGND_c_310_n A_411_47# 0.00236501f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
