* NGSPICE file created from sky130_fd_sc_hdll__inv_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__inv_1 A VGND VNB VPB VPWR Y
M1000 Y A VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=2.015e+11p ps=1.92e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=2.7e+11p ps=2.54e+06u
.ends

