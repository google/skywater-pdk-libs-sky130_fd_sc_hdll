* File: sky130_fd_sc_hdll__o21ba_2.pex.spice
* Created: Thu Aug 27 19:19:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%B1_N 1 3 4 6 7 8 20
r34 20 21 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.715 $Y2=1.16
r35 14 21 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.715 $Y=1.325
+ $X2=0.715 $Y2=1.16
r36 13 20 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=0.53 $Y=1.16 $X2=0.69
+ $Y2=1.16
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.53
+ $Y=1.16 $X2=0.53 $Y2=1.16
r38 8 14 10.7387 $w=2.18e-07 $l=2.05e-07 $layer=LI1_cond $X=0.715 $Y=1.53
+ $X2=0.715 $Y2=1.325
r39 7 21 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=0.74 $Y=1.16
+ $X2=0.715 $Y2=1.16
r40 4 12 49.2447 $w=2.79e-07 $l=2.73861e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.545 $Y2=1.16
r41 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
r42 1 12 38.7444 $w=2.79e-07 $l=1.98997e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.545 $Y2=1.16
r43 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%A_186_21# 1 2 7 9 10 12 13 15 16 18 21 24
+ 25 28 31 34 37 39 45
c105 34 0 4.88489e-20 $X=2.305 $Y=0.74
c106 21 0 1.78374e-19 $X=1.49 $Y=1.16
r107 45 46 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=1.525 $Y=1.202
+ $X2=1.55 $Y2=1.202
r108 42 43 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.03 $Y2=1.202
r109 37 39 0.371197 $w=5.78e-07 $l=1.8e-08 $layer=LI1_cond $X=2.762 $Y=1.745
+ $X2=2.78 $Y2=1.745
r110 35 37 8.24882 $w=5.78e-07 $l=4e-07 $layer=LI1_cond $X=2.362 $Y=1.745
+ $X2=2.762 $Y2=1.745
r111 31 35 6.62809 $w=2.15e-07 $l=2.9e-07 $layer=LI1_cond $X=2.362 $Y=1.455
+ $X2=2.362 $Y2=1.745
r112 30 34 3.43356 $w=2.72e-07 $l=1.09864e-07 $layer=LI1_cond $X=2.362 $Y=0.825
+ $X2=2.305 $Y2=0.74
r113 30 31 33.7693 $w=2.13e-07 $l=6.3e-07 $layer=LI1_cond $X=2.362 $Y=0.825
+ $X2=2.362 $Y2=1.455
r114 26 34 3.43356 $w=2.72e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.655
+ $X2=2.305 $Y2=0.74
r115 26 28 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.305 $Y=0.655
+ $X2=2.305 $Y2=0.38
r116 24 34 3.08518 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.14 $Y=0.74
+ $X2=2.305 $Y2=0.74
r117 24 25 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.14 $Y=0.74
+ $X2=1.575 $Y2=0.74
r118 22 45 4.46296 $w=3.78e-07 $l=3.5e-08 $layer=POLY_cond $X=1.49 $Y=1.202
+ $X2=1.525 $Y2=1.202
r119 22 43 58.6561 $w=3.78e-07 $l=4.6e-07 $layer=POLY_cond $X=1.49 $Y=1.202
+ $X2=1.03 $Y2=1.202
r120 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.49
+ $Y=1.16 $X2=1.49 $Y2=1.16
r121 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.575 $Y2=0.74
r122 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.49 $Y=0.825
+ $X2=1.49 $Y2=1.16
r123 16 46 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.55 $Y=0.995
+ $X2=1.55 $Y2=1.202
r124 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.55 $Y=0.995
+ $X2=1.55 $Y2=0.56
r125 13 45 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.525 $Y=1.41
+ $X2=1.525 $Y2=1.202
r126 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.525 $Y=1.41
+ $X2=1.525 $Y2=1.985
r127 10 43 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r128 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.985
r129 7 42 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=1.202
r130 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r131 2 39 300 $w=1.7e-07 $l=5.66238e-07 $layer=licon1_PDIFF $count=2 $X=2.58
+ $Y=1.485 $X2=2.78 $Y2=1.96
r132 2 39 600 $w=1.7e-07 $l=2.58844e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=1.485 $X2=2.78 $Y2=1.62
r133 1 28 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=2.18
+ $Y=0.235 $X2=2.305 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%A_27_93# 1 2 7 9 10 12 13 14 17 20 21 22
+ 25 31 33
r74 28 31 2.62582 $w=3.93e-07 $l=9e-08 $layer=LI1_cond $X=0.17 $Y=0.627 $X2=0.26
+ $Y2=0.627
r75 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=1.16
+ $X2=2 $Y2=1.16
r76 23 25 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2 $Y=1.865 $X2=2
+ $Y2=1.16
r77 21 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.915 $Y=1.95
+ $X2=2 $Y2=1.865
r78 21 22 99.1658 $w=1.68e-07 $l=1.52e-06 $layer=LI1_cond $X=1.915 $Y=1.95
+ $X2=0.395 $Y2=1.95
r79 18 22 7.59919 $w=1.7e-07 $l=1.92873e-07 $layer=LI1_cond $X=0.24 $Y=1.865
+ $X2=0.395 $Y2=1.95
r80 18 20 7.62099 $w=3.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.24 $Y=1.865
+ $X2=0.24 $Y2=1.66
r81 17 33 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=0.24 $Y=1.65
+ $X2=0.24 $Y2=1.495
r82 17 20 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=0.24 $Y=1.65 $X2=0.24
+ $Y2=1.66
r83 15 28 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=0.627
r84 15 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=0.17 $Y=0.825
+ $X2=0.17 $Y2=1.495
r85 13 26 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=2.39 $Y=1.16 $X2=2
+ $Y2=1.16
r86 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.39 $Y=1.16
+ $X2=2.49 $Y2=1.202
r87 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.49 $Y2=1.202
r88 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=0.56
r89 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.49 $Y=1.41
+ $X2=2.49 $Y2=1.202
r90 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.49 $Y=1.41 $X2=2.49
+ $Y2=1.985
r91 2 20 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r92 1 31 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%A2 1 3 4 6 7 15
c30 4 0 4.88489e-20 $X=3.04 $Y=0.995
r31 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r32 7 15 8.71429 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=2.73 $Y=1.18
+ $X2=2.895 $Y2=1.18
r33 4 10 38.6072 $w=2.91e-07 $l=2.02287e-07 $layer=POLY_cond $X=3.04 $Y=0.995
+ $X2=2.957 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.04 $Y=0.995 $X2=3.04
+ $Y2=0.56
r35 1 10 48.3784 $w=2.91e-07 $l=2.77489e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=2.957 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%A1 1 3 4 6 7 8 13
r23 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.515
+ $Y=1.16 $X2=3.515 $Y2=1.16
r24 7 8 7.46177 $w=5.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.622 $Y=1.19
+ $X2=3.622 $Y2=1.53
r25 7 13 0.658392 $w=5.43e-07 $l=3e-08 $layer=LI1_cond $X=3.622 $Y=1.19
+ $X2=3.622 $Y2=1.16
r26 4 12 38.8967 $w=3.59e-07 $l=1.96914e-07 $layer=POLY_cond $X=3.46 $Y=0.995
+ $X2=3.53 $Y2=1.16
r27 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.46 $Y=0.995 $X2=3.46
+ $Y2=0.56
r28 1 12 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=3.43 $Y=1.41
+ $X2=3.53 $Y2=1.16
r29 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.43 $Y=1.41 $X2=3.43
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%VPWR 1 2 3 12 14 16 26 33 34 37 46 49 51
r54 51 52 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 48 49 10.1561 $w=5.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.215 $Y=2.505
+ $X2=2.38 $Y2=2.505
r56 44 48 2.89052 $w=5.98e-07 $l=1.45e-07 $layer=LI1_cond $X=2.07 $Y=2.505
+ $X2=2.215 $Y2=2.505
r57 44 46 17.8309 $w=5.98e-07 $l=5.5e-07 $layer=LI1_cond $X=2.07 $Y=2.505
+ $X2=1.52 $Y2=2.505
r58 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r59 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 37 40 11.2625 $w=4.38e-07 $l=4.3e-07 $layer=LI1_cond $X=0.74 $Y=2.29
+ $X2=0.74 $Y2=2.72
r61 34 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 31 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.83 $Y=2.72 $X2=3.64
+ $Y2=2.72
r64 31 33 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=3.83 $Y=2.72 $X2=3.91
+ $Y2=2.72
r65 30 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 30 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r67 29 49 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.53 $Y=2.72 $X2=2.38
+ $Y2=2.72
r68 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 26 51 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.45 $Y=2.72 $X2=3.64
+ $Y2=2.72
r70 26 29 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 25 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 25 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 24 46 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.15 $Y=2.72 $X2=1.52
+ $Y2=2.72
r74 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r75 22 40 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.96 $Y=2.72 $X2=0.74
+ $Y2=2.72
r76 22 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.96 $Y=2.72
+ $X2=1.15 $Y2=2.72
r77 16 40 6.36164 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.52 $Y=2.72 $X2=0.74
+ $Y2=2.72
r78 16 18 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r79 14 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 14 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 10 51 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.64 $Y=2.635
+ $X2=3.64 $Y2=2.72
r82 10 12 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.64 $Y=2.635
+ $X2=3.64 $Y2=1.96
r83 3 12 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.52
+ $Y=1.485 $X2=3.665 $Y2=1.96
r84 2 48 300 $w=1.7e-07 $l=1.0635e-06 $layer=licon1_PDIFF $count=2 $X=1.615
+ $Y=1.485 $X2=2.215 $Y2=2.29
r85 1 37 600 $w=1.7e-07 $l=9.03922e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.795 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%X 1 2 11 13 18 23
r33 13 23 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=1.115 $Y=0.38
+ $X2=1.215 $Y2=0.38
r34 13 18 0.960369 $w=2.38e-07 $l=2e-08 $layer=LI1_cond $X=1.115 $Y=0.53
+ $X2=1.115 $Y2=0.51
r35 13 18 2.16083 $w=2.38e-07 $l=4.5e-08 $layer=LI1_cond $X=1.115 $Y=0.465
+ $X2=1.115 $Y2=0.51
r36 8 13 46.3378 $w=2.38e-07 $l=9.65e-07 $layer=LI1_cond $X=1.115 $Y=1.495
+ $X2=1.115 $Y2=0.53
r37 8 11 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.115 $Y=1.595
+ $X2=1.265 $Y2=1.595
r38 2 11 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.12
+ $Y=1.485 $X2=1.265 $Y2=1.61
r39 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.215 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%VGND 1 2 3 14 16 20 24 27 28 29 39 40 43
+ 46
r62 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r63 44 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r64 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r65 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r66 37 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r67 36 37 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r68 34 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r69 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r70 33 36 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r71 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r72 31 46 9.23004 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=1.742
+ $Y2=0
r73 31 33 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.925 $Y=0 $X2=2.07
+ $Y2=0
r74 29 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r75 27 36 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.165 $Y=0 $X2=2.99
+ $Y2=0
r76 27 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.25
+ $Y2=0
r77 26 39 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.91
+ $Y2=0
r78 26 28 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.335 $Y=0 $X2=3.25
+ $Y2=0
r79 22 28 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0
r80 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.25 $Y=0.085
+ $X2=3.25 $Y2=0.39
r81 18 46 1.2012 $w=3.65e-07 $l=8.5e-08 $layer=LI1_cond $X=1.742 $Y=0.085
+ $X2=1.742 $Y2=0
r82 18 20 9.31427 $w=3.63e-07 $l=2.95e-07 $layer=LI1_cond $X=1.742 $Y=0.085
+ $X2=1.742 $Y2=0.38
r83 17 43 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=0.825 $Y=0 $X2=0.735
+ $Y2=0
r84 16 46 9.23004 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=1.742
+ $Y2=0
r85 16 17 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.56 $Y=0 $X2=0.825
+ $Y2=0
r86 12 43 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r87 12 14 35.4293 $w=1.78e-07 $l=5.75e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.66
r88 3 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.25 $Y2=0.39
r89 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.625
+ $Y=0.235 $X2=1.76 $Y2=0.38
r90 1 14 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.465 $X2=0.73 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BA_2%A_518_47# 1 2 9 11 12 15
r28 13 15 11.8684 $w=3.33e-07 $l=3.45e-07 $layer=LI1_cond $X=3.722 $Y=0.735
+ $X2=3.722 $Y2=0.39
r29 11 13 7.80856 $w=1.7e-07 $l=2.05144e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=3.722 $Y2=0.735
r30 11 12 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.555 $Y=0.82
+ $X2=2.945 $Y2=0.82
r31 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.82 $Y=0.735
+ $X2=2.945 $Y2=0.82
r32 7 9 7.14515 $w=2.48e-07 $l=1.55e-07 $layer=LI1_cond $X=2.82 $Y=0.735
+ $X2=2.82 $Y2=0.58
r33 2 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.535
+ $Y=0.235 $X2=3.72 $Y2=0.39
r34 1 9 182 $w=1.7e-07 $l=4.29622e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.235 $X2=2.78 $Y2=0.58
.ends

