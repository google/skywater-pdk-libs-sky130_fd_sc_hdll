# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a32oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a32oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 1.075000 3.255000 1.625000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.720000 1.075000 4.575000 1.625000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.075000 6.320000 1.625000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.795000 1.285000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 1.075000 0.875000 1.285000 ;
        RECT 0.145000 1.285000 0.325000 1.625000 ;
    END
  END B2
  PIN VGND
    ANTENNADIFFAREA  0.646750 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.195000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  2.080000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.455000 2.195000 1.625000 ;
        RECT 0.565000 1.625000 0.895000 2.125000 ;
        RECT 1.455000 0.655000 3.245000 0.825000 ;
        RECT 1.585000 1.625000 1.755000 2.125000 ;
        RECT 1.965000 0.825000 2.195000 1.455000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.095000  0.295000 0.425000 0.715000 ;
      RECT 0.095000  0.715000 1.285000 0.885000 ;
      RECT 0.175000  1.795000 0.345000 2.295000 ;
      RECT 0.175000  2.295000 2.225000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.545000 ;
      RECT 1.035000  0.295000 2.305000 0.465000 ;
      RECT 1.035000  0.465000 1.285000 0.715000 ;
      RECT 1.115000  1.795000 1.285000 2.295000 ;
      RECT 2.055000  1.795000 6.265000 1.965000 ;
      RECT 2.055000  1.965000 2.225000 2.295000 ;
      RECT 2.445000  2.255000 3.165000 2.635000 ;
      RECT 2.495000  0.295000 4.605000 0.465000 ;
      RECT 3.415000  1.965000 3.585000 2.465000 ;
      RECT 3.755000  0.635000 5.800000 0.805000 ;
      RECT 3.770000  2.255000 4.525000 2.635000 ;
      RECT 4.695000  1.965000 4.865000 2.465000 ;
      RECT 4.865000  0.085000 5.250000 0.465000 ;
      RECT 5.125000  2.255000 5.845000 2.635000 ;
      RECT 5.420000  0.275000 5.800000 0.635000 ;
      RECT 6.095000  0.085000 6.265000 0.885000 ;
      RECT 6.095000  1.965000 6.265000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a32oi_2
END LIBRARY
