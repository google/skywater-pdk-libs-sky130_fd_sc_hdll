* File: sky130_fd_sc_hdll__or2b_2.pex.spice
* Created: Wed Sep  2 08:48:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%B_N 1 3 6 8 13 16
r26 13 14 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r27 11 13 31.1181 $w=3.64e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r28 8 16 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r29 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r30 4 14 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r31 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r32 1 13 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r33 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%A_27_53# 1 2 9 11 13 16 18 19 22 26
r43 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.16 $X2=1.265 $Y2=1.16
r44 24 32 8.85254 $w=2.43e-07 $l=1.65e-07 $layer=LI1_cond $X=0.767 $Y=1.16
+ $X2=0.767 $Y2=1.325
r45 24 26 13.0959 $w=3.28e-07 $l=3.75e-07 $layer=LI1_cond $X=0.89 $Y=1.16
+ $X2=1.265 $Y2=1.16
r46 22 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=1.63
+ $X2=0.73 $Y2=1.325
r47 18 24 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=0.767 $Y=0.82
+ $X2=0.767 $Y2=1.16
r48 18 19 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=0.645 $Y=0.82
+ $X2=0.42 $Y2=0.82
r49 14 19 7.64049 $w=1.7e-07 $l=1.95944e-07 $layer=LI1_cond $X=0.262 $Y=0.735
+ $X2=0.42 $Y2=0.82
r50 14 16 10.6098 $w=3.13e-07 $l=2.9e-07 $layer=LI1_cond $X=0.262 $Y=0.735
+ $X2=0.262 $Y2=0.445
r51 11 27 44.7829 $w=4.14e-07 $l=3.10242e-07 $layer=POLY_cond $X=1.5 $Y=1.41
+ $X2=1.365 $Y2=1.16
r52 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.5 $Y=1.41 $X2=1.5
+ $Y2=1.695
r53 7 27 39.8702 $w=4.14e-07 $l=2.09105e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.365 $Y2=1.16
r54 7 9 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=0.475
r55 2 22 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r56 1 16 182 $w=1.7e-07 $l=2.34307e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%A 1 5 7 8 9 12 14 16 22 26
c48 8 0 8.49032e-20 $X=1.91 $Y=1.31
r49 20 26 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=1.055 $Y=2.25
+ $X2=1.15 $Y2=2.25
r50 19 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.055 $Y=2.28
+ $X2=1.22 $Y2=2.28
r51 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.055
+ $Y=2.28 $X2=1.055 $Y2=2.28
r52 16 26 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=2.25 $X2=1.15
+ $Y2=2.25
r53 10 14 101.939 $w=2e-07 $l=3.05e-07 $layer=POLY_cond $X=1.91 $Y=2.035
+ $X2=1.91 $Y2=2.34
r54 10 12 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.91 $Y=2.035
+ $X2=1.91 $Y2=1.695
r55 9 12 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.91 $Y=1.41
+ $X2=1.91 $Y2=1.695
r56 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.91 $Y=1.31 $X2=1.91
+ $Y2=1.41
r57 7 13 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.91 $Y=1.06 $X2=1.91
+ $Y2=0.96
r58 7 8 82.8943 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=1.91 $Y=1.06 $X2=1.91
+ $Y2=1.31
r59 5 13 248.691 $w=1.5e-07 $l=4.85e-07 $layer=POLY_cond $X=1.885 $Y=0.475
+ $X2=1.885 $Y2=0.96
r60 1 14 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.81 $Y=2.34 $X2=1.91
+ $Y2=2.34
r61 1 22 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=1.81 $Y=2.34 $X2=1.22
+ $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%A_228_297# 1 2 7 9 10 12 13 14 15 17 18 20
+ 21 22 26 28 29 33 35
c76 33 0 1.12758e-19 $X=2.355 $Y=1.16
r77 41 42 3.16273 $w=3.81e-07 $l=2.5e-08 $layer=POLY_cond $X=2.45 $Y=1.202
+ $X2=2.475 $Y2=1.202
r78 35 38 2.88111 $w=4.18e-07 $l=1.05e-07 $layer=LI1_cond $X=1.245 $Y=1.58
+ $X2=1.245 $Y2=1.685
r79 34 41 12.0184 $w=3.81e-07 $l=9.5e-08 $layer=POLY_cond $X=2.355 $Y=1.202
+ $X2=2.45 $Y2=1.202
r80 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.355
+ $Y=1.16 $X2=2.355 $Y2=1.16
r81 31 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.355 $Y=1.495
+ $X2=2.355 $Y2=1.16
r82 30 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.355 $Y=0.825
+ $X2=2.355 $Y2=1.16
r83 28 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.27 $Y=0.74
+ $X2=2.355 $Y2=0.825
r84 28 29 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.27 $Y=0.74
+ $X2=1.76 $Y2=0.74
r85 24 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.675 $Y=0.655
+ $X2=1.76 $Y2=0.74
r86 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.675 $Y=0.655
+ $X2=1.675 $Y2=0.47
r87 23 35 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.245 $Y2=1.58
r88 22 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.27 $Y=1.58
+ $X2=2.355 $Y2=1.495
r89 22 23 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=2.27 $Y=1.58
+ $X2=1.455 $Y2=1.58
r90 18 21 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.135 $Y=0.995
+ $X2=3.11 $Y2=1.202
r91 18 20 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.135 $Y=0.995
+ $X2=3.135 $Y2=0.56
r92 15 21 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.11 $Y=1.41
+ $X2=3.11 $Y2=1.202
r93 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.11 $Y=1.41
+ $X2=3.11 $Y2=1.985
r94 14 42 10.4828 $w=3.81e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.55 $Y=1.16
+ $X2=2.475 $Y2=1.202
r95 13 21 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=3.11 $Y2=1.202
r96 13 14 80.4362 $w=3.3e-07 $l=4.6e-07 $layer=POLY_cond $X=3.01 $Y=1.16
+ $X2=2.55 $Y2=1.16
r97 10 42 24.6764 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.475 $Y=0.995
+ $X2=2.475 $Y2=1.202
r98 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.475 $Y=0.995
+ $X2=2.475 $Y2=0.56
r99 7 41 20.3063 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.45 $Y2=1.202
r100 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.45 $Y=1.41
+ $X2=2.45 $Y2=1.985
r101 2 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.14
+ $Y=1.485 $X2=1.265 $Y2=1.685
r102 1 26 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.265 $X2=1.675 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%VPWR 1 2 3 10 12 16 18 20 24 26 31 40 44
c40 2 0 1.12758e-19 $X=2 $Y=1.485
r41 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r42 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 35 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 35 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r45 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 32 40 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.34 $Y=2.72 $X2=2.2
+ $Y2=2.72
r47 32 34 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.34 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 31 43 3.83517 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=3.482 $Y2=2.72
r49 31 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.285 $Y=2.72
+ $X2=2.99 $Y2=2.72
r50 30 41 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r51 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r52 27 37 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r53 27 29 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r54 26 40 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.06 $Y=2.72 $X2=2.2
+ $Y2=2.72
r55 26 29 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 24 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 24 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 20 23 33.3473 $w=2.33e-07 $l=6.8e-07 $layer=LI1_cond $X=3.402 $Y=1.65
+ $X2=3.402 $Y2=2.33
r59 18 43 3.2122 $w=2.35e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.402 $Y=2.635
+ $X2=3.482 $Y2=2.72
r60 18 23 14.9572 $w=2.33e-07 $l=3.05e-07 $layer=LI1_cond $X=3.402 $Y=2.635
+ $X2=3.402 $Y2=2.33
r61 14 40 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.2 $Y=2.635 $X2=2.2
+ $Y2=2.72
r62 14 16 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.2 $Y=2.635
+ $X2=2.2 $Y2=2
r63 10 37 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r64 10 12 43.2166 $w=2.58e-07 $l=9.75e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.66
r65 3 23 400 $w=1.7e-07 $l=9.26107e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.485 $X2=3.37 $Y2=2.33
r66 3 20 400 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_PDIFF $count=1 $X=3.2
+ $Y=1.485 $X2=3.37 $Y2=1.65
r67 2 16 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.485 $X2=2.21 $Y2=2
r68 1 12 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%X 1 2 7 10
r20 10 13 45.1974 $w=3.18e-07 $l=1.255e-06 $layer=LI1_cond $X=2.95 $Y=0.59
+ $X2=2.95 $Y2=1.845
r21 7 13 0.900346 $w=3.18e-07 $l=2.5e-08 $layer=LI1_cond $X=2.95 $Y=1.87
+ $X2=2.95 $Y2=1.845
r22 2 13 300 $w=1.7e-07 $l=5.002e-07 $layer=licon1_PDIFF $count=2 $X=2.54
+ $Y=1.485 $X2=2.875 $Y2=1.845
r23 1 10 182 $w=1.7e-07 $l=4.91325e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.235 $X2=2.875 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2B_2%VGND 1 2 3 12 16 18 20 22 24 30 38 40 44
r45 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r46 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r47 37 38 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.205 $Y=0.24
+ $X2=1.37 $Y2=0.24
r48 35 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r49 34 37 1.01207 $w=6.48e-07 $l=5.5e-08 $layer=LI1_cond $X=1.15 $Y=0.24
+ $X2=1.205 $Y2=0.24
r50 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r51 31 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r52 30 34 8.46455 $w=6.48e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.24
+ $X2=1.15 $Y2=0.24
r53 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 28 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r55 28 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r56 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r57 25 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.195
+ $Y2=0
r58 25 27 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.36 $Y=0 $X2=2.99
+ $Y2=0
r59 24 43 3.83517 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=3.482
+ $Y2=0
r60 24 27 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.285 $Y=0 $X2=2.99
+ $Y2=0
r61 22 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r62 18 43 3.2122 $w=2.35e-07 $l=1.18427e-07 $layer=LI1_cond $X=3.402 $Y=0.085
+ $X2=3.482 $Y2=0
r63 18 20 14.712 $w=2.33e-07 $l=3e-07 $layer=LI1_cond $X=3.402 $Y=0.085
+ $X2=3.402 $Y2=0.385
r64 14 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0
r65 14 16 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.195 $Y=0.085
+ $X2=2.195 $Y2=0.4
r66 12 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=2.195
+ $Y2=0
r67 12 38 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.03 $Y=0 $X2=1.37
+ $Y2=0
r68 3 20 91 $w=1.7e-07 $l=2.22711e-07 $layer=licon1_NDIFF $count=2 $X=3.21
+ $Y=0.235 $X2=3.37 $Y2=0.385
r69 2 16 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=1.96
+ $Y=0.265 $X2=2.195 $Y2=0.4
r70 1 37 91 $w=1.7e-07 $l=6.74129e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.265 $X2=1.205 $Y2=0.4
.ends

