* File: sky130_fd_sc_hdll__and4bb_2.pxi.spice
* Created: Wed Sep  2 08:23:41 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%A_N N_A_N_c_95_n N_A_N_c_96_n N_A_N_M1002_g
+ N_A_N_M1011_g A_N A_N N_A_N_c_94_n PM_SKY130_FD_SC_HDLL__AND4BB_2%A_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%A_184_21# N_A_184_21#_M1000_s
+ N_A_184_21#_M1008_d N_A_184_21#_M1003_d N_A_184_21#_c_124_n
+ N_A_184_21#_M1012_g N_A_184_21#_c_131_n N_A_184_21#_M1010_g
+ N_A_184_21#_c_125_n N_A_184_21#_M1013_g N_A_184_21#_c_132_n
+ N_A_184_21#_M1015_g N_A_184_21#_c_126_n N_A_184_21#_c_127_n
+ N_A_184_21#_c_218_p N_A_184_21#_c_220_p N_A_184_21#_c_128_n
+ N_A_184_21#_c_129_n N_A_184_21#_c_144_p N_A_184_21#_c_135_n
+ N_A_184_21#_c_136_n N_A_184_21#_c_181_p N_A_184_21#_c_130_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_2%A_184_21#
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%A_27_47# N_A_27_47#_M1011_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_242_n N_A_27_47#_c_243_n N_A_27_47#_M1008_g N_A_27_47#_M1000_g
+ N_A_27_47#_c_250_n N_A_27_47#_c_244_n N_A_27_47#_c_238_n N_A_27_47#_c_239_n
+ N_A_27_47#_c_273_n N_A_27_47#_c_246_n N_A_27_47#_c_247_n N_A_27_47#_c_240_n
+ N_A_27_47#_c_241_n PM_SKY130_FD_SC_HDLL__AND4BB_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%A_545_280# N_A_545_280#_M1014_d
+ N_A_545_280#_M1007_d N_A_545_280#_c_335_n N_A_545_280#_c_336_n
+ N_A_545_280#_M1009_g N_A_545_280#_M1004_g N_A_545_280#_c_338_n
+ N_A_545_280#_c_339_n N_A_545_280#_c_340_n N_A_545_280#_c_352_n
+ N_A_545_280#_c_341_n N_A_545_280#_c_333_n N_A_545_280#_c_343_n
+ N_A_545_280#_c_344_n N_A_545_280#_c_334_n N_A_545_280#_c_345_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_2%A_545_280#
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%C N_C_c_406_n N_C_c_411_n N_C_M1003_g
+ N_C_M1006_g C C C N_C_c_408_n N_C_c_409_n PM_SKY130_FD_SC_HDLL__AND4BB_2%C
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%D N_D_M1005_g N_D_c_449_n N_D_c_450_n
+ N_D_M1001_g D D D N_D_c_448_n PM_SKY130_FD_SC_HDLL__AND4BB_2%D
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%B_N N_B_N_c_493_n N_B_N_c_498_n N_B_N_M1007_g
+ N_B_N_M1014_g B_N B_N N_B_N_c_495_n N_B_N_c_496_n B_N
+ PM_SKY130_FD_SC_HDLL__AND4BB_2%B_N
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%VPWR N_VPWR_M1002_d N_VPWR_M1015_d
+ N_VPWR_M1009_d N_VPWR_M1001_d N_VPWR_c_529_n N_VPWR_c_530_n N_VPWR_c_531_n
+ N_VPWR_c_532_n VPWR N_VPWR_c_533_n N_VPWR_c_534_n N_VPWR_c_528_n
+ N_VPWR_c_536_n N_VPWR_c_537_n N_VPWR_c_538_n N_VPWR_c_539_n
+ PM_SKY130_FD_SC_HDLL__AND4BB_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%X N_X_M1012_s N_X_M1010_s X X X N_X_c_608_n X
+ PM_SKY130_FD_SC_HDLL__AND4BB_2%X
x_PM_SKY130_FD_SC_HDLL__AND4BB_2%VGND N_VGND_M1011_d N_VGND_M1013_d
+ N_VGND_M1005_d N_VGND_c_631_n N_VGND_c_632_n N_VGND_c_633_n VGND
+ N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n PM_SKY130_FD_SC_HDLL__AND4BB_2%VGND
cc_1 VNB N_A_N_M1011_g 0.0366941f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.0024619f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_94_n 0.0476084f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_184_21#_c_124_n 0.0167243f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_5 VNB N_A_184_21#_c_125_n 0.0194832f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_6 VNB N_A_184_21#_c_126_n 0.00126655f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.53
cc_7 VNB N_A_184_21#_c_127_n 0.00929626f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_184_21#_c_128_n 0.00396616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_184_21#_c_129_n 0.00545721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_184_21#_c_130_n 0.0488871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_M1000_g 0.0344412f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_12 VNB N_A_27_47#_c_238_n 0.00871067f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.53
cc_13 VNB N_A_27_47#_c_239_n 0.00348446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_240_n 0.0027408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_241_n 0.0349739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_545_280#_M1004_g 0.0472855f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_17 VNB N_A_545_280#_c_333_n 0.0335361f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_545_280#_c_334_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_C_c_406_n 0.00984718f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.89
cc_20 VNB C 0.00764007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_C_c_408_n 0.025027f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_22 VNB N_C_c_409_n 0.0162171f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_23 VNB N_D_M1005_g 0.0314793f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_24 VNB D 0.00761073f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_25 VNB N_D_c_448_n 0.0187436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_B_N_c_493_n 0.0126372f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.89
cc_27 VNB B_N 0.00618481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_B_N_c_495_n 0.0310032f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_29 VNB N_B_N_c_496_n 0.0215191f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_30 VNB N_VPWR_c_528_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_608_n 6.41148e-19 $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_32 VNB N_VGND_c_631_n 0.00518f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_632_n 0.0651889f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_34 VNB N_VGND_c_633_n 0.00478242f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_35 VNB N_VGND_c_634_n 0.0151529f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_36 VNB N_VGND_c_635_n 0.0158181f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.53
cc_37 VNB N_VGND_c_636_n 0.0195874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_637_n 0.263393f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_638_n 0.00794401f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_639_n 0.0120591f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VPB N_A_N_c_95_n 0.0395156f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_42 VPB N_A_N_c_96_n 0.0263918f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_43 VPB A_N 0.0159685f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_44 VPB N_A_N_c_94_n 0.0119448f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_45 VPB N_A_184_21#_c_131_n 0.0164808f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_184_21#_c_132_n 0.0193829f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_47 VPB N_A_184_21#_c_126_n 0.00227696f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.53
cc_48 VPB N_A_184_21#_c_129_n 0.00509073f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_184_21#_c_135_n 0.00603654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_184_21#_c_136_n 0.00479883f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_184_21#_c_130_n 0.0254581f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_47#_c_242_n 0.0321384f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_53 VPB N_A_27_47#_c_243_n 0.0260709f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_244_n 9.28565e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_239_n 0.00161481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_246_n 0.0114947f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_247_n 0.00309144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_240_n 3.69208e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_27_47#_c_241_n 0.0162144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_545_280#_c_335_n 0.00938267f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_61 VPB N_A_545_280#_c_336_n 0.0212533f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_545_280#_M1004_g 0.00531358f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_63 VPB N_A_545_280#_c_338_n 0.0261302f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_64 VPB N_A_545_280#_c_339_n 0.00158592f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_65 VPB N_A_545_280#_c_340_n 0.00819307f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_545_280#_c_341_n 0.0147617f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.53
cc_67 VPB N_A_545_280#_c_333_n 0.0299179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_545_280#_c_343_n 0.00267539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_545_280#_c_344_n 0.0288152f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_545_280#_c_345_n 0.0112142f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_C_c_406_n 0.0326647f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_72 VPB N_C_c_411_n 0.0211659f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_73 VPB N_D_c_449_n 0.0284578f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_74 VPB N_D_c_450_n 0.0237727f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_75 VPB D 0.00197901f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_76 VPB N_D_c_448_n 0.00830225f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B_N_c_493_n 0.0397583f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_78 VPB N_B_N_c_498_n 0.0276075f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_79 VPB B_N 0.00376338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_529_n 0.0154753f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_530_n 0.00287347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_531_n 0.020191f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_532_n 0.00513086f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.16
cc_84 VPB N_VPWR_c_533_n 0.015197f $X=-0.19 $Y=1.305 $X2=0.24 $Y2=1.53
cc_85 VPB N_VPWR_c_534_n 0.0175722f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_528_n 0.0479122f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_536_n 0.00870752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_537_n 0.0205616f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_538_n 0.0198385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_539_n 0.00560816f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_X_c_608_n 0.00144092f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_92 N_A_N_M1011_g N_A_184_21#_c_124_n 0.0172714f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_93 N_A_N_c_95_n N_A_184_21#_c_131_n 0.0191578f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_94 N_A_N_c_96_n N_A_184_21#_c_131_n 0.015502f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_95 N_A_N_c_94_n N_A_184_21#_c_130_n 0.0172714f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_N_M1011_g N_A_27_47#_c_250_n 0.00407642f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_N_c_96_n N_A_27_47#_c_244_n 0.00548009f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_98 N_A_N_M1011_g N_A_27_47#_c_238_n 0.0124225f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_99 A_N N_A_27_47#_c_238_n 0.0112557f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A_N_c_94_n N_A_27_47#_c_238_n 0.00551734f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_N_c_95_n N_A_27_47#_c_239_n 0.0218972f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_102 N_A_N_M1011_g N_A_27_47#_c_239_n 0.0106834f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_103 A_N N_A_27_47#_c_239_n 0.0455797f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A_N_c_94_n N_A_27_47#_c_239_n 0.0100507f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_N_c_95_n N_A_27_47#_c_246_n 0.00504117f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_106 N_A_N_c_96_n N_A_27_47#_c_246_n 0.0121785f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_107 A_N N_A_27_47#_c_246_n 0.00987856f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A_N_c_94_n N_A_27_47#_c_246_n 0.00220498f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_N_c_96_n N_VPWR_c_533_n 0.00318288f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_110 N_A_N_c_96_n N_VPWR_c_528_n 0.00467603f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_111 N_A_N_c_96_n N_VPWR_c_536_n 0.0110746f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_112 N_A_N_c_94_n X 4.06861e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_113 N_A_N_M1011_g N_X_c_608_n 0.00110555f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_114 N_A_N_M1011_g N_VGND_c_634_n 0.00198377f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_N_M1011_g N_VGND_c_637_n 0.00358947f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_116 N_A_N_M1011_g N_VGND_c_638_n 0.0112293f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_117 N_A_184_21#_c_129_n N_A_27_47#_c_242_n 0.0156306f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_118 N_A_184_21#_c_129_n N_A_27_47#_c_243_n 0.00113113f $X=2.495 $Y=1.915
+ $X2=0 $Y2=0
cc_119 N_A_184_21#_c_144_p N_A_27_47#_c_243_n 0.00418243f $X=2.68 $Y=2.3 $X2=0
+ $Y2=0
cc_120 N_A_184_21#_c_136_n N_A_27_47#_c_243_n 0.0101117f $X=2.765 $Y=2 $X2=0
+ $Y2=0
cc_121 N_A_184_21#_c_126_n N_A_27_47#_M1000_g 0.00262779f $X=1.6 $Y=1.16 $X2=0
+ $Y2=0
cc_122 N_A_184_21#_c_128_n N_A_27_47#_M1000_g 0.0124031f $X=2.495 $Y=0.805 $X2=0
+ $Y2=0
cc_123 N_A_184_21#_c_129_n N_A_27_47#_M1000_g 0.0072739f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_124 N_A_184_21#_c_124_n N_A_27_47#_c_238_n 0.00146411f $X=0.995 $Y=0.995
+ $X2=0 $Y2=0
cc_125 N_A_184_21#_c_124_n N_A_27_47#_c_239_n 0.00521458f $X=0.995 $Y=0.995
+ $X2=0 $Y2=0
cc_126 N_A_184_21#_c_131_n N_A_27_47#_c_239_n 0.00602919f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_184_21#_c_131_n N_A_27_47#_c_273_n 0.0180938f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_184_21#_c_132_n N_A_27_47#_c_273_n 0.0191971f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_184_21#_c_126_n N_A_27_47#_c_273_n 0.00570971f $X=1.6 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_184_21#_c_129_n N_A_27_47#_c_273_n 0.00149775f $X=2.495 $Y=1.915
+ $X2=0 $Y2=0
cc_131 N_A_184_21#_c_136_n N_A_27_47#_c_273_n 0.00760817f $X=2.765 $Y=2 $X2=0
+ $Y2=0
cc_132 N_A_184_21#_c_130_n N_A_27_47#_c_273_n 0.00125481f $X=1.49 $Y=1.202 $X2=0
+ $Y2=0
cc_133 N_A_184_21#_c_132_n N_A_27_47#_c_247_n 0.010906f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_184_21#_c_129_n N_A_27_47#_c_247_n 0.0254709f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_135 N_A_184_21#_c_130_n N_A_27_47#_c_247_n 0.00172208f $X=1.49 $Y=1.202 $X2=0
+ $Y2=0
cc_136 N_A_184_21#_c_126_n N_A_27_47#_c_240_n 0.0252121f $X=1.6 $Y=1.16 $X2=0
+ $Y2=0
cc_137 N_A_184_21#_c_127_n N_A_27_47#_c_240_n 0.0217712f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_138 N_A_184_21#_c_129_n N_A_27_47#_c_240_n 0.0238805f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_139 N_A_184_21#_c_130_n N_A_27_47#_c_240_n 0.00229343f $X=1.49 $Y=1.202 $X2=0
+ $Y2=0
cc_140 N_A_184_21#_c_126_n N_A_27_47#_c_241_n 3.51933e-19 $X=1.6 $Y=1.16 $X2=0
+ $Y2=0
cc_141 N_A_184_21#_c_127_n N_A_27_47#_c_241_n 0.010574f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_142 N_A_184_21#_c_129_n N_A_27_47#_c_241_n 0.0107911f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_143 N_A_184_21#_c_130_n N_A_27_47#_c_241_n 0.0166636f $X=1.49 $Y=1.202 $X2=0
+ $Y2=0
cc_144 N_A_184_21#_c_129_n N_A_545_280#_c_335_n 0.00363775f $X=2.495 $Y=1.915
+ $X2=0 $Y2=0
cc_145 N_A_184_21#_c_144_p N_A_545_280#_c_336_n 0.00399826f $X=2.68 $Y=2.3 $X2=0
+ $Y2=0
cc_146 N_A_184_21#_c_135_n N_A_545_280#_c_336_n 0.0136067f $X=3.545 $Y=2 $X2=0
+ $Y2=0
cc_147 N_A_184_21#_c_128_n N_A_545_280#_M1004_g 0.00199899f $X=2.495 $Y=0.805
+ $X2=0 $Y2=0
cc_148 N_A_184_21#_c_129_n N_A_545_280#_M1004_g 0.00716103f $X=2.495 $Y=1.915
+ $X2=0 $Y2=0
cc_149 N_A_184_21#_c_135_n N_A_545_280#_c_338_n 0.0524799f $X=3.545 $Y=2 $X2=0
+ $Y2=0
cc_150 N_A_184_21#_c_135_n N_A_545_280#_c_352_n 0.0150771f $X=3.545 $Y=2 $X2=0
+ $Y2=0
cc_151 N_A_184_21#_c_129_n N_A_545_280#_c_343_n 0.02367f $X=2.495 $Y=1.915 $X2=0
+ $Y2=0
cc_152 N_A_184_21#_c_135_n N_A_545_280#_c_343_n 0.015855f $X=3.545 $Y=2 $X2=0
+ $Y2=0
cc_153 N_A_184_21#_c_129_n N_A_545_280#_c_344_n 0.00203181f $X=2.495 $Y=1.915
+ $X2=0 $Y2=0
cc_154 N_A_184_21#_c_136_n N_A_545_280#_c_344_n 0.00260732f $X=2.765 $Y=2 $X2=0
+ $Y2=0
cc_155 N_A_184_21#_c_135_n N_C_c_411_n 0.0134879f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_156 N_A_184_21#_c_181_p N_C_c_411_n 0.00412276f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_157 N_A_184_21#_c_128_n C 0.00538925f $X=2.495 $Y=0.805 $X2=0 $Y2=0
cc_158 N_A_184_21#_c_129_n C 0.0130988f $X=2.495 $Y=1.915 $X2=0 $Y2=0
cc_159 N_A_184_21#_c_135_n N_D_c_450_n 0.0014042f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_160 N_A_184_21#_c_181_p N_D_c_450_n 0.00459241f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_161 N_A_184_21#_c_135_n N_VPWR_M1009_d 0.00190219f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_162 N_A_184_21#_c_144_p N_VPWR_c_529_n 0.0113299f $X=2.68 $Y=2.3 $X2=0 $Y2=0
cc_163 N_A_184_21#_c_136_n N_VPWR_c_529_n 0.00552107f $X=2.765 $Y=2 $X2=0 $Y2=0
cc_164 N_A_184_21#_c_181_p N_VPWR_c_530_n 0.0086977f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_165 N_A_184_21#_c_135_n N_VPWR_c_531_n 0.00320526f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_166 N_A_184_21#_c_181_p N_VPWR_c_531_n 0.0116326f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_167 N_A_184_21#_M1008_d N_VPWR_c_528_n 0.00310074f $X=2.505 $Y=2.065 $X2=0
+ $Y2=0
cc_168 N_A_184_21#_M1003_d N_VPWR_c_528_n 0.00439382f $X=3.485 $Y=2.065 $X2=0
+ $Y2=0
cc_169 N_A_184_21#_c_131_n N_VPWR_c_528_n 0.00692453f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_170 N_A_184_21#_c_132_n N_VPWR_c_528_n 0.00816029f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_184_21#_c_144_p N_VPWR_c_528_n 0.00637602f $X=2.68 $Y=2.3 $X2=0 $Y2=0
cc_172 N_A_184_21#_c_135_n N_VPWR_c_528_n 0.00709978f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_173 N_A_184_21#_c_136_n N_VPWR_c_528_n 0.00960989f $X=2.765 $Y=2 $X2=0 $Y2=0
cc_174 N_A_184_21#_c_181_p N_VPWR_c_528_n 0.00643448f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_175 N_A_184_21#_c_131_n N_VPWR_c_536_n 0.00438976f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_184_21#_c_131_n N_VPWR_c_537_n 0.00515358f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_184_21#_c_132_n N_VPWR_c_537_n 0.00515358f $X=1.49 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A_184_21#_c_132_n N_VPWR_c_538_n 0.0153776f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_184_21#_c_144_p N_VPWR_c_539_n 0.0157096f $X=2.68 $Y=2.3 $X2=0 $Y2=0
cc_180 N_A_184_21#_c_135_n N_VPWR_c_539_n 0.0203937f $X=3.545 $Y=2 $X2=0 $Y2=0
cc_181 N_A_184_21#_c_181_p N_VPWR_c_539_n 0.0128798f $X=3.63 $Y=2.3 $X2=0 $Y2=0
cc_182 N_A_184_21#_c_131_n X 0.00339678f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_184_21#_c_132_n X 0.00424556f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_184_21#_c_130_n X 0.00119575f $X=1.49 $Y=1.202 $X2=0 $Y2=0
cc_185 N_A_184_21#_c_124_n N_X_c_608_n 0.0134531f $X=0.995 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_184_21#_c_131_n N_X_c_608_n 0.00286192f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_184_21#_c_125_n N_X_c_608_n 0.00216197f $X=1.465 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_184_21#_c_132_n N_X_c_608_n 0.00148219f $X=1.49 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_184_21#_c_126_n N_X_c_608_n 0.0339317f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_184_21#_c_130_n N_X_c_608_n 0.0288149f $X=1.49 $Y=1.202 $X2=0 $Y2=0
cc_191 N_A_184_21#_c_126_n N_VGND_M1013_d 0.00134422f $X=1.6 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_184_21#_c_127_n N_VGND_M1013_d 0.00571044f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_193 N_A_184_21#_c_218_p N_VGND_M1013_d 0.00160022f $X=1.735 $Y=0.72 $X2=0
+ $Y2=0
cc_194 N_A_184_21#_c_127_n N_VGND_c_632_n 0.00872817f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_195 N_A_184_21#_c_220_p N_VGND_c_632_n 0.0111381f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_196 N_A_184_21#_c_124_n N_VGND_c_635_n 0.00579312f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_197 N_A_184_21#_c_125_n N_VGND_c_635_n 0.00468308f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_198 N_A_184_21#_M1000_s N_VGND_c_637_n 0.00242518f $X=2.105 $Y=0.235 $X2=0
+ $Y2=0
cc_199 N_A_184_21#_c_124_n N_VGND_c_637_n 0.0106199f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_200 N_A_184_21#_c_125_n N_VGND_c_637_n 0.00801881f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_184_21#_c_127_n N_VGND_c_637_n 0.0154255f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_202 N_A_184_21#_c_218_p N_VGND_c_637_n 0.00110018f $X=1.735 $Y=0.72 $X2=0
+ $Y2=0
cc_203 N_A_184_21#_c_220_p N_VGND_c_637_n 0.00637602f $X=2.23 $Y=0.42 $X2=0
+ $Y2=0
cc_204 N_A_184_21#_c_124_n N_VGND_c_638_n 0.00169113f $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_184_21#_c_124_n N_VGND_c_639_n 4.64464e-19 $X=0.995 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_184_21#_c_125_n N_VGND_c_639_n 0.0080434f $X=1.465 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_184_21#_c_127_n N_VGND_c_639_n 0.0118732f $X=2.145 $Y=0.72 $X2=0
+ $Y2=0
cc_208 N_A_184_21#_c_218_p N_VGND_c_639_n 0.0135801f $X=1.735 $Y=0.72 $X2=0
+ $Y2=0
cc_209 N_A_184_21#_c_220_p N_VGND_c_639_n 0.0123915f $X=2.23 $Y=0.42 $X2=0 $Y2=0
cc_210 N_A_184_21#_c_130_n N_VGND_c_639_n 6.20318e-19 $X=1.49 $Y=1.202 $X2=0
+ $Y2=0
cc_211 N_A_184_21#_c_128_n A_503_47# 8.81158e-19 $X=2.495 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_212 N_A_27_47#_c_242_n N_A_545_280#_c_335_n 0.00507307f $X=2.415 $Y=1.89
+ $X2=0 $Y2=0
cc_213 N_A_27_47#_c_243_n N_A_545_280#_c_336_n 0.0149149f $X=2.415 $Y=1.99 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_M1000_g N_A_545_280#_M1004_g 0.0440605f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_215 N_A_27_47#_c_242_n N_A_545_280#_c_343_n 3.57603e-19 $X=2.415 $Y=1.89
+ $X2=0 $Y2=0
cc_216 N_A_27_47#_c_242_n N_A_545_280#_c_344_n 0.0202467f $X=2.415 $Y=1.89 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_239_n N_VPWR_M1002_d 0.0048752f $X=0.61 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_27_47#_c_273_n N_VPWR_M1002_d 0.0074704f $X=1.905 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_27_47#_c_246_n N_VPWR_M1002_d 6.83486e-19 $X=0.72 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_220 N_A_27_47#_c_273_n N_VPWR_M1015_d 0.0177908f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_247_n N_VPWR_M1015_d 0.0133969f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_243_n N_VPWR_c_529_n 0.00598209f $X=2.415 $Y=1.99 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_244_n N_VPWR_c_533_n 0.0113907f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_246_n N_VPWR_c_533_n 0.00274481f $X=0.72 $Y=1.97 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1002_s N_VPWR_c_528_n 0.00380082f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_243_n N_VPWR_c_528_n 0.010102f $X=2.415 $Y=1.99 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_244_n N_VPWR_c_528_n 0.00638769f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_273_n N_VPWR_c_528_n 0.0208938f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_246_n N_VPWR_c_528_n 0.00587866f $X=0.72 $Y=1.97 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_244_n N_VPWR_c_536_n 0.0156776f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_246_n N_VPWR_c_536_n 0.0212706f $X=0.72 $Y=1.97 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_273_n N_VPWR_c_537_n 0.0102899f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_243_n N_VPWR_c_538_n 0.00359305f $X=2.415 $Y=1.99 $X2=0
+ $Y2=0
cc_234 N_A_27_47#_c_273_n N_VPWR_c_538_n 0.0299059f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_243_n N_VPWR_c_539_n 5.39753e-19 $X=2.415 $Y=1.99 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_273_n N_X_M1010_s 0.00475732f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_273_n X 0.0188647f $X=1.905 $Y=1.97 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_247_n X 0.00558816f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_238_n N_X_c_608_n 0.00780848f $X=0.61 $Y=0.805 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_239_n N_X_c_608_n 0.0402216f $X=0.61 $Y=1.885 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_247_n N_X_c_608_n 0.00720448f $X=1.99 $Y=1.885 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_238_n N_VGND_M1011_d 0.00281405f $X=0.61 $Y=0.805 $X2=-0.19
+ $Y2=-0.24
cc_243 N_A_27_47#_c_239_n N_VGND_M1011_d 0.00105765f $X=0.61 $Y=1.885 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_M1000_g N_VGND_c_632_n 0.00425094f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_250_n N_VGND_c_634_n 0.0113299f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_238_n N_VGND_c_634_n 0.00249084f $X=0.61 $Y=0.805 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_M1011_s N_VGND_c_637_n 0.00427389f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_M1000_g N_VGND_c_637_n 0.0073684f $X=2.44 $Y=0.445 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_250_n N_VGND_c_637_n 0.00637602f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_238_n N_VGND_c_637_n 0.00539404f $X=0.61 $Y=0.805 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_250_n N_VGND_c_638_n 0.0156777f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_238_n N_VGND_c_638_n 0.0107888f $X=0.61 $Y=0.805 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1000_g N_VGND_c_639_n 0.00289666f $X=2.44 $Y=0.445 $X2=0
+ $Y2=0
cc_254 N_A_545_280#_M1004_g N_C_c_406_n 0.0124783f $X=2.935 $Y=0.445 $X2=0 $Y2=0
cc_255 N_A_545_280#_c_338_n N_C_c_406_n 0.0134954f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_256 N_A_545_280#_c_339_n N_C_c_406_n 8.59234e-19 $X=3.995 $Y=1.915 $X2=0
+ $Y2=0
cc_257 N_A_545_280#_c_343_n N_C_c_406_n 0.00125138f $X=2.88 $Y=1.565 $X2=0 $Y2=0
cc_258 N_A_545_280#_c_344_n N_C_c_406_n 0.0139511f $X=2.88 $Y=1.565 $X2=0 $Y2=0
cc_259 N_A_545_280#_c_335_n N_C_c_411_n 0.0139511f $X=2.915 $Y=1.89 $X2=0 $Y2=0
cc_260 N_A_545_280#_c_336_n N_C_c_411_n 0.0116808f $X=2.915 $Y=1.99 $X2=0 $Y2=0
cc_261 N_A_545_280#_M1004_g C 0.00869038f $X=2.935 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_545_280#_c_338_n C 0.0132358f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_263 N_A_545_280#_M1004_g N_C_c_408_n 0.0196338f $X=2.935 $Y=0.445 $X2=0 $Y2=0
cc_264 N_A_545_280#_c_338_n N_C_c_408_n 0.00136896f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_265 N_A_545_280#_M1004_g N_C_c_409_n 0.0248325f $X=2.935 $Y=0.445 $X2=0 $Y2=0
cc_266 N_A_545_280#_c_338_n N_D_c_449_n 0.0148143f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_267 N_A_545_280#_c_339_n N_D_c_449_n 0.00470465f $X=3.995 $Y=1.915 $X2=0
+ $Y2=0
cc_268 N_A_545_280#_c_339_n N_D_c_450_n 7.89591e-19 $X=3.995 $Y=1.915 $X2=0
+ $Y2=0
cc_269 N_A_545_280#_c_352_n N_D_c_450_n 0.007018f $X=4.105 $Y=2 $X2=0 $Y2=0
cc_270 N_A_545_280#_c_338_n D 0.0241169f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_271 N_A_545_280#_c_338_n N_D_c_448_n 0.00162068f $X=3.885 $Y=1.66 $X2=0 $Y2=0
cc_272 N_A_545_280#_c_338_n N_B_N_c_493_n 0.00199883f $X=3.885 $Y=1.66 $X2=0
+ $Y2=0
cc_273 N_A_545_280#_c_339_n N_B_N_c_493_n 0.00167318f $X=3.995 $Y=1.915 $X2=0
+ $Y2=0
cc_274 N_A_545_280#_c_340_n N_B_N_c_498_n 0.0202368f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_275 N_A_545_280#_c_341_n N_B_N_c_498_n 0.00484502f $X=4.74 $Y=2.3 $X2=0 $Y2=0
cc_276 N_A_545_280#_c_340_n B_N 0.0108555f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_277 N_A_545_280#_c_333_n B_N 0.0335659f $X=4.83 $Y=1.915 $X2=0 $Y2=0
cc_278 N_A_545_280#_c_333_n N_B_N_c_496_n 0.0367088f $X=4.83 $Y=1.915 $X2=0
+ $Y2=0
cc_279 N_A_545_280#_c_340_n N_VPWR_M1001_d 0.0026613f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_280 N_A_545_280#_c_352_n N_VPWR_M1001_d 0.00168336f $X=4.105 $Y=2 $X2=0 $Y2=0
cc_281 N_A_545_280#_c_336_n N_VPWR_c_529_n 0.00315022f $X=2.915 $Y=1.99 $X2=0
+ $Y2=0
cc_282 N_A_545_280#_c_340_n N_VPWR_c_530_n 0.0205428f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_283 N_A_545_280#_c_341_n N_VPWR_c_530_n 0.0131278f $X=4.74 $Y=2.3 $X2=0 $Y2=0
cc_284 N_A_545_280#_c_352_n N_VPWR_c_531_n 0.0035426f $X=4.105 $Y=2 $X2=0 $Y2=0
cc_285 N_A_545_280#_c_340_n N_VPWR_c_534_n 0.00319548f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_286 N_A_545_280#_c_341_n N_VPWR_c_534_n 0.018114f $X=4.74 $Y=2.3 $X2=0 $Y2=0
cc_287 N_A_545_280#_M1007_d N_VPWR_c_528_n 0.00238238f $X=4.595 $Y=2.065 $X2=0
+ $Y2=0
cc_288 N_A_545_280#_c_336_n N_VPWR_c_528_n 0.00380608f $X=2.915 $Y=1.99 $X2=0
+ $Y2=0
cc_289 N_A_545_280#_c_340_n N_VPWR_c_528_n 0.00685901f $X=4.655 $Y=2 $X2=0 $Y2=0
cc_290 N_A_545_280#_c_352_n N_VPWR_c_528_n 0.00617483f $X=4.105 $Y=2 $X2=0 $Y2=0
cc_291 N_A_545_280#_c_341_n N_VPWR_c_528_n 0.00991723f $X=4.74 $Y=2.3 $X2=0
+ $Y2=0
cc_292 N_A_545_280#_c_336_n N_VPWR_c_539_n 0.00959326f $X=2.915 $Y=1.99 $X2=0
+ $Y2=0
cc_293 N_A_545_280#_M1004_g N_VGND_c_632_n 0.00585385f $X=2.935 $Y=0.445 $X2=0
+ $Y2=0
cc_294 N_A_545_280#_c_334_n N_VGND_c_636_n 0.0170867f $X=4.83 $Y=0.42 $X2=0
+ $Y2=0
cc_295 N_A_545_280#_M1014_d N_VGND_c_637_n 0.00379446f $X=4.605 $Y=0.235 $X2=0
+ $Y2=0
cc_296 N_A_545_280#_M1004_g N_VGND_c_637_n 0.0112057f $X=2.935 $Y=0.445 $X2=0
+ $Y2=0
cc_297 N_A_545_280#_c_334_n N_VGND_c_637_n 0.00982816f $X=4.83 $Y=0.42 $X2=0
+ $Y2=0
cc_298 C N_D_M1005_g 0.00197219f $X=3.27 $Y=0.425 $X2=0 $Y2=0
cc_299 N_C_c_409_n N_D_M1005_g 0.0227355f $X=3.36 $Y=0.775 $X2=0 $Y2=0
cc_300 N_C_c_406_n N_D_c_449_n 0.0227355f $X=3.395 $Y=1.89 $X2=0 $Y2=0
cc_301 N_C_c_411_n N_D_c_450_n 0.0333858f $X=3.395 $Y=1.99 $X2=0 $Y2=0
cc_302 N_C_c_406_n D 0.00287595f $X=3.395 $Y=1.89 $X2=0 $Y2=0
cc_303 C D 0.0594526f $X=3.27 $Y=0.425 $X2=0 $Y2=0
cc_304 N_C_c_409_n D 0.00264451f $X=3.36 $Y=0.775 $X2=0 $Y2=0
cc_305 N_C_c_408_n N_D_c_448_n 0.0227355f $X=3.36 $Y=0.94 $X2=0 $Y2=0
cc_306 N_C_c_411_n N_VPWR_c_531_n 0.00456711f $X=3.395 $Y=1.99 $X2=0 $Y2=0
cc_307 N_C_c_411_n N_VPWR_c_528_n 0.00516277f $X=3.395 $Y=1.99 $X2=0 $Y2=0
cc_308 N_C_c_411_n N_VPWR_c_539_n 0.00786257f $X=3.395 $Y=1.99 $X2=0 $Y2=0
cc_309 C N_VGND_c_632_n 0.00712416f $X=3.27 $Y=0.425 $X2=0 $Y2=0
cc_310 N_C_c_408_n N_VGND_c_632_n 9.83499e-19 $X=3.36 $Y=0.94 $X2=0 $Y2=0
cc_311 N_C_c_409_n N_VGND_c_632_n 0.0038979f $X=3.36 $Y=0.775 $X2=0 $Y2=0
cc_312 C N_VGND_c_637_n 0.00846732f $X=3.27 $Y=0.425 $X2=0 $Y2=0
cc_313 N_C_c_408_n N_VGND_c_637_n 0.00107677f $X=3.36 $Y=0.94 $X2=0 $Y2=0
cc_314 N_C_c_409_n N_VGND_c_637_n 0.00563436f $X=3.36 $Y=0.775 $X2=0 $Y2=0
cc_315 C A_602_47# 0.0033564f $X=3.27 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_316 N_D_c_449_n N_B_N_c_493_n 0.00768321f $X=3.865 $Y=1.89 $X2=0 $Y2=0
cc_317 D N_B_N_c_493_n 7.57099e-19 $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_318 N_D_c_448_n N_B_N_c_493_n 0.00957091f $X=3.9 $Y=1.24 $X2=0 $Y2=0
cc_319 N_D_c_450_n N_B_N_c_498_n 0.0189196f $X=3.865 $Y=1.99 $X2=0 $Y2=0
cc_320 N_D_M1005_g B_N 9.63354e-19 $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_321 D B_N 0.0439013f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_322 N_D_c_448_n B_N 0.00179693f $X=3.9 $Y=1.24 $X2=0 $Y2=0
cc_323 N_D_M1005_g N_B_N_c_495_n 0.00892162f $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_324 D N_B_N_c_495_n 8.73602e-19 $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_325 N_D_c_448_n N_B_N_c_495_n 8.85797e-19 $X=3.9 $Y=1.24 $X2=0 $Y2=0
cc_326 N_D_M1005_g N_B_N_c_496_n 0.00833793f $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_327 D N_B_N_c_496_n 0.00343003f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_328 N_D_c_450_n N_VPWR_c_530_n 0.00539424f $X=3.865 $Y=1.99 $X2=0 $Y2=0
cc_329 N_D_c_450_n N_VPWR_c_531_n 0.00651568f $X=3.865 $Y=1.99 $X2=0 $Y2=0
cc_330 N_D_c_450_n N_VPWR_c_528_n 0.0110541f $X=3.865 $Y=1.99 $X2=0 $Y2=0
cc_331 N_D_c_450_n N_VPWR_c_539_n 0.00107401f $X=3.865 $Y=1.99 $X2=0 $Y2=0
cc_332 D N_VGND_M1005_d 0.00308014f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_333 N_D_M1005_g N_VGND_c_631_n 0.00663019f $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_334 D N_VGND_c_631_n 0.011963f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_335 N_D_M1005_g N_VGND_c_632_n 0.00390689f $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_336 D N_VGND_c_632_n 0.0078617f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_337 N_D_M1005_g N_VGND_c_637_n 0.00603312f $X=3.84 $Y=0.445 $X2=0 $Y2=0
cc_338 D N_VGND_c_637_n 0.00964347f $X=3.785 $Y=0.425 $X2=0 $Y2=0
cc_339 D A_699_47# 0.001987f $X=3.785 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_340 N_B_N_c_498_n N_VPWR_c_530_n 0.0085817f $X=4.505 $Y=1.99 $X2=0 $Y2=0
cc_341 N_B_N_c_498_n N_VPWR_c_534_n 0.00456002f $X=4.505 $Y=1.99 $X2=0 $Y2=0
cc_342 N_B_N_c_498_n N_VPWR_c_528_n 0.00610017f $X=4.505 $Y=1.99 $X2=0 $Y2=0
cc_343 B_N N_VGND_c_631_n 0.0185899f $X=4.175 $Y=0.765 $X2=0 $Y2=0
cc_344 N_B_N_c_495_n N_VGND_c_631_n 8.93205e-19 $X=4.44 $Y=0.93 $X2=0 $Y2=0
cc_345 N_B_N_c_496_n N_VGND_c_631_n 0.00335421f $X=4.455 $Y=0.765 $X2=0 $Y2=0
cc_346 N_B_N_c_496_n N_VGND_c_636_n 0.00585385f $X=4.455 $Y=0.765 $X2=0 $Y2=0
cc_347 B_N N_VGND_c_637_n 0.00436117f $X=4.175 $Y=0.765 $X2=0 $Y2=0
cc_348 N_B_N_c_496_n N_VGND_c_637_n 0.00993123f $X=4.455 $Y=0.765 $X2=0 $Y2=0
cc_349 N_VPWR_c_528_n N_X_M1010_s 0.00351307f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_350 N_X_c_608_n N_VGND_c_635_n 0.0169614f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_351 N_X_M1012_s N_VGND_c_637_n 0.00428929f $X=1.07 $Y=0.235 $X2=0 $Y2=0
cc_352 N_X_c_608_n N_VGND_c_637_n 0.010423f $X=1.255 $Y=0.42 $X2=0 $Y2=0
cc_353 N_VGND_c_637_n A_503_47# 0.0119395f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_354 N_VGND_c_637_n A_602_47# 0.0107664f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_355 N_VGND_c_637_n A_699_47# 0.00823311f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
