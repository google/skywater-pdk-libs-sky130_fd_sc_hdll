* File: sky130_fd_sc_hdll__einvn_1.spice
* Created: Thu Aug 27 19:07:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__einvn_1.pex.spice"
.subckt sky130_fd_sc_hdll__einvn_1  VNB VPB TE_B A VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* A	A
* TE_B	TE_B
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_TE_B_M1002_g N_A_27_47#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.206271 AS=0.1302 PD=1.16579 PS=1.46 NRD=15.708 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75002 A=0.063 P=1.14 MULT=1
MM1000 A_316_47# N_A_27_47#_M1000_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.190125 AS=0.319229 PD=1.235 PS=1.80421 NRD=43.836 NRS=29.532 M=1
+ R=4.33333 SA=75001 SB=75001 A=0.0975 P=1.6 MULT=1
MM1005 N_Z_M1005_d N_A_M1005_g A_316_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.190125 PD=1.92 PS=1.235 NRD=8.304 NRS=43.836 M=1 R=4.33333 SA=75001.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_TE_B_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=9.2196 NRS=1.5366 M=1
+ R=3.55556 SA=90000.2 SB=90001.9 A=0.1152 P=1.64 MULT=1
MM1004 A_222_297# N_TE_B_M1004_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1 AD=0.5325
+ AS=0.191707 PD=2.065 PS=1.64024 NRD=94.0478 NRS=6.8753 M=1 R=5.55556
+ SA=90000.5 SB=90001.4 A=0.18 P=2.36 MULT=1
MM1003 N_Z_M1003_d N_A_M1003_g A_222_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.5325 PD=2.54 PS=2.065 NRD=0.9653 NRS=94.0478 M=1 R=5.55556 SA=90001.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX7_noxref noxref_11 Z Z PROBETYPE=1
pX8_noxref noxref_12 Z Z PROBETYPE=1
*
.include "sky130_fd_sc_hdll__einvn_1.pxi.spice"
*
.ends
*
*
