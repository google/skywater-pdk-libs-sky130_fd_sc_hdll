* NGSPICE file created from sky130_fd_sc_hdll__and4bb_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
M1000 a_606_47# D VGND VNB nshort w=650000u l=150000u
+  ad=2.6975e+11p pd=2.13e+06u as=8.552e+11p ps=7.75e+06u
M1001 a_912_21# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=1.9814e+12p ps=1.503e+07u
M1002 VPWR B_N a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_184_21# a_912_21# a_836_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=2.47e+11p ps=2.06e+06u
M1004 a_184_21# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=7.35e+11p pd=5.47e+06u as=0p ps=0u
M1005 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=4.16e+11p ps=3.88e+06u
M1006 VPWR C a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1009 a_836_47# a_27_47# a_719_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.8275e+11p ps=2.17e+06u
M1010 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_184_21# D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_912_21# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=0p ps=0u
M1013 VPWR a_184_21# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND B_N a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1015 VGND a_184_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 X a_184_21# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_719_47# C a_606_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VPWR a_912_21# a_184_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1019 X a_184_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

