* File: sky130_fd_sc_hdll__o21ai_1.pex.spice
* Created: Thu Aug 27 19:19:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%A1 1 3 4 6 7 11
r22 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.325
+ $Y=1.16 $X2=0.325 $Y2=1.16
r23 7 11 3.31764 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.325 $Y2=1.16
r24 4 10 38.952 $w=3.63e-07 $l=2.19875e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.392 $Y2=1.16
r25 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r26 1 10 45.4477 $w=3.63e-07 $l=2.97069e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.392 $Y2=1.16
r27 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%A2 1 3 4 6 7 8 9 10 17
r37 18 29 2.26808 $w=2.55e-07 $l=1.65e-07 $layer=LI1_cond $X=0.707 $Y=1.325
+ $X2=0.707 $Y2=1.16
r38 17 29 8.13695 $w=3.28e-07 $l=2.33e-07 $layer=LI1_cond $X=0.94 $Y=1.16
+ $X2=0.707 $Y2=1.16
r39 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r40 9 10 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.707 $Y=1.87
+ $X2=0.707 $Y2=2.21
r41 8 9 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=0.707 $Y=1.53
+ $X2=0.707 $Y2=1.87
r42 8 18 9.26474 $w=2.53e-07 $l=2.05e-07 $layer=LI1_cond $X=0.707 $Y=1.53
+ $X2=0.707 $Y2=1.325
r43 7 29 0.593683 $w=3.28e-07 $l=1.7e-08 $layer=LI1_cond $X=0.69 $Y=1.16
+ $X2=0.707 $Y2=1.16
r44 4 16 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=1.06 $Y=0.995
+ $X2=0.97 $Y2=1.16
r45 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.06 $Y=0.995 $X2=1.06
+ $Y2=0.56
r46 1 16 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.97 $Y2=1.16
r47 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.905 $Y=1.41
+ $X2=0.905 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%B1 3 5 7 8 11
r30 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.46 $X2=1.75 $Y2=1.46
r31 11 13 32.3534 $w=3.65e-07 $l=2.45e-07 $layer=POLY_cond $X=1.505 $Y=1.502
+ $X2=1.75 $Y2=1.502
r32 10 11 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.48 $Y=1.502
+ $X2=1.505 $Y2=1.502
r33 8 14 10.2439 $w=3.58e-07 $l=3.2e-07 $layer=LI1_cond $X=2.07 $Y=1.475
+ $X2=1.75 $Y2=1.475
r34 5 11 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.505 $Y=1.71
+ $X2=1.505 $Y2=1.502
r35 5 7 113.806 $w=1.8e-07 $l=4.25e-07 $layer=POLY_cond $X=1.505 $Y=1.71
+ $X2=1.505 $Y2=2.135
r36 1 10 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=1.295
+ $X2=1.48 $Y2=1.502
r37 1 3 376.883 $w=1.5e-07 $l=7.35e-07 $layer=POLY_cond $X=1.48 $Y=1.295
+ $X2=1.48 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%VPWR 1 2 7 9 13 15 17 19 32
r26 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r27 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r28 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r29 23 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r30 22 25 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r31 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r32 20 28 4.70099 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=0.205 $Y2=2.72
r33 20 22 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=0.41 $Y=2.72
+ $X2=0.69 $Y2=2.72
r34 19 31 5.76191 $w=1.7e-07 $l=3.27e-07 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.972 $Y2=2.72
r35 19 25 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=1.645 $Y=2.72
+ $X2=1.61 $Y2=2.72
r36 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r37 17 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r38 13 31 3.17169 $w=4.65e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.877 $Y=2.635
+ $X2=1.972 $Y2=2.72
r39 13 15 16.3335 $w=4.63e-07 $l=6.35e-07 $layer=LI1_cond $X=1.877 $Y=2.635
+ $X2=1.877 $Y2=2
r40 9 12 24.4894 $w=3.18e-07 $l=6.8e-07 $layer=LI1_cond $X=0.25 $Y=1.66 $X2=0.25
+ $Y2=2.34
r41 7 28 2.98112 $w=3.2e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.205 $Y2=2.72
r42 7 12 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.25 $Y=2.635
+ $X2=0.25 $Y2=2.34
r43 2 15 300 $w=1.7e-07 $l=3.82688e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.785 $X2=1.885 $Y2=2
r44 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r45 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%Y 1 2 9 10 13 15 16 17 18
r33 18 24 5.90276 $w=4.08e-07 $l=2.1e-07 $layer=LI1_cond $X=1.21 $Y=2.21
+ $X2=1.21 $Y2=2
r34 17 24 3.65409 $w=4.08e-07 $l=1.3e-07 $layer=LI1_cond $X=1.21 $Y=1.87
+ $X2=1.21 $Y2=2
r35 15 17 4.49734 $w=4.08e-07 $l=1.6e-07 $layer=LI1_cond $X=1.21 $Y=1.71
+ $X2=1.21 $Y2=1.87
r36 15 16 9.81506 $w=4.08e-07 $l=2.05e-07 $layer=LI1_cond $X=1.21 $Y=1.71
+ $X2=1.21 $Y2=1.505
r37 11 13 15.3047 $w=4.63e-07 $l=5.95e-07 $layer=LI1_cond $X=1.877 $Y=0.955
+ $X2=1.877 $Y2=0.36
r38 9 11 8.93361 $w=1.7e-07 $l=2.7119e-07 $layer=LI1_cond $X=1.645 $Y=1.04
+ $X2=1.877 $Y2=0.955
r39 9 10 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.645 $Y=1.04
+ $X2=1.415 $Y2=1.04
r40 7 10 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.33 $Y=1.125
+ $X2=1.415 $Y2=1.04
r41 7 16 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.33 $Y=1.125
+ $X2=1.33 $Y2=1.505
r42 2 24 300 $w=1.7e-07 $l=6.2149e-07 $layer=licon1_PDIFF $count=2 $X=0.995
+ $Y=1.485 $X2=1.23 $Y2=2
r43 1 13 91 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_NDIFF $count=2 $X=1.555
+ $Y=0.235 $X2=1.885 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%A_27_47# 1 2 9 11 12 15
r24 13 15 7.01487 $w=2.28e-07 $l=1.4e-07 $layer=LI1_cond $X=1.29 $Y=0.615
+ $X2=1.29 $Y2=0.475
r25 11 13 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=1.175 $Y=0.7
+ $X2=1.29 $Y2=0.615
r26 11 12 51.8663 $w=1.68e-07 $l=7.95e-07 $layer=LI1_cond $X=1.175 $Y=0.7
+ $X2=0.38 $Y2=0.7
r27 7 12 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=0.235 $Y=0.615
+ $X2=0.38 $Y2=0.7
r28 7 9 7.35179 $w=2.88e-07 $l=1.85e-07 $layer=LI1_cond $X=0.235 $Y=0.615
+ $X2=0.235 $Y2=0.43
r29 2 15 182 $w=1.7e-07 $l=3e-07 $layer=licon1_NDIFF $count=1 $X=1.135 $Y=0.235
+ $X2=1.27 $Y2=0.475
r30 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_1%VGND 1 6 13 14 18 24
r25 18 21 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.815
+ $Y2=0.36
r26 18 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r27 13 14 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r28 11 14 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r29 11 19 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r30 10 13 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r31 10 11 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r32 8 18 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=0.815
+ $Y2=0
r33 8 10 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=1.005 $Y=0 $X2=1.15
+ $Y2=0
r34 6 19 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.69
+ $Y2=0
r35 6 24 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r36 1 21 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.79 $Y2=0.36
.ends

