* File: sky130_fd_sc_hdll__clkinv_16.pex.spice
* Created: Wed Sep  2 08:26:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_16%A 1 3 4 6 7 9 10 12 15 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 47 50 52 54 57 59 61 62 63 66 68 70 73 75 77 80 82 84 87
+ 89 91 94 96 98 101 103 105 108 110 112 115 117 119 122 124 126 127 129 130 132
+ 133 135 136 138 139 141 146 147 148 150 202 203
c296 124 0 1.08667e-19 $X=9.82 $Y=1.41
c297 117 0 1.08667e-19 $X=9.34 $Y=1.41
c298 110 0 1.08667e-19 $X=8.86 $Y=1.41
c299 103 0 1.08667e-19 $X=8.38 $Y=1.41
c300 96 0 1.08667e-19 $X=7.9 $Y=1.41
c301 89 0 1.08667e-19 $X=7.42 $Y=1.41
c302 82 0 1.08667e-19 $X=6.94 $Y=1.41
c303 75 0 1.08667e-19 $X=6.46 $Y=1.41
c304 68 0 1.14801e-19 $X=5.98 $Y=1.41
c305 59 0 1.24926e-19 $X=5.345 $Y=1.41
c306 52 0 1.0646e-19 $X=4.83 $Y=1.41
c307 45 0 1.07837e-19 $X=4.35 $Y=1.41
c308 38 0 1.09776e-19 $X=3.87 $Y=1.41
c309 31 0 1.09072e-19 $X=3.39 $Y=1.41
c310 24 0 1.0723e-19 $X=2.91 $Y=1.41
c311 17 0 1.02518e-19 $X=2.43 $Y=1.41
r312 202 204 16.2332 $w=3.86e-07 $l=1.3e-07 $layer=POLY_cond $X=11.61 $Y=1.2
+ $X2=11.74 $Y2=1.2
r313 202 203 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=11.61
+ $Y=1.16 $X2=11.61 $Y2=1.16
r314 200 202 43.7047 $w=3.86e-07 $l=3.5e-07 $layer=POLY_cond $X=11.26 $Y=1.2
+ $X2=11.61 $Y2=1.2
r315 199 200 59.9378 $w=3.86e-07 $l=4.8e-07 $layer=POLY_cond $X=10.78 $Y=1.2
+ $X2=11.26 $Y2=1.2
r316 198 199 59.9378 $w=3.86e-07 $l=4.8e-07 $layer=POLY_cond $X=10.3 $Y=1.2
+ $X2=10.78 $Y2=1.2
r317 196 198 24.9741 $w=3.86e-07 $l=2e-07 $layer=POLY_cond $X=10.1 $Y=1.2
+ $X2=10.3 $Y2=1.2
r318 196 197 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=10.1
+ $Y=1.16 $X2=10.1 $Y2=1.16
r319 194 196 34.9637 $w=3.86e-07 $l=2.8e-07 $layer=POLY_cond $X=9.82 $Y=1.2
+ $X2=10.1 $Y2=1.2
r320 193 194 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=9.795 $Y=1.2
+ $X2=9.82 $Y2=1.2
r321 192 193 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=9.34 $Y=1.2
+ $X2=9.795 $Y2=1.2
r322 191 192 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=9.315 $Y=1.2
+ $X2=9.34 $Y2=1.2
r323 190 191 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=8.86 $Y=1.2
+ $X2=9.315 $Y2=1.2
r324 189 190 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=8.835 $Y=1.2
+ $X2=8.86 $Y2=1.2
r325 188 189 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=8.38 $Y=1.2
+ $X2=8.835 $Y2=1.2
r326 187 188 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=8.355 $Y=1.2
+ $X2=8.38 $Y2=1.2
r327 186 187 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=7.9 $Y=1.2
+ $X2=8.355 $Y2=1.2
r328 185 186 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=7.875 $Y=1.2
+ $X2=7.9 $Y2=1.2
r329 184 185 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=7.42 $Y=1.2
+ $X2=7.875 $Y2=1.2
r330 183 184 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=7.395 $Y=1.2
+ $X2=7.42 $Y2=1.2
r331 182 183 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=6.94 $Y=1.2
+ $X2=7.395 $Y2=1.2
r332 181 182 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=6.915 $Y=1.2
+ $X2=6.94 $Y2=1.2
r333 180 181 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=6.46 $Y=1.2
+ $X2=6.915 $Y2=1.2
r334 179 180 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=6.435 $Y=1.2
+ $X2=6.46 $Y2=1.2
r335 178 179 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=5.98 $Y=1.2
+ $X2=6.435 $Y2=1.2
r336 177 178 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=5.955 $Y=1.2
+ $X2=5.98 $Y2=1.2
r337 175 176 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=5.32 $Y=1.2
+ $X2=5.345 $Y2=1.2
r338 174 175 61.1865 $w=3.86e-07 $l=4.9e-07 $layer=POLY_cond $X=4.83 $Y=1.2
+ $X2=5.32 $Y2=1.2
r339 173 174 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=4.805 $Y=1.2
+ $X2=4.83 $Y2=1.2
r340 172 173 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=4.35 $Y=1.2
+ $X2=4.805 $Y2=1.2
r341 171 172 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=4.325 $Y=1.2
+ $X2=4.35 $Y2=1.2
r342 170 171 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=3.87 $Y=1.2
+ $X2=4.325 $Y2=1.2
r343 169 170 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=3.845 $Y=1.2
+ $X2=3.87 $Y2=1.2
r344 168 169 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=3.39 $Y=1.2
+ $X2=3.845 $Y2=1.2
r345 167 168 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=3.365 $Y=1.2
+ $X2=3.39 $Y2=1.2
r346 166 167 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=2.91 $Y=1.2
+ $X2=3.365 $Y2=1.2
r347 165 166 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=2.885 $Y=1.2
+ $X2=2.91 $Y2=1.2
r348 164 165 56.8161 $w=3.86e-07 $l=4.55e-07 $layer=POLY_cond $X=2.43 $Y=1.2
+ $X2=2.885 $Y2=1.2
r349 163 164 3.12176 $w=3.86e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.2
+ $X2=2.43 $Y2=1.2
r350 161 163 31.842 $w=3.86e-07 $l=2.55e-07 $layer=POLY_cond $X=2.15 $Y=1.2
+ $X2=2.405 $Y2=1.2
r351 159 161 24.9741 $w=3.86e-07 $l=2e-07 $layer=POLY_cond $X=1.95 $Y=1.2
+ $X2=2.15 $Y2=1.2
r352 158 159 59.9378 $w=3.86e-07 $l=4.8e-07 $layer=POLY_cond $X=1.47 $Y=1.2
+ $X2=1.95 $Y2=1.2
r353 157 158 59.9378 $w=3.86e-07 $l=4.8e-07 $layer=POLY_cond $X=0.99 $Y=1.2
+ $X2=1.47 $Y2=1.2
r354 155 157 49.9482 $w=3.86e-07 $l=4e-07 $layer=POLY_cond $X=0.59 $Y=1.2
+ $X2=0.99 $Y2=1.2
r355 155 156 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.59
+ $Y=1.16 $X2=0.59 $Y2=1.16
r356 153 155 9.98964 $w=3.86e-07 $l=8e-08 $layer=POLY_cond $X=0.51 $Y=1.2
+ $X2=0.59 $Y2=1.2
r357 151 203 18.803 $w=3.78e-07 $l=6.2e-07 $layer=LI1_cond $X=10.99 $Y=1.085
+ $X2=11.61 $Y2=1.085
r358 151 197 26.9914 $w=3.78e-07 $l=8.9e-07 $layer=LI1_cond $X=10.99 $Y=1.085
+ $X2=10.1 $Y2=1.085
r359 150 151 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.99 $Y=1.19
+ $X2=10.99 $Y2=1.19
r360 148 150 0.378547 $w=2.3e-07 $l=5.9e-07 $layer=MET1_cond $X=10.4 $Y=1.19
+ $X2=10.99 $Y2=1.19
r361 146 148 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=10.285 $Y=1.19
+ $X2=10.4 $Y2=1.19
r362 146 147 9.74008 $w=1.4e-07 $l=7.87e-06 $layer=MET1_cond $X=10.285 $Y=1.19
+ $X2=2.415 $Y2=1.19
r363 141 147 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=2.3 $Y=1.19
+ $X2=2.415 $Y2=1.19
r364 141 143 0.0192481 $w=2.3e-07 $l=3e-08 $layer=MET1_cond $X=2.3 $Y=1.19
+ $X2=2.27 $Y2=1.19
r365 139 156 44.8846 $w=3.78e-07 $l=1.48e-06 $layer=LI1_cond $X=2.07 $Y=1.085
+ $X2=0.59 $Y2=1.085
r366 139 161 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r367 139 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.27 $Y=1.19
+ $X2=2.27 $Y2=1.19
r368 136 204 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=11.74 $Y=1.41
+ $X2=11.74 $Y2=1.2
r369 136 138 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.74 $Y=1.41
+ $X2=11.74 $Y2=1.985
r370 133 200 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=11.26 $Y=1.41
+ $X2=11.26 $Y2=1.2
r371 133 135 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.26 $Y=1.41
+ $X2=11.26 $Y2=1.985
r372 130 199 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=10.78 $Y=1.41
+ $X2=10.78 $Y2=1.2
r373 130 132 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.78 $Y=1.41
+ $X2=10.78 $Y2=1.985
r374 127 198 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=10.3 $Y=1.41
+ $X2=10.3 $Y2=1.2
r375 127 129 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.3 $Y=1.41
+ $X2=10.3 $Y2=1.985
r376 124 194 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=9.82 $Y=1.41
+ $X2=9.82 $Y2=1.2
r377 124 126 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.82 $Y=1.41
+ $X2=9.82 $Y2=1.985
r378 120 193 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.795 $Y=0.99
+ $X2=9.795 $Y2=1.2
r379 120 122 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=9.795 $Y=0.99
+ $X2=9.795 $Y2=0.445
r380 117 192 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=9.34 $Y=1.41
+ $X2=9.34 $Y2=1.2
r381 117 119 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.34 $Y=1.41
+ $X2=9.34 $Y2=1.985
r382 113 191 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=9.315 $Y=0.99
+ $X2=9.315 $Y2=1.2
r383 113 115 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=9.315 $Y=0.99
+ $X2=9.315 $Y2=0.445
r384 110 190 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.86 $Y=1.41
+ $X2=8.86 $Y2=1.2
r385 110 112 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.86 $Y=1.41
+ $X2=8.86 $Y2=1.985
r386 106 189 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.835 $Y=0.99
+ $X2=8.835 $Y2=1.2
r387 106 108 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.835 $Y=0.99
+ $X2=8.835 $Y2=0.445
r388 103 188 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=8.38 $Y=1.41
+ $X2=8.38 $Y2=1.2
r389 103 105 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.38 $Y=1.41
+ $X2=8.38 $Y2=1.985
r390 99 187 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=8.355 $Y=0.99
+ $X2=8.355 $Y2=1.2
r391 99 101 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=8.355 $Y=0.99
+ $X2=8.355 $Y2=0.445
r392 96 186 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=7.9 $Y=1.41
+ $X2=7.9 $Y2=1.2
r393 96 98 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.9 $Y=1.41
+ $X2=7.9 $Y2=1.985
r394 92 185 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.875 $Y=0.99
+ $X2=7.875 $Y2=1.2
r395 92 94 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.875 $Y=0.99
+ $X2=7.875 $Y2=0.445
r396 89 184 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=7.42 $Y=1.41
+ $X2=7.42 $Y2=1.2
r397 89 91 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.42 $Y=1.41
+ $X2=7.42 $Y2=1.985
r398 85 183 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=7.395 $Y=0.99
+ $X2=7.395 $Y2=1.2
r399 85 87 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=7.395 $Y=0.99
+ $X2=7.395 $Y2=0.445
r400 82 182 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=6.94 $Y=1.41
+ $X2=6.94 $Y2=1.2
r401 82 84 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.94 $Y=1.41
+ $X2=6.94 $Y2=1.985
r402 78 181 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.915 $Y=0.99
+ $X2=6.915 $Y2=1.2
r403 78 80 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.915 $Y=0.99
+ $X2=6.915 $Y2=0.445
r404 75 180 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=6.46 $Y=1.41
+ $X2=6.46 $Y2=1.2
r405 75 77 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.46 $Y=1.41
+ $X2=6.46 $Y2=1.985
r406 71 179 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=6.435 $Y=0.99
+ $X2=6.435 $Y2=1.2
r407 71 73 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=6.435 $Y=0.99
+ $X2=6.435 $Y2=0.445
r408 68 178 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.98 $Y=1.41
+ $X2=5.98 $Y2=1.2
r409 68 70 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.98 $Y=1.41
+ $X2=5.98 $Y2=1.985
r410 64 177 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.955 $Y=0.99
+ $X2=5.955 $Y2=1.2
r411 64 66 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.955 $Y=0.99
+ $X2=5.955 $Y2=0.445
r412 63 176 12.7749 $w=3.86e-07 $l=1.14018e-07 $layer=POLY_cond $X=5.445 $Y=1.17
+ $X2=5.345 $Y2=1.2
r413 62 177 9.65311 $w=3.86e-07 $l=8.87412e-08 $layer=POLY_cond $X=5.88 $Y=1.17
+ $X2=5.955 $Y2=1.2
r414 62 63 69.7259 $w=3.6e-07 $l=4.35e-07 $layer=POLY_cond $X=5.88 $Y=1.17
+ $X2=5.445 $Y2=1.17
r415 59 176 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=5.345 $Y=1.41
+ $X2=5.345 $Y2=1.2
r416 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.345 $Y=1.41
+ $X2=5.345 $Y2=1.985
r417 55 175 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=5.32 $Y=0.99
+ $X2=5.32 $Y2=1.2
r418 55 57 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=5.32 $Y=0.99
+ $X2=5.32 $Y2=0.445
r419 52 174 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.83 $Y=1.41
+ $X2=4.83 $Y2=1.2
r420 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.83 $Y=1.41
+ $X2=4.83 $Y2=1.985
r421 48 173 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.805 $Y=0.99
+ $X2=4.805 $Y2=1.2
r422 48 50 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.805 $Y=0.99
+ $X2=4.805 $Y2=0.445
r423 45 172 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=4.35 $Y=1.41
+ $X2=4.35 $Y2=1.2
r424 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.35 $Y=1.41
+ $X2=4.35 $Y2=1.985
r425 41 171 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=4.325 $Y=0.99
+ $X2=4.325 $Y2=1.2
r426 41 43 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=4.325 $Y=0.99
+ $X2=4.325 $Y2=0.445
r427 38 170 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.87 $Y=1.41
+ $X2=3.87 $Y2=1.2
r428 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.87 $Y=1.41
+ $X2=3.87 $Y2=1.985
r429 34 169 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.845 $Y=0.99
+ $X2=3.845 $Y2=1.2
r430 34 36 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.845 $Y=0.99
+ $X2=3.845 $Y2=0.445
r431 31 168 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=3.39 $Y=1.41
+ $X2=3.39 $Y2=1.2
r432 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.39 $Y=1.41
+ $X2=3.39 $Y2=1.985
r433 27 167 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.365 $Y=0.99
+ $X2=3.365 $Y2=1.2
r434 27 29 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=3.365 $Y=0.99
+ $X2=3.365 $Y2=0.445
r435 24 166 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.2
r436 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.91 $Y=1.41
+ $X2=2.91 $Y2=1.985
r437 20 165 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.885 $Y=0.99
+ $X2=2.885 $Y2=1.2
r438 20 22 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.885 $Y=0.99
+ $X2=2.885 $Y2=0.445
r439 17 164 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.2
r440 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.985
r441 13 163 24.9932 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.405 $Y=0.99
+ $X2=2.405 $Y2=1.2
r442 13 15 279.457 $w=1.5e-07 $l=5.45e-07 $layer=POLY_cond $X=2.405 $Y=0.99
+ $X2=2.405 $Y2=0.445
r443 10 159 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.95 $Y=1.41
+ $X2=1.95 $Y2=1.2
r444 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.95 $Y=1.41
+ $X2=1.95 $Y2=1.985
r445 7 158 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.47 $Y2=1.2
r446 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.47 $Y2=1.985
r447 4 157 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.2
r448 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.985
r449 1 153 20.6153 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.2
r450 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.51 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 46 50 52 56 60 64 68 72 77 78 82 84 88 92 96 100 104 107 108 110 111 113 114
+ 117 118 120 121 123 124 126 127 128 140 158 159 165 168 171 174 177
r173 177 178 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r174 175 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r175 174 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r176 172 175 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r177 171 172 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r178 168 169 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r179 166 169 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r180 165 166 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r181 158 159 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r182 156 159 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r183 155 156 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r184 153 156 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r185 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r186 150 153 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r187 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r188 147 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r189 147 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.05 $Y2=2.72
r190 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r191 144 177 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=8.27 $Y=2.72
+ $X2=8.142 $Y2=2.72
r192 144 146 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.27 $Y=2.72
+ $X2=8.97 $Y2=2.72
r193 143 172 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r194 142 143 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r195 140 171 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=6.22 $Y2=2.72
r196 140 142 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=2.72
+ $X2=5.75 $Y2=2.72
r197 139 143 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r198 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r199 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r200 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r201 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r202 133 169 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r203 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r204 130 168 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=2.32 $Y=2.72
+ $X2=2.192 $Y2=2.72
r205 130 132 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.32 $Y=2.72
+ $X2=2.99 $Y2=2.72
r206 128 166 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r207 128 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r208 126 155 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=11.85 $Y=2.72
+ $X2=11.73 $Y2=2.72
r209 126 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.85 $Y=2.72
+ $X2=11.98 $Y2=2.72
r210 125 158 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=12.11 $Y=2.72
+ $X2=12.19 $Y2=2.72
r211 125 127 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=12.11 $Y=2.72
+ $X2=11.98 $Y2=2.72
r212 123 152 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.895 $Y=2.72
+ $X2=10.81 $Y2=2.72
r213 123 124 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.895 $Y=2.72
+ $X2=11.022 $Y2=2.72
r214 122 155 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=11.15 $Y=2.72
+ $X2=11.73 $Y2=2.72
r215 122 124 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=11.15 $Y=2.72
+ $X2=11.022 $Y2=2.72
r216 120 149 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=9.89 $Y2=2.72
r217 120 121 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=9.935 $Y=2.72
+ $X2=10.062 $Y2=2.72
r218 119 152 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=10.81 $Y2=2.72
r219 119 121 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.19 $Y=2.72
+ $X2=10.062 $Y2=2.72
r220 117 146 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=8.975 $Y=2.72
+ $X2=8.97 $Y2=2.72
r221 117 118 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.975 $Y=2.72
+ $X2=9.102 $Y2=2.72
r222 116 149 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=9.23 $Y=2.72
+ $X2=9.89 $Y2=2.72
r223 116 118 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=9.23 $Y=2.72
+ $X2=9.102 $Y2=2.72
r224 113 138 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=4.83 $Y2=2.72
r225 113 114 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.965 $Y=2.72
+ $X2=5.092 $Y2=2.72
r226 112 142 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.75 $Y2=2.72
r227 112 114 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=5.22 $Y=2.72
+ $X2=5.092 $Y2=2.72
r228 110 135 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=3.91 $Y2=2.72
r229 110 111 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=4.112 $Y2=2.72
r230 109 138 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.24 $Y=2.72
+ $X2=4.83 $Y2=2.72
r231 109 111 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=4.24 $Y=2.72
+ $X2=4.112 $Y2=2.72
r232 107 132 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=2.99 $Y2=2.72
r233 107 108 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=3.15 $Y2=2.72
r234 106 135 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=3.28 $Y=2.72
+ $X2=3.91 $Y2=2.72
r235 106 108 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.28 $Y=2.72
+ $X2=3.15 $Y2=2.72
r236 102 127 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=11.98 $Y=2.635
+ $X2=11.98 $Y2=2.72
r237 102 104 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=11.98 $Y=2.635
+ $X2=11.98 $Y2=2
r238 98 124 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=11.022 $Y=2.635
+ $X2=11.022 $Y2=2.72
r239 98 100 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=11.022 $Y=2.635
+ $X2=11.022 $Y2=2
r240 94 121 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.062 $Y=2.635
+ $X2=10.062 $Y2=2.72
r241 94 96 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=10.062 $Y=2.635
+ $X2=10.062 $Y2=2
r242 90 118 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.102 $Y=2.635
+ $X2=9.102 $Y2=2.72
r243 90 92 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=9.102 $Y=2.635
+ $X2=9.102 $Y2=2
r244 86 177 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=8.142 $Y=2.635
+ $X2=8.142 $Y2=2.72
r245 86 88 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=8.142 $Y=2.635
+ $X2=8.142 $Y2=2
r246 85 174 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=7.31 $Y=2.72
+ $X2=7.182 $Y2=2.72
r247 84 177 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=8.015 $Y=2.72
+ $X2=8.142 $Y2=2.72
r248 84 85 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=8.015 $Y=2.72
+ $X2=7.31 $Y2=2.72
r249 80 174 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=7.182 $Y=2.635
+ $X2=7.182 $Y2=2.72
r250 80 82 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=7.182 $Y=2.635
+ $X2=7.182 $Y2=2
r251 79 171 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.35 $Y=2.72
+ $X2=6.22 $Y2=2.72
r252 78 174 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=7.182 $Y2=2.72
r253 78 79 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=7.055 $Y=2.72
+ $X2=6.35 $Y2=2.72
r254 75 171 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.72
r255 75 77 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=6.22 $Y=2.635
+ $X2=6.22 $Y2=2.34
r256 74 115 5.76222 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=6.22 $Y=2.25
+ $X2=6.22 $Y2=2.12
r257 74 77 3.98923 $w=2.58e-07 $l=9e-08 $layer=LI1_cond $X=6.22 $Y=2.25 $X2=6.22
+ $Y2=2.34
r258 72 115 5.42326 $w=2.53e-07 $l=1.2e-07 $layer=LI1_cond $X=6.217 $Y=2
+ $X2=6.217 $Y2=2.12
r259 66 114 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=5.092 $Y=2.635
+ $X2=5.092 $Y2=2.72
r260 66 68 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=5.092 $Y=2.635
+ $X2=5.092 $Y2=2
r261 62 111 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.112 $Y=2.635
+ $X2=4.112 $Y2=2.72
r262 62 64 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=4.112 $Y=2.635
+ $X2=4.112 $Y2=2
r263 58 108 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.15 $Y=2.635
+ $X2=3.15 $Y2=2.72
r264 58 60 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=3.15 $Y=2.635
+ $X2=3.15 $Y2=2
r265 54 168 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=2.192 $Y=2.635
+ $X2=2.192 $Y2=2.72
r266 54 56 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=2.192 $Y=2.635
+ $X2=2.192 $Y2=2
r267 53 165 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.36 $Y=2.72
+ $X2=1.23 $Y2=2.72
r268 52 168 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.192 $Y2=2.72
r269 52 53 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.36 $Y2=2.72
r270 48 165 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2.72
r271 48 50 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=1.23 $Y=2.635
+ $X2=1.23 $Y2=2
r272 47 162 4.10994 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r273 46 165 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.1 $Y=2.72
+ $X2=1.23 $Y2=2.72
r274 46 47 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.1 $Y=2.72
+ $X2=0.405 $Y2=2.72
r275 42 45 29.5721 $w=2.63e-07 $l=6.8e-07 $layer=LI1_cond $X=0.272 $Y=1.66
+ $X2=0.272 $Y2=2.34
r276 40 162 3.13813 $w=2.65e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.272 $Y=2.635
+ $X2=0.202 $Y2=2.72
r277 40 45 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=0.272 $Y=2.635
+ $X2=0.272 $Y2=2.34
r278 13 104 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=11.83
+ $Y=1.485 $X2=11.975 $Y2=2
r279 12 100 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=10.87
+ $Y=1.485 $X2=11.02 $Y2=2
r280 11 96 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=9.91
+ $Y=1.485 $X2=10.06 $Y2=2
r281 10 92 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=8.95
+ $Y=1.485 $X2=9.1 $Y2=2
r282 9 88 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=7.99
+ $Y=1.485 $X2=8.14 $Y2=2
r283 8 82 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=7.03
+ $Y=1.485 $X2=7.18 $Y2=2
r284 7 77 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.215 $Y2=2.34
r285 7 72 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=6.07
+ $Y=1.485 $X2=6.215 $Y2=2
r286 6 68 300 $w=1.7e-07 $l=5.93949e-07 $layer=licon1_PDIFF $count=2 $X=4.92
+ $Y=1.485 $X2=5.09 $Y2=2
r287 5 64 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=3.96
+ $Y=1.485 $X2=4.11 $Y2=2
r288 4 60 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=3
+ $Y=1.485 $X2=3.15 $Y2=2
r289 3 56 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.04
+ $Y=1.485 $X2=2.19 $Y2=2
r290 2 50 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.08
+ $Y=1.485 $X2=1.23 $Y2=2
r291 1 45 400 $w=1.7e-07 $l=9.22348e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=2.34
r292 1 42 400 $w=1.7e-07 $l=2.34787e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.275 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_16%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 19 20 61 63 65 69 73 77 81 85 89 93 96 100 106 110 114 118 122 126 130
+ 134 138 145 147 149 151 152 154 156 158 160 162 164 165
c222 165 0 8.51807e-20 $X=5.675 $Y=1.445
c223 130 0 2.17334e-19 $X=9.58 $Y=0.445
c224 122 0 2.17334e-19 $X=8.62 $Y=0.445
c225 114 0 2.17334e-19 $X=7.66 $Y=0.445
c226 106 0 2.17334e-19 $X=6.7 $Y=0.445
c227 100 0 2.39727e-19 $X=5.615 $Y=0.445
c228 89 0 2.14296e-19 $X=4.59 $Y=0.445
c229 81 0 2.18848e-19 $X=3.63 $Y=0.445
c230 73 0 2.09748e-19 $X=2.67 $Y=0.445
r231 165 168 4.25218 $w=2.5e-07 $l=1.88e-07 $layer=LI1_cond $X=5.642 $Y=1.54
+ $X2=5.83 $Y2=1.54
r232 165 168 0.322684 $w=2.48e-07 $l=7e-09 $layer=LI1_cond $X=5.837 $Y=1.54
+ $X2=5.83 $Y2=1.54
r233 152 165 34.0201 $w=2.48e-07 $l=7.38e-07 $layer=LI1_cond $X=6.575 $Y=1.54
+ $X2=5.837 $Y2=1.54
r234 152 154 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.575 $Y=1.54 $X2=6.7
+ $Y2=1.54
r235 139 162 5.7647 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=10.655 $Y=1.56
+ $X2=10.535 $Y2=1.56
r236 138 164 3.77708 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=11.375 $Y=1.56
+ $X2=11.502 $Y2=1.56
r237 138 139 38.026 $w=2.08e-07 $l=7.2e-07 $layer=LI1_cond $X=11.375 $Y=1.56
+ $X2=10.655 $Y2=1.56
r238 135 160 3.30809 $w=2.1e-07 $l=1.34629e-07 $layer=LI1_cond $X=9.705 $Y=1.56
+ $X2=9.58 $Y2=1.54
r239 134 162 5.7647 $w=2.1e-07 $l=1.2e-07 $layer=LI1_cond $X=10.415 $Y=1.56
+ $X2=10.535 $Y2=1.56
r240 134 135 37.4978 $w=2.08e-07 $l=7.1e-07 $layer=LI1_cond $X=10.415 $Y=1.56
+ $X2=9.705 $Y2=1.56
r241 128 160 2.79962 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=9.58 $Y=1.415
+ $X2=9.58 $Y2=1.54
r242 128 130 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=9.58 $Y=1.415
+ $X2=9.58 $Y2=0.445
r243 127 158 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.745 $Y=1.54
+ $X2=8.62 $Y2=1.54
r244 126 160 3.30809 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=9.455 $Y=1.54
+ $X2=9.58 $Y2=1.54
r245 126 127 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=9.455 $Y=1.54
+ $X2=8.745 $Y2=1.54
r246 120 158 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.62 $Y=1.415
+ $X2=8.62 $Y2=1.54
r247 120 122 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=8.62 $Y=1.415
+ $X2=8.62 $Y2=0.445
r248 119 156 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.785 $Y=1.54
+ $X2=7.66 $Y2=1.54
r249 118 158 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=8.495 $Y=1.54
+ $X2=8.62 $Y2=1.54
r250 118 119 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=8.495 $Y=1.54
+ $X2=7.785 $Y2=1.54
r251 112 156 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.66 $Y=1.415
+ $X2=7.66 $Y2=1.54
r252 112 114 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=7.66 $Y=1.415
+ $X2=7.66 $Y2=0.445
r253 111 154 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.825 $Y=1.54 $X2=6.7
+ $Y2=1.54
r254 110 156 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=7.535 $Y=1.54
+ $X2=7.66 $Y2=1.54
r255 110 111 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=7.535 $Y=1.54
+ $X2=6.825 $Y2=1.54
r256 104 154 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=6.7 $Y=1.415 $X2=6.7
+ $Y2=1.54
r257 104 106 44.7148 $w=2.48e-07 $l=9.7e-07 $layer=LI1_cond $X=6.7 $Y=1.415
+ $X2=6.7 $Y2=0.445
r258 98 165 1.99954 $w=3.5e-07 $l=1.30863e-07 $layer=LI1_cond $X=5.63 $Y=1.415
+ $X2=5.642 $Y2=1.54
r259 98 100 31.9391 $w=3.48e-07 $l=9.7e-07 $layer=LI1_cond $X=5.63 $Y=1.415
+ $X2=5.63 $Y2=0.445
r260 94 151 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.705 $Y=1.54
+ $X2=4.585 $Y2=1.54
r261 94 96 26.9672 $w=2.48e-07 $l=5.85e-07 $layer=LI1_cond $X=4.705 $Y=1.54
+ $X2=5.29 $Y2=1.54
r262 93 165 4.25218 $w=2.5e-07 $l=1.87e-07 $layer=LI1_cond $X=5.455 $Y=1.54
+ $X2=5.642 $Y2=1.54
r263 93 96 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.455 $Y=1.54
+ $X2=5.29 $Y2=1.54
r264 87 151 6.35417 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=4.585 $Y=1.415
+ $X2=4.585 $Y2=1.54
r265 87 89 46.5779 $w=2.38e-07 $l=9.7e-07 $layer=LI1_cond $X=4.585 $Y=1.415
+ $X2=4.585 $Y2=0.445
r266 86 149 6.1976 $w=2.5e-07 $l=1.28e-07 $layer=LI1_cond $X=3.76 $Y=1.54
+ $X2=3.632 $Y2=1.54
r267 85 151 5.856 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=4.465 $Y=1.54
+ $X2=4.585 $Y2=1.54
r268 85 86 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=4.465 $Y=1.54
+ $X2=3.76 $Y2=1.54
r269 79 149 5.98039 $w=2.55e-07 $l=1.25e-07 $layer=LI1_cond $X=3.632 $Y=1.415
+ $X2=3.632 $Y2=1.54
r270 79 81 43.838 $w=2.53e-07 $l=9.7e-07 $layer=LI1_cond $X=3.632 $Y=1.415
+ $X2=3.632 $Y2=0.445
r271 78 147 2.98324 $w=2.5e-07 $l=1.13e-07 $layer=LI1_cond $X=2.8 $Y=1.54
+ $X2=2.687 $Y2=1.54
r272 77 149 6.1976 $w=2.5e-07 $l=1.27e-07 $layer=LI1_cond $X=3.505 $Y=1.54
+ $X2=3.632 $Y2=1.54
r273 77 78 32.4989 $w=2.48e-07 $l=7.05e-07 $layer=LI1_cond $X=3.505 $Y=1.54
+ $X2=2.8 $Y2=1.54
r274 71 147 3.11731 $w=2.25e-07 $l=1.25e-07 $layer=LI1_cond $X=2.687 $Y=1.415
+ $X2=2.687 $Y2=1.54
r275 71 73 49.6831 $w=2.23e-07 $l=9.7e-07 $layer=LI1_cond $X=2.687 $Y=1.415
+ $X2=2.687 $Y2=0.445
r276 70 145 6.05271 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=1.84 $Y=1.56
+ $X2=1.712 $Y2=1.56
r277 69 147 2.98324 $w=2.1e-07 $l=1.21589e-07 $layer=LI1_cond $X=2.575 $Y=1.56
+ $X2=2.687 $Y2=1.54
r278 69 70 38.8182 $w=2.08e-07 $l=7.35e-07 $layer=LI1_cond $X=2.575 $Y=1.56
+ $X2=1.84 $Y2=1.56
r279 66 143 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.88 $Y=1.56
+ $X2=0.752 $Y2=1.56
r280 65 145 6.05271 $w=2.1e-07 $l=1.27e-07 $layer=LI1_cond $X=1.585 $Y=1.56
+ $X2=1.712 $Y2=1.56
r281 65 66 37.2338 $w=2.08e-07 $l=7.05e-07 $layer=LI1_cond $X=1.585 $Y=1.56
+ $X2=0.88 $Y2=1.56
r282 61 143 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.752 $Y=1.665
+ $X2=0.752 $Y2=1.56
r283 61 63 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.752 $Y=1.665
+ $X2=0.752 $Y2=2.3
r284 20 164 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=11.35
+ $Y=1.485 $X2=11.5 $Y2=1.62
r285 19 162 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=10.39
+ $Y=1.485 $X2=10.54 $Y2=1.62
r286 18 160 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=9.43
+ $Y=1.485 $X2=9.58 $Y2=1.62
r287 17 158 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=8.47
+ $Y=1.485 $X2=8.62 $Y2=1.62
r288 16 156 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=7.51
+ $Y=1.485 $X2=7.66 $Y2=1.62
r289 15 154 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=6.55
+ $Y=1.485 $X2=6.7 $Y2=1.62
r290 14 165 300 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_PDIFF $count=2 $X=5.435
+ $Y=1.485 $X2=5.715 $Y2=1.62
r291 13 151 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=4.44
+ $Y=1.485 $X2=4.59 $Y2=1.62
r292 12 149 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=3.48
+ $Y=1.485 $X2=3.63 $Y2=1.62
r293 11 147 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=1.485 $X2=2.67 $Y2=1.62
r294 10 145 300 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=2 $X=1.56
+ $Y=1.485 $X2=1.71 $Y2=1.62
r295 9 143 400 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.75 $Y2=1.62
r296 9 63 400 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=0.6
+ $Y=1.485 $X2=0.75 $Y2=2.3
r297 8 130 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=9.39
+ $Y=0.235 $X2=9.58 $Y2=0.445
r298 7 122 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=8.43
+ $Y=0.235 $X2=8.62 $Y2=0.445
r299 6 114 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=7.47
+ $Y=0.235 $X2=7.66 $Y2=0.445
r300 5 106 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=6.51
+ $Y=0.235 $X2=6.7 $Y2=0.445
r301 4 100 182 $w=1.7e-07 $l=3.07571e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.615 $Y2=0.445
r302 3 89 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.4
+ $Y=0.235 $X2=4.59 $Y2=0.445
r303 2 81 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.44
+ $Y=0.235 $X2=3.63 $Y2=0.445
r304 1 73 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.67 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_16%VGND 1 2 3 4 5 6 7 8 9 30 34 38 42 46 48
+ 52 54 58 60 64 68 71 72 74 75 77 78 80 81 82 84 99 111 112 115 118 121 124 127
r122 127 128 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r123 125 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r124 124 125 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r125 122 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r126 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r127 119 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r128 118 119 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r129 115 116 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r130 111 112 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r131 109 112 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=12.19 $Y2=0
r132 108 111 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=10.35 $Y=0
+ $X2=12.19 $Y2=0
r133 108 109 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r134 106 109 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r135 106 128 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=8.97 $Y2=0
r136 105 106 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r137 103 127 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=9.102 $Y2=0
r138 103 105 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=9.235 $Y=0
+ $X2=9.89 $Y2=0
r139 102 119 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r140 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r141 99 118 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=6.09 $Y=0
+ $X2=6.222 $Y2=0
r142 99 101 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.09 $Y=0 $X2=5.75
+ $Y2=0
r143 98 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r144 97 98 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r145 95 98 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r146 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r147 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r148 92 116 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r149 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r150 89 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.325 $Y=0
+ $X2=2.19 $Y2=0
r151 89 91 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=2.325 $Y=0 $X2=2.99
+ $Y2=0
r152 84 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=2.19 $Y2=0
r153 84 86 119.064 $w=1.68e-07 $l=1.825e-06 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=0.23 $Y2=0
r154 82 116 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=2.07 $Y2=0
r155 82 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r156 80 105 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=9.93 $Y=0 $X2=9.89
+ $Y2=0
r157 80 81 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=9.93 $Y=0
+ $X2=10.062 $Y2=0
r158 79 108 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.35 $Y2=0
r159 79 81 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.062 $Y2=0
r160 77 97 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.965 $Y=0
+ $X2=4.83 $Y2=0
r161 77 78 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=4.965 $Y=0
+ $X2=5.097 $Y2=0
r162 76 101 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.75
+ $Y2=0
r163 76 78 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=5.23 $Y=0 $X2=5.097
+ $Y2=0
r164 74 94 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.98 $Y=0 $X2=3.91
+ $Y2=0
r165 74 75 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.98 $Y=0 $X2=4.112
+ $Y2=0
r166 73 97 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=4.245 $Y=0
+ $X2=4.83 $Y2=0
r167 73 75 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=4.245 $Y=0
+ $X2=4.112 $Y2=0
r168 71 91 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.99
+ $Y2=0
r169 71 72 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.152
+ $Y2=0
r170 70 94 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.91 $Y2=0
r171 70 72 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=3.285 $Y=0
+ $X2=3.152 $Y2=0
r172 66 81 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=10.062 $Y=0.085
+ $X2=10.062 $Y2=0
r173 66 68 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=10.062 $Y=0.085
+ $X2=10.062 $Y2=0.445
r174 62 127 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=9.102 $Y=0.085
+ $X2=9.102 $Y2=0
r175 62 64 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=9.102 $Y=0.085
+ $X2=9.102 $Y2=0.445
r176 61 124 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=8.275 $Y=0
+ $X2=8.142 $Y2=0
r177 60 127 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=9.102 $Y2=0
r178 60 61 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=8.97 $Y=0
+ $X2=8.275 $Y2=0
r179 56 124 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=8.142 $Y=0.085
+ $X2=8.142 $Y2=0
r180 56 58 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=8.142 $Y=0.085
+ $X2=8.142 $Y2=0.445
r181 55 121 6.47928 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.162 $Y2=0
r182 54 124 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=8.01 $Y=0
+ $X2=8.142 $Y2=0
r183 54 55 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=8.01 $Y=0
+ $X2=7.275 $Y2=0
r184 50 121 0.355529 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=7.162 $Y=0.085
+ $X2=7.162 $Y2=0
r185 50 52 18.4391 $w=2.23e-07 $l=3.6e-07 $layer=LI1_cond $X=7.162 $Y=0.085
+ $X2=7.162 $Y2=0.445
r186 49 118 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=6.355 $Y=0
+ $X2=6.222 $Y2=0
r187 48 121 6.47928 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=7.05 $Y=0
+ $X2=7.162 $Y2=0
r188 48 49 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=7.05 $Y=0
+ $X2=6.355 $Y2=0
r189 44 118 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=6.222 $Y=0.085
+ $X2=6.222 $Y2=0
r190 44 46 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=6.222 $Y=0.085
+ $X2=6.222 $Y2=0.445
r191 40 78 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=5.097 $Y=0.085
+ $X2=5.097 $Y2=0
r192 40 42 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=5.097 $Y=0.085
+ $X2=5.097 $Y2=0.445
r193 36 75 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=4.112 $Y=0.085
+ $X2=4.112 $Y2=0
r194 36 38 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=4.112 $Y=0.085
+ $X2=4.112 $Y2=0.445
r195 32 72 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=3.152 $Y=0.085
+ $X2=3.152 $Y2=0
r196 32 34 15.6558 $w=2.63e-07 $l=3.6e-07 $layer=LI1_cond $X=3.152 $Y=0.085
+ $X2=3.152 $Y2=0.445
r197 28 115 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r198 28 30 15.3659 $w=2.68e-07 $l=3.6e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.445
r199 9 68 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=9.87
+ $Y=0.235 $X2=10.06 $Y2=0.445
r200 8 64 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=8.91
+ $Y=0.235 $X2=9.1 $Y2=0.445
r201 7 58 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=7.95
+ $Y=0.235 $X2=8.14 $Y2=0.445
r202 6 52 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=6.99
+ $Y=0.235 $X2=7.18 $Y2=0.445
r203 5 46 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=6.03
+ $Y=0.235 $X2=6.22 $Y2=0.445
r204 4 42 182 $w=1.7e-07 $l=3.02283e-07 $layer=licon1_NDIFF $count=1 $X=4.88
+ $Y=0.235 $X2=5.095 $Y2=0.445
r205 3 38 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.92
+ $Y=0.235 $X2=4.11 $Y2=0.445
r206 2 34 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.96
+ $Y=0.235 $X2=3.15 $Y2=0.445
r207 1 30 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.235 $X2=2.19 $Y2=0.445
.ends

