* NGSPICE file created from sky130_fd_sc_hdll__sdlclkp_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__sdlclkp_2 CLK GATE SCE VGND VNB VPB VPWR GCLK
M1000 a_484_315# a_299_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.6654e+12p ps=1.474e+07u
M1001 a_269_21# CLK VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1002 a_27_47# GATE a_117_369# VPB phighvt w=640000u l=180000u
+  ad=2.021e+11p pd=1.97e+06u as=1.472e+11p ps=1.74e+06u
M1003 VPWR a_1093_47# GCLK VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1004 a_1185_47# a_484_315# a_1093_47# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.302e+11p ps=1.46e+06u
M1005 VGND CLK a_1185_47# VNB nshort w=420000u l=150000u
+  ad=9.4605e+11p pd=9.05e+06u as=0p ps=0u
M1006 a_484_315# a_299_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1007 a_117_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_415_47# a_266_243# a_299_47# VNB nshort w=360000u l=150000u
+  ad=1.977e+11p pd=1.85e+06u as=1.548e+11p ps=1.58e+06u
M1009 a_410_413# a_269_21# a_299_47# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=1.47e+11p ps=1.54e+06u
M1010 VPWR a_484_315# a_410_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 GCLK a_1093_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_1093_47# GCLK VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.08e+11p ps=1.94e+06u
M1013 VPWR CLK a_1093_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.856e+11p ps=1.86e+06u
M1014 GCLK a_1093_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND a_484_315# a_415_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_269_21# CLK VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1017 VGND a_269_21# a_266_243# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1018 a_299_47# a_269_21# a_27_47# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=2.622e+11p ps=2.95e+06u
M1019 a_1093_47# a_484_315# VPWR VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VGND SCE a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_299_47# a_266_243# a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VPWR a_269_21# a_266_243# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1023 a_27_47# GATE VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

