* File: sky130_fd_sc_hdll__decap_4.pex.spice
* Created: Wed Sep  2 08:27:39 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DECAP_4%VGND 1 7 10 13 24 27
r9 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r10 24 26 0.338889 $w=1.08e-06 $l=3e-08 $layer=LI1_cond $X=1.58 $Y=0.645
+ $X2=1.61 $Y2=0.645
r11 22 27 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r12 21 24 10.0537 $w=1.08e-06 $l=8.9e-07 $layer=LI1_cond $X=0.69 $Y=0.645
+ $X2=1.58 $Y2=0.645
r13 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r14 15 18 0.338889 $w=1.08e-06 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.645
+ $X2=0.26 $Y2=0.645
r15 11 21 4.74444 $w=1.08e-06 $l=4.2e-07 $layer=LI1_cond $X=0.27 $Y=0.645
+ $X2=0.69 $Y2=0.645
r16 11 18 0.112963 $w=1.08e-06 $l=1e-08 $layer=LI1_cond $X=0.27 $Y=0.645
+ $X2=0.26 $Y2=0.645
r17 10 13 41.1323 $w=9.62e-07 $l=7.6e-07 $layer=POLY_cond $X=0.775 $Y=1.29
+ $X2=0.775 $Y2=2.05
r18 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.29 $X2=0.27 $Y2=1.29
r19 7 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r20 7 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r21 1 24 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=1.58 $Y2=0.51
r22 1 18 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.445
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DECAP_4%VPWR 1 7 10 19 22
r9 19 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r10 16 19 7.66267 $w=1.417e-06 $l=8.9e-07 $layer=LI1_cond $X=0.92 $Y=1.83
+ $X2=0.92 $Y2=2.72
r11 13 16 6.19901 $w=1.417e-06 $l=9.93177e-07 $layer=LI1_cond $X=1.57 $Y=1.11
+ $X2=0.92 $Y2=1.83
r12 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.11 $X2=1.57 $Y2=1.11
r13 10 12 38.6501 $w=8.18e-07 $l=8.33966e-07 $layer=POLY_cond $X=0.92 $Y=0.69
+ $X2=1.57 $Y2=1.11
r14 7 22 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r15 7 19 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r16 1 16 300 $w=1.7e-07 $l=2.74317e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.615 $X2=1.58 $Y2=1.83
r17 1 16 300 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_PDIFF $count=2 $X=1.445
+ $Y=1.615 $X2=0.26 $Y2=1.83
.ends

