* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkmux2_4 A0 A1 S VGND VNB VPB VPWR X
X0 VPWR S a_523_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X1 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 a_523_309# A0 a_79_199# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X3 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X4 a_79_199# A0 a_754_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_79_199# A1 a_875_309# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X7 a_754_47# a_925_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR a_79_199# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 X a_79_199# VGND VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X11 VGND S a_525_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_875_309# a_925_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X13 VGND a_79_199# X VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X14 X a_79_199# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VPWR S a_925_21# VPB sky130_fd_pr__pfet_01v8_hvt w=940000u l=180000u
X16 a_525_47# A1 a_79_199# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 VGND S a_925_21# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
.ends
