* File: sky130_fd_sc_hdll__clkbuf_8.pxi.spice
* Created: Thu Aug 27 19:02:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_8%A N_A_c_87_n N_A_M1004_g N_A_M1001_g N_A_c_88_n
+ N_A_M1013_g N_A_M1002_g A A N_A_c_86_n PM_SKY130_FD_SC_HDLL__CLKBUF_8%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_8%A_118_297# N_A_118_297#_M1001_d
+ N_A_118_297#_M1004_d N_A_118_297#_M1000_g N_A_118_297#_c_133_n
+ N_A_118_297#_M1003_g N_A_118_297#_M1007_g N_A_118_297#_c_134_n
+ N_A_118_297#_M1005_g N_A_118_297#_M1008_g N_A_118_297#_c_135_n
+ N_A_118_297#_M1006_g N_A_118_297#_M1009_g N_A_118_297#_c_136_n
+ N_A_118_297#_M1010_g N_A_118_297#_M1012_g N_A_118_297#_c_137_n
+ N_A_118_297#_M1011_g N_A_118_297#_M1014_g N_A_118_297#_c_138_n
+ N_A_118_297#_M1015_g N_A_118_297#_M1016_g N_A_118_297#_c_139_n
+ N_A_118_297#_M1017_g N_A_118_297#_c_140_n N_A_118_297#_M1019_g
+ N_A_118_297#_M1018_g N_A_118_297#_c_130_n N_A_118_297#_c_141_n
+ N_A_118_297#_c_131_n N_A_118_297#_c_154_n N_A_118_297#_c_132_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_8%A_118_297#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_8%VPWR N_VPWR_M1004_s N_VPWR_M1013_s
+ N_VPWR_M1005_d N_VPWR_M1010_d N_VPWR_M1015_d N_VPWR_M1019_d N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_272_n N_VPWR_c_273_n
+ N_VPWR_c_274_n N_VPWR_c_275_n N_VPWR_c_276_n N_VPWR_c_277_n N_VPWR_c_278_n
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n VPWR
+ N_VPWR_c_283_n N_VPWR_c_267_n N_VPWR_c_285_n N_VPWR_c_286_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_8%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_8%X N_X_M1000_s N_X_M1008_s N_X_M1012_s
+ N_X_M1016_s N_X_M1003_s N_X_M1006_s N_X_M1011_s N_X_M1017_s N_X_c_346_n
+ N_X_c_347_n N_X_c_348_n N_X_c_368_n N_X_c_349_n N_X_c_350_n N_X_c_378_n
+ N_X_c_351_n N_X_c_352_n N_X_c_387_n N_X_c_353_n N_X_c_392_n N_X_c_354_n
+ N_X_c_396_n N_X_c_355_n N_X_c_400_n X X X PM_SKY130_FD_SC_HDLL__CLKBUF_8%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_8%VGND N_VGND_M1001_s N_VGND_M1002_s
+ N_VGND_M1007_d N_VGND_M1009_d N_VGND_M1014_d N_VGND_M1018_d N_VGND_c_461_n
+ N_VGND_c_462_n N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n N_VGND_c_466_n
+ N_VGND_c_467_n N_VGND_c_468_n N_VGND_c_469_n N_VGND_c_470_n N_VGND_c_471_n
+ N_VGND_c_472_n N_VGND_c_473_n N_VGND_c_474_n N_VGND_c_475_n VGND
+ N_VGND_c_476_n N_VGND_c_477_n N_VGND_c_478_n N_VGND_c_479_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_8%VGND
cc_1 VNB N_A_M1001_g 0.0288268f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.445
cc_2 VNB N_A_M1002_g 0.0241662f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=0.445
cc_3 VNB A 0.0261816f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_4 VNB N_A_c_86_n 0.0755189f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.155
cc_5 VNB N_A_118_297#_M1000_g 0.0268891f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.985
cc_6 VNB N_A_118_297#_M1007_g 0.0258077f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_A_118_297#_M1008_g 0.0258075f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.155
cc_8 VNB N_A_118_297#_M1009_g 0.0258077f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_118_297#_M1012_g 0.0258075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_118_297#_M1014_g 0.0257771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_118_297#_M1016_g 0.0261623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_118_297#_M1018_g 0.0336194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_118_297#_c_130_n 0.00465316f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_118_297#_c_131_n 0.00442652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_118_297#_c_132_n 0.176502f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VPWR_c_267_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_X_c_346_n 0.0017582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_347_n 0.00733625f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.16
cc_19 VNB N_X_c_348_n 0.00426583f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_349_n 0.00149815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_350_n 0.00733625f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_351_n 0.00149815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_352_n 0.0048892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_353_n 0.0015723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_354_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_355_n 0.0018976f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB X 0.0317353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_461_n 0.0112866f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.155
cc_29 VNB N_VGND_c_462_n 0.005166f $X=-0.19 $Y=-0.24 $X2=0.27 $Y2=1.16
cc_30 VNB N_VGND_c_463_n 0.0198934f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.155
cc_31 VNB N_VGND_c_464_n 0.00522139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_465_n 0.0190904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_466_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_467_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_468_n 0.00523594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_469_n 0.018338f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_470_n 0.0182806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_471_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_472_n 0.0182806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_473_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_474_n 0.0182774f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_475_n 0.00574315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_476_n 0.0113717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_477_n 0.283434f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_478_n 0.00497572f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_479_n 0.00497395f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VPB N_A_c_87_n 0.0211429f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_48 VPB N_A_c_88_n 0.0165782f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_49 VPB A 0.00123221f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_50 VPB N_A_c_86_n 0.0301893f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.155
cc_51 VPB N_A_118_297#_c_133_n 0.0166021f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=0.9
cc_52 VPB N_A_118_297#_c_134_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_118_297#_c_135_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.155
cc_54 VPB N_A_118_297#_c_136_n 0.0164285f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_118_297#_c_137_n 0.0164277f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_118_297#_c_138_n 0.0164107f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_118_297#_c_139_n 0.0157624f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_118_297#_c_140_n 0.0193677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_118_297#_c_141_n 0.00140153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_118_297#_c_131_n 0.00331269f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_118_297#_c_132_n 0.102242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_268_n 0.0108797f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.155
cc_63 VPB N_VPWR_c_269_n 0.0422667f $X=-0.19 $Y=1.305 $X2=0.27 $Y2=1.16
cc_64 VPB N_VPWR_c_270_n 0.0199013f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.155
cc_65 VPB N_VPWR_c_271_n 0.00522213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_272_n 0.0198082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_273_n 0.00522213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_274_n 0.00522213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_275_n 0.00522213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_276_n 0.0278366f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_277_n 0.0198082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_278_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_279_n 0.0198082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_280_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_281_n 0.0198082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_282_n 0.00564836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_283_n 0.0114539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_267_n 0.0516179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_285_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_286_n 0.00497514f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB X 0.0104376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB X 0.0107432f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_A_118_297#_M1000_g 0.0220403f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_84 N_A_c_88_n N_A_118_297#_c_133_n 0.0166985f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_M1001_g N_A_118_297#_c_130_n 0.00343385f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_M1002_g N_A_118_297#_c_130_n 0.00875058f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_87 A N_A_118_297#_c_130_n 0.0229331f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_c_86_n N_A_118_297#_c_130_n 0.0133594f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_89 N_A_c_87_n N_A_118_297#_c_141_n 0.00295477f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_88_n N_A_118_297#_c_141_n 0.00300089f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_86_n N_A_118_297#_c_141_n 0.0100729f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_92 N_A_c_86_n N_A_118_297#_c_131_n 0.027109f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_93 A N_A_118_297#_c_154_n 0.0161665f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_94 N_A_c_86_n N_A_118_297#_c_154_n 0.0100412f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_95 N_A_c_86_n N_A_118_297#_c_132_n 0.0220403f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_96 N_A_c_87_n N_VPWR_c_269_n 0.00918636f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_97 A N_VPWR_c_269_n 0.0210616f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A_c_86_n N_VPWR_c_269_n 0.00771804f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_99 N_A_c_87_n N_VPWR_c_270_n 0.00702461f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_88_n N_VPWR_c_270_n 0.00702461f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_88_n N_VPWR_c_271_n 0.00408512f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_87_n N_VPWR_c_267_n 0.0135424f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_88_n N_VPWR_c_267_n 0.0126419f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_104 A N_VGND_c_461_n 0.00101698f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_M1001_g N_VGND_c_462_n 0.00609576f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_106 A N_VGND_c_462_n 0.0211866f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_107 N_A_c_86_n N_VGND_c_462_n 0.00122559f $X=1.005 $Y=1.155 $X2=0 $Y2=0
cc_108 N_A_M1001_g N_VGND_c_463_n 0.00585385f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_M1002_g N_VGND_c_463_n 0.00585385f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_110 N_A_M1002_g N_VGND_c_464_n 0.00311641f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_M1001_g N_VGND_c_477_n 0.0117978f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_112 N_A_M1002_g N_VGND_c_477_n 0.0107987f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_113 A N_VGND_c_477_n 0.00306056f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_114 N_A_118_297#_c_141_n N_VPWR_c_270_n 0.0148098f $X=0.74 $Y=1.69 $X2=0
+ $Y2=0
cc_115 N_A_118_297#_c_133_n N_VPWR_c_271_n 0.00408512f $X=1.46 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_A_118_297#_c_131_n N_VPWR_c_271_n 0.0166171f $X=3.595 $Y=1.16 $X2=0
+ $Y2=0
cc_117 N_A_118_297#_c_133_n N_VPWR_c_272_n 0.00702461f $X=1.46 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_118_297#_c_134_n N_VPWR_c_272_n 0.00702461f $X=1.94 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_118_297#_c_134_n N_VPWR_c_273_n 0.00398486f $X=1.94 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_118_297#_c_135_n N_VPWR_c_273_n 0.00398486f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_121 N_A_118_297#_c_136_n N_VPWR_c_274_n 0.00398486f $X=2.9 $Y=1.41 $X2=0
+ $Y2=0
cc_122 N_A_118_297#_c_137_n N_VPWR_c_274_n 0.00398486f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A_118_297#_c_138_n N_VPWR_c_275_n 0.00398486f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_118_297#_c_139_n N_VPWR_c_275_n 0.00398486f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_125 N_A_118_297#_c_132_n N_VPWR_c_275_n 4.17622e-19 $X=4.82 $Y=1.18 $X2=0
+ $Y2=0
cc_126 N_A_118_297#_c_140_n N_VPWR_c_276_n 0.00877126f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_127 N_A_118_297#_c_135_n N_VPWR_c_277_n 0.00702461f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_118_297#_c_136_n N_VPWR_c_277_n 0.00702461f $X=2.9 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_118_297#_c_137_n N_VPWR_c_279_n 0.00702461f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_118_297#_c_138_n N_VPWR_c_279_n 0.00702461f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_118_297#_c_139_n N_VPWR_c_281_n 0.00702461f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_132 N_A_118_297#_c_140_n N_VPWR_c_281_n 0.00702461f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A_118_297#_M1004_d N_VPWR_c_267_n 0.00421554f $X=0.59 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_A_118_297#_c_133_n N_VPWR_c_267_n 0.0126419f $X=1.46 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_118_297#_c_134_n N_VPWR_c_267_n 0.0126174f $X=1.94 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_118_297#_c_135_n N_VPWR_c_267_n 0.0126174f $X=2.42 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_118_297#_c_136_n N_VPWR_c_267_n 0.0126174f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_118_297#_c_137_n N_VPWR_c_267_n 0.0126174f $X=3.38 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_118_297#_c_138_n N_VPWR_c_267_n 0.0126174f $X=3.86 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_118_297#_c_139_n N_VPWR_c_267_n 0.0126174f $X=4.34 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_118_297#_c_140_n N_VPWR_c_267_n 0.0136856f $X=4.82 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_118_297#_c_141_n N_VPWR_c_267_n 0.00952853f $X=0.74 $Y=1.69 $X2=0
+ $Y2=0
cc_143 N_A_118_297#_M1000_g N_X_c_346_n 0.00439403f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_A_118_297#_M1007_g N_X_c_346_n 0.00228345f $X=1.915 $Y=0.445 $X2=0
+ $Y2=0
cc_145 N_A_118_297#_M1007_g N_X_c_347_n 0.0124132f $X=1.915 $Y=0.445 $X2=0 $Y2=0
cc_146 N_A_118_297#_M1008_g N_X_c_347_n 0.0128559f $X=2.395 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_118_297#_c_131_n N_X_c_347_n 0.0503195f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A_118_297#_c_132_n N_X_c_347_n 0.00400618f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_149 N_A_118_297#_M1000_g N_X_c_348_n 0.00545572f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_A_118_297#_c_131_n N_X_c_348_n 0.021367f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_118_297#_c_132_n N_X_c_348_n 0.00415703f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_152 N_A_118_297#_c_134_n N_X_c_368_n 0.017751f $X=1.94 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_118_297#_c_135_n N_X_c_368_n 0.017751f $X=2.42 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_118_297#_c_131_n N_X_c_368_n 0.0450774f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_118_297#_c_132_n N_X_c_368_n 0.00670724f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_156 N_A_118_297#_M1008_g N_X_c_349_n 0.00519179f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_157 N_A_118_297#_M1009_g N_X_c_349_n 0.00228345f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_158 N_A_118_297#_M1009_g N_X_c_350_n 0.0128559f $X=2.875 $Y=0.445 $X2=0 $Y2=0
cc_159 N_A_118_297#_M1012_g N_X_c_350_n 0.0128559f $X=3.355 $Y=0.445 $X2=0 $Y2=0
cc_160 N_A_118_297#_c_131_n N_X_c_350_n 0.0503195f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_118_297#_c_132_n N_X_c_350_n 0.00400618f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_162 N_A_118_297#_c_136_n N_X_c_378_n 0.017751f $X=2.9 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_118_297#_c_137_n N_X_c_378_n 0.017751f $X=3.38 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_118_297#_c_131_n N_X_c_378_n 0.0450774f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_118_297#_c_132_n N_X_c_378_n 0.00670724f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_166 N_A_118_297#_M1012_g N_X_c_351_n 0.00519179f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_167 N_A_118_297#_M1014_g N_X_c_351_n 0.00228345f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_168 N_A_118_297#_M1014_g N_X_c_352_n 0.0128559f $X=3.835 $Y=0.445 $X2=0 $Y2=0
cc_169 N_A_118_297#_c_131_n N_X_c_352_n 0.0170647f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_170 N_A_118_297#_c_132_n N_X_c_352_n 0.00480754f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_171 N_A_118_297#_c_138_n N_X_c_387_n 0.017751f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_118_297#_c_131_n N_X_c_387_n 0.0150268f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_173 N_A_118_297#_c_132_n N_X_c_387_n 0.00539432f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_174 N_A_118_297#_M1016_g N_X_c_353_n 0.00525012f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_175 N_A_118_297#_M1018_g N_X_c_353_n 0.00525012f $X=4.845 $Y=0.445 $X2=0
+ $Y2=0
cc_176 N_A_118_297#_c_131_n N_X_c_392_n 0.0177415f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_177 N_A_118_297#_c_132_n N_X_c_392_n 0.00635512f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_178 N_A_118_297#_c_131_n N_X_c_354_n 0.021367f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_118_297#_c_132_n N_X_c_354_n 0.00415703f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_180 N_A_118_297#_c_131_n N_X_c_396_n 0.0177415f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_118_297#_c_132_n N_X_c_396_n 0.00635512f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_182 N_A_118_297#_c_131_n N_X_c_355_n 0.021367f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_183 N_A_118_297#_c_132_n N_X_c_355_n 0.00415703f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_184 N_A_118_297#_c_131_n N_X_c_400_n 0.0177415f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_118_297#_c_132_n N_X_c_400_n 0.00635512f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_186 N_A_118_297#_M1014_g X 0.00112182f $X=3.835 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_118_297#_c_138_n X 0.0022323f $X=3.86 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_118_297#_M1016_g X 0.0126798f $X=4.315 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_118_297#_c_139_n X 0.00297541f $X=4.34 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_118_297#_c_140_n X 0.00412953f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_118_297#_M1018_g X 0.0143761f $X=4.845 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_118_297#_c_131_n X 0.0208936f $X=3.595 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_118_297#_c_132_n X 0.068352f $X=4.82 $Y=1.18 $X2=0 $Y2=0
cc_194 N_A_118_297#_c_139_n X 0.0163761f $X=4.34 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_118_297#_c_140_n X 0.018241f $X=4.82 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_118_297#_c_130_n N_VGND_c_463_n 0.0152148f $X=0.74 $Y=0.445 $X2=0
+ $Y2=0
cc_197 N_A_118_297#_M1000_g N_VGND_c_464_n 0.00311641f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_198 N_A_118_297#_c_131_n N_VGND_c_464_n 0.00869033f $X=3.595 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_118_297#_M1000_g N_VGND_c_465_n 0.00585385f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_200 N_A_118_297#_M1007_g N_VGND_c_465_n 0.00439206f $X=1.915 $Y=0.445 $X2=0
+ $Y2=0
cc_201 N_A_118_297#_M1007_g N_VGND_c_466_n 0.00484691f $X=1.915 $Y=0.445 $X2=0
+ $Y2=0
cc_202 N_A_118_297#_M1008_g N_VGND_c_466_n 0.00313102f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_203 N_A_118_297#_M1009_g N_VGND_c_467_n 0.00484691f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_204 N_A_118_297#_M1012_g N_VGND_c_467_n 0.00313102f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_205 N_A_118_297#_M1014_g N_VGND_c_468_n 0.00484691f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_206 N_A_118_297#_M1016_g N_VGND_c_468_n 0.00313102f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_207 N_A_118_297#_M1018_g N_VGND_c_469_n 0.00488085f $X=4.845 $Y=0.445 $X2=0
+ $Y2=0
cc_208 N_A_118_297#_M1008_g N_VGND_c_470_n 0.00439206f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_209 N_A_118_297#_M1009_g N_VGND_c_470_n 0.00439206f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_210 N_A_118_297#_M1012_g N_VGND_c_472_n 0.00439206f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_211 N_A_118_297#_M1014_g N_VGND_c_472_n 0.00439206f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_212 N_A_118_297#_M1016_g N_VGND_c_474_n 0.00439071f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_213 N_A_118_297#_M1018_g N_VGND_c_474_n 0.00439071f $X=4.845 $Y=0.445 $X2=0
+ $Y2=0
cc_214 N_A_118_297#_M1001_d N_VGND_c_477_n 0.00549964f $X=0.6 $Y=0.235 $X2=0
+ $Y2=0
cc_215 N_A_118_297#_M1000_g N_VGND_c_477_n 0.0107987f $X=1.435 $Y=0.445 $X2=0
+ $Y2=0
cc_216 N_A_118_297#_M1007_g N_VGND_c_477_n 0.00628867f $X=1.915 $Y=0.445 $X2=0
+ $Y2=0
cc_217 N_A_118_297#_M1008_g N_VGND_c_477_n 0.00616322f $X=2.395 $Y=0.445 $X2=0
+ $Y2=0
cc_218 N_A_118_297#_M1009_g N_VGND_c_477_n 0.00628867f $X=2.875 $Y=0.445 $X2=0
+ $Y2=0
cc_219 N_A_118_297#_M1012_g N_VGND_c_477_n 0.00616322f $X=3.355 $Y=0.445 $X2=0
+ $Y2=0
cc_220 N_A_118_297#_M1014_g N_VGND_c_477_n 0.00628867f $X=3.835 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_118_297#_M1016_g N_VGND_c_477_n 0.00627824f $X=4.315 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_118_297#_M1018_g N_VGND_c_477_n 0.00722843f $X=4.845 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_118_297#_c_130_n N_VGND_c_477_n 0.00950576f $X=0.74 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_VPWR_c_267_n N_X_M1003_s 0.00386843f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_267_n N_X_M1006_s 0.00386843f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_267_n N_X_M1011_s 0.00386843f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_c_267_n N_X_M1017_s 0.00386843f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_228 N_VPWR_M1005_d N_X_c_368_n 0.00357164f $X=2.03 $Y=1.485 $X2=0 $Y2=0
cc_229 N_VPWR_c_273_n N_X_c_368_n 0.0154924f $X=2.18 $Y=2.22 $X2=0 $Y2=0
cc_230 N_VPWR_M1010_d N_X_c_378_n 0.00357164f $X=2.99 $Y=1.485 $X2=0 $Y2=0
cc_231 N_VPWR_c_274_n N_X_c_378_n 0.0154924f $X=3.14 $Y=2.22 $X2=0 $Y2=0
cc_232 N_VPWR_M1015_d N_X_c_387_n 0.00363829f $X=3.95 $Y=1.485 $X2=0 $Y2=0
cc_233 N_VPWR_c_275_n N_X_c_387_n 0.0127053f $X=4.1 $Y=2.22 $X2=0 $Y2=0
cc_234 N_VPWR_c_272_n N_X_c_392_n 0.0151544f $X=2.05 $Y=2.72 $X2=0 $Y2=0
cc_235 N_VPWR_c_267_n N_X_c_392_n 0.00991274f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_236 N_VPWR_c_277_n N_X_c_396_n 0.0151544f $X=3.01 $Y=2.72 $X2=0 $Y2=0
cc_237 N_VPWR_c_267_n N_X_c_396_n 0.00991274f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_238 N_VPWR_c_279_n N_X_c_400_n 0.0151544f $X=3.97 $Y=2.72 $X2=0 $Y2=0
cc_239 N_VPWR_c_267_n N_X_c_400_n 0.00991274f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_240 N_VPWR_M1015_d X 3.5412e-19 $X=3.95 $Y=1.485 $X2=0 $Y2=0
cc_241 N_VPWR_M1019_d X 0.00362185f $X=4.91 $Y=1.485 $X2=0 $Y2=0
cc_242 N_VPWR_c_275_n X 0.00293026f $X=4.1 $Y=2.22 $X2=0 $Y2=0
cc_243 N_VPWR_c_276_n X 0.0233095f $X=5.06 $Y=2.22 $X2=0 $Y2=0
cc_244 N_VPWR_c_281_n X 0.0151544f $X=4.93 $Y=2.72 $X2=0 $Y2=0
cc_245 N_VPWR_c_267_n X 0.00991274f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_246 N_X_c_346_n N_VGND_c_465_n 0.0141875f $X=1.7 $Y=0.445 $X2=0 $Y2=0
cc_247 N_X_c_347_n N_VGND_c_465_n 0.00299761f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_248 N_X_c_347_n N_VGND_c_466_n 0.0185136f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_249 N_X_c_350_n N_VGND_c_467_n 0.0185136f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_250 N_X_c_352_n N_VGND_c_468_n 0.0150295f $X=4.16 $Y=0.82 $X2=0 $Y2=0
cc_251 X N_VGND_c_468_n 0.00403581f $X=4.28 $Y=0.765 $X2=0 $Y2=0
cc_252 X N_VGND_c_469_n 0.0243348f $X=4.28 $Y=0.765 $X2=0 $Y2=0
cc_253 N_X_c_347_n N_VGND_c_470_n 0.00299761f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_254 N_X_c_349_n N_VGND_c_470_n 0.0141875f $X=2.66 $Y=0.445 $X2=0 $Y2=0
cc_255 N_X_c_350_n N_VGND_c_470_n 0.00299761f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_256 N_X_c_350_n N_VGND_c_472_n 0.00299761f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_257 N_X_c_351_n N_VGND_c_472_n 0.0141875f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_258 N_X_c_352_n N_VGND_c_472_n 0.00299761f $X=4.16 $Y=0.82 $X2=0 $Y2=0
cc_259 N_X_c_353_n N_VGND_c_474_n 0.0156284f $X=4.58 $Y=0.445 $X2=0 $Y2=0
cc_260 X N_VGND_c_474_n 0.00665978f $X=4.28 $Y=0.765 $X2=0 $Y2=0
cc_261 N_X_M1000_s N_VGND_c_477_n 0.00482172f $X=1.51 $Y=0.235 $X2=0 $Y2=0
cc_262 N_X_M1008_s N_VGND_c_477_n 0.00300326f $X=2.47 $Y=0.235 $X2=0 $Y2=0
cc_263 N_X_M1012_s N_VGND_c_477_n 0.00300326f $X=3.43 $Y=0.235 $X2=0 $Y2=0
cc_264 N_X_M1016_s N_VGND_c_477_n 0.00365899f $X=4.39 $Y=0.235 $X2=0 $Y2=0
cc_265 N_X_c_346_n N_VGND_c_477_n 0.00979224f $X=1.7 $Y=0.445 $X2=0 $Y2=0
cc_266 N_X_c_347_n N_VGND_c_477_n 0.0109571f $X=2.53 $Y=0.82 $X2=0 $Y2=0
cc_267 N_X_c_349_n N_VGND_c_477_n 0.00979224f $X=2.66 $Y=0.445 $X2=0 $Y2=0
cc_268 N_X_c_350_n N_VGND_c_477_n 0.0109571f $X=3.49 $Y=0.82 $X2=0 $Y2=0
cc_269 N_X_c_351_n N_VGND_c_477_n 0.00979224f $X=3.62 $Y=0.445 $X2=0 $Y2=0
cc_270 N_X_c_352_n N_VGND_c_477_n 0.00572224f $X=4.16 $Y=0.82 $X2=0 $Y2=0
cc_271 N_X_c_353_n N_VGND_c_477_n 0.00981584f $X=4.58 $Y=0.445 $X2=0 $Y2=0
cc_272 X N_VGND_c_477_n 0.0122417f $X=4.28 $Y=0.765 $X2=0 $Y2=0
