* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_326_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.65e+11p pd=5.13e+06u as=6.834e+11p ps=6.52e+06u
M1001 a_412_47# A1 a_235_297# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=1.755e+11p ps=1.84e+06u
M1002 VPWR B1_N a_27_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.134e+11p ps=1.38e+06u
M1003 a_235_297# a_27_413# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=9.0705e+11p ps=5.49e+06u
M1004 VGND B1_N a_27_413# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.323e+11p ps=1.47e+06u
M1005 X a_235_297# VGND VNB nshort w=650000u l=150000u
+  ad=2.4375e+11p pd=2.05e+06u as=0p ps=0u
M1006 VGND A2 a_412_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR A1 a_326_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_326_297# a_27_413# a_235_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.75e+11p ps=2.55e+06u
M1009 X a_235_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.85e+11p pd=2.77e+06u as=0p ps=0u
.ends
