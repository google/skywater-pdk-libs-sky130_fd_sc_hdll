* File: sky130_fd_sc_hdll__o22ai_2.pex.spice
* Created: Wed Sep  2 08:45:44 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%B1 1 3 4 6 7 9 10 12 13 19 20 23
r38 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 18 20 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=0.95 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.95
+ $Y=1.16 $X2=0.95 $Y2=1.16
r41 16 18 55.1763 $w=3.8e-07 $l=4.35e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.95 $Y2=1.202
r42 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r43 13 19 10.8268 $w=2.08e-07 $l=2.05e-07 $layer=LI1_cond $X=0.745 $Y=1.18
+ $X2=0.95 $Y2=1.18
r44 13 23 2.64069 $w=2.08e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.18
+ $X2=0.695 $Y2=1.18
r45 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r46 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r47 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r48 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r49 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r51 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%B2 1 3 4 6 7 9 10 12 13 19 20 23
r41 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r42 18 20 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=1.88 $Y=1.202
+ $X2=1.925 $Y2=1.202
r43 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r44 16 18 53.9079 $w=3.8e-07 $l=4.25e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.88 $Y2=1.202
r45 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r46 13 19 6.37727 $w=1.98e-07 $l=1.15e-07 $layer=LI1_cond $X=1.765 $Y=1.175
+ $X2=1.88 $Y2=1.175
r47 13 23 8.31818 $w=1.98e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.175
+ $X2=1.615 $Y2=1.175
r48 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r49 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r50 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r51 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r52 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r53 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r54 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r55 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%A2 1 3 4 6 7 9 10 12 13 19 20 23
r51 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.425 $Y=1.202
+ $X2=3.45 $Y2=1.202
r52 18 20 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=3.39 $Y=1.202
+ $X2=3.425 $Y2=1.202
r53 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.39
+ $Y=1.16 $X2=3.39 $Y2=1.16
r54 16 18 55.1763 $w=3.8e-07 $l=4.35e-07 $layer=POLY_cond $X=2.955 $Y=1.202
+ $X2=3.39 $Y2=1.202
r55 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.93 $Y=1.202
+ $X2=2.955 $Y2=1.202
r56 13 19 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=3.265 $Y=1.175
+ $X2=3.39 $Y2=1.175
r57 13 23 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=3.265 $Y=1.175
+ $X2=3.015 $Y2=1.175
r58 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=1.202
r59 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.45 $Y2=0.56
r60 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.202
r61 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.425 $Y=1.41
+ $X2=3.425 $Y2=1.985
r62 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.202
r63 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.955 $Y=1.41
+ $X2=2.955 $Y2=1.985
r64 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.93 $Y=0.995
+ $X2=2.93 $Y2=1.202
r65 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.93 $Y=0.995 $X2=2.93
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%A1 1 3 4 6 7 9 10 12 13 20 23
r41 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.365 $Y=1.202
+ $X2=4.39 $Y2=1.202
r42 18 20 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=4.32 $Y=1.202
+ $X2=4.365 $Y2=1.202
r43 16 18 53.9079 $w=3.8e-07 $l=4.25e-07 $layer=POLY_cond $X=3.895 $Y=1.202
+ $X2=4.32 $Y2=1.202
r44 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.87 $Y=1.202
+ $X2=3.895 $Y2=1.202
r45 13 23 18.4848 $w=2.08e-07 $l=3.5e-07 $layer=LI1_cond $X=4.285 $Y=1.18
+ $X2=3.935 $Y2=1.18
r46 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.32
+ $Y=1.16 $X2=4.32 $Y2=1.16
r47 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.39 $Y=0.995
+ $X2=4.39 $Y2=1.202
r48 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.39 $Y=0.995
+ $X2=4.39 $Y2=0.56
r49 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.202
r50 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.365 $Y=1.41
+ $X2=4.365 $Y2=1.985
r51 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.202
r52 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.895 $Y=1.41
+ $X2=3.895 $Y2=1.985
r53 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.87 $Y=0.995
+ $X2=3.87 $Y2=1.202
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.87 $Y=0.995 $X2=3.87
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_297# 1 2 3 10 12 14 16 17 18 22
r34 20 22 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.16 $Y=2.295
+ $X2=2.16 $Y2=1.96
r35 19 29 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.38
+ $X2=1.22 $Y2=2.38
r36 18 20 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=2.16 $Y2=2.295
r37 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=2.38
+ $X2=1.345 $Y2=2.38
r38 17 29 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.295
+ $X2=1.22 $Y2=2.38
r39 16 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r40 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.295
r41 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r42 14 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r43 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r44 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r45 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r46 3 22 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.96
r47 2 29 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r48 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r49 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r50 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%VPWR 1 2 11 15 18 19 20 30 31 34
r54 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r55 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r56 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r57 27 28 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 25 28 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r59 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r60 24 27 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 24 25 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r62 22 34 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r63 22 24 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 18 27 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=3.91 $Y2=2.72
r66 18 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.005 $Y=2.72
+ $X2=4.13 $Y2=2.72
r67 17 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.83 $Y2=2.72
r68 17 19 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.255 $Y=2.72
+ $X2=4.13 $Y2=2.72
r69 13 19 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=2.635
+ $X2=4.13 $Y2=2.72
r70 13 15 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=4.13 $Y=2.635
+ $X2=4.13 $Y2=1.96
r71 9 34 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r72 9 11 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=1.96
r73 2 15 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.985
+ $Y=1.485 $X2=4.13 $Y2=1.96
r74 1 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%Y 1 2 3 4 13 22 23 29 30 31 33 34
r64 30 34 8.0101 $w=1.78e-07 $l=1.3e-07 $layer=LI1_cond $X=2.405 $Y=1.535
+ $X2=2.275 $Y2=1.535
r65 30 31 6.51676 $w=1.8e-07 $l=1.2e-07 $layer=LI1_cond $X=2.405 $Y=1.535
+ $X2=2.525 $Y2=1.535
r66 27 34 28.3434 $w=1.78e-07 $l=4.6e-07 $layer=LI1_cond $X=1.815 $Y=1.535
+ $X2=2.275 $Y2=1.535
r67 27 29 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=1.815 $Y=1.535
+ $X2=1.69 $Y2=1.535
r68 24 31 6.51676 $w=1.8e-07 $l=1.2e-07 $layer=LI1_cond $X=2.645 $Y=1.535
+ $X2=2.525 $Y2=1.535
r69 23 33 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.065 $Y=1.535
+ $X2=3.19 $Y2=1.535
r70 23 24 25.8788 $w=1.78e-07 $l=4.2e-07 $layer=LI1_cond $X=3.065 $Y=1.535
+ $X2=2.645 $Y2=1.535
r71 22 31 0.330231 $w=2.4e-07 $l=9e-08 $layer=LI1_cond $X=2.525 $Y=1.445
+ $X2=2.525 $Y2=1.535
r72 21 22 25.93 $w=2.38e-07 $l=5.4e-07 $layer=LI1_cond $X=2.525 $Y=0.905
+ $X2=2.525 $Y2=1.445
r73 15 18 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=0.75 $Y=0.775
+ $X2=1.69 $Y2=0.775
r74 13 21 6.83069 $w=2.6e-07 $l=1.80278e-07 $layer=LI1_cond $X=2.405 $Y=0.775
+ $X2=2.525 $Y2=0.905
r75 13 18 31.6922 $w=2.58e-07 $l=7.15e-07 $layer=LI1_cond $X=2.405 $Y=0.775
+ $X2=1.69 $Y2=0.775
r76 4 33 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.045
+ $Y=1.485 $X2=3.19 $Y2=1.62
r77 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.62
r78 2 18 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.73
r79 1 15 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%A_515_297# 1 2 3 12 14 15 16 17 18 20 22
r38 20 29 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=4.602 $Y=1.625
+ $X2=4.602 $Y2=1.54
r39 20 22 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=4.602 $Y=1.625
+ $X2=4.602 $Y2=2.3
r40 19 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.785 $Y=1.54
+ $X2=3.66 $Y2=1.54
r41 18 29 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=4.475 $Y=1.54
+ $X2=4.602 $Y2=1.54
r42 18 19 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.475 $Y=1.54
+ $X2=3.785 $Y2=1.54
r43 17 27 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=2.295
+ $X2=3.66 $Y2=2.38
r44 16 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.66 $Y=1.625
+ $X2=3.66 $Y2=1.54
r45 16 17 30.8855 $w=2.48e-07 $l=6.7e-07 $layer=LI1_cond $X=3.66 $Y=1.625
+ $X2=3.66 $Y2=2.295
r46 14 27 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.535 $Y=2.38
+ $X2=3.66 $Y2=2.38
r47 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.535 $Y=2.38
+ $X2=2.845 $Y2=2.38
r48 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.72 $Y=2.295
+ $X2=2.845 $Y2=2.38
r49 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.72 $Y=2.295
+ $X2=2.72 $Y2=1.96
r50 3 29 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.485 $X2=4.6 $Y2=1.62
r51 3 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.455
+ $Y=1.485 $X2=4.6 $Y2=2.3
r52 2 27 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=2.3
r53 2 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.515
+ $Y=1.485 $X2=3.66 $Y2=1.62
r54 1 12 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.575
+ $Y=1.485 $X2=2.72 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%A_27_47# 1 2 3 4 5 16 18 20 27 28 29 32 34
+ 38 42
r75 36 38 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.575 $Y=0.725
+ $X2=4.575 $Y2=0.39
r76 35 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.825 $Y=0.815
+ $X2=3.66 $Y2=0.815
r77 34 36 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=4.385 $Y=0.815
+ $X2=4.575 $Y2=0.725
r78 34 35 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.385 $Y=0.815
+ $X2=3.825 $Y2=0.815
r79 30 42 0.718145 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=3.66 $Y=0.725 $X2=3.66
+ $Y2=0.815
r80 30 32 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.66 $Y=0.725
+ $X2=3.66 $Y2=0.39
r81 28 42 8.26956 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=3.495 $Y=0.815
+ $X2=3.66 $Y2=0.815
r82 28 29 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=3.495 $Y=0.815
+ $X2=2.985 $Y2=0.815
r83 27 29 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.9 $Y=0.725
+ $X2=2.985 $Y2=0.815
r84 26 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=2.9 $Y=0.475 $X2=2.9
+ $Y2=0.725
r85 23 25 97.5348 $w=1.68e-07 $l=1.495e-06 $layer=LI1_cond $X=1.22 $Y=0.39
+ $X2=2.715 $Y2=0.39
r86 21 41 4.53113 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=0.365 $Y=0.39
+ $X2=0.227 $Y2=0.39
r87 21 23 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.365 $Y=0.39
+ $X2=1.22 $Y2=0.39
r88 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.815 $Y=0.39
+ $X2=2.9 $Y2=0.475
r89 20 25 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.815 $Y=0.39
+ $X2=2.715 $Y2=0.39
r90 16 41 2.79091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.227 $Y=0.475
+ $X2=0.227 $Y2=0.39
r91 16 18 10.6863 $w=2.73e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=0.475
+ $X2=0.227 $Y2=0.73
r92 5 38 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=4.465
+ $Y=0.235 $X2=4.6 $Y2=0.39
r93 4 32 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=3.525
+ $Y=0.235 $X2=3.66 $Y2=0.39
r94 3 25 91 $w=1.7e-07 $l=7.63577e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.235 $X2=2.715 $Y2=0.39
r95 2 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r96 1 41 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
r97 1 18 182 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22AI_2%VGND 1 2 9 13 16 17 19 20 21 34 35
r57 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r58 32 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r59 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r60 29 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r61 28 29 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r62 24 28 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.99
+ $Y2=0
r63 21 29 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.99
+ $Y2=0
r64 21 24 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r65 19 31 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=4.045 $Y=0 $X2=3.91
+ $Y2=0
r66 19 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.045 $Y=0 $X2=4.13
+ $Y2=0
r67 18 34 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.83
+ $Y2=0
r68 18 20 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0 $X2=4.13
+ $Y2=0
r69 16 28 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=0 $X2=2.99
+ $Y2=0
r70 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=0 $X2=3.24
+ $Y2=0
r71 15 31 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.325 $Y=0 $X2=3.91
+ $Y2=0
r72 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=0 $X2=3.24
+ $Y2=0
r73 11 20 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0
r74 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.13 $Y=0.085
+ $X2=4.13 $Y2=0.39
r75 7 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=0.085 $X2=3.24
+ $Y2=0
r76 7 9 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.24 $Y=0.085
+ $X2=3.24 $Y2=0.39
r77 2 13 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.945
+ $Y=0.235 $X2=4.13 $Y2=0.39
r78 1 9 182 $w=1.7e-07 $l=3.02738e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.24 $Y2=0.39
.ends

