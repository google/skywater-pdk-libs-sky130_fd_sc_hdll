# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xnor2_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xnor2_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.075000 2.905000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.485000 1.075000 1.010000 1.285000 ;
        RECT 0.840000 1.285000 1.010000 1.445000 ;
        RECT 0.840000 1.445000 3.350000 1.615000 ;
        RECT 3.180000 1.075000 4.305000 1.285000 ;
        RECT 3.180000 1.285000 3.350000 1.445000 ;
    END
  END B
  PIN Y
    ANTENNADIFFAREA  0.953000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.075000 1.795000 5.745000 1.965000 ;
        RECT 4.075000 1.965000 4.285000 2.125000 ;
        RECT 4.985000 0.305000 6.340000 0.475000 ;
        RECT 5.495000 1.415000 6.340000 1.625000 ;
        RECT 5.495000 1.625000 5.745000 1.795000 ;
        RECT 5.495000 1.965000 5.745000 2.125000 ;
        RECT 5.950000 0.475000 6.340000 1.415000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.645000 0.910000 0.895000 ;
      RECT 0.085000  0.895000 0.315000 1.785000 ;
      RECT 0.085000  1.785000 3.780000 1.955000 ;
      RECT 0.085000  1.955000 2.280000 1.965000 ;
      RECT 0.085000  1.965000 0.400000 2.465000 ;
      RECT 0.105000  0.255000 1.380000 0.475000 ;
      RECT 0.620000  2.135000 0.870000 2.635000 ;
      RECT 1.090000  1.965000 1.340000 2.465000 ;
      RECT 1.130000  0.475000 1.380000 0.725000 ;
      RECT 1.130000  0.725000 2.320000 0.905000 ;
      RECT 1.560000  2.135000 1.810000 2.635000 ;
      RECT 1.600000  0.085000 1.770000 0.555000 ;
      RECT 1.940000  0.255000 2.320000 0.725000 ;
      RECT 2.030000  1.965000 2.280000 2.465000 ;
      RECT 2.590000  2.125000 2.840000 2.465000 ;
      RECT 2.630000  0.085000 2.800000 0.905000 ;
      RECT 2.970000  0.255000 3.350000 0.725000 ;
      RECT 2.970000  0.725000 5.755000 0.905000 ;
      RECT 3.060000  2.135000 3.310000 2.635000 ;
      RECT 3.530000  2.125000 3.855000 2.295000 ;
      RECT 3.530000  2.295000 4.755000 2.465000 ;
      RECT 3.570000  0.085000 3.740000 0.555000 ;
      RECT 3.610000  1.455000 5.205000 1.625000 ;
      RECT 3.610000  1.625000 3.780000 1.785000 ;
      RECT 3.910000  0.255000 4.325000 0.725000 ;
      RECT 4.505000  2.135000 4.755000 2.295000 ;
      RECT 4.545000  0.085000 4.715000 0.555000 ;
      RECT 5.025000  2.135000 5.275000 2.635000 ;
      RECT 5.035000  1.075000 5.745000 1.245000 ;
      RECT 5.035000  1.245000 5.205000 1.455000 ;
      RECT 5.405000  0.645000 5.755000 0.725000 ;
      RECT 5.965000  1.795000 6.340000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.665000  2.125000 2.835000 2.295000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.685000  2.125000 3.855000 2.295000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
    LAYER met1 ;
      RECT 2.605000 2.095000 2.895000 2.140000 ;
      RECT 2.605000 2.140000 3.915000 2.280000 ;
      RECT 2.605000 2.280000 2.895000 2.325000 ;
      RECT 3.625000 2.095000 3.915000 2.140000 ;
      RECT 3.625000 2.280000 3.915000 2.325000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xnor2_2
END LIBRARY
