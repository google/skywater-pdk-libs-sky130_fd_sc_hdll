* File: sky130_fd_sc_hdll__a31oi_1.spice
* Created: Wed Sep  2 08:20:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a31oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a31oi_1  VNB VPB A3 A2 A1 B1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B1	B1
* A1	A1
* A2	A2
* A3	A3
* VPB	VPB
* VNB	VNB
MM1005 A_119_47# N_A3_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.2015 PD=0.92 PS=1.92 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1002 A_203_47# N_A2_M1002_g A_119_47# VNB NSHORT L=0.15 W=0.65 AD=0.115375
+ AS=0.08775 PD=1.005 PS=0.92 NRD=22.608 NRS=14.76 M=1 R=4.33333 SA=75000.7
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g A_203_47# VNB NSHORT L=0.15 W=0.65 AD=0.121875
+ AS=0.115375 PD=1.025 PS=1.005 NRD=8.304 NRS=22.608 M=1 R=4.33333 SA=75001.2
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1003 N_VGND_M1003_d N_B1_M1003_g N_Y_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.3185 AS=0.121875 PD=2.28 PS=1.025 NRD=41.532 NRS=9.228 M=1 R=4.33333
+ SA=75001.7 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_117_297#_M1004_d N_A3_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A2_M1000_g N_A_117_297#_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.145 PD=1.325 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_A_117_297#_M1001_d N_A1_M1001_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1725 AS=0.1625 PD=1.345 PS=1.325 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90001.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_117_297#_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.28 AS=0.1725 PD=2.56 PS=1.345 NRD=2.9353 NRS=11.8003 M=1 R=5.55556
+ SA=90001.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_13 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a31oi_1.pxi.spice"
*
.ends
*
*
