* File: sky130_fd_sc_hdll__o21ba_2.pxi.spice
* Created: Thu Aug 27 19:19:41 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BA_2%B1_N N_B1_N_c_70_n N_B1_N_M1011_g N_B1_N_c_71_n
+ N_B1_N_M1005_g B1_N B1_N B1_N PM_SKY130_FD_SC_HDLL__O21BA_2%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BA_2%A_186_21# N_A_186_21#_M1004_s
+ N_A_186_21#_M1001_d N_A_186_21#_c_104_n N_A_186_21#_M1002_g
+ N_A_186_21#_c_112_n N_A_186_21#_M1000_g N_A_186_21#_c_113_n
+ N_A_186_21#_M1008_g N_A_186_21#_c_105_n N_A_186_21#_M1003_g
+ N_A_186_21#_c_106_n N_A_186_21#_c_107_n N_A_186_21#_c_172_p
+ N_A_186_21#_c_108_n N_A_186_21#_c_109_n N_A_186_21#_c_110_n
+ N_A_186_21#_c_155_p N_A_186_21#_c_115_n N_A_186_21#_c_111_n
+ PM_SKY130_FD_SC_HDLL__O21BA_2%A_186_21#
x_PM_SKY130_FD_SC_HDLL__O21BA_2%A_27_93# N_A_27_93#_M1011_s N_A_27_93#_M1005_s
+ N_A_27_93#_c_215_n N_A_27_93#_M1001_g N_A_27_93#_c_209_n N_A_27_93#_M1004_g
+ N_A_27_93#_c_210_n N_A_27_93#_c_211_n N_A_27_93#_c_218_n N_A_27_93#_c_219_n
+ N_A_27_93#_c_220_n N_A_27_93#_c_221_n N_A_27_93#_c_212_n N_A_27_93#_c_213_n
+ N_A_27_93#_c_214_n PM_SKY130_FD_SC_HDLL__O21BA_2%A_27_93#
x_PM_SKY130_FD_SC_HDLL__O21BA_2%A2 N_A2_c_283_n N_A2_M1010_g N_A2_c_284_n
+ N_A2_M1006_g A2 A2 PM_SKY130_FD_SC_HDLL__O21BA_2%A2
x_PM_SKY130_FD_SC_HDLL__O21BA_2%A1 N_A1_c_313_n N_A1_M1009_g N_A1_c_314_n
+ N_A1_M1007_g A1 A1 N_A1_c_315_n PM_SKY130_FD_SC_HDLL__O21BA_2%A1
x_PM_SKY130_FD_SC_HDLL__O21BA_2%VPWR N_VPWR_M1005_d N_VPWR_M1008_d
+ N_VPWR_M1009_d N_VPWR_c_337_n VPWR N_VPWR_c_338_n N_VPWR_c_339_n
+ N_VPWR_c_340_n N_VPWR_c_336_n N_VPWR_c_342_n N_VPWR_c_343_n N_VPWR_c_344_n
+ N_VPWR_c_345_n PM_SKY130_FD_SC_HDLL__O21BA_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BA_2%X N_X_M1002_s N_X_M1000_s N_X_c_392_n X X
+ N_X_c_410_n PM_SKY130_FD_SC_HDLL__O21BA_2%X
x_PM_SKY130_FD_SC_HDLL__O21BA_2%VGND N_VGND_M1011_d N_VGND_M1003_d
+ N_VGND_M1006_d N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n
+ N_VGND_c_428_n N_VGND_c_429_n VGND N_VGND_c_430_n N_VGND_c_431_n
+ N_VGND_c_432_n N_VGND_c_433_n PM_SKY130_FD_SC_HDLL__O21BA_2%VGND
x_PM_SKY130_FD_SC_HDLL__O21BA_2%A_518_47# N_A_518_47#_M1004_d
+ N_A_518_47#_M1007_d N_A_518_47#_c_489_n N_A_518_47#_c_486_n
+ N_A_518_47#_c_487_n N_A_518_47#_c_488_n
+ PM_SKY130_FD_SC_HDLL__O21BA_2%A_518_47#
cc_1 VNB N_B1_N_c_70_n 0.0209348f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B1_N_c_71_n 0.027205f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB B1_N 0.00303026f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_4 VNB N_A_186_21#_c_104_n 0.0199684f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_5 VNB N_A_186_21#_c_105_n 0.0197339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_186_21#_c_106_n 7.17385e-19 $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.16
cc_7 VNB N_A_186_21#_c_107_n 0.00648759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_186_21#_c_108_n 0.00517942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_186_21#_c_109_n 0.00162459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_186_21#_c_110_n 6.70754e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_186_21#_c_111_n 0.0407142f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_93#_c_209_n 0.0210882f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_93#_c_210_n 0.0368755f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_14 VNB N_A_27_93#_c_211_n 0.0132651f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.325
cc_15 VNB N_A_27_93#_c_212_n 0.0015776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_93#_c_213_n 0.0181339f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_93#_c_214_n 0.0220784f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_283_n 0.021993f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_19 VNB N_A2_c_284_n 0.0171353f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_20 VNB A2 0.00954676f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.53
cc_21 VNB N_A1_c_313_n 0.0350549f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_22 VNB N_A1_c_314_n 0.0217065f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_23 VNB N_A1_c_315_n 0.0106083f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_24 VNB N_VPWR_c_336_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 6.88344e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_424_n 0.00944581f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.325
cc_27 VNB N_VGND_c_425_n 0.0182728f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_426_n 0.0053872f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.19
cc_29 VNB N_VGND_c_427_n 0.00471543f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_428_n 0.0325632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_429_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_430_n 0.0239079f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_431_n 0.23903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_432_n 0.0243983f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_433_n 0.00553701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_518_47#_c_486_n 0.0161236f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_37 VNB N_A_518_47#_c_487_n 0.00199567f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_38 VNB N_A_518_47#_c_488_n 0.0184083f $X=-0.19 $Y=-0.24 $X2=0.715 $Y2=1.53
cc_39 VPB N_B1_N_c_71_n 0.0289456f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_40 VPB B1_N 4.81078e-19 $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.105
cc_41 VPB B1_N 0.00248918f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.445
cc_42 VPB N_A_186_21#_c_112_n 0.0181519f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_186_21#_c_113_n 0.0182975f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_44 VPB N_A_186_21#_c_109_n 0.00140353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_186_21#_c_115_n 0.00513521f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_186_21#_c_111_n 0.0212717f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_93#_c_215_n 0.0199904f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=1.105
cc_48 VPB N_A_27_93#_c_210_n 0.0204344f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_49 VPB N_A_27_93#_c_211_n 0.00732488f $X=-0.19 $Y=1.305 $X2=0.715 $Y2=1.325
cc_50 VPB N_A_27_93#_c_218_n 0.00601347f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_51 VPB N_A_27_93#_c_219_n 0.00826367f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.19
cc_52 VPB N_A_27_93#_c_220_n 8.35915e-19 $X=-0.19 $Y=1.305 $X2=0.715 $Y2=1.16
cc_53 VPB N_A_27_93#_c_221_n 0.0119905f $X=-0.19 $Y=1.305 $X2=0.74 $Y2=1.16
cc_54 VPB N_A_27_93#_c_212_n 0.00272572f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_93#_c_214_n 0.00889791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A2_c_283_n 0.0261803f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_57 VPB N_A1_c_313_n 0.0321553f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_58 VPB N_A1_c_315_n 0.0158381f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_59 VPB N_VPWR_c_337_n 0.0265149f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_60 VPB N_VPWR_c_338_n 0.0169571f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_339_n 0.0290028f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_340_n 0.0120081f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_336_n 0.0571187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_342_n 0.0240464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_343_n 0.0134349f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_344_n 0.0202127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_345_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB X 0.00163045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 N_B1_N_c_70_n N_A_186_21#_c_104_n 0.0112421f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_70 N_B1_N_c_71_n N_A_186_21#_c_112_n 0.0191956f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_71 B1_N N_A_186_21#_c_112_n 0.0021295f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_72 N_B1_N_c_71_n N_A_186_21#_c_111_n 0.0211063f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 B1_N N_A_186_21#_c_111_n 0.00251163f $X=0.655 $Y=1.105 $X2=0 $Y2=0
cc_74 B1_N N_A_186_21#_c_111_n 6.29384e-19 $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_75 N_B1_N_c_71_n N_A_27_93#_c_220_n 0.0159082f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_76 B1_N N_A_27_93#_c_220_n 0.00476922f $X=0.655 $Y=1.105 $X2=0 $Y2=0
cc_77 B1_N N_A_27_93#_c_220_n 0.0141022f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_78 N_B1_N_c_70_n N_A_27_93#_c_213_n 8.2544e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B1_N_c_70_n N_A_27_93#_c_214_n 0.0149764f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_N_c_71_n N_A_27_93#_c_214_n 0.00169815f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_81 B1_N N_A_27_93#_c_214_n 0.0251396f $X=0.655 $Y=1.105 $X2=0 $Y2=0
cc_82 B1_N N_A_27_93#_c_214_n 0.00759904f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_83 B1_N N_VPWR_M1005_d 0.00544716f $X=0.655 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_84 N_B1_N_c_71_n N_VPWR_c_338_n 0.00198707f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B1_N_c_71_n N_VPWR_c_336_n 0.00322858f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B1_N_c_71_n N_VPWR_c_342_n 0.00173541f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_87 B1_N N_X_c_392_n 0.0153654f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_88 N_B1_N_c_70_n X 8.85961e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_N_c_71_n X 2.94934e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 B1_N X 0.025897f $X=0.655 $Y=1.105 $X2=0 $Y2=0
cc_91 B1_N X 0.0126777f $X=0.655 $Y=1.445 $X2=0 $Y2=0
cc_92 N_B1_N_c_70_n N_VGND_c_424_n 0.00416861f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_93 N_B1_N_c_71_n N_VGND_c_424_n 0.00114149f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 B1_N N_VGND_c_424_n 0.0152296f $X=0.655 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B1_N_c_70_n N_VGND_c_431_n 0.00512902f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_N_c_70_n N_VGND_c_432_n 0.00510437f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_186_21#_c_109_n N_A_27_93#_c_215_n 0.00196289f $X=2.362 $Y=1.455 $X2=0
+ $Y2=0
cc_98 N_A_186_21#_c_115_n N_A_27_93#_c_215_n 0.0380026f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_99 N_A_186_21#_c_108_n N_A_27_93#_c_209_n 0.00588332f $X=2.305 $Y=0.38 $X2=0
+ $Y2=0
cc_100 N_A_186_21#_c_109_n N_A_27_93#_c_209_n 0.00459865f $X=2.362 $Y=1.455
+ $X2=0 $Y2=0
cc_101 N_A_186_21#_c_110_n N_A_27_93#_c_209_n 0.00201891f $X=2.305 $Y=0.74 $X2=0
+ $Y2=0
cc_102 N_A_186_21#_c_106_n N_A_27_93#_c_210_n 0.0013398f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_186_21#_c_107_n N_A_27_93#_c_210_n 0.00518656f $X=2.14 $Y=0.74 $X2=0
+ $Y2=0
cc_104 N_A_186_21#_c_109_n N_A_27_93#_c_210_n 0.0140884f $X=2.362 $Y=1.455 $X2=0
+ $Y2=0
cc_105 N_A_186_21#_c_110_n N_A_27_93#_c_210_n 0.00496762f $X=2.305 $Y=0.74 $X2=0
+ $Y2=0
cc_106 N_A_186_21#_c_115_n N_A_27_93#_c_210_n 7.55821e-19 $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_107 N_A_186_21#_c_111_n N_A_27_93#_c_210_n 0.0195819f $X=1.525 $Y=1.202 $X2=0
+ $Y2=0
cc_108 N_A_186_21#_c_109_n N_A_27_93#_c_211_n 0.0106435f $X=2.362 $Y=1.455 $X2=0
+ $Y2=0
cc_109 N_A_186_21#_c_115_n N_A_27_93#_c_211_n 6.36461e-19 $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_110 N_A_186_21#_c_112_n N_A_27_93#_c_220_n 0.0157047f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_111 N_A_186_21#_c_113_n N_A_27_93#_c_220_n 0.0173078f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_112 N_A_186_21#_c_106_n N_A_27_93#_c_220_n 0.0034991f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_113 N_A_186_21#_c_115_n N_A_27_93#_c_220_n 0.0152206f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_114 N_A_186_21#_c_113_n N_A_27_93#_c_212_n 0.0116452f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_A_186_21#_c_106_n N_A_27_93#_c_212_n 0.0128323f $X=1.49 $Y=1.16 $X2=0
+ $Y2=0
cc_116 N_A_186_21#_c_107_n N_A_27_93#_c_212_n 0.0134259f $X=2.14 $Y=0.74 $X2=0
+ $Y2=0
cc_117 N_A_186_21#_c_109_n N_A_27_93#_c_212_n 0.032745f $X=2.362 $Y=1.455 $X2=0
+ $Y2=0
cc_118 N_A_186_21#_c_115_n N_A_27_93#_c_212_n 0.0332884f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_119 N_A_186_21#_c_111_n N_A_27_93#_c_212_n 0.00397638f $X=1.525 $Y=1.202
+ $X2=0 $Y2=0
cc_120 N_A_186_21#_c_109_n N_A2_c_283_n 0.00147351f $X=2.362 $Y=1.455 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_186_21#_c_115_n N_A2_c_283_n 0.00352021f $X=2.78 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_186_21#_c_108_n N_A2_c_284_n 6.02205e-19 $X=2.305 $Y=0.38 $X2=0 $Y2=0
cc_123 N_A_186_21#_c_109_n N_A2_c_284_n 4.84066e-19 $X=2.362 $Y=1.455 $X2=0
+ $Y2=0
cc_124 N_A_186_21#_c_109_n A2 0.0163359f $X=2.362 $Y=1.455 $X2=0 $Y2=0
cc_125 N_A_186_21#_c_115_n A2 0.0230937f $X=2.78 $Y=1.62 $X2=0 $Y2=0
cc_126 N_A_186_21#_c_115_n N_A1_c_313_n 0.00110855f $X=2.78 $Y=1.62 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_186_21#_c_115_n N_A1_c_315_n 0.00729904f $X=2.78 $Y=1.62 $X2=0 $Y2=0
cc_128 N_A_186_21#_c_115_n N_VPWR_M1008_d 0.00655021f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_129 N_A_186_21#_c_155_p N_VPWR_c_337_n 0.0146307f $X=2.762 $Y=1.745 $X2=0
+ $Y2=0
cc_130 N_A_186_21#_c_115_n N_VPWR_c_337_n 0.00579884f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_131 N_A_186_21#_c_155_p N_VPWR_c_339_n 0.0189795f $X=2.762 $Y=1.745 $X2=0
+ $Y2=0
cc_132 N_A_186_21#_c_115_n N_VPWR_c_339_n 0.00320582f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_133 N_A_186_21#_M1001_d N_VPWR_c_336_n 0.00285422f $X=2.58 $Y=1.485 $X2=0
+ $Y2=0
cc_134 N_A_186_21#_c_112_n N_VPWR_c_336_n 0.00537865f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_186_21#_c_113_n N_VPWR_c_336_n 0.00319897f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_186_21#_c_155_p N_VPWR_c_336_n 0.0122953f $X=2.762 $Y=1.745 $X2=0
+ $Y2=0
cc_137 N_A_186_21#_c_115_n N_VPWR_c_336_n 0.00594575f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_138 N_A_186_21#_c_112_n N_VPWR_c_342_n 0.0103547f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_186_21#_c_113_n N_VPWR_c_342_n 0.00120895f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_186_21#_c_112_n N_VPWR_c_343_n 0.00461133f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_186_21#_c_113_n N_VPWR_c_343_n 0.0024422f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_186_21#_c_112_n N_VPWR_c_344_n 0.00142269f $X=1.03 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_186_21#_c_113_n N_VPWR_c_344_n 0.0152894f $X=1.525 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_186_21#_c_115_n N_VPWR_c_344_n 0.00736638f $X=2.78 $Y=1.62 $X2=0
+ $Y2=0
cc_145 N_A_186_21#_c_106_n N_X_M1002_s 5.2422e-19 $X=1.49 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_186_21#_c_172_p N_X_M1002_s 0.00179652f $X=1.575 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_186_21#_c_112_n N_X_c_392_n 0.00559747f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_186_21#_c_113_n N_X_c_392_n 0.00415118f $X=1.525 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_186_21#_c_106_n N_X_c_392_n 0.00272279f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_150 N_A_186_21#_c_111_n N_X_c_392_n 0.00665725f $X=1.525 $Y=1.202 $X2=0 $Y2=0
cc_151 N_A_186_21#_c_104_n X 0.0138252f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_186_21#_c_112_n X 0.00241341f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_186_21#_c_113_n X 0.00181494f $X=1.525 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_186_21#_c_105_n X 0.00510892f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_186_21#_c_106_n X 0.0359176f $X=1.49 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_186_21#_c_172_p X 0.0141595f $X=1.575 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_186_21#_c_111_n X 0.0213925f $X=1.525 $Y=1.202 $X2=0 $Y2=0
cc_158 N_A_186_21#_c_104_n N_X_c_410_n 0.00355546f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_186_21#_c_105_n N_X_c_410_n 0.00142386f $X=1.55 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_186_21#_c_111_n N_X_c_410_n 0.00390339f $X=1.525 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_186_21#_c_107_n N_VGND_M1003_d 0.0100985f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_162 N_A_186_21#_c_104_n N_VGND_c_424_n 0.0107061f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_186_21#_c_104_n N_VGND_c_425_n 0.0046113f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_186_21#_c_105_n N_VGND_c_425_n 0.00241736f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_165 N_A_186_21#_c_172_p N_VGND_c_425_n 0.00221971f $X=1.575 $Y=0.74 $X2=0
+ $Y2=0
cc_166 N_A_186_21#_c_104_n N_VGND_c_426_n 0.00109216f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_186_21#_c_105_n N_VGND_c_426_n 0.0115488f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_186_21#_c_107_n N_VGND_c_426_n 0.0201152f $X=2.14 $Y=0.74 $X2=0 $Y2=0
cc_169 N_A_186_21#_c_172_p N_VGND_c_426_n 0.00100003f $X=1.575 $Y=0.74 $X2=0
+ $Y2=0
cc_170 N_A_186_21#_c_108_n N_VGND_c_426_n 0.0149491f $X=2.305 $Y=0.38 $X2=0
+ $Y2=0
cc_171 N_A_186_21#_c_107_n N_VGND_c_428_n 0.00375027f $X=2.14 $Y=0.74 $X2=0
+ $Y2=0
cc_172 N_A_186_21#_c_108_n N_VGND_c_428_n 0.0209337f $X=2.305 $Y=0.38 $X2=0
+ $Y2=0
cc_173 N_A_186_21#_M1004_s N_VGND_c_431_n 0.00209319f $X=2.18 $Y=0.235 $X2=0
+ $Y2=0
cc_174 N_A_186_21#_c_104_n N_VGND_c_431_n 0.00930138f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_175 N_A_186_21#_c_105_n N_VGND_c_431_n 0.00335745f $X=1.55 $Y=0.995 $X2=0
+ $Y2=0
cc_176 N_A_186_21#_c_107_n N_VGND_c_431_n 0.00757744f $X=2.14 $Y=0.74 $X2=0
+ $Y2=0
cc_177 N_A_186_21#_c_172_p N_VGND_c_431_n 0.00425962f $X=1.575 $Y=0.74 $X2=0
+ $Y2=0
cc_178 N_A_186_21#_c_108_n N_VGND_c_431_n 0.0124067f $X=2.305 $Y=0.38 $X2=0
+ $Y2=0
cc_179 N_A_186_21#_c_108_n N_A_518_47#_c_489_n 0.0177367f $X=2.305 $Y=0.38 $X2=0
+ $Y2=0
cc_180 N_A_186_21#_c_110_n N_A_518_47#_c_489_n 0.00516904f $X=2.305 $Y=0.74
+ $X2=0 $Y2=0
cc_181 N_A_186_21#_c_109_n N_A_518_47#_c_487_n 0.00517819f $X=2.362 $Y=1.455
+ $X2=0 $Y2=0
cc_182 N_A_186_21#_c_110_n N_A_518_47#_c_487_n 0.00632777f $X=2.305 $Y=0.74
+ $X2=0 $Y2=0
cc_183 N_A_27_93#_c_215_n N_A2_c_283_n 0.0234215f $X=2.49 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_184 N_A_27_93#_c_211_n N_A2_c_283_n 0.0260283f $X=2.49 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_185 N_A_27_93#_c_209_n N_A2_c_284_n 0.0155366f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_27_93#_c_211_n A2 0.00174008f $X=2.49 $Y=1.202 $X2=0 $Y2=0
cc_187 N_A_27_93#_c_220_n N_VPWR_M1005_d 0.00628812f $X=1.915 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_188 N_A_27_93#_c_220_n N_VPWR_M1008_d 0.0167146f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_189 N_A_27_93#_c_212_n N_VPWR_M1008_d 0.0116695f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_93#_c_220_n N_VPWR_c_338_n 0.00183693f $X=1.915 $Y=1.95 $X2=0
+ $Y2=0
cc_191 N_A_27_93#_c_221_n N_VPWR_c_338_n 0.00563795f $X=0.395 $Y=1.95 $X2=0
+ $Y2=0
cc_192 N_A_27_93#_c_215_n N_VPWR_c_339_n 0.00518775f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_27_93#_c_215_n N_VPWR_c_336_n 0.00818019f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_27_93#_c_220_n N_VPWR_c_336_n 0.0214921f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_195 N_A_27_93#_c_221_n N_VPWR_c_336_n 0.00893864f $X=0.395 $Y=1.95 $X2=0
+ $Y2=0
cc_196 N_A_27_93#_c_220_n N_VPWR_c_342_n 0.0295864f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_197 N_A_27_93#_c_220_n N_VPWR_c_343_n 0.00770957f $X=1.915 $Y=1.95 $X2=0
+ $Y2=0
cc_198 N_A_27_93#_c_215_n N_VPWR_c_344_n 0.00514457f $X=2.49 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_27_93#_c_220_n N_VPWR_c_344_n 0.0398773f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_200 N_A_27_93#_c_220_n N_X_M1000_s 0.00563172f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_201 N_A_27_93#_c_220_n N_X_c_392_n 0.0246277f $X=1.915 $Y=1.95 $X2=0 $Y2=0
cc_202 N_A_27_93#_c_212_n N_X_c_392_n 0.00694472f $X=2 $Y=1.16 $X2=0 $Y2=0
cc_203 N_A_27_93#_c_213_n N_VGND_c_424_n 0.0104422f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_204 N_A_27_93#_c_209_n N_VGND_c_426_n 0.00227117f $X=2.515 $Y=0.995 $X2=0
+ $Y2=0
cc_205 N_A_27_93#_c_209_n N_VGND_c_428_n 0.00541359f $X=2.515 $Y=0.995 $X2=0
+ $Y2=0
cc_206 N_A_27_93#_c_209_n N_VGND_c_431_n 0.0113f $X=2.515 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_27_93#_c_213_n N_VGND_c_431_n 0.00885431f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_208 N_A_27_93#_c_213_n N_VGND_c_432_n 0.00842023f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_209 N_A_27_93#_c_209_n N_A_518_47#_c_489_n 0.0013994f $X=2.515 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_27_93#_c_209_n N_A_518_47#_c_487_n 0.00140025f $X=2.515 $Y=0.995
+ $X2=0 $Y2=0
cc_211 N_A2_c_283_n N_A1_c_313_n 0.0913309f $X=3.015 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_212 A2 N_A1_c_313_n 0.00132953f $X=2.895 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_213 N_A2_c_284_n N_A1_c_314_n 0.0259631f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A2_c_283_n N_A1_c_315_n 0.00193657f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_215 A2 N_A1_c_315_n 0.0178225f $X=2.895 $Y=1.19 $X2=0 $Y2=0
cc_216 N_A2_c_283_n N_VPWR_c_337_n 0.0030306f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A2_c_283_n N_VPWR_c_339_n 0.00702461f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A2_c_283_n N_VPWR_c_336_n 0.012718f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A2_c_284_n N_VGND_c_427_n 0.00268723f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_220 N_A2_c_284_n N_VGND_c_428_n 0.00439206f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A2_c_284_n N_VGND_c_431_n 0.00625689f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A2_c_283_n N_A_518_47#_c_486_n 5.76324e-19 $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A2_c_284_n N_A_518_47#_c_486_n 0.0116761f $X=3.04 $Y=0.995 $X2=0 $Y2=0
cc_224 A2 N_A_518_47#_c_486_n 0.0167245f $X=2.895 $Y=1.19 $X2=0 $Y2=0
cc_225 N_A2_c_283_n N_A_518_47#_c_487_n 0.00378812f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_226 A2 N_A_518_47#_c_487_n 0.0204648f $X=2.895 $Y=1.19 $X2=0 $Y2=0
cc_227 N_A1_c_315_n N_VPWR_M1009_d 0.00373249f $X=3.515 $Y=1.16 $X2=0 $Y2=0
cc_228 N_A1_c_313_n N_VPWR_c_337_n 0.0219598f $X=3.43 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A1_c_315_n N_VPWR_c_337_n 0.021035f $X=3.515 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A1_c_313_n N_VPWR_c_339_n 0.00427505f $X=3.43 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A1_c_313_n N_VPWR_c_336_n 0.00729026f $X=3.43 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A1_c_314_n N_VGND_c_427_n 0.00268723f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A1_c_314_n N_VGND_c_430_n 0.00439206f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A1_c_314_n N_VGND_c_431_n 0.00704219f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A1_c_313_n N_A_518_47#_c_486_n 0.00686583f $X=3.43 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A1_c_314_n N_A_518_47#_c_486_n 0.0104968f $X=3.46 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A1_c_315_n N_A_518_47#_c_486_n 0.0453921f $X=3.515 $Y=1.16 $X2=0 $Y2=0
cc_238 N_VPWR_c_336_n N_X_M1000_s 0.00392867f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_239 N_VPWR_c_336_n A_621_297# 0.0100452f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_240 X N_VGND_c_424_n 0.0260503f $X=1.12 $Y=0.51 $X2=0 $Y2=0
cc_241 N_X_c_410_n N_VGND_c_424_n 0.0126705f $X=1.215 $Y=0.38 $X2=0 $Y2=0
cc_242 N_X_c_410_n N_VGND_c_425_n 0.0180504f $X=1.215 $Y=0.38 $X2=0 $Y2=0
cc_243 N_X_c_410_n N_VGND_c_426_n 0.0127818f $X=1.215 $Y=0.38 $X2=0 $Y2=0
cc_244 N_X_M1002_s N_VGND_c_431_n 0.00436704f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_245 N_X_c_410_n N_VGND_c_431_n 0.0135275f $X=1.215 $Y=0.38 $X2=0 $Y2=0
cc_246 N_VGND_c_431_n N_A_518_47#_M1004_d 0.00690006f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_247 N_VGND_c_431_n N_A_518_47#_M1007_d 0.00259842f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_248 N_VGND_c_428_n N_A_518_47#_c_489_n 0.009328f $X=3.165 $Y=0 $X2=0 $Y2=0
cc_249 N_VGND_c_431_n N_A_518_47#_c_489_n 0.00892163f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_250 N_VGND_M1006_d N_A_518_47#_c_486_n 0.00165819f $X=3.115 $Y=0.235 $X2=0
+ $Y2=0
cc_251 N_VGND_c_427_n N_A_518_47#_c_486_n 0.0116529f $X=3.25 $Y=0.39 $X2=0 $Y2=0
cc_252 N_VGND_c_428_n N_A_518_47#_c_486_n 0.00248202f $X=3.165 $Y=0 $X2=0 $Y2=0
cc_253 N_VGND_c_430_n N_A_518_47#_c_486_n 0.00248202f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_254 N_VGND_c_431_n N_A_518_47#_c_486_n 0.0105368f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_255 N_VGND_c_430_n N_A_518_47#_c_488_n 0.0201871f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_256 N_VGND_c_431_n N_A_518_47#_c_488_n 0.0127086f $X=3.91 $Y=0 $X2=0 $Y2=0
