* File: sky130_fd_sc_hdll__a21o_4.pex.spice
* Created: Thu Aug 27 18:52:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21O_4%A_84_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 43 44 45 48 52 54 59 71
r125 70 71 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.935 $Y=1.202
+ $X2=1.96 $Y2=1.202
r126 69 70 59.5951 $w=3.68e-07 $l=4.55e-07 $layer=POLY_cond $X=1.48 $Y=1.202
+ $X2=1.935 $Y2=1.202
r127 68 69 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r128 65 66 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.975 $Y=1.202
+ $X2=1 $Y2=1.202
r129 64 65 59.5951 $w=3.68e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.975 $Y2=1.202
r130 63 64 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r131 59 61 7.61436 $w=2.78e-07 $l=1.85e-07 $layer=LI1_cond $X=4.625 $Y=0.57
+ $X2=4.625 $Y2=0.755
r132 55 57 3.05 $w=1.7e-07 $l=9.80051e-08 $layer=LI1_cond $X=3.295 $Y=0.755
+ $X2=3.21 $Y2=0.727
r133 54 61 3.65648 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.485 $Y=0.755
+ $X2=4.625 $Y2=0.755
r134 54 55 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=4.485 $Y=0.755
+ $X2=3.295 $Y2=0.755
r135 50 57 3.05 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=3.21 $Y=0.84 $X2=3.21
+ $Y2=0.727
r136 50 52 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.21 $Y=0.84
+ $X2=3.21 $Y2=1.62
r137 46 57 3.05 $w=1.7e-07 $l=1.12e-07 $layer=LI1_cond $X=3.21 $Y=0.615 $X2=3.21
+ $Y2=0.727
r138 46 48 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.21 $Y=0.615
+ $X2=3.21 $Y2=0.42
r139 44 57 3.05 $w=1.7e-07 $l=9.75705e-08 $layer=LI1_cond $X=3.125 $Y=0.7
+ $X2=3.21 $Y2=0.727
r140 44 45 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.125 $Y=0.7
+ $X2=2.3 $Y2=0.7
r141 42 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=0.785
+ $X2=2.3 $Y2=0.7
r142 42 43 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.215 $Y=0.785
+ $X2=2.215 $Y2=0.995
r143 41 71 3.92935 $w=3.68e-07 $l=3e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=1.96 $Y2=1.202
r144 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.99
+ $Y=1.16 $X2=1.99 $Y2=1.16
r145 37 68 25.5408 $w=3.68e-07 $l=1.95e-07 $layer=POLY_cond $X=1.26 $Y=1.202
+ $X2=1.455 $Y2=1.202
r146 37 66 34.0543 $w=3.68e-07 $l=2.6e-07 $layer=POLY_cond $X=1.26 $Y=1.202
+ $X2=1 $Y2=1.202
r147 36 40 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=1.26 $Y=1.16
+ $X2=1.99 $Y2=1.16
r148 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.26
+ $Y=1.16 $X2=1.26 $Y2=1.16
r149 34 43 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.13 $Y=1.16
+ $X2=2.215 $Y2=0.995
r150 34 40 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.13 $Y=1.16
+ $X2=1.99 $Y2=1.16
r151 31 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.202
r152 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.985
r153 28 70 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.935 $Y=0.995
+ $X2=1.935 $Y2=1.202
r154 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.935 $Y=0.995
+ $X2=1.935 $Y2=0.56
r155 25 69 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.48 $Y=1.41
+ $X2=1.48 $Y2=1.202
r156 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.48 $Y=1.41
+ $X2=1.48 $Y2=1.985
r157 22 68 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.455 $Y=0.995
+ $X2=1.455 $Y2=1.202
r158 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.455 $Y=0.995
+ $X2=1.455 $Y2=0.56
r159 19 66 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.202
r160 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1 $Y=1.41 $X2=1
+ $Y2=1.985
r161 16 65 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=1.202
r162 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.975 $Y=0.995
+ $X2=0.975 $Y2=0.56
r163 13 64 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.202
r164 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.52 $Y=1.41
+ $X2=0.52 $Y2=1.985
r165 10 63 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=1.202
r166 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.495 $Y=0.995
+ $X2=0.495 $Y2=0.56
r167 3 52 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.065
+ $Y=1.485 $X2=3.21 $Y2=1.62
r168 2 59 182 $w=1.7e-07 $l=4.17373e-07 $layer=licon1_NDIFF $count=1 $X=4.435
+ $Y=0.235 $X2=4.62 $Y2=0.57
r169 1 57 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.235 $X2=3.21 $Y2=0.76
r170 1 48 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=3.025
+ $Y=0.235 $X2=3.21 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%B1 1 3 4 6 7 9 10 12 13 20 23
c50 7 0 1.28785e-19 $X=3.445 $Y=1.41
r51 20 21 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=3.445 $Y=1.202
+ $X2=3.47 $Y2=1.202
r52 19 20 61.393 $w=3.69e-07 $l=4.7e-07 $layer=POLY_cond $X=2.975 $Y=1.202
+ $X2=3.445 $Y2=1.202
r53 18 19 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=2.95 $Y=1.202
+ $X2=2.975 $Y2=1.202
r54 16 18 16.981 $w=3.69e-07 $l=1.3e-07 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.95 $Y2=1.202
r55 13 23 4.5135 $w=5.28e-07 $l=2e-07 $layer=LI1_cond $X=2.75 $Y=1.26 $X2=2.55
+ $Y2=1.26
r56 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.82
+ $Y=1.16 $X2=2.82 $Y2=1.16
r57 10 21 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.47 $Y=0.995
+ $X2=3.47 $Y2=1.202
r58 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.47 $Y=0.995
+ $X2=3.47 $Y2=0.56
r59 7 20 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.445 $Y=1.41
+ $X2=3.445 $Y2=1.202
r60 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.445 $Y=1.41
+ $X2=3.445 $Y2=1.985
r61 4 19 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.202
r62 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.975 $Y=1.41
+ $X2=2.975 $Y2=1.985
r63 1 18 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.95 $Y=0.995
+ $X2=2.95 $Y2=1.202
r64 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.95 $Y=0.995 $X2=2.95
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%A2 1 3 4 6 7 9 10 12 14 15 16 18 24 30 33
+ 38
c84 14 0 1.28785e-19 $X=4.057 $Y=1.51
r85 33 38 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.285 $Y=1.595
+ $X2=5.285 $Y2=1.51
r86 33 38 1.26769 $w=2.98e-07 $l=3.3e-08 $layer=LI1_cond $X=5.285 $Y=1.477
+ $X2=5.285 $Y2=1.51
r87 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.36
+ $Y=1.16 $X2=5.36 $Y2=1.16
r88 27 33 7.18356 $w=2.98e-07 $l=1.87e-07 $layer=LI1_cond $X=5.285 $Y=1.29
+ $X2=5.285 $Y2=1.477
r89 27 30 3.67801 $w=2.33e-07 $l=7.5e-08 $layer=LI1_cond $X=5.285 $Y=1.172
+ $X2=5.36 $Y2=1.172
r90 21 24 7.26257 $w=2.63e-07 $l=1.67e-07 $layer=LI1_cond $X=3.89 $Y=1.142
+ $X2=4.057 $Y2=1.142
r91 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.89
+ $Y=1.16 $X2=3.89 $Y2=1.16
r92 16 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.17 $Y=1.595
+ $X2=4.85 $Y2=1.595
r93 15 33 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.135 $Y=1.595
+ $X2=5.285 $Y2=1.595
r94 15 18 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=5.135 $Y=1.595
+ $X2=4.85 $Y2=1.595
r95 14 16 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=4.057 $Y=1.51
+ $X2=4.17 $Y2=1.595
r96 13 24 1.71951 $w=2.25e-07 $l=1.33e-07 $layer=LI1_cond $X=4.057 $Y=1.275
+ $X2=4.057 $Y2=1.142
r97 13 14 12.0366 $w=2.23e-07 $l=2.35e-07 $layer=LI1_cond $X=4.057 $Y=1.275
+ $X2=4.057 $Y2=1.51
r98 10 31 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.325 $Y=1.41
+ $X2=5.385 $Y2=1.16
r99 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.325 $Y=1.41
+ $X2=5.325 $Y2=1.985
r100 7 31 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=5.3 $Y=0.995
+ $X2=5.385 $Y2=1.16
r101 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.3 $Y=0.995 $X2=5.3
+ $Y2=0.56
r102 4 22 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.915 $Y2=1.16
r103 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.93 $Y=0.995
+ $X2=3.93 $Y2=0.56
r104 1 22 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.915 $Y=1.41
+ $X2=3.915 $Y2=1.16
r105 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.915 $Y=1.41
+ $X2=3.915 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%A1 1 3 4 6 7 9 10 12 13 20 23
r46 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.855 $Y=1.202
+ $X2=4.88 $Y2=1.202
r47 19 23 8.69768 $w=2.63e-07 $l=2e-07 $layer=LI1_cond $X=4.59 $Y=1.142 $X2=4.39
+ $Y2=1.142
r48 18 20 33.6132 $w=3.8e-07 $l=2.65e-07 $layer=POLY_cond $X=4.59 $Y=1.202
+ $X2=4.855 $Y2=1.202
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.59
+ $Y=1.16 $X2=4.59 $Y2=1.16
r50 16 18 26.0026 $w=3.8e-07 $l=2.05e-07 $layer=POLY_cond $X=4.385 $Y=1.202
+ $X2=4.59 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.36 $Y=1.202
+ $X2=4.385 $Y2=1.202
r52 13 19 10.6547 $w=2.63e-07 $l=2.45e-07 $layer=LI1_cond $X=4.835 $Y=1.142
+ $X2=4.59 $Y2=1.142
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.88 $Y=0.995
+ $X2=4.88 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.88 $Y=0.995
+ $X2=4.88 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.855 $Y=1.41
+ $X2=4.855 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.855 $Y=1.41
+ $X2=4.855 $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.385 $Y=1.41
+ $X2=4.385 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.385 $Y=1.41
+ $X2=4.385 $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.36 $Y=0.995
+ $X2=4.36 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.36 $Y=0.995 $X2=4.36
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%VPWR 1 2 3 4 5 16 18 22 24 28 33 36 40 43
+ 46 48 64 65 71 74
r102 74 75 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r103 72 75 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r104 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r105 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r107 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r108 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r109 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r110 56 59 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r111 56 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 55 58 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r114 53 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.19 $Y2=2.72
r115 53 55 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.315 $Y=2.72
+ $X2=2.53 $Y2=2.72
r116 52 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r118 49 68 4.73185 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.222 $Y2=2.72
r119 49 51 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=2.72
+ $X2=0.69 $Y2=2.72
r120 48 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=1.215 $Y2=2.72
r121 48 51 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 46 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 46 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 44 64 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.255 $Y=2.72
+ $X2=5.75 $Y2=2.72
r125 43 61 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 42 44 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=5.255 $Y2=2.72
r127 42 43 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.065 $Y=2.72
+ $X2=4.875 $Y2=2.72
r128 40 42 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.065 $Y=2.36
+ $X2=5.065 $Y2=2.72
r129 37 61 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.315 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 36 58 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r131 35 37 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=4.315 $Y2=2.72
r132 35 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.125 $Y=2.72
+ $X2=3.935 $Y2=2.72
r133 33 35 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.125 $Y=2.36
+ $X2=4.125 $Y2=2.72
r134 28 31 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=2.19 $Y=1.68
+ $X2=2.19 $Y2=2.36
r135 26 74 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r136 26 31 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.36
r137 25 71 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.405 $Y=2.72
+ $X2=1.215 $Y2=2.72
r138 24 74 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=2.19 $Y2=2.72
r139 24 25 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=2.065 $Y=2.72
+ $X2=1.405 $Y2=2.72
r140 20 71 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=2.72
r141 20 22 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=1.215 $Y=2.635
+ $X2=1.215 $Y2=2.02
r142 16 68 3.03433 $w=3.3e-07 $l=1.1025e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.222 $Y2=2.72
r143 16 18 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=0.28 $Y=2.635
+ $X2=0.28 $Y2=2.02
r144 5 40 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.945
+ $Y=1.485 $X2=5.09 $Y2=2.36
r145 4 33 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=4.005
+ $Y=1.485 $X2=4.15 $Y2=2.36
r146 3 31 400 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.485 $X2=2.2 $Y2=2.36
r147 3 28 400 $w=1.7e-07 $l=2.59374e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.485 $X2=2.2 $Y2=1.68
r148 2 22 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=1.09
+ $Y=1.485 $X2=1.24 $Y2=2.02
r149 1 18 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%X 1 2 3 4 15 17 21 23 25 27 32 38
r48 35 38 1.22961 $w=5.33e-07 $l=5.5e-08 $layer=LI1_cond $X=0.412 $Y=1.585
+ $X2=0.412 $Y2=1.53
r49 32 35 2.71818 $w=3.52e-07 $l=1.19499e-07 $layer=LI1_cond $X=0.495 $Y=1.67
+ $X2=0.412 $Y2=1.585
r50 32 38 0.335349 $w=5.33e-07 $l=1.5e-08 $layer=LI1_cond $X=0.412 $Y=1.515
+ $X2=0.412 $Y2=1.53
r51 29 32 16.3203 $w=5.33e-07 $l=7.3e-07 $layer=LI1_cond $X=0.412 $Y=0.785
+ $X2=0.412 $Y2=1.515
r52 25 31 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=1.755
+ $X2=1.76 $Y2=1.67
r53 25 27 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=1.76 $Y=1.755
+ $X2=1.76 $Y2=2.02
r54 24 32 4.06059 $w=1.7e-07 $l=3.5e-07 $layer=LI1_cond $X=0.845 $Y=1.67
+ $X2=0.495 $Y2=1.67
r55 23 31 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.635 $Y=1.67
+ $X2=1.76 $Y2=1.67
r56 23 24 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=1.635 $Y=1.67
+ $X2=0.845 $Y2=1.67
r57 19 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=0.76 $Y=0.7 $X2=1.72
+ $Y2=0.7
r58 17 29 9.52189 $w=1.7e-07 $l=3.07578e-07 $layer=LI1_cond $X=0.68 $Y=0.7
+ $X2=0.412 $Y2=0.785
r59 17 19 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=0.68 $Y=0.7 $X2=0.76
+ $Y2=0.7
r60 13 32 2.71818 $w=3.52e-07 $l=3.04549e-07 $layer=LI1_cond $X=0.76 $Y=1.755
+ $X2=0.495 $Y2=1.67
r61 13 15 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.76 $Y=1.755
+ $X2=0.76 $Y2=2.02
r62 4 31 600 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.485 $X2=1.72 $Y2=1.67
r63 4 27 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=1.57
+ $Y=1.485 $X2=1.72 $Y2=2.02
r64 3 32 600 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.485 $X2=0.76 $Y2=1.67
r65 3 15 600 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=1 $X=0.61
+ $Y=1.485 $X2=0.76 $Y2=2.02
r66 2 21 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=1.53
+ $Y=0.235 $X2=1.72 $Y2=0.7
r67 1 19 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=0.57
+ $Y=0.235 $X2=0.76 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%A_523_297# 1 2 3 4 15 17 18 21 26 27 31 33
+ 39 43 45
r66 37 45 3.22182 $w=2.92e-07 $l=1.01833e-07 $layer=LI1_cond $X=5.732 $Y=1.85
+ $X2=5.695 $Y2=1.935
r67 37 39 9.94265 $w=2.53e-07 $l=2.2e-07 $layer=LI1_cond $X=5.732 $Y=1.85
+ $X2=5.732 $Y2=1.63
r68 34 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.705 $Y=1.935
+ $X2=4.62 $Y2=1.935
r69 33 45 3.35233 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.53 $Y=1.935
+ $X2=5.695 $Y2=1.935
r70 33 34 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.53 $Y=1.935
+ $X2=4.705 $Y2=1.935
r71 29 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.62 $Y=2.02 $X2=4.62
+ $Y2=1.935
r72 29 31 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=4.62 $Y=2.02
+ $X2=4.62 $Y2=2.3
r73 28 41 1.54918 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=3.765 $Y=1.935
+ $X2=3.675 $Y2=1.935
r74 27 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.535 $Y=1.935
+ $X2=4.62 $Y2=1.935
r75 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.535 $Y=1.935
+ $X2=3.765 $Y2=1.935
r76 24 26 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=3.675 $Y=2.295
+ $X2=3.675 $Y2=2.055
r77 23 41 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=2.02
+ $X2=3.675 $Y2=1.935
r78 23 26 2.15657 $w=1.78e-07 $l=3.5e-08 $layer=LI1_cond $X=3.675 $Y=2.02
+ $X2=3.675 $Y2=2.055
r79 19 41 4.92476 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.85
+ $X2=3.675 $Y2=1.935
r80 19 21 14.7879 $w=1.78e-07 $l=2.4e-07 $layer=LI1_cond $X=3.675 $Y=1.85
+ $X2=3.675 $Y2=1.61
r81 17 24 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=3.585 $Y=2.38
+ $X2=3.675 $Y2=2.295
r82 17 18 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=3.585 $Y=2.38
+ $X2=2.825 $Y2=2.38
r83 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.74 $Y=2.295
+ $X2=2.825 $Y2=2.38
r84 13 15 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.74 $Y=2.295
+ $X2=2.74 $Y2=1.86
r85 4 45 300 $w=1.7e-07 $l=6.09118e-07 $layer=licon1_PDIFF $count=2 $X=5.415
+ $Y=1.485 $X2=5.695 $Y2=1.97
r86 4 39 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=5.415
+ $Y=1.485 $X2=5.695 $Y2=1.63
r87 3 43 600 $w=1.7e-07 $l=5.17446e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.62 $Y2=1.935
r88 3 31 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.62 $Y2=2.3
r89 2 26 600 $w=1.7e-07 $l=6.38396e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=1.485 $X2=3.68 $Y2=2.055
r90 2 21 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.535
+ $Y=1.485 $X2=3.68 $Y2=1.61
r91 1 15 300 $w=1.7e-07 $l=4.33013e-07 $layer=licon1_PDIFF $count=2 $X=2.615
+ $Y=1.485 $X2=2.74 $Y2=1.86
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21O_4%VGND 1 2 3 4 5 16 18 22 24 26 29 30 31 33
+ 47 59 67 70 73
r85 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r86 69 70 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.72 $Y=0.18
+ $X2=2.885 $Y2=0.18
r87 65 69 4.28783 $w=5.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.72 $Y2=0.18
r88 65 67 15.4591 $w=5.28e-07 $l=4.2e-07 $layer=LI1_cond $X=2.53 $Y=0.18
+ $X2=2.11 $Y2=0.18
r89 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r90 59 62 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.215 $Y=0 $X2=1.215
+ $Y2=0.36
r91 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r92 53 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r93 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r94 50 53 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r95 49 52 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r96 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r97 47 72 4.10258 $w=1.7e-07 $l=2.67e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=5.712
+ $Y2=0
r98 47 52 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.445 $Y=0 $X2=5.29
+ $Y2=0
r99 46 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r100 46 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r101 45 70 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.885
+ $Y2=0
r102 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r103 42 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r104 42 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r105 41 67 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.11
+ $Y2=0
r106 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r107 39 59 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=1.215
+ $Y2=0
r108 39 41 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.405 $Y=0 $X2=2.07
+ $Y2=0
r109 37 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r110 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r111 34 55 4.84988 $w=1.7e-07 $l=2.23e-07 $layer=LI1_cond $X=0.445 $Y=0
+ $X2=0.222 $Y2=0
r112 34 36 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.445 $Y=0 $X2=0.69
+ $Y2=0
r113 33 59 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.215
+ $Y2=0
r114 33 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0
+ $X2=0.69 $Y2=0
r115 31 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r116 31 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r117 29 45 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.555 $Y=0
+ $X2=3.45 $Y2=0
r118 29 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0 $X2=3.72
+ $Y2=0
r119 28 49 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.91
+ $Y2=0
r120 28 30 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0 $X2=3.72
+ $Y2=0
r121 24 72 3.25748 $w=2.8e-07 $l=1.64085e-07 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.712 $Y2=0
r122 24 26 12.1418 $w=2.78e-07 $l=2.95e-07 $layer=LI1_cond $X=5.585 $Y=0.085
+ $X2=5.585 $Y2=0.38
r123 20 30 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0
r124 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.72 $Y=0.085
+ $X2=3.72 $Y2=0.36
r125 16 55 3.00127 $w=3.4e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.222 $Y2=0
r126 16 18 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.36
r127 5 26 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=5.375
+ $Y=0.235 $X2=5.56 $Y2=0.38
r128 4 22 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=3.545
+ $Y=0.235 $X2=3.72 $Y2=0.36
r129 3 69 91 $w=1.7e-07 $l=7.69968e-07 $layer=licon1_NDIFF $count=2 $X=2.01
+ $Y=0.235 $X2=2.72 $Y2=0.36
r130 2 62 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.05
+ $Y=0.235 $X2=1.24 $Y2=0.36
r131 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

