* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
X0 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 VGND B2 a_616_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_616_47# B2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_96_21# A1 a_1008_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 X a_96_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_96_21# B1 a_616_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VPWR A2 a_524_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_96_21# B2 a_524_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_524_297# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_524_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_524_297# B1 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 VGND A2 a_1008_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_1008_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_1008_47# A1 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VPWR A1 a_524_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND a_96_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 X a_96_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_96_21# B1 a_524_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 a_616_47# B1 a_96_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VPWR a_96_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_524_297# B2 a_96_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
