* File: sky130_fd_sc_hdll__and4_1.spice
* Created: Wed Sep  2 08:22:53 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4_1.pex.spice"
.subckt sky130_fd_sc_hdll__and4_1  VNB VPB A B C D VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* D	D
* C	C
* B	B
* A	A
* VPB	VPB
* VNB	VNB
MM1007 A_119_47# N_A_M1007_g N_A_27_47#_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=22.848 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1002 A_203_47# N_B_M1002_g A_119_47# VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0567 PD=0.75 PS=0.69 NRD=31.428 NRS=22.848 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1006 A_299_47# N_C_M1006_g A_203_47# VNB NSHORT L=0.15 W=0.42 AD=0.0714
+ AS=0.0693 PD=0.76 PS=0.75 NRD=32.856 NRS=31.428 M=1 R=2.8 SA=75001.1
+ SB=75001.5 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1000_d N_D_M1000_g A_299_47# VNB NSHORT L=0.15 W=0.42 AD=0.108042
+ AS=0.0714 PD=0.863551 PS=0.76 NRD=14.28 NRS=32.856 M=1 R=2.8 SA=75001.6
+ SB=75001 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_27_47#_M1005_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2925 AS=0.167208 PD=2.2 PS=1.33645 NRD=34.152 NRS=22.152 M=1 R=4.33333
+ SA=75001.5 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1001 N_A_27_47#_M1001_d N_A_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0609 AS=0.1134 PD=0.71 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1008_d N_B_M1008_g N_A_27_47#_M1001_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.063 AS=0.0609 PD=0.72 PS=0.71 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.6 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1004 N_A_27_47#_M1004_d N_C_M1004_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0651 AS=0.063 PD=0.73 PS=0.72 NRD=4.6886 NRS=7.0329 M=1 R=2.33333
+ SA=90001.1 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1009 N_VPWR_M1009_d N_D_M1009_g N_A_27_47#_M1004_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0948549 AS=0.0651 PD=0.810423 PS=0.73 NRD=41.0351 NRS=9.3772 M=1
+ R=2.33333 SA=90001.6 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.46 AS=0.225845 PD=2.92 PS=1.92958 NRD=38.3953 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.4 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX11_noxref noxref_14 B B PROBETYPE=1
pX12_noxref noxref_15 B B PROBETYPE=1
pX13_noxref noxref_16 C C PROBETYPE=1
pX14_noxref noxref_17 C C PROBETYPE=1
pX15_noxref noxref_18 C C PROBETYPE=1
pX16_noxref noxref_19 D D PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and4_1.pxi.spice"
*
.ends
*
*
