* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4bb_1 A_N B_N C D VGND VNB VPB VPWR Y
M1000 VPWR B_N a_27_93# VPB phighvt w=420000u l=180000u
+  ad=1.1325e+12p pd=8.99e+06u as=1.134e+11p ps=1.38e+06u
M1001 VPWR a_500_21# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=7e+11p ps=5.4e+06u
M1002 a_434_47# a_27_93# a_334_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=2.275e+11p ps=2e+06u
M1003 Y D VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_334_47# C a_218_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.795e+11p ps=2.16e+06u
M1005 VPWR C Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y a_500_21# a_434_47# VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1007 a_218_47# D VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=3.372e+11p ps=3.45e+06u
M1008 a_500_21# A_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1009 Y a_27_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_500_21# A_N VGND VNB nshort w=420000u l=150000u
+  ad=1.533e+11p pd=1.57e+06u as=0p ps=0u
M1011 VGND B_N a_27_93# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.092e+11p ps=1.36e+06u
.ends
