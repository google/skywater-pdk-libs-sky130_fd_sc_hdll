* File: sky130_fd_sc_hdll__and3b_4.pex.spice
* Created: Thu Aug 27 18:58:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%A_98_199# 1 2 7 9 10 12 14 15 16 21 27
c75 16 0 7.42278e-20 $X=0.865 $Y=1.99
c76 7 0 1.60824e-19 $X=0.71 $Y=1.41
r77 24 27 5.13361 $w=3.28e-07 $l=1.47e-07 $layer=LI1_cond $X=0.625 $Y=1.16
+ $X2=0.772 $Y2=1.16
r78 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.625
+ $Y=1.16 $X2=0.625 $Y2=1.16
r79 19 21 52.8889 $w=2.78e-07 $l=1.285e-06 $layer=LI1_cond $X=4.765 $Y=1.875
+ $X2=4.765 $Y2=0.59
r80 16 18 186.145 $w=2.28e-07 $l=3.715e-06 $layer=LI1_cond $X=0.865 $Y=1.99
+ $X2=4.58 $Y2=1.99
r81 15 19 6.90206 $w=2.3e-07 $l=1.88944e-07 $layer=LI1_cond $X=4.625 $Y=1.99
+ $X2=4.765 $Y2=1.875
r82 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.625 $Y=1.99
+ $X2=4.58 $Y2=1.99
r83 14 16 6.92126 $w=2.3e-07 $l=1.54661e-07 $layer=LI1_cond $X=0.772 $Y=1.875
+ $X2=0.865 $Y2=1.99
r84 13 27 4.14273 $w=1.85e-07 $l=1.65e-07 $layer=LI1_cond $X=0.772 $Y=1.325
+ $X2=0.772 $Y2=1.16
r85 13 14 32.973 $w=1.83e-07 $l=5.5e-07 $layer=LI1_cond $X=0.772 $Y=1.325
+ $X2=0.772 $Y2=1.875
r86 10 25 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.735 $Y=0.995
+ $X2=0.65 $Y2=1.16
r87 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.735 $Y=0.995
+ $X2=0.735 $Y2=0.56
r88 7 25 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.71 $Y=1.41
+ $X2=0.65 $Y2=1.16
r89 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.71 $Y=1.41 $X2=0.71
+ $Y2=1.985
r90 2 18 600 $w=1.7e-07 $l=3.62319e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.725 $X2=4.58 $Y2=2.02
r91 1 21 182 $w=1.7e-07 $l=3.26573e-07 $layer=licon1_NDIFF $count=1 $X=4.44
+ $Y=0.465 $X2=4.71 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%B 1 3 4 6 7 8
r34 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.155
+ $Y=1.16 $X2=1.155 $Y2=1.16
r35 7 8 14.2903 $w=2.48e-07 $l=3.1e-07 $layer=LI1_cond $X=1.16 $Y=0.85 $X2=1.16
+ $Y2=1.16
r36 4 12 38.6069 $w=3.31e-07 $l=2.12238e-07 $layer=POLY_cond $X=1.31 $Y=0.995
+ $X2=1.202 $Y2=1.16
r37 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.31 $Y=0.995 $X2=1.31
+ $Y2=0.56
r38 1 12 46.3664 $w=3.31e-07 $l=2.88531e-07 $layer=POLY_cond $X=1.285 $Y=1.41
+ $X2=1.202 $Y2=1.16
r39 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.285 $Y=1.41
+ $X2=1.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%C 1 3 4 6 7 13
c39 4 0 1.52606e-19 $X=1.785 $Y=1.41
r40 7 13 3.34041 $w=3.43e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=1.167 $X2=1.61
+ $Y2=1.167
r41 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r42 4 10 48.1208 $w=2.95e-07 $l=2.64575e-07 $layer=POLY_cond $X=1.785 $Y=1.41
+ $X2=1.755 $Y2=1.16
r43 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.785 $Y=1.41
+ $X2=1.785 $Y2=1.985
r44 1 10 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=1.74 $Y=0.995
+ $X2=1.755 $Y2=1.16
r45 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.74 $Y=0.995 $X2=1.74
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%A_56_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 38 40 44 47 49 55 59 64 65 66 70 79
c148 44 0 8.37355e-20 $X=2.035 $Y=0.71
c149 40 0 1.60824e-19 $X=2.035 $Y=1.61
r150 79 80 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.78 $Y=1.202
+ $X2=3.805 $Y2=1.202
r151 78 79 62.3612 $w=3.71e-07 $l=4.8e-07 $layer=POLY_cond $X=3.3 $Y=1.202
+ $X2=3.78 $Y2=1.202
r152 77 78 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.275 $Y=1.202
+ $X2=3.3 $Y2=1.202
r153 74 75 4.54717 $w=3.71e-07 $l=3.5e-08 $layer=POLY_cond $X=2.795 $Y=1.202
+ $X2=2.83 $Y2=1.202
r154 71 72 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.315 $Y=1.202
+ $X2=2.34 $Y2=1.202
r155 66 68 16.0202 $w=1.78e-07 $l=2.6e-07 $layer=LI1_cond $X=1.61 $Y=0.45
+ $X2=1.61 $Y2=0.71
r156 64 65 7.01282 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.33 $Y=1.66
+ $X2=0.33 $Y2=1.495
r157 62 65 36.1448 $w=2.18e-07 $l=6.9e-07 $layer=LI1_cond $X=0.26 $Y=0.805
+ $X2=0.26 $Y2=1.495
r158 61 62 12.3665 $w=4.83e-07 $l=3.55e-07 $layer=LI1_cond $X=0.392 $Y=0.45
+ $X2=0.392 $Y2=0.805
r159 59 61 1.7263 $w=4.83e-07 $l=7e-08 $layer=LI1_cond $X=0.392 $Y=0.38
+ $X2=0.392 $Y2=0.45
r160 56 77 11.6927 $w=3.71e-07 $l=9e-08 $layer=POLY_cond $X=3.185 $Y=1.202
+ $X2=3.275 $Y2=1.202
r161 56 75 46.1213 $w=3.71e-07 $l=3.55e-07 $layer=POLY_cond $X=3.185 $Y=1.202
+ $X2=2.83 $Y2=1.202
r162 55 56 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.185
+ $Y=1.16 $X2=3.185 $Y2=1.16
r163 53 74 50.6685 $w=3.71e-07 $l=3.9e-07 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.795 $Y2=1.202
r164 53 72 8.44474 $w=3.71e-07 $l=6.5e-08 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.34 $Y2=1.202
r165 52 55 26.833 $w=3.33e-07 $l=7.8e-07 $layer=LI1_cond $X=2.405 $Y=1.187
+ $X2=3.185 $Y2=1.187
r166 52 53 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.405
+ $Y=1.16 $X2=2.405 $Y2=1.16
r167 50 70 0.43014 $w=3.35e-07 $l=1.15e-07 $layer=LI1_cond $X=2.265 $Y=1.187
+ $X2=2.15 $Y2=1.187
r168 50 52 4.81618 $w=3.33e-07 $l=1.4e-07 $layer=LI1_cond $X=2.265 $Y=1.187
+ $X2=2.405 $Y2=1.187
r169 48 70 7.74634 $w=2e-07 $l=1.82384e-07 $layer=LI1_cond $X=2.12 $Y=1.355
+ $X2=2.15 $Y2=1.187
r170 48 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.12 $Y=1.355
+ $X2=2.12 $Y2=1.525
r171 47 70 7.74634 $w=2e-07 $l=1.67e-07 $layer=LI1_cond $X=2.15 $Y=1.02 $X2=2.15
+ $Y2=1.187
r172 46 47 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=2.15 $Y=0.805
+ $X2=2.15 $Y2=1.02
r173 45 68 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.7 $Y=0.71 $X2=1.61
+ $Y2=0.71
r174 44 46 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=2.035 $Y=0.71
+ $X2=2.15 $Y2=0.805
r175 44 45 19.555 $w=1.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.035 $Y=0.71
+ $X2=1.7 $Y2=0.71
r176 40 49 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.035 $Y=1.61
+ $X2=2.12 $Y2=1.525
r177 40 42 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=2.035 $Y=1.61
+ $X2=1.545 $Y2=1.61
r178 39 61 6.27638 $w=1.9e-07 $l=2.43e-07 $layer=LI1_cond $X=0.635 $Y=0.45
+ $X2=0.392 $Y2=0.45
r179 38 66 0.384081 $w=1.9e-07 $l=9e-08 $layer=LI1_cond $X=1.52 $Y=0.45 $X2=1.61
+ $Y2=0.45
r180 38 39 51.6603 $w=1.88e-07 $l=8.85e-07 $layer=LI1_cond $X=1.52 $Y=0.45
+ $X2=0.635 $Y2=0.45
r181 31 80 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.805 $Y=0.995
+ $X2=3.805 $Y2=1.202
r182 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.805 $Y=0.995
+ $X2=3.805 $Y2=0.56
r183 28 79 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.78 $Y=1.41
+ $X2=3.78 $Y2=1.202
r184 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.78 $Y=1.41
+ $X2=3.78 $Y2=1.985
r185 25 78 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.3 $Y=1.41
+ $X2=3.3 $Y2=1.202
r186 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.3 $Y=1.41
+ $X2=3.3 $Y2=1.985
r187 22 77 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.275 $Y=0.995
+ $X2=3.275 $Y2=1.202
r188 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.275 $Y=0.995
+ $X2=3.275 $Y2=0.56
r189 19 75 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.83 $Y=1.41
+ $X2=2.83 $Y2=1.202
r190 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.83 $Y=1.41
+ $X2=2.83 $Y2=1.985
r191 16 74 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.795 $Y=0.995
+ $X2=2.795 $Y2=1.202
r192 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.795 $Y=0.995
+ $X2=2.795 $Y2=0.56
r193 13 72 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.34 $Y=1.41
+ $X2=2.34 $Y2=1.202
r194 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.34 $Y=1.41
+ $X2=2.34 $Y2=1.985
r195 10 71 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=1.202
r196 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.315 $Y=0.995
+ $X2=2.315 $Y2=0.56
r197 3 42 600 $w=1.7e-07 $l=2.23942e-07 $layer=licon1_PDIFF $count=1 $X=1.375
+ $Y=1.485 $X2=1.545 $Y2=1.61
r198 2 64 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.28
+ $Y=1.485 $X2=0.425 $Y2=1.66
r199 1 59 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=0.305
+ $Y=0.235 $X2=0.47 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%A_N 2 3 6 9 11 12 16 18
c41 6 0 1.92207e-19 $X=4.34 $Y=1.935
r42 16 19 37.7763 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.277 $Y=1.16
+ $X2=4.277 $Y2=1.325
r43 16 18 46.1766 $w=3.25e-07 $l=1.65e-07 $layer=POLY_cond $X=4.277 $Y=1.16
+ $X2=4.277 $Y2=0.995
r44 11 12 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=4.31 $Y=1.16
+ $X2=4.31 $Y2=1.53
r45 11 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=1.16 $X2=4.25 $Y2=1.16
r46 9 18 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=4.365 $Y=0.675
+ $X2=4.365 $Y2=0.995
r47 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.34 $Y=1.65 $X2=4.34
+ $Y2=1.935
r48 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.34 $Y=1.55 $X2=4.34
+ $Y2=1.65
r49 2 19 74.6049 $w=2e-07 $l=2.25e-07 $layer=POLY_cond $X=4.34 $Y=1.55 $X2=4.34
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%VPWR 1 2 3 4 15 17 19 24 29 34 41 42 45 52
+ 55 62
c68 1 0 7.42278e-20 $X=0.8 $Y=1.485
r69 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r70 62 65 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.995 $Y=2.36
+ $X2=3.995 $Y2=2.72
r71 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r73 45 48 8.61176 $w=4.98e-07 $l=3.6e-07 $layer=LI1_cond $X=0.98 $Y=2.36
+ $X2=0.98 $Y2=2.72
r74 42 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r75 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 39 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=3.995 $Y2=2.72
r77 39 41 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.83 $Y2=2.72
r78 38 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r79 38 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r80 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r81 35 37 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=3.23 $Y=2.72
+ $X2=3.45 $Y2=2.72
r82 34 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.995 $Y2=2.72
r83 34 37 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=2.72
+ $X2=3.45 $Y2=2.72
r84 33 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r85 33 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r87 30 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.06 $Y2=2.72
r88 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.53 $Y2=2.72
r89 29 35 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=3.037 $Y=2.72
+ $X2=3.23 $Y2=2.72
r90 29 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r91 29 55 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=3.037 $Y=2.72
+ $X2=3.037 $Y2=2.36
r92 29 32 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=2.72
+ $X2=2.53 $Y2=2.72
r93 28 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r94 28 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r96 25 48 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=1.23 $Y=2.72 $X2=0.98
+ $Y2=2.72
r97 25 27 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r98 24 52 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.06 $Y2=2.72
r99 24 27 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r100 22 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r101 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r102 19 48 7.15667 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=0.73 $Y=2.72
+ $X2=0.98 $Y2=2.72
r103 19 21 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=0.73 $Y=2.72 $X2=0.69
+ $Y2=2.72
r104 17 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r105 13 52 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2.72
r106 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.06 $Y=2.635
+ $X2=2.06 $Y2=2.36
r107 4 62 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.87
+ $Y=1.485 $X2=4.02 $Y2=2.36
r108 3 55 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.92
+ $Y=1.485 $X2=3.065 $Y2=2.36
r109 2 15 600 $w=1.7e-07 $l=9.63068e-07 $layer=licon1_PDIFF $count=1 $X=1.875
+ $Y=1.485 $X2=2.06 $Y2=2.36
r110 1 45 600 $w=1.7e-07 $l=9.76601e-07 $layer=licon1_PDIFF $count=1 $X=0.8
+ $Y=1.485 $X2=1.015 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%X 1 2 3 4 13 19 23 28 30 35
c56 13 0 3.44813e-19 $X=3.57 $Y=1.62
r57 33 35 0.135582 $w=4.23e-07 $l=5e-09 $layer=LI1_cond $X=3.782 $Y=0.845
+ $X2=3.782 $Y2=0.85
r58 30 33 3.61955 $w=3.47e-07 $l=1.57972e-07 $layer=LI1_cond $X=3.68 $Y=0.73
+ $X2=3.782 $Y2=0.845
r59 30 35 1.08465 $w=4.23e-07 $l=4e-08 $layer=LI1_cond $X=3.782 $Y=0.89
+ $X2=3.782 $Y2=0.85
r60 29 30 17.49 $w=4.23e-07 $l=6.45e-07 $layer=LI1_cond $X=3.782 $Y=1.535
+ $X2=3.782 $Y2=0.89
r61 26 28 4.38803 $w=3.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.58 $Y=0.68
+ $X2=2.675 $Y2=0.68
r62 21 30 3.61955 $w=3.47e-07 $l=2.30434e-07 $layer=LI1_cond $X=3.5 $Y=0.615
+ $X2=3.68 $Y2=0.73
r63 21 23 8.3232 $w=2.68e-07 $l=1.95e-07 $layer=LI1_cond $X=3.5 $Y=0.615 $X2=3.5
+ $Y2=0.42
r64 19 30 2.86291 $w=2.3e-07 $l=3.15e-07 $layer=LI1_cond $X=3.365 $Y=0.73
+ $X2=3.68 $Y2=0.73
r65 19 28 34.5733 $w=2.28e-07 $l=6.9e-07 $layer=LI1_cond $X=3.365 $Y=0.73
+ $X2=2.675 $Y2=0.73
r66 15 18 61.9786 $w=1.68e-07 $l=9.5e-07 $layer=LI1_cond $X=2.59 $Y=1.62
+ $X2=3.54 $Y2=1.62
r67 13 29 8.58847 $w=1.7e-07 $l=2.50926e-07 $layer=LI1_cond $X=3.57 $Y=1.62
+ $X2=3.782 $Y2=1.535
r68 13 18 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=3.57 $Y=1.62 $X2=3.54
+ $Y2=1.62
r69 4 18 600 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=3.39
+ $Y=1.485 $X2=3.54 $Y2=1.62
r70 3 15 600 $w=1.7e-07 $l=2.17256e-07 $layer=licon1_PDIFF $count=1 $X=2.43
+ $Y=1.485 $X2=2.59 $Y2=1.62
r71 2 30 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.235 $X2=3.54 $Y2=0.76
r72 2 23 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=3.35
+ $Y=0.235 $X2=3.54 $Y2=0.42
r73 1 26 182 $w=1.7e-07 $l=5.31578e-07 $layer=licon1_NDIFF $count=1 $X=2.39
+ $Y=0.235 $X2=2.58 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_4%VGND 1 2 3 12 16 18 20 28 33 40 41 44 47
+ 51
c75 28 0 8.37355e-20 $X=2.845 $Y=0
r76 51 54 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.995 $Y=0 $X2=3.995
+ $Y2=0.36
r77 51 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r78 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r79 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r80 41 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=3.91
+ $Y2=0
r81 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r82 38 51 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=3.995
+ $Y2=0
r83 38 40 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.83
+ $Y2=0
r84 37 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r85 37 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r86 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r87 34 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=3.195 $Y=0 $X2=3.02
+ $Y2=0
r88 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.195 $Y=0 $X2=3.45
+ $Y2=0
r89 33 51 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.995
+ $Y2=0
r90 33 36 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=3.805 $Y=0 $X2=3.45
+ $Y2=0
r91 32 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r92 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r93 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r94 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.095
+ $Y2=0
r95 29 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=2.26 $Y=0 $X2=2.53
+ $Y2=0
r96 28 47 8.9695 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=3.02
+ $Y2=0
r97 28 31 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.845 $Y=0 $X2=2.53
+ $Y2=0
r98 27 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r99 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r100 22 26 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=1.61
+ $Y2=0
r101 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=2.095
+ $Y2=0
r102 20 26 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=1.93 $Y=0 $X2=1.61
+ $Y2=0
r103 18 27 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.61 $Y2=0
r104 18 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r105 14 47 1.07557 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.02 $Y=0.085
+ $X2=3.02 $Y2=0
r106 14 16 9.05491 $w=3.48e-07 $l=2.75e-07 $layer=LI1_cond $X=3.02 $Y=0.085
+ $X2=3.02 $Y2=0.36
r107 10 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0
r108 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.095 $Y=0.085
+ $X2=2.095 $Y2=0.36
r109 3 54 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.88
+ $Y=0.235 $X2=4.02 $Y2=0.36
r110 2 16 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=2.87
+ $Y=0.235 $X2=3.03 $Y2=0.36
r111 1 12 182 $w=1.7e-07 $l=3.36749e-07 $layer=licon1_NDIFF $count=1 $X=1.815
+ $Y=0.235 $X2=2.095 $Y2=0.36
.ends

