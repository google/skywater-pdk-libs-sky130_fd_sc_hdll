* File: sky130_fd_sc_hdll__probec_p_8.pex.spice
* Created: Wed Sep  2 08:50:19 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A 1 3 6 8 10 13 17 19 21 22 32 34
c86 34 0 4.1351e-20 $X=1.41 $Y=1.212
c87 13 0 5.2712e-21 $X=0.99 $Y=0.56
c88 8 0 8.78971e-21 $X=0.965 $Y=1.41
r89 34 35 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.212
+ $X2=1.435 $Y2=1.212
r90 33 34 62.4815 $w=3.24e-07 $l=4.2e-07 $layer=POLY_cond $X=0.99 $Y=1.212
+ $X2=1.41 $Y2=1.212
r91 31 33 0.743827 $w=3.24e-07 $l=5e-09 $layer=POLY_cond $X=0.985 $Y=1.212
+ $X2=0.99 $Y2=1.212
r92 31 32 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r93 29 31 2.97531 $w=3.24e-07 $l=2e-08 $layer=POLY_cond $X=0.965 $Y=1.212
+ $X2=0.985 $Y2=1.212
r94 28 29 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.212
+ $X2=0.965 $Y2=1.212
r95 27 28 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r96 25 27 28.2654 $w=3.24e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.212
+ $X2=0.495 $Y2=1.212
r97 25 26 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=0.305
+ $Y=1.16 $X2=0.305 $Y2=1.16
r98 22 32 16.0818 $w=1.98e-07 $l=2.9e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.985 $Y2=1.175
r99 22 26 21.6273 $w=1.98e-07 $l=3.9e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=0.305 $Y2=1.175
r100 19 35 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r101 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r102 15 34 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.212
r103 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r104 11 33 20.7868 $w=1.5e-07 $l=1.87e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=1.212
r105 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.99 $Y=1.025
+ $X2=0.99 $Y2=0.56
r106 8 29 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.212
r107 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r108 4 28 20.7868 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r109 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r110 1 27 16.5046 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r111 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_27_47# 1 2 3 4 13 15 18 22 24 26 27
+ 29 32 36 38 40 41 43 46 50 52 54 55 57 60 64 66 68 71 77 79 80 81 82 85 91 94
+ 96 102 106 109 111 128
c288 128 0 6.43277e-20 $X=5.17 $Y=1.217
c289 106 0 2.87386e-20 $X=1.507 $Y=1.53
c290 55 0 8.5977e-20 $X=4.725 $Y=1.41
c291 38 0 1.23615e-19 $X=3.315 $Y=1.41
c292 24 0 2.00692e-20 $X=2.375 $Y=1.41
c293 22 0 4.02009e-21 $X=2.35 $Y=0.56
c294 13 0 2.00692e-20 $X=1.905 $Y=1.41
r295 128 129 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r296 127 128 62.8696 $w=3.22e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.217
+ $X2=5.17 $Y2=1.217
r297 126 127 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.217
+ $X2=4.75 $Y2=1.217
r298 125 126 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.725 $Y2=1.217
r299 124 125 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r300 121 122 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=3.81 $Y2=1.217
r301 120 121 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=3.315 $Y=1.217
+ $X2=3.785 $Y2=1.217
r302 119 120 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r303 118 119 62.8696 $w=3.22e-07 $l=4.2e-07 $layer=POLY_cond $X=2.87 $Y=1.217
+ $X2=3.29 $Y2=1.217
r304 117 118 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=2.87 $Y2=1.217
r305 116 117 70.354 $w=3.22e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.845 $Y2=1.217
r306 115 116 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r307 112 113 3.74224 $w=3.22e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r308 103 124 52.3913 $w=3.22e-07 $l=3.5e-07 $layer=POLY_cond $X=3.88 $Y=1.217
+ $X2=4.23 $Y2=1.217
r309 103 122 10.4783 $w=3.22e-07 $l=7e-08 $layer=POLY_cond $X=3.88 $Y=1.217
+ $X2=3.81 $Y2=1.217
r310 102 103 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r311 100 115 25.4472 $w=3.22e-07 $l=1.7e-07 $layer=POLY_cond $X=2.18 $Y=1.217
+ $X2=2.35 $Y2=1.217
r312 100 113 37.4224 $w=3.22e-07 $l=2.5e-07 $layer=POLY_cond $X=2.18 $Y=1.217
+ $X2=1.93 $Y2=1.217
r313 99 102 110.909 $w=1.68e-07 $l=1.7e-06 $layer=LI1_cond $X=2.18 $Y=1.16
+ $X2=3.88 $Y2=1.16
r314 99 100 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.18
+ $Y=1.16 $X2=2.18 $Y2=1.16
r315 97 111 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=1.507 $Y2=1.16
r316 97 99 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=1.595 $Y=1.16
+ $X2=2.18 $Y2=1.16
r317 96 106 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.445
+ $X2=1.507 $Y2=1.53
r318 95 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.16
r319 95 96 12.6753 $w=1.73e-07 $l=2e-07 $layer=LI1_cond $X=1.507 $Y=1.245
+ $X2=1.507 $Y2=1.445
r320 94 111 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=1.075
+ $X2=1.507 $Y2=1.16
r321 93 109 0.574824 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=0.82
r322 93 94 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=1.507 $Y=0.905
+ $X2=1.507 $Y2=1.075
r323 89 109 20.0289 $w=1.68e-07 $l=3.07e-07 $layer=LI1_cond $X=1.2 $Y=0.82
+ $X2=1.507 $Y2=0.82
r324 89 91 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=0.735
+ $X2=1.2 $Y2=0.42
r325 85 87 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=1.2 $Y=1.63 $X2=1.2
+ $Y2=2.31
r326 83 106 20.0289 $w=1.68e-07 $l=3.07e-07 $layer=LI1_cond $X=1.2 $Y=1.53
+ $X2=1.507 $Y2=1.53
r327 83 85 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.2 $Y=1.615
+ $X2=1.2 $Y2=1.63
r328 81 89 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=1.2 $Y2=0.82
r329 81 82 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.065 $Y=0.82
+ $X2=0.445 $Y2=0.82
r330 79 83 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=1.2 $Y2=1.53
r331 79 80 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=1.53
+ $X2=0.425 $Y2=1.53
r332 75 82 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=0.295 $Y=0.735
+ $X2=0.445 $Y2=0.82
r333 75 77 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=0.295 $Y=0.735
+ $X2=0.295 $Y2=0.42
r334 71 73 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.63
+ $X2=0.26 $Y2=2.31
r335 69 80 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.425 $Y2=1.53
r336 69 71 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=0.26 $Y=1.615
+ $X2=0.26 $Y2=1.63
r337 66 129 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r338 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r339 62 128 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r340 62 64 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r341 58 127 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=1.217
r342 58 60 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.75 $Y=1.025
+ $X2=4.75 $Y2=0.56
r343 55 126 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r344 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r345 52 125 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r346 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r347 48 124 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r348 48 50 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
r349 44 122 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r350 44 46 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r351 41 121 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r352 41 43 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r353 38 120 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r354 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r355 34 119 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r356 34 36 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r357 30 118 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r358 30 32 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r359 27 117 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r360 27 29 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r361 24 116 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r362 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r363 20 115 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r364 20 22 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r365 16 113 20.6399 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r366 16 18 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r367 13 112 16.3606 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r368 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r369 4 87 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.31
r370 4 85 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r371 3 73 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.31
r372 3 71 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.63
r373 2 91 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.42
r374 1 77 91 $w=1.7e-07 $l=2.5807e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VPWR 1 2 3 4 5 6 21 23 27 29 33 35 39
+ 41 45 49 54 55 56 58 61 69 74 85 89 92 95 98 101 113
c125 69 0 6.43277e-20 $X=4.46 $Y=2.875
c126 61 0 2.5603e-19 $X=5.72 $Y=2.72
c127 2 0 1.8139e-19 $X=1.525 $Y=1.485
r128 113 114 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=5.68 $Y=2.72
+ $X2=5.68 $Y2=2.72
r129 101 102 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r130 99 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r131 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r132 96 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r133 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r134 93 96 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r135 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r136 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r137 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r138 85 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r139 83 113 0.110971 $w=4.8e-07 $l=3.9e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.68 $Y2=2.72
r140 83 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r141 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r142 80 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=4.49 $Y2=2.72
r143 80 82 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=2.72
+ $X2=5.29 $Y2=2.72
r144 74 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.73 $Y2=2.72
r145 66 69 0.0160563 $w=1.704e-06 $l=9.6e-07 $layer=MET5_cond $X=5.52 $Y=3.025
+ $X2=4.56 $Y2=3.025
r146 65 66 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=5.52 $Y=3.025
+ $X2=5.52 $Y2=3.025
r147 62 114 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=5.72 $Y=2.72
+ $X2=5.72 $Y2=2.72
r148 61 65 0.0123962 $w=1.18e-06 $l=3.05e-07 $layer=MET4_cond $X=5.52 $Y=2.72
+ $X2=5.52 $Y2=3.025
r149 61 62 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=5.72 $Y=2.72
+ $X2=5.72 $Y2=2.72
r150 58 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 56 74 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.595 $Y2=2.72
r152 56 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r153 54 82 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.29 $Y2=2.72
r154 54 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.295 $Y=2.72
+ $X2=5.445 $Y2=2.72
r155 53 85 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.75 $Y2=2.72
r156 53 55 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.595 $Y=2.72
+ $X2=5.445 $Y2=2.72
r157 49 52 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=5.445 $Y=1.66
+ $X2=5.445 $Y2=2.34
r158 47 55 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.72
r159 47 52 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.445 $Y=2.635
+ $X2=5.445 $Y2=2.34
r160 43 101 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2.72
r161 43 45 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.49 $Y=2.635
+ $X2=4.49 $Y2=2
r162 42 98 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=2.72
+ $X2=3.55 $Y2=2.72
r163 41 101 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=4.49 $Y2=2.72
r164 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=2.72
+ $X2=3.685 $Y2=2.72
r165 37 98 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2.72
r166 37 39 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.55 $Y=2.635
+ $X2=3.55 $Y2=2
r167 36 95 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=2.72
+ $X2=2.61 $Y2=2.72
r168 35 98 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=3.55 $Y2=2.72
r169 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=2.72
+ $X2=2.745 $Y2=2.72
r170 31 95 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2.72
r171 31 33 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.61 $Y=2.635
+ $X2=2.61 $Y2=2
r172 30 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=2.72
+ $X2=1.67 $Y2=2.72
r173 29 95 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=2.61 $Y2=2.72
r174 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=2.72
+ $X2=1.805 $Y2=2.72
r175 25 92 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2.72
r176 25 27 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.67 $Y=2.635
+ $X2=1.67 $Y2=2
r177 24 89 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=2.72
+ $X2=0.73 $Y2=2.72
r178 23 92 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=1.67 $Y2=2.72
r179 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=2.72
+ $X2=0.865 $Y2=2.72
r180 19 89 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r181 19 21 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2
r182 6 52 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r183 6 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r184 5 45 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2
r185 4 39 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2
r186 3 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2
r187 2 27 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2
r188 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%A_399_297# 1 2 3 4 5 6 7 8 27 31 33 34
+ 35 36 39 43 45 47 51 55 59 63 65 66 67 68 69 71 74 76 77 80 82 87 93
c239 93 0 1.32773e-19 $X=2.475 $Y=1.19
c240 80 0 1.1937e-20 $X=2.475 $Y=1.19
c241 77 0 1.67773e-19 $X=2.05 $Y=1.36
c242 76 0 1.95451e-19 $X=2.05 $Y=1.36
c243 74 0 1.42241e-19 $X=2.53 $Y=1.19
c244 68 0 1.26775e-19 $X=2.66 $Y=1.19
c245 8 0 1.70053e-19 $X=4.815 $Y=1.485
c246 4 0 1.70053e-19 $X=4.825 $Y=0.235
r247 89 93 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=2.5 $Y=1.19 $X2=2.5
+ $Y2=1.19
r248 80 93 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=2.475 $Y=1.19
+ $X2=2.475 $Y2=1.19
r249 77 82 0.0191979 $w=4.93e-06 $l=8.9e-07 $layer=MET5_cond $X=2.05 $Y=1.36
+ $X2=1.16 $Y2=1.36
r250 76 80 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=2.475 $Y=1.19
+ $X2=2.475 $Y2=1.19
r251 76 77 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=2.05 $Y=1.36
+ $X2=2.05 $Y2=1.36
r252 74 89 0.0170272 $w=2.6e-07 $l=3e-08 $layer=MET1_cond $X=2.53 $Y=1.19
+ $X2=2.5 $Y2=1.19
r253 72 87 3.68633 $w=6.95e-07 $l=2.1e-07 $layer=LI1_cond $X=4.75 $Y=1.175
+ $X2=4.96 $Y2=1.175
r254 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.75 $Y=1.19
+ $X2=4.75 $Y2=1.19
r255 69 71 0.250226 $w=2.3e-07 $l=3.9e-07 $layer=MET1_cond $X=4.36 $Y=1.19
+ $X2=4.75 $Y2=1.19
r256 68 74 0.089401 $w=2.6e-07 $l=1.3e-07 $layer=MET1_cond $X=2.66 $Y=1.19
+ $X2=2.53 $Y2=1.19
r257 67 69 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=4.245 $Y=1.19
+ $X2=4.36 $Y2=1.19
r258 67 68 1.96163 $w=1.4e-07 $l=1.585e-06 $layer=MET1_cond $X=4.245 $Y=1.19
+ $X2=2.66 $Y2=1.19
r259 61 87 5.10968 $w=3.3e-07 $l=4.4e-07 $layer=LI1_cond $X=4.96 $Y=1.615
+ $X2=4.96 $Y2=1.175
r260 61 63 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.96 $Y=1.615
+ $X2=4.96 $Y2=1.755
r261 57 87 5.10968 $w=3.3e-07 $l=4.4e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.96 $Y2=1.175
r262 57 59 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.96 $Y=0.735
+ $X2=4.96 $Y2=0.42
r263 53 55 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=4.02 $Y=1.615
+ $X2=4.02 $Y2=1.755
r264 49 72 12.8144 $w=6.95e-07 $l=9.24175e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.75 $Y2=1.175
r265 49 53 5.10968 $w=3.3e-07 $l=8.8e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=1.615
r266 49 51 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.02 $Y=0.735
+ $X2=4.02 $Y2=0.42
r267 48 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=1.53
+ $X2=3.08 $Y2=1.53
r268 47 49 6.53734 $w=3.47e-07 $l=8.73613e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=4.02 $Y2=0.735
r269 47 48 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=1.53
+ $X2=3.245 $Y2=1.53
r270 46 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0.82
+ $X2=3.08 $Y2=0.82
r271 45 49 6.53734 $w=3.47e-07 $l=2.03101e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=4.02 $Y2=0.735
r272 45 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0.82
+ $X2=3.245 $Y2=0.82
r273 41 66 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.53
r274 41 43 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=3.08 $Y=1.615
+ $X2=3.08 $Y2=1.755
r275 37 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.82
r276 37 39 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=3.08 $Y=0.735
+ $X2=3.08 $Y2=0.42
r277 35 66 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=1.53
+ $X2=3.08 $Y2=1.53
r278 35 36 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=1.53
+ $X2=2.305 $Y2=1.53
r279 33 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=3.08 $Y2=0.82
r280 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.82
+ $X2=2.305 $Y2=0.82
r281 29 36 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.305 $Y2=1.53
r282 29 31 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=2.14 $Y=1.615
+ $X2=2.14 $Y2=1.755
r283 25 34 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.305 $Y2=0.82
r284 25 27 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.14 $Y2=0.42
r285 8 63 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.755
r286 7 55 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.755
r287 6 43 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.755
r288 5 31 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.755
r289 4 59 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.42
r290 3 51 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.42
r291 2 39 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.42
r292 1 27 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%VGND 1 2 3 4 5 6 21 25 27 31 33 37 39
+ 43 47 50 51 52 54 57 64 69 79 82 84 87 90 93 96 99 103 114
c140 57 0 1.70053e-19 $X=5.52 $Y=-0.304
r141 114 115 2.25 $w=1.5e-07 $l=3e-07 $layer=via $count=2 $X=5.68 $Y=0 $X2=5.68
+ $Y2=0
r142 96 97 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r143 94 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r144 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r145 91 94 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r146 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r147 88 91 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r148 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r149 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r150 82 84 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.615 $Y=0 $X2=0.755
+ $Y2=0
r151 79 114 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r152 77 114 0.110971 $w=4.8e-07 $l=3.9e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.68 $Y2=0
r153 77 97 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r154 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r155 74 96 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.49
+ $Y2=0
r156 74 76 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r157 73 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r158 73 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r159 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r160 70 84 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.755
+ $Y2=0
r161 70 72 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r162 69 87 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.655
+ $Y2=0
r163 69 72 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.505 $Y=0
+ $X2=1.15 $Y2=0
r164 61 115 1.705 $w=2e-07 $l=4e-07 $layer=via2 $count=2 $X=5.72 $Y=0 $X2=5.72
+ $Y2=0
r165 58 64 0.0160563 $w=1.704e-06 $l=9.6e-07 $layer=MET5_cond $X=5.52 $Y=-0.305
+ $X2=4.56 $Y2=-0.305
r166 57 61 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=5.72 $Y=0
+ $X2=5.72 $Y2=0
r167 57 58 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=5.52
+ $Y=-0.304 $X2=5.52 $Y2=-0.304
r168 54 85 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r169 54 103 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r170 52 82 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=0.235 $Y=0
+ $X2=0.615 $Y2=0
r171 52 99 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r172 50 76 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.29
+ $Y2=0
r173 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.42
+ $Y2=0
r174 49 79 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.75 $Y2=0
r175 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.545 $Y=0 $X2=5.42
+ $Y2=0
r176 45 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0
r177 45 47 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.42 $Y=0.085
+ $X2=5.42 $Y2=0.38
r178 41 96 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r179 41 43 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.4
r180 40 93 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.55
+ $Y2=0
r181 39 96 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.49
+ $Y2=0
r182 39 40 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=3.685 $Y2=0
r183 35 93 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r184 35 37 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.4
r185 34 90 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.61
+ $Y2=0
r186 33 93 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.55
+ $Y2=0
r187 33 34 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=2.745 $Y2=0
r188 29 90 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r189 29 31 13.4452 $w=2.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.4
r190 28 87 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.655
+ $Y2=0
r191 27 90 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.61
+ $Y2=0
r192 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.805 $Y2=0
r193 23 87 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0
r194 23 25 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=1.655 $Y=0.085
+ $X2=1.655 $Y2=0.4
r195 19 84 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0
r196 19 21 12.965 $w=2.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.755 $Y=0.085
+ $X2=0.755 $Y2=0.4
r197 6 47 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.245
+ $Y=0.235 $X2=5.38 $Y2=0.38
r198 5 43 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.4
r199 4 37 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
r200 3 31 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r201 2 25 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.4
r202 1 21 182 $w=1.7e-07 $l=2.33345e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.76 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__PROBEC_P_8%X 1 4 8 10
c37 10 0 2.87386e-20 $X=1.06 $Y=1.36
r38 5 10 0.0302819 $w=1.6e-06 $l=1.609e-06 $layer=MET5_cond $X=-0.549 $Y=1.36
+ $X2=1.06 $Y2=1.36
r39 4 8 1.705 $w=2e-07 $l=4e-07 $layer=via3_notcapm $count=2 $X=-0.124 $Y=1.19
+ $X2=-0.124 $Y2=1.19
r40 4 5 0.38 $w=8e-07 $l=8e-07 $layer=via4_notcap2m $count=1 $X=-0.549 $Y=1.36
+ $X2=-0.549 $Y2=1.36
r41 1 8 0.033007 $w=3.2e-07 $l=2.06e-07 $layer=MET3_cond $X=-0.33 $Y=1.19
+ $X2=-0.124 $Y2=1.19
.ends

