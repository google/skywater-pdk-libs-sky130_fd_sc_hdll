* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 a_276_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=1.95e+11p pd=1.9e+06u as=6.045e+11p ps=4.46e+06u
M1001 VPWR a_93_21# X VPB phighvt w=1e+06u l=180000u
+  ad=9.75e+11p pd=5.95e+06u as=3.4e+11p ps=2.68e+06u
M1002 a_93_21# B1 a_268_297# VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=1.015e+12p ps=8.03e+06u
M1003 a_93_21# A1 a_366_47# VNB nshort w=650000u l=150000u
+  ad=3.185e+11p pd=2.28e+06u as=3.575e+11p ps=2.4e+06u
M1004 a_366_47# A2 a_276_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_93_21# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.145e+11p ps=1.96e+06u
M1006 a_634_47# B1 a_93_21# VNB nshort w=650000u l=150000u
+  ad=1.365e+11p pd=1.72e+06u as=0p ps=0u
M1007 VPWR A2 a_268_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_268_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_268_297# A3 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_268_297# B2 a_93_21# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND B2 a_634_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
