* File: sky130_fd_sc_hdll__or3_1.pxi.spice
* Created: Thu Aug 27 19:24:05 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR3_1%C N_C_c_56_n N_C_M1002_g N_C_M1001_g C N_C_c_55_n
+ PM_SKY130_FD_SC_HDLL__OR3_1%C
x_PM_SKY130_FD_SC_HDLL__OR3_1%B N_B_c_81_n N_B_c_82_n N_B_c_84_n N_B_c_85_n
+ N_B_M1006_g N_B_M1007_g N_B_c_83_n B B N_B_c_87_n B
+ PM_SKY130_FD_SC_HDLL__OR3_1%B
x_PM_SKY130_FD_SC_HDLL__OR3_1%A N_A_c_123_n N_A_M1003_g N_A_M1005_g A A A
+ N_A_c_125_n N_A_c_126_n A PM_SKY130_FD_SC_HDLL__OR3_1%A
x_PM_SKY130_FD_SC_HDLL__OR3_1%A_29_53# N_A_29_53#_M1001_s N_A_29_53#_M1007_d
+ N_A_29_53#_M1002_s N_A_29_53#_c_173_n N_A_29_53#_M1000_g N_A_29_53#_c_174_n
+ N_A_29_53#_M1004_g N_A_29_53#_c_175_n N_A_29_53#_c_176_n N_A_29_53#_c_177_n
+ N_A_29_53#_c_182_n N_A_29_53#_c_247_p N_A_29_53#_c_178_n N_A_29_53#_c_215_n
+ N_A_29_53#_c_179_n N_A_29_53#_c_184_n N_A_29_53#_c_180_n N_A_29_53#_c_185_n
+ PM_SKY130_FD_SC_HDLL__OR3_1%A_29_53#
x_PM_SKY130_FD_SC_HDLL__OR3_1%VPWR N_VPWR_M1003_d N_VPWR_c_269_n VPWR
+ N_VPWR_c_270_n N_VPWR_c_271_n N_VPWR_c_268_n N_VPWR_c_273_n VPWR
+ PM_SKY130_FD_SC_HDLL__OR3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR3_1%X N_X_M1004_d N_X_M1000_d N_X_c_292_n N_X_c_294_n
+ N_X_c_293_n X PM_SKY130_FD_SC_HDLL__OR3_1%X
x_PM_SKY130_FD_SC_HDLL__OR3_1%VGND N_VGND_M1001_d N_VGND_M1005_d N_VGND_c_311_n
+ VGND N_VGND_c_312_n N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n
+ N_VGND_c_316_n N_VGND_c_317_n VGND PM_SKY130_FD_SC_HDLL__OR3_1%VGND
cc_1 VNB N_C_M1001_g 0.0344462f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.475
cc_2 VNB C 0.0123316f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_C_c_55_n 0.0362629f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_4 VNB N_B_c_81_n 0.00672106f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_5 VNB N_B_c_82_n 0.0216796f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.695
cc_6 VNB N_B_c_83_n 0.0143238f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_7 VNB N_A_c_123_n 0.0209385f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.41
cc_8 VNB N_A_M1005_g 0.0285191f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.475
cc_9 VNB N_A_c_125_n 0.00227398f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_126_n 0.00244293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_29_53#_c_173_n 0.0294189f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.202
cc_12 VNB N_A_29_53#_c_174_n 0.0207304f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_13 VNB N_A_29_53#_c_175_n 0.0135183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_29_53#_c_176_n 0.00360508f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_29_53#_c_177_n 0.00942926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_29_53#_c_178_n 0.00172906f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_29_53#_c_179_n 0.00113231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_29_53#_c_180_n 0.00154117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_268_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_292_n 0.013635f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_21 VNB N_X_c_293_n 0.025699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_311_n 0.0010436f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_312_n 0.0151077f $X=-0.19 $Y=-0.24 $X2=0.505 $Y2=1.202
cc_24 VNB N_VGND_c_313_n 0.0129653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_314_n 0.0274657f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_315_n 0.171023f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_316_n 0.00544933f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_317_n 0.0102719f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_C_c_56_n 0.0204874f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_30 VPB C 0.00162495f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_31 VPB N_C_c_55_n 0.0165533f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.202
cc_32 VPB N_B_c_84_n 0.0056146f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.695
cc_33 VPB N_B_c_85_n 0.0482502f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_34 VPB N_B_M1006_g 0.0107354f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.475
cc_35 VPB N_B_c_87_n 0.0377963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_c_123_n 0.0273735f $X=-0.19 $Y=1.305 $X2=0.505 $Y2=1.41
cc_37 VPB A 0.00169108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_c_125_n 0.00313301f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_29_53#_c_173_n 0.0331655f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_40 VPB N_A_29_53#_c_182_n 0.0033481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_29_53#_c_179_n 0.00165371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_29_53#_c_184_n 0.0209087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_29_53#_c_185_n 0.00139636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_269_n 0.0129433f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.475
cc_45 VPB N_VPWR_c_270_n 0.0419151f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.202
cc_46 VPB N_VPWR_c_271_n 0.0277375f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_268_n 0.061976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_273_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_X_c_294_n 0.00521594f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.202
cc_50 VPB N_X_c_293_n 0.00936334f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB X 0.0319967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 N_C_M1001_g N_B_c_81_n 0.0199009f $X=0.53 $Y=0.475 $X2=-0.19 $Y2=-0.24
cc_53 C N_B_c_82_n 2.18655e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_54 N_C_c_55_n N_B_c_82_n 0.0199009f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_55 N_C_c_56_n N_B_M1006_g 0.033095f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_56 N_C_M1001_g N_B_c_83_n 0.0137274f $X=0.53 $Y=0.475 $X2=0 $Y2=0
cc_57 N_C_c_56_n N_B_c_87_n 0.00528921f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_58 N_C_c_56_n A 0.00251338f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_59 N_C_c_55_n A 0.00224594f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_60 C N_A_c_126_n 0.0257891f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_61 N_C_c_55_n N_A_c_126_n 0.00316301f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_62 N_C_M1001_g N_A_29_53#_c_176_n 0.0167603f $X=0.53 $Y=0.475 $X2=0 $Y2=0
cc_63 C N_A_29_53#_c_176_n 0.00559912f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_64 N_C_c_55_n N_A_29_53#_c_176_n 0.00278696f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_65 C N_A_29_53#_c_177_n 0.0211211f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_66 N_C_c_55_n N_A_29_53#_c_177_n 0.00542346f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_67 N_C_c_56_n N_A_29_53#_c_182_n 0.0133471f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_68 N_C_c_56_n N_A_29_53#_c_184_n 0.00674133f $X=0.505 $Y=1.41 $X2=0 $Y2=0
cc_69 C N_A_29_53#_c_184_n 0.023487f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_70 N_C_c_55_n N_A_29_53#_c_184_n 0.00642559f $X=0.505 $Y=1.202 $X2=0 $Y2=0
cc_71 N_C_M1001_g N_VGND_c_311_n 0.0124902f $X=0.53 $Y=0.475 $X2=0 $Y2=0
cc_72 N_C_M1001_g N_VGND_c_312_n 0.00187556f $X=0.53 $Y=0.475 $X2=0 $Y2=0
cc_73 N_C_M1001_g N_VGND_c_315_n 0.00330947f $X=0.53 $Y=0.475 $X2=0 $Y2=0
cc_74 N_B_c_82_n N_A_c_123_n 0.0176216f $X=0.925 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_75 N_B_c_84_n N_A_c_123_n 0.00357417f $X=0.925 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_76 N_B_M1006_g N_A_c_123_n 0.0215164f $X=0.925 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_77 N_B_c_87_n N_A_c_123_n 6.03833e-19 $X=0.99 $Y=2.28 $X2=-0.19 $Y2=-0.24
cc_78 N_B_c_83_n N_A_M1005_g 0.0166388f $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_79 N_B_c_84_n A 0.00236103f $X=0.925 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B_M1006_g A 0.00502076f $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_81 N_B_c_82_n N_A_c_125_n 0.0110177f $X=0.925 $Y=1.31 $X2=0 $Y2=0
cc_82 N_B_c_84_n N_A_c_125_n 0.00464961f $X=0.925 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_82_n N_A_c_126_n 0.0037757f $X=0.925 $Y=1.31 $X2=0 $Y2=0
cc_84 N_B_c_81_n N_A_29_53#_c_176_n 0.00629366f $X=0.925 $Y=0.86 $X2=0 $Y2=0
cc_85 N_B_c_83_n N_A_29_53#_c_176_n 0.00713678f $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_86 N_B_c_85_n N_A_29_53#_c_182_n 0.00111426f $X=0.925 $Y=2.035 $X2=0 $Y2=0
cc_87 N_B_M1006_g N_A_29_53#_c_182_n 0.0127838f $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_88 N_B_c_87_n N_A_29_53#_c_182_n 0.0569078f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_89 N_B_M1006_g N_A_29_53#_c_184_n 9.46988e-19 $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_90 N_B_c_87_n N_A_29_53#_c_184_n 0.026488f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_91 N_B_M1006_g N_A_29_53#_c_185_n 0.00473678f $X=0.925 $Y=1.695 $X2=0 $Y2=0
cc_92 N_B_c_87_n N_A_29_53#_c_185_n 0.0137296f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_93 N_B_c_85_n N_VPWR_c_269_n 0.00350614f $X=0.925 $Y=2.035 $X2=0 $Y2=0
cc_94 N_B_c_87_n N_VPWR_c_269_n 0.0210032f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_95 N_B_c_85_n N_VPWR_c_270_n 0.00753055f $X=0.925 $Y=2.035 $X2=0 $Y2=0
cc_96 N_B_c_87_n N_VPWR_c_270_n 0.0647515f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_97 N_B_c_85_n N_VPWR_c_268_n 0.0107919f $X=0.925 $Y=2.035 $X2=0 $Y2=0
cc_98 N_B_c_87_n N_VPWR_c_268_n 0.0469974f $X=0.99 $Y=2.28 $X2=0 $Y2=0
cc_99 N_B_c_83_n N_VGND_c_311_n 0.00720367f $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_100 N_B_c_83_n N_VGND_c_313_n 0.00322006f $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_101 N_B_c_83_n N_VGND_c_315_n 0.00408297f $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_102 N_B_c_83_n N_VGND_c_317_n 5.53035e-19 $X=0.925 $Y=0.76 $X2=0 $Y2=0
cc_103 N_A_c_123_n N_A_29_53#_c_173_n 0.0392073f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_125_n N_A_29_53#_c_173_n 0.00108448f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_M1005_g N_A_29_53#_c_174_n 0.0191905f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_106 N_A_c_125_n N_A_29_53#_c_176_n 0.0207076f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A_c_126_n N_A_29_53#_c_176_n 0.0199527f $X=0.725 $Y=1.325 $X2=0 $Y2=0
cc_108 N_A_c_123_n N_A_29_53#_c_182_n 2.17268e-19 $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_109 A N_A_29_53#_c_182_n 0.0108545f $X=0.65 $Y=1.445 $X2=0 $Y2=0
cc_110 N_A_c_125_n N_A_29_53#_c_182_n 0.0116476f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_c_123_n N_A_29_53#_c_178_n 0.00240831f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_M1005_g N_A_29_53#_c_178_n 0.0127189f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_113 N_A_c_125_n N_A_29_53#_c_178_n 0.0142622f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_c_123_n N_A_29_53#_c_215_n 0.0147956f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_c_125_n N_A_29_53#_c_215_n 0.00821244f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_116 N_A_c_123_n N_A_29_53#_c_179_n 0.00433378f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_M1005_g N_A_29_53#_c_179_n 0.00329784f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_118 N_A_c_125_n N_A_29_53#_c_179_n 0.015218f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_119 N_A_c_123_n N_A_29_53#_c_180_n 5.77159e-19 $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_c_125_n N_A_29_53#_c_180_n 0.0146254f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_c_123_n N_A_29_53#_c_185_n 0.0113899f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_122 A N_A_29_53#_c_185_n 0.00485635f $X=0.65 $Y=1.445 $X2=0 $Y2=0
cc_123 N_A_c_125_n N_A_29_53#_c_185_n 0.0112473f $X=1.405 $Y=1.16 $X2=0 $Y2=0
cc_124 A A_119_297# 0.00139384f $X=0.65 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_125 N_A_c_123_n N_VPWR_c_269_n 0.00330158f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_c_123_n N_VPWR_c_270_n 0.00351268f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_c_123_n N_VPWR_c_268_n 0.00445321f $X=1.445 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_VGND_c_311_n 5.02092e-19 $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_129 N_A_M1005_g N_VGND_c_313_n 0.00188229f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_130 N_A_M1005_g N_VGND_c_315_n 0.00270076f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_131 N_A_M1005_g N_VGND_c_317_n 0.01011f $X=1.47 $Y=0.475 $X2=0 $Y2=0
cc_132 N_A_29_53#_c_182_n A_119_297# 0.0013394f $X=1.205 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_29_53#_c_182_n A_203_297# 0.00258366f $X=1.205 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_134 N_A_29_53#_c_185_n A_203_297# 0.00459651f $X=1.29 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_29_53#_c_215_n N_VPWR_M1003_d 0.00651861f $X=1.805 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_136 N_A_29_53#_c_173_n N_VPWR_c_269_n 0.00512739f $X=1.985 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_29_53#_c_215_n N_VPWR_c_269_n 0.0198977f $X=1.805 $Y=1.58 $X2=0 $Y2=0
cc_138 N_A_29_53#_c_185_n N_VPWR_c_269_n 0.00726621f $X=1.29 $Y=1.58 $X2=0 $Y2=0
cc_139 N_A_29_53#_c_173_n N_VPWR_c_271_n 0.00702461f $X=1.985 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_29_53#_c_173_n N_VPWR_c_268_n 0.0148987f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_29_53#_c_174_n N_X_c_292_n 0.00907889f $X=2.01 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_29_53#_c_178_n N_X_c_292_n 0.00469632f $X=1.805 $Y=0.74 $X2=0 $Y2=0
cc_143 N_A_29_53#_c_173_n N_X_c_294_n 0.0222372f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_29_53#_c_215_n N_X_c_294_n 0.00756186f $X=1.805 $Y=1.58 $X2=0 $Y2=0
cc_145 N_A_29_53#_c_173_n N_X_c_293_n 0.001511f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_29_53#_c_174_n N_X_c_293_n 0.0124142f $X=2.01 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_29_53#_c_178_n N_X_c_293_n 0.00230974f $X=1.805 $Y=0.74 $X2=0 $Y2=0
cc_148 N_A_29_53#_c_179_n N_X_c_293_n 0.0222238f $X=1.89 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_29_53#_c_176_n N_VGND_M1001_d 0.00160115f $X=1.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_150 N_A_29_53#_c_178_n N_VGND_M1005_d 0.00650959f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_29_53#_c_179_n N_VGND_M1005_d 7.32946e-19 $X=1.89 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_29_53#_c_175_n N_VGND_c_311_n 0.0138472f $X=0.27 $Y=0.47 $X2=0 $Y2=0
cc_153 N_A_29_53#_c_176_n N_VGND_c_311_n 0.0196541f $X=1.125 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_29_53#_c_247_p N_VGND_c_311_n 0.0110177f $X=1.21 $Y=0.47 $X2=0 $Y2=0
cc_155 N_A_29_53#_c_175_n N_VGND_c_312_n 0.0132481f $X=0.27 $Y=0.47 $X2=0 $Y2=0
cc_156 N_A_29_53#_c_176_n N_VGND_c_312_n 0.0023206f $X=1.125 $Y=0.74 $X2=0 $Y2=0
cc_157 N_A_29_53#_c_176_n N_VGND_c_313_n 0.00310196f $X=1.125 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_A_29_53#_c_247_p N_VGND_c_313_n 0.00876148f $X=1.21 $Y=0.47 $X2=0 $Y2=0
cc_159 N_A_29_53#_c_178_n N_VGND_c_313_n 0.00232988f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_29_53#_c_174_n N_VGND_c_314_n 0.00543382f $X=2.01 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_A_29_53#_c_178_n N_VGND_c_314_n 0.00105918f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_162 N_A_29_53#_c_174_n N_VGND_c_315_n 0.0110827f $X=2.01 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_29_53#_c_175_n N_VGND_c_315_n 0.00942308f $X=0.27 $Y=0.47 $X2=0 $Y2=0
cc_164 N_A_29_53#_c_176_n N_VGND_c_315_n 0.0115456f $X=1.125 $Y=0.74 $X2=0 $Y2=0
cc_165 N_A_29_53#_c_247_p N_VGND_c_315_n 0.00625722f $X=1.21 $Y=0.47 $X2=0 $Y2=0
cc_166 N_A_29_53#_c_178_n N_VGND_c_315_n 0.00843284f $X=1.805 $Y=0.74 $X2=0
+ $Y2=0
cc_167 N_A_29_53#_c_173_n N_VGND_c_317_n 4.00709e-19 $X=1.985 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_29_53#_c_174_n N_VGND_c_317_n 0.00498808f $X=2.01 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_29_53#_c_247_p N_VGND_c_317_n 0.0135697f $X=1.21 $Y=0.47 $X2=0 $Y2=0
cc_170 N_A_29_53#_c_178_n N_VGND_c_317_n 0.0273767f $X=1.805 $Y=0.74 $X2=0 $Y2=0
cc_171 N_VPWR_c_268_n N_X_M1000_d 0.0132621f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_172 N_VPWR_c_271_n X 0.019258f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_173 N_VPWR_c_268_n X 0.0105137f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_174 N_X_c_292_n N_VGND_c_314_n 0.00902248f $X=2.53 $Y=0.587 $X2=0 $Y2=0
cc_175 N_X_M1004_d N_VGND_c_315_n 0.0130032f $X=2.085 $Y=0.235 $X2=0 $Y2=0
cc_176 N_X_c_292_n N_VGND_c_315_n 0.00941771f $X=2.53 $Y=0.587 $X2=0 $Y2=0
