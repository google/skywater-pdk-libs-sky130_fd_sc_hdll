* File: sky130_fd_sc_hdll__o21a_4.spice
* Created: Thu Aug 27 19:19:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21a_4.pex.spice"
.subckt sky130_fd_sc_hdll__o21a_4  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_X_M1005_d N_A_80_21#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.17225 PD=0.98 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1005_d N_A_80_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_A_80_21#_M1009_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1018 N_X_M1009_d N_A_80_21#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_A_525_47#_M1013_d N_B1_M1013_g N_A_80_21#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1015 N_A_525_47#_M1015_d N_B1_M1015_g N_A_80_21#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.147875 AS=0.08775 PD=1.105 PS=0.92 NRD=23.076 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1012 N_A_525_47#_M1015_d N_A1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.147875 AS=0.10075 PD=1.105 PS=0.96 NRD=9.228 NRS=3.684 M=1 R=4.33333
+ SA=75001.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 N_A_525_47#_M1003_d N_A2_M1003_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10075 PD=0.98 PS=0.96 NRD=9.228 NRS=1.836 M=1 R=4.33333
+ SA=75001.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_525_47#_M1003_d N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75002.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1016 N_A_525_47#_M1016_d N_A1_M1016_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.20475 AS=0.10725 PD=1.93 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_A_80_21#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.325 PD=1.3 PS=2.65 NRD=1.9503 NRS=11.8003 M=1 R=5.55556
+ SA=90000.2 SB=90004.8 A=0.18 P=2.36 MULT=1
MM1002 N_X_M1000_d N_A_80_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90004.3 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1010_d N_A_80_21#_M1010_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90003.8 A=0.18 P=2.36 MULT=1
MM1017 N_X_M1010_d N_A_80_21#_M1017_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=1.9503 NRS=5.8903 M=1 R=5.55556 SA=90001.7
+ SB=90003.3 A=0.18 P=2.36 MULT=1
MM1001 N_A_80_21#_M1001_d N_B1_M1001_g N_VPWR_M1017_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.16 PD=1.35 PS=1.32 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90002.2 SB=90002.8 A=0.18 P=2.36 MULT=1
MM1011 N_A_80_21#_M1001_d N_B1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.26 PD=1.35 PS=1.52 NRD=11.8003 NRS=21.67 M=1 R=5.55556
+ SA=90002.7 SB=90002.3 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1011_s N_A1_M1014_g A_826_297# VPB PHIGHVT L=0.18 W=1 AD=0.26
+ AS=0.125 PD=1.52 PS=1.25 NRD=25.5903 NRS=13.7703 M=1 R=5.55556 SA=90003.4
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 A_826_297# N_A2_M1004_g N_A_80_21#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.125 AS=0.15 PD=1.25 PS=1.3 NRD=13.7703 NRS=1.9503 M=1 R=5.55556
+ SA=90003.8 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1019 A_1008_297# N_A2_M1019_g N_A_80_21#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=18.6953 NRS=1.9503 M=1 R=5.55556 SA=90004.3
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A1_M1008_g A_1008_297# VPB PHIGHVT L=0.18 W=1 AD=0.295
+ AS=0.15 PD=2.59 PS=1.3 NRD=1.9503 NRS=18.6953 M=1 R=5.55556 SA=90004.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
c_78 VPB 0 1.79518e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__o21a_4.pxi.spice"
*
.ends
*
*
