* File: sky130_fd_sc_hdll__a32o_2.pex.spice
* Created: Thu Aug 27 18:56:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32O_2%A_21_199# 1 2 7 9 10 12 13 15 16 18 21 24
+ 25 27 28 31 32 33 36 42 48
r97 48 49 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r98 45 46 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r99 42 43 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.03
+ $X2=2.19 $Y2=1.945
r100 34 36 6.33844 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=2.555 $Y=0.675
+ $X2=2.555 $Y2=0.51
r101 32 34 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=2.405 $Y=0.76
+ $X2=2.555 $Y2=0.675
r102 32 33 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=2.405 $Y=0.76
+ $X2=2.04 $Y2=0.76
r103 31 43 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=2.15 $Y=1.63
+ $X2=2.15 $Y2=1.945
r104 28 31 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=2.15 $Y=1.615
+ $X2=2.15 $Y2=1.63
r105 27 28 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.92 $Y=1.53
+ $X2=2.15 $Y2=1.53
r106 26 33 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=1.92 $Y=0.845
+ $X2=2.04 $Y2=0.76
r107 26 27 28.8111 $w=2.38e-07 $l=6e-07 $layer=LI1_cond $X=1.92 $Y=0.845
+ $X2=1.92 $Y2=1.445
r108 24 27 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.8 $Y=1.53
+ $X2=1.92 $Y2=1.53
r109 24 25 68.1765 $w=1.68e-07 $l=1.045e-06 $layer=LI1_cond $X=1.8 $Y=1.53
+ $X2=0.755 $Y2=1.53
r110 22 48 45.5589 $w=3.65e-07 $l=3.45e-07 $layer=POLY_cond $X=0.62 $Y=1.202
+ $X2=0.965 $Y2=1.202
r111 22 46 13.2055 $w=3.65e-07 $l=1e-07 $layer=POLY_cond $X=0.62 $Y=1.202
+ $X2=0.52 $Y2=1.202
r112 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r113 19 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.645 $Y=1.445
+ $X2=0.755 $Y2=1.53
r114 19 21 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=0.645 $Y=1.445
+ $X2=0.645 $Y2=1.16
r115 16 49 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r116 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r117 13 48 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r118 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r119 10 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r120 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r121 7 45 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r122 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r123 2 42 600 $w=1.7e-07 $l=6.13229e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2.03
r124 2 31 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=1.63
r125 1 36 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.235 $X2=2.62 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%B2 1 3 4 6 8 9 10
r37 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.465
+ $Y=1.16 $X2=1.465 $Y2=1.16
r38 10 15 0.635086 $w=5.63e-07 $l=3e-08 $layer=LI1_cond $X=1.347 $Y=1.19
+ $X2=1.347 $Y2=1.16
r39 9 15 6.56255 $w=5.63e-07 $l=3.1e-07 $layer=LI1_cond $X=1.347 $Y=0.85
+ $X2=1.347 $Y2=1.16
r40 8 14 51.5841 $w=3.3e-07 $l=2.95e-07 $layer=POLY_cond $X=1.76 $Y=1.16
+ $X2=1.465 $Y2=1.16
r41 4 8 49.5676 $w=2.75e-07 $l=2.72947e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.907 $Y2=1.16
r42 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r43 1 8 38.8084 $w=2.75e-07 $l=1.9775e-07 $layer=POLY_cond $X=1.835 $Y=0.995
+ $X2=1.907 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.835 $Y=0.995
+ $X2=1.835 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%B1 1 3 4 6 12 14
c40 12 0 3.53479e-20 $X=2.557 $Y=1.245
c41 4 0 4.20925e-20 $X=2.425 $Y=1.41
r42 12 14 14.5976 $w=2.23e-07 $l=2.85e-07 $layer=LI1_cond $X=2.557 $Y=1.245
+ $X2=2.557 $Y2=1.53
r43 8 12 10.2428 $w=1.68e-07 $l=1.57e-07 $layer=LI1_cond $X=2.4 $Y=1.16
+ $X2=2.557 $Y2=1.16
r44 8 9 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4 $Y=1.16
+ $X2=2.4 $Y2=1.16
r45 4 9 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.16
r46 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r47 1 9 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.34 $Y=0.995
+ $X2=2.425 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.34 $Y=0.995 $X2=2.34
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%A1 1 3 4 6 7
r34 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=1.16 $X2=2.97 $Y2=1.16
r35 7 11 27.744 $w=2.68e-07 $l=6.5e-07 $layer=LI1_cond $X=3.01 $Y=0.51 $X2=3.01
+ $Y2=1.16
r36 4 10 46.5183 $w=3.27e-07 $l=2.87228e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.975 $Y2=1.16
r37 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r38 1 10 38.5818 $w=3.27e-07 $l=2.11069e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.975 $Y2=1.16
r39 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995 $X2=2.87
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%A2 1 3 4 6 7 8 9 10
r35 9 10 12.7285 $w=3.33e-07 $l=3.7e-07 $layer=LI1_cond $X=3.482 $Y=1.16
+ $X2=3.482 $Y2=1.53
r36 9 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.5 $Y=1.16
+ $X2=3.5 $Y2=1.16
r37 8 9 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=3.482 $Y=0.85
+ $X2=3.482 $Y2=1.16
r38 7 8 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=3.482 $Y=0.51
+ $X2=3.482 $Y2=0.85
r39 4 16 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.55 $Y=0.995
+ $X2=3.525 $Y2=1.16
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.55 $Y=0.995 $X2=3.55
+ $Y2=0.56
r41 1 16 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.525 $Y=1.41
+ $X2=3.525 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%A3 1 3 4 6 7 8 12
r25 12 14 33.7665 $w=3.64e-07 $l=2.55e-07 $layer=POLY_cond $X=3.995 $Y=1.202
+ $X2=4.25 $Y2=1.202
r26 11 12 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=3.97 $Y=1.202
+ $X2=3.995 $Y2=1.202
r27 7 8 12.5413 $w=3.38e-07 $l=3.7e-07 $layer=LI1_cond $X=4.335 $Y=1.16
+ $X2=4.335 $Y2=1.53
r28 7 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.25
+ $Y=1.16 $X2=4.25 $Y2=1.16
r29 4 12 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.202
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.995 $Y=1.41
+ $X2=3.995 $Y2=1.985
r31 1 11 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.97 $Y=0.995
+ $X2=3.97 $Y2=1.202
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.97 $Y=0.995 $X2=3.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%X 1 2 3 12 14 19 20 21 22 23 24 33 36
r42 33 36 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=0.24 $Y=0.825
+ $X2=0.24 $Y2=0.85
r43 23 24 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=1.955
+ $X2=0.24 $Y2=2.21
r44 22 23 10.0225 $w=3.78e-07 $l=2.55e-07 $layer=LI1_cond $X=0.24 $Y=1.53
+ $X2=0.24 $Y2=1.785
r45 21 22 17.9567 $w=2.08e-07 $l=3.4e-07 $layer=LI1_cond $X=0.24 $Y=1.19
+ $X2=0.24 $Y2=1.53
r46 20 33 3.09364 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=0.24 $Y=0.74 $X2=0.24
+ $Y2=0.825
r47 20 21 16.3723 $w=2.08e-07 $l=3.1e-07 $layer=LI1_cond $X=0.24 $Y=0.88
+ $X2=0.24 $Y2=1.19
r48 20 36 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=0.24 $Y=0.88 $X2=0.24
+ $Y2=0.85
r49 15 23 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.345 $Y=1.87
+ $X2=0.24 $Y2=1.87
r50 14 19 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=1.87 $X2=1.2
+ $Y2=1.87
r51 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=1.87
+ $X2=0.345 $Y2=1.87
r52 10 20 3.82155 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.24 $Y2=0.74
r53 10 12 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.73 $Y2=0.74
r54 3 19 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.95
r55 2 23 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.95
r56 1 12 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%VPWR 1 2 3 12 16 18 20 22 24 29 34 40 43 47
r68 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r69 43 44 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r71 38 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r72 38 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r74 35 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.105 $Y2=2.72
r75 35 37 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.295 $Y=2.72
+ $X2=3.91 $Y2=2.72
r76 34 46 5.04433 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=4.307 $Y2=2.72
r77 34 37 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=2.72
+ $X2=3.91 $Y2=2.72
r78 33 44 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 33 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r81 30 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r82 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r83 29 43 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.105 $Y2=2.72
r84 29 32 115.15 $w=1.68e-07 $l=1.765e-06 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 24 40 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r86 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r87 22 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r88 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r89 18 46 3.19589 $w=3.85e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.207 $Y=2.635
+ $X2=4.307 $Y2=2.72
r90 18 20 19.0078 $w=3.83e-07 $l=6.35e-07 $layer=LI1_cond $X=4.207 $Y=2.635
+ $X2=4.207 $Y2=2
r91 14 43 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.105 $Y=2.635
+ $X2=3.105 $Y2=2.72
r92 14 16 12.4343 $w=3.78e-07 $l=4.1e-07 $layer=LI1_cond $X=3.105 $Y=2.635
+ $X2=3.105 $Y2=2.225
r93 10 40 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r94 10 12 12.8892 $w=3.78e-07 $l=4.25e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.21
r95 3 20 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.085
+ $Y=1.485 $X2=4.23 $Y2=2
r96 2 16 600 $w=1.7e-07 $l=8.09259e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.225
r97 1 12 600 $w=1.7e-07 $l=7.94198e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%A_319_297# 1 2 3 12 14 15 16 17 18 25
c37 16 0 7.74404e-20 $X=2.66 $Y=1.965
r38 19 23 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.745 $Y=1.88
+ $X2=2.66 $Y2=1.88
r39 18 25 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.675 $Y=1.88
+ $X2=3.76 $Y2=1.88
r40 18 19 60.6738 $w=1.68e-07 $l=9.3e-07 $layer=LI1_cond $X=3.675 $Y=1.88
+ $X2=2.745 $Y2=1.88
r41 16 23 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.66 $Y=1.965
+ $X2=2.66 $Y2=1.88
r42 16 17 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.66 $Y=1.965
+ $X2=2.66 $Y2=2.295
r43 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.575 $Y=2.38
+ $X2=2.66 $Y2=2.295
r44 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.575 $Y=2.38
+ $X2=1.805 $Y2=2.38
r45 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.72 $Y=2.295
+ $X2=1.805 $Y2=2.38
r46 10 12 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.72 $Y=2.295
+ $X2=1.72 $Y2=1.95
r47 3 25 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.615
+ $Y=1.485 $X2=3.76 $Y2=1.96
r48 2 23 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.96
r49 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32O_2%VGND 1 2 3 10 12 14 16 18 25 39 45 48
r58 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r59 43 45 8.91451 $w=5.28e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=0.18
+ $X2=1.74 $Y2=0.18
r60 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r61 41 43 0.789863 $w=5.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.575 $Y=0.18
+ $X2=1.61 $Y2=0.18
r62 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r63 37 41 9.5912 $w=5.28e-07 $l=4.25e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=1.575 $Y2=0.18
r64 37 39 9.70437 $w=5.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.15 $Y=0.18
+ $X2=0.985 $Y2=0.18
r65 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r66 32 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r67 31 32 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r68 29 32 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r69 29 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r70 28 31 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.91
+ $Y2=0
r71 28 45 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.07 $Y=0 $X2=1.74
+ $Y2=0
r72 28 29 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 25 47 5.04433 $w=1.7e-07 $l=2.92e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.307
+ $Y2=0
r74 25 31 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=3.91
+ $Y2=0
r75 24 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r76 23 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=0.985
+ $Y2=0
r77 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r78 21 34 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r79 21 23 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r80 18 24 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r81 18 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r82 14 47 3.19589 $w=3.85e-07 $l=1.36015e-07 $layer=LI1_cond $X=4.207 $Y=0.085
+ $X2=4.307 $Y2=0
r83 14 16 8.83041 $w=3.83e-07 $l=2.95e-07 $layer=LI1_cond $X=4.207 $Y=0.085
+ $X2=4.207 $Y2=0.38
r84 10 34 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r85 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.38
r86 3 16 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.045
+ $Y=0.235 $X2=4.23 $Y2=0.38
r87 2 41 91 $w=1.7e-07 $l=5.69078e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.575 $Y2=0.36
r88 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

