* File: sky130_fd_sc_hdll__clkbuf_6.spice
* Created: Wed Sep  2 08:25:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkbuf_6.pex.spice"
.subckt sky130_fd_sc_hdll__clkbuf_6  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_117_297#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0567 PD=1.46 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75003.5 A=0.063 P=1.14 MULT=1
MM1010 N_VGND_M1010_d N_A_M1010_g N_A_117_297#_M1004_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75003.1 A=0.063 P=1.14 MULT=1
MM1005 N_X_M1005_d N_A_117_297#_M1005_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.2
+ SB=75002.5 A=0.063 P=1.14 MULT=1
MM1007 N_X_M1005_d N_A_117_297#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.07665 PD=0.69 PS=0.785 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.6
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1011 N_X_M1011_d N_A_117_297#_M1011_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.07665 PD=0.695 PS=0.785 NRD=0 NRS=11.424 M=1 R=2.8 SA=75002.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1013 N_X_M1011_d N_A_117_297#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.05775 AS=0.0777 PD=0.695 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75002.5
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1014 N_X_M1014_d N_A_117_297#_M1014_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75003.1
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1015 N_X_M1014_d N_A_117_297#_M1015_g N_VGND_M1015_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.1302 PD=0.69 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75003.5
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1006_d N_A_117_297#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A_117_297#_M1002_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1002_d N_A_117_297#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_117_297#_M1008_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1008_d N_A_117_297#_M1009_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_117_297#_M1012_g N_X_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=7.9929 P=13.17
*
.include "sky130_fd_sc_hdll__clkbuf_6.pxi.spice"
*
.ends
*
*
