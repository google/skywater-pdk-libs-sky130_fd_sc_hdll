* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0

.SUBCKT sky130_fd_sc_hdll__or3b_1 A B C_N VGND VNB VPB VPWR X
*.PININFO A:I B:I C_N:I VGND:I VNB:I VPB:I VPWR:I X:O
MMP0 VPWR A VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP1 sndPA B VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMP2 sndPB C VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP2 C C_N VPB pfet_01v8_hvt m=1 w=0.42 l=0.18 mult=1 sa=0.265
+ sb=0.265 sd=0.28 topography=normal area=0.063 perim=1.14
MMIP3 X y VPB pfet_01v8_hvt m=1 w=1.0 l=0.18 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN0 y A VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN1 y B VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMN2 y C VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN2 C C_N VNB nfet_01v8 m=1 w=0.42 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
MMIN3 X y VNB nfet_01v8 m=1 w=0.65 l=0.15 mult=1 sa=0.265 sb=0.265
+ sd=0.28 topography=normal area=0.063 perim=1.14
.ENDS sky130_fd_sc_hdll__or3b_1
