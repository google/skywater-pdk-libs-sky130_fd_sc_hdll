* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_225_47# B a_693_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_693_47# C a_1081_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_1081_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND D a_1081_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 a_225_47# B a_693_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_693_47# C a_1081_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_27_47# A_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 Y a_27_47# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_1081_47# C a_693_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_1081_47# C a_693_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 VGND D a_1081_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_27_47# A_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 Y a_27_47# a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_1081_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_693_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_225_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 a_693_47# B a_225_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X32 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_225_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
