* File: sky130_fd_sc_hdll__clkbuf_1.pex.spice
* Created: Thu Aug 27 19:01:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_1%A_75_212# 1 2 7 9 12 15 17 18 19 20 21 24
+ 28 34
r65 31 34 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=0.51 $Y=1.225
+ $X2=0.65 $Y2=1.225
r66 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.51
+ $Y=1.225 $X2=0.51 $Y2=1.225
r67 26 28 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.58 $Y=1.705
+ $X2=1.58 $Y2=1.96
r68 22 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=1.54 $Y=0.635
+ $X2=1.54 $Y2=0.445
r69 20 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.495 $Y=1.62
+ $X2=1.58 $Y2=1.705
r70 20 21 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.495 $Y=1.62
+ $X2=0.76 $Y2=1.62
r71 18 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.455 $Y=0.72
+ $X2=1.54 $Y2=0.635
r72 18 19 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.455 $Y=0.72
+ $X2=0.76 $Y2=0.72
r73 17 21 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.65 $Y=1.535
+ $X2=0.76 $Y2=1.62
r74 16 34 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=1.39
+ $X2=0.65 $Y2=1.225
r75 16 17 7.59565 $w=2.18e-07 $l=1.45e-07 $layer=LI1_cond $X=0.65 $Y=1.39
+ $X2=0.65 $Y2=1.535
r76 15 34 3.11056 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=0.65 $Y=1.06
+ $X2=0.65 $Y2=1.225
r77 14 19 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.65 $Y=0.805
+ $X2=0.76 $Y2=0.72
r78 14 15 13.3579 $w=2.18e-07 $l=2.55e-07 $layer=LI1_cond $X=0.65 $Y=0.805
+ $X2=0.65 $Y2=1.06
r79 10 32 38.9026 $w=2.7e-07 $l=1.72337e-07 $layer=POLY_cond $X=0.52 $Y=1.06
+ $X2=0.535 $Y2=1.225
r80 10 12 289.713 $w=1.5e-07 $l=5.65e-07 $layer=POLY_cond $X=0.52 $Y=1.06
+ $X2=0.52 $Y2=0.495
r81 7 32 75.8829 $w=2.7e-07 $l=4.14518e-07 $layer=POLY_cond $X=0.495 $Y=1.62
+ $X2=0.535 $Y2=1.225
r82 7 9 125.856 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=0.495 $Y=1.62
+ $X2=0.495 $Y2=2.09
r83 2 28 300 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=2 $X=1.435
+ $Y=1.695 $X2=1.58 $Y2=1.96
r84 1 24 182 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_NDIFF $count=1 $X=1.395
+ $Y=0.235 $X2=1.54 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_1%A 3 6 7 9 10 16 22
r30 16 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.58
+ $Y=1.16 $X2=1.58 $Y2=1.16
r31 14 16 41.0924 $w=3.3e-07 $l=2.35e-07 $layer=POLY_cond $X=1.345 $Y=1.16
+ $X2=1.58 $Y2=1.16
r32 12 14 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=1.32 $Y=1.16
+ $X2=1.345 $Y2=1.16
r33 10 22 0.155736 $w=3.68e-07 $l=5e-09 $layer=LI1_cond $X=1.515 $Y=1.17
+ $X2=1.52 $Y2=1.17
r34 7 9 125.856 $w=1.8e-07 $l=4.7e-07 $layer=POLY_cond $X=1.345 $Y=1.62
+ $X2=1.345 $Y2=2.09
r35 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.345 $Y=1.52 $X2=1.345
+ $Y2=1.62
r36 5 14 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=1.16
r37 5 6 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=1.345 $Y=1.325
+ $X2=1.345 $Y2=1.52
r38 1 12 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.32 $Y=0.995
+ $X2=1.32 $Y2=1.16
r39 1 3 256.383 $w=1.5e-07 $l=5e-07 $layer=POLY_cond $X=1.32 $Y=0.995 $X2=1.32
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_1%X 1 2 10 11 12 13 14 15
r24 14 15 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=1.87
+ $X2=0.22 $Y2=2.21
r25 11 14 7.46954 $w=2.68e-07 $l=1.75e-07 $layer=LI1_cond $X=0.22 $Y=1.695
+ $X2=0.22 $Y2=1.87
r26 11 12 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=0.22 $Y=1.695
+ $X2=0.22 $Y2=1.56
r27 10 12 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=0.17 $Y=0.76 $X2=0.17
+ $Y2=1.56
r28 9 13 5.31897 $w=2.58e-07 $l=1.2e-07 $layer=LI1_cond $X=0.215 $Y=0.63
+ $X2=0.215 $Y2=0.51
r29 9 10 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=0.215 $Y=0.63
+ $X2=0.215 $Y2=0.76
r30 2 14 300 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.695 $X2=0.26 $Y2=1.895
r31 1 13 182 $w=1.7e-07 $l=3.51994e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_1%VPWR 1 6 8 10 17 18 21 26
r24 21 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r25 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r26 15 21 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=0.9 $Y2=2.72
r27 15 17 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.275 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 13 26 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 12 13 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 10 21 14.1623 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.9 $Y2=2.72
r31 10 12 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r32 8 18 0.102435 $w=4.8e-07 $l=3.6e-07 $layer=MET1_cond $X=1.25 $Y=2.72
+ $X2=1.61 $Y2=2.72
r33 8 26 0.0284542 $w=4.8e-07 $l=1e-07 $layer=MET1_cond $X=1.25 $Y=2.72 $X2=1.15
+ $Y2=2.72
r34 4 21 3.00456 $w=7.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=2.635 $X2=0.9
+ $Y2=2.72
r35 4 6 10.7647 $w=7.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.9 $Y=2.635 $X2=0.9
+ $Y2=1.96
r36 1 6 150 $w=1.7e-07 $l=6.13351e-07 $layer=licon1_PDIFF $count=4 $X=0.585
+ $Y=1.695 $X2=1.08 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_1%VGND 1 4 13 14 19 25 30
r27 23 25 8.96211 $w=5.48e-07 $l=1.25e-07 $layer=LI1_cond $X=1.15 $Y=0.19
+ $X2=1.275 $Y2=0.19
r28 23 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r29 21 23 1.52228 $w=5.48e-07 $l=7e-08 $layer=LI1_cond $X=1.08 $Y=0.19 $X2=1.15
+ $Y2=0.19
r30 18 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r31 17 21 8.48128 $w=5.48e-07 $l=3.9e-07 $layer=LI1_cond $X=0.69 $Y=0.19
+ $X2=1.08 $Y2=0.19
r32 17 19 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=0.69 $Y=0.19
+ $X2=0.525 $Y2=0.19
r33 17 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r34 13 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.275
+ $Y2=0
r35 13 14 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r36 9 18 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r37 8 19 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.23 $Y=0 $X2=0.525
+ $Y2=0
r38 8 9 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r39 4 14 0.102435 $w=4.8e-07 $l=3.6e-07 $layer=MET1_cond $X=1.25 $Y=0 $X2=1.61
+ $Y2=0
r40 4 30 0.0284542 $w=4.8e-07 $l=1e-07 $layer=MET1_cond $X=1.25 $Y=0 $X2=1.15
+ $Y2=0
r41 1 21 91 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_NDIFF $count=2 $X=0.595
+ $Y=0.235 $X2=1.08 $Y2=0.38
.ends

