* File: sky130_fd_sc_hdll__ebufn_4.pxi.spice
* Created: Wed Sep  2 08:30:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%A N_A_c_95_n N_A_M1018_g N_A_c_96_n N_A_M1007_g
+ A A PM_SKY130_FD_SC_HDLL__EBUFN_4%A
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%TE_B N_TE_B_M1009_g N_TE_B_c_130_n
+ N_TE_B_M1017_g N_TE_B_c_131_n N_TE_B_c_128_n N_TE_B_c_133_n N_TE_B_M1005_g
+ N_TE_B_c_134_n N_TE_B_c_135_n N_TE_B_M1008_g N_TE_B_c_136_n N_TE_B_c_137_n
+ N_TE_B_M1012_g N_TE_B_c_138_n N_TE_B_c_139_n N_TE_B_M1016_g N_TE_B_c_140_n
+ N_TE_B_c_141_n N_TE_B_c_142_n TE_B PM_SKY130_FD_SC_HDLL__EBUFN_4%TE_B
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%A_224_47# N_A_224_47#_M1009_d
+ N_A_224_47#_M1017_d N_A_224_47#_c_214_n N_A_224_47#_M1002_g
+ N_A_224_47#_c_215_n N_A_224_47#_c_216_n N_A_224_47#_c_217_n
+ N_A_224_47#_M1006_g N_A_224_47#_c_218_n N_A_224_47#_c_219_n
+ N_A_224_47#_M1014_g N_A_224_47#_c_220_n N_A_224_47#_M1015_g
+ N_A_224_47#_c_221_n N_A_224_47#_c_222_n N_A_224_47#_c_223_n
+ N_A_224_47#_c_230_n N_A_224_47#_c_224_n N_A_224_47#_c_225_n
+ N_A_224_47#_c_226_n N_A_224_47#_c_227_n N_A_224_47#_c_228_n
+ N_A_224_47#_c_229_n PM_SKY130_FD_SC_HDLL__EBUFN_4%A_224_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%A_27_47# N_A_27_47#_M1018_s N_A_27_47#_M1007_s
+ N_A_27_47#_M1001_g N_A_27_47#_c_319_n N_A_27_47#_M1000_g N_A_27_47#_M1003_g
+ N_A_27_47#_c_320_n N_A_27_47#_M1004_g N_A_27_47#_M1010_g N_A_27_47#_c_321_n
+ N_A_27_47#_M1011_g N_A_27_47#_c_322_n N_A_27_47#_M1013_g N_A_27_47#_M1019_g
+ N_A_27_47#_c_323_n N_A_27_47#_c_324_n N_A_27_47#_c_313_n N_A_27_47#_c_314_n
+ N_A_27_47#_c_315_n N_A_27_47#_c_327_n N_A_27_47#_c_316_n N_A_27_47#_c_317_n
+ N_A_27_47#_c_318_n PM_SKY130_FD_SC_HDLL__EBUFN_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%VPWR N_VPWR_M1007_d N_VPWR_M1005_s
+ N_VPWR_M1012_s N_VPWR_c_408_n N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n VPWR N_VPWR_c_414_n N_VPWR_c_415_n
+ N_VPWR_c_407_n N_VPWR_c_417_n PM_SKY130_FD_SC_HDLL__EBUFN_4%VPWR
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%A_340_309# N_A_340_309#_M1005_d
+ N_A_340_309#_M1008_d N_A_340_309#_M1016_d N_A_340_309#_M1004_d
+ N_A_340_309#_M1013_d N_A_340_309#_c_485_n N_A_340_309#_c_514_n
+ N_A_340_309#_c_486_n N_A_340_309#_c_493_n N_A_340_309#_c_487_n
+ N_A_340_309#_c_494_n PM_SKY130_FD_SC_HDLL__EBUFN_4%A_340_309#
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%Z N_Z_M1001_d N_Z_M1010_d N_Z_M1000_s
+ N_Z_M1011_s N_Z_c_561_n Z Z Z Z Z Z Z Z Z Z N_Z_c_545_n Z Z Z Z Z Z Z
+ N_Z_c_542_n PM_SKY130_FD_SC_HDLL__EBUFN_4%Z
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%VGND N_VGND_M1018_d N_VGND_M1002_s
+ N_VGND_M1014_s N_VGND_c_606_n N_VGND_c_607_n N_VGND_c_608_n N_VGND_c_609_n
+ VGND N_VGND_c_610_n N_VGND_c_611_n N_VGND_c_612_n N_VGND_c_613_n
+ N_VGND_c_614_n N_VGND_c_615_n N_VGND_c_616_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_4%VGND
x_PM_SKY130_FD_SC_HDLL__EBUFN_4%A_413_47# N_A_413_47#_M1002_d
+ N_A_413_47#_M1006_d N_A_413_47#_M1015_d N_A_413_47#_M1003_s
+ N_A_413_47#_M1019_s N_A_413_47#_c_685_n N_A_413_47#_c_690_n
+ N_A_413_47#_c_686_n N_A_413_47#_c_696_n N_A_413_47#_c_697_n
+ N_A_413_47#_c_743_n N_A_413_47#_c_687_n N_A_413_47#_c_703_n
+ PM_SKY130_FD_SC_HDLL__EBUFN_4%A_413_47#
cc_1 VNB N_A_c_95_n 0.0197693f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_c_96_n 0.0300357f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB A 0.00216056f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_4 VNB N_TE_B_M1009_g 0.0230541f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_5 VNB N_TE_B_c_128_n 0.0431218f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB TE_B 0.00130409f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_224_47#_c_214_n 0.0184073f $X=-0.19 $Y=-0.24 $X2=0.61 $Y2=0.765
cc_8 VNB N_A_224_47#_c_215_n 0.0137076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_224_47#_c_216_n 0.00853733f $X=-0.19 $Y=-0.24 $X2=0.577 $Y2=1.16
cc_10 VNB N_A_224_47#_c_217_n 0.0154576f $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_11 VNB N_A_224_47#_c_218_n 0.0113204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_224_47#_c_219_n 0.0145707f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.16
cc_13 VNB N_A_224_47#_c_220_n 0.0137381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_224_47#_c_221_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_224_47#_c_222_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_224_47#_c_223_n 0.0112749f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_224_47#_c_224_n 0.0125344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_224_47#_c_225_n 3.72754e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_224_47#_c_226_n 0.0208019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_224_47#_c_227_n 0.00171924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_224_47#_c_228_n 0.0398595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_224_47#_c_229_n 0.0157353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_M1001_g 0.0190941f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_M1003_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_M1010_g 0.0190914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_M1019_g 0.0219052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_313_n 0.0150059f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_27_47#_c_314_n 0.023363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_27_47#_c_315_n 0.0113098f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_27_47#_c_316_n 0.00524072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_27_47#_c_317_n 0.0020849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_27_47#_c_318_n 0.0916105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_407_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB Z 0.0222703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Z_c_542_n 0.0112101f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_606_n 8.48704e-19 $X=-0.19 $Y=-0.24 $X2=0.575 $Y2=1.16
cc_37 VNB N_VGND_c_607_n 0.00241972f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_608_n 0.0135077f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.53
cc_39 VNB N_VGND_c_609_n 0.00272154f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_610_n 0.0151734f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_611_n 0.0363596f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_612_n 0.0627984f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_613_n 0.326404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_614_n 0.00655113f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_615_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_616_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_413_47#_c_685_n 0.00522107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_413_47#_c_686_n 0.00282551f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_413_47#_c_687_n 0.00812227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_A_c_96_n 0.0312312f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB A 0.00133979f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=0.765
cc_52 VPB N_TE_B_c_130_n 0.0199329f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_53 VPB N_TE_B_c_131_n 0.0187253f $X=-0.19 $Y=1.305 $X2=0.61 $Y2=1.445
cc_54 VPB N_TE_B_c_128_n 0.0277413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_TE_B_c_133_n 0.0184062f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_TE_B_c_134_n 0.0139927f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_57 VPB N_TE_B_c_135_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_TE_B_c_136_n 0.0125186f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.53
cc_59 VPB N_TE_B_c_137_n 0.0154273f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_TE_B_c_138_n 0.0266127f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_TE_B_c_139_n 0.0191144f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_TE_B_c_140_n 0.00735165f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_TE_B_c_141_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_TE_B_c_142_n 0.00590532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB TE_B 0.00338357f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_224_47#_c_230_n 0.00719229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_224_47#_c_225_n 0.0124082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_319_n 0.0201091f $X=-0.19 $Y=1.305 $X2=0.577 $Y2=1.16
cc_69 VPB N_A_27_47#_c_320_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.53
cc_70 VPB N_A_27_47#_c_321_n 0.0158725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_47#_c_322_n 0.0191865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_47#_c_323_n 0.00494099f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_47#_c_324_n 0.0219831f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_47#_c_314_n 0.0194654f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_315_n 0.00158633f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_47#_c_327_n 0.00136192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_316_n 0.0206984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_318_n 0.0290885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_408_n 0.00333285f $X=-0.19 $Y=1.305 $X2=0.575 $Y2=1.16
cc_80 VPB N_VPWR_c_409_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_410_n 0.00547148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_411_n 0.028693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_412_n 0.0138823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_413_n 0.00436029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_414_n 0.0150576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_415_n 0.0712237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_407_n 0.056778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_417_n 0.00743881f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_340_309#_c_485_n 0.0034756f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.53
cc_90 VPB N_A_340_309#_c_486_n 0.00180023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_340_309#_c_487_n 0.023886f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB Z 0.0144748f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB Z 0.0072218f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Z_c_545_n 0.0124309f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 N_A_c_95_n N_TE_B_M1009_g 0.0185669f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_c_96_n N_TE_B_M1009_g 0.0215233f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_97 A N_TE_B_M1009_g 0.00439489f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A_c_96_n N_TE_B_c_130_n 0.0222862f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 A N_TE_B_c_130_n 0.00530706f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A_c_96_n N_TE_B_c_128_n 0.00255013f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_96_n TE_B 5.03739e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_102 A TE_B 0.0510354f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_103 N_A_c_95_n N_A_27_47#_c_314_n 0.0184886f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_96_n N_A_27_47#_c_314_n 0.00940857f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_105 A N_A_27_47#_c_314_n 0.0674439f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_106 N_A_c_96_n N_A_27_47#_c_315_n 0.00269146f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_107 A N_A_27_47#_c_315_n 0.00275793f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_108 N_A_c_96_n N_A_27_47#_c_316_n 0.00959072f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_109 A N_A_27_47#_c_316_n 0.0221286f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_110 A N_VPWR_M1007_d 0.00488784f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_111 N_A_c_96_n N_VPWR_c_408_n 0.0177792f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_112 A N_VPWR_c_408_n 0.0219873f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_113 N_A_c_96_n N_VPWR_c_414_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_96_n N_VPWR_c_407_n 0.0082412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 A N_VGND_M1018_d 0.00372716f $X=0.61 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_116 N_A_c_95_n N_VGND_c_606_n 0.0118659f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_c_96_n N_VGND_c_606_n 8.9449e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_118 A N_VGND_c_606_n 0.0215942f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_119 N_A_c_95_n N_VGND_c_610_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_95_n N_VGND_c_613_n 0.00818925f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_121 A N_VGND_c_613_n 0.00210925f $X=0.61 $Y=0.765 $X2=0 $Y2=0
cc_122 TE_B N_A_224_47#_M1009_d 0.00411646f $X=1.075 $Y=0.765 $X2=-0.19
+ $Y2=-0.24
cc_123 N_TE_B_c_141_n N_A_224_47#_c_215_n 0.0152647f $X=2.53 $Y=1.395 $X2=0
+ $Y2=0
cc_124 N_TE_B_c_134_n N_A_224_47#_c_216_n 0.0152647f $X=2.44 $Y=1.395 $X2=0
+ $Y2=0
cc_125 N_TE_B_c_142_n N_A_224_47#_c_218_n 0.0152647f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_126 N_TE_B_c_136_n N_A_224_47#_c_221_n 0.0152647f $X=2.91 $Y=1.395 $X2=0
+ $Y2=0
cc_127 N_TE_B_c_138_n N_A_224_47#_c_222_n 0.0152647f $X=3.38 $Y=1.395 $X2=0
+ $Y2=0
cc_128 N_TE_B_c_128_n N_A_224_47#_c_223_n 0.00402323f $X=1.695 $Y=1.395 $X2=0
+ $Y2=0
cc_129 TE_B N_A_224_47#_c_223_n 0.0143413f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_130 N_TE_B_c_133_n N_A_224_47#_c_230_n 0.00460224f $X=2.06 $Y=1.47 $X2=0
+ $Y2=0
cc_131 N_TE_B_M1009_g N_A_224_47#_c_224_n 0.00535911f $X=1.045 $Y=0.56 $X2=0
+ $Y2=0
cc_132 TE_B N_A_224_47#_c_224_n 0.0213591f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_133 N_TE_B_c_130_n N_A_224_47#_c_225_n 0.00392628f $X=1.07 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_TE_B_c_131_n N_A_224_47#_c_225_n 0.0132701f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_135 N_TE_B_c_128_n N_A_224_47#_c_225_n 0.0170621f $X=1.695 $Y=1.395 $X2=0
+ $Y2=0
cc_136 N_TE_B_c_133_n N_A_224_47#_c_225_n 0.00696587f $X=2.06 $Y=1.47 $X2=0
+ $Y2=0
cc_137 TE_B N_A_224_47#_c_225_n 0.0243642f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_138 N_TE_B_c_131_n N_A_224_47#_c_226_n 0.0237476f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_139 N_TE_B_c_128_n N_A_224_47#_c_227_n 0.00943564f $X=1.695 $Y=1.395 $X2=0
+ $Y2=0
cc_140 TE_B N_A_224_47#_c_227_n 0.019555f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_141 N_TE_B_c_131_n N_A_27_47#_c_316_n 0.0323665f $X=1.97 $Y=1.395 $X2=0 $Y2=0
cc_142 N_TE_B_c_128_n N_A_27_47#_c_316_n 0.00750138f $X=1.695 $Y=1.395 $X2=0
+ $Y2=0
cc_143 TE_B N_A_27_47#_c_316_n 0.0325489f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_144 N_TE_B_c_130_n N_VPWR_c_408_n 0.00772308f $X=1.07 $Y=1.41 $X2=0 $Y2=0
cc_145 N_TE_B_c_135_n N_VPWR_c_409_n 4.96664e-19 $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_146 N_TE_B_c_137_n N_VPWR_c_409_n 0.00666322f $X=3 $Y=1.47 $X2=0 $Y2=0
cc_147 N_TE_B_c_139_n N_VPWR_c_409_n 0.00813391f $X=3.47 $Y=1.47 $X2=0 $Y2=0
cc_148 N_TE_B_c_133_n N_VPWR_c_410_n 0.0107351f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_149 N_TE_B_c_135_n N_VPWR_c_410_n 0.00666244f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_150 N_TE_B_c_137_n N_VPWR_c_410_n 4.99599e-19 $X=3 $Y=1.47 $X2=0 $Y2=0
cc_151 N_TE_B_c_130_n N_VPWR_c_411_n 0.00700684f $X=1.07 $Y=1.41 $X2=0 $Y2=0
cc_152 N_TE_B_c_133_n N_VPWR_c_411_n 0.00309439f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_153 N_TE_B_c_135_n N_VPWR_c_412_n 0.00450093f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_154 N_TE_B_c_137_n N_VPWR_c_412_n 0.00449565f $X=3 $Y=1.47 $X2=0 $Y2=0
cc_155 N_TE_B_c_139_n N_VPWR_c_415_n 0.00449565f $X=3.47 $Y=1.47 $X2=0 $Y2=0
cc_156 N_TE_B_c_130_n N_VPWR_c_407_n 0.0139825f $X=1.07 $Y=1.41 $X2=0 $Y2=0
cc_157 N_TE_B_c_133_n N_VPWR_c_407_n 0.00495648f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_158 N_TE_B_c_135_n N_VPWR_c_407_n 0.00508383f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_159 N_TE_B_c_137_n N_VPWR_c_407_n 0.00508633f $X=3 $Y=1.47 $X2=0 $Y2=0
cc_160 N_TE_B_c_139_n N_VPWR_c_407_n 0.00646266f $X=3.47 $Y=1.47 $X2=0 $Y2=0
cc_161 N_TE_B_c_131_n N_A_340_309#_c_486_n 0.00228495f $X=1.97 $Y=1.395 $X2=0
+ $Y2=0
cc_162 N_TE_B_c_133_n N_A_340_309#_c_486_n 0.01623f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_163 N_TE_B_c_134_n N_A_340_309#_c_486_n 4.50429e-19 $X=2.44 $Y=1.395 $X2=0
+ $Y2=0
cc_164 N_TE_B_c_135_n N_A_340_309#_c_486_n 0.0149975f $X=2.53 $Y=1.47 $X2=0
+ $Y2=0
cc_165 N_TE_B_c_136_n N_A_340_309#_c_486_n 4.9053e-19 $X=2.91 $Y=1.395 $X2=0
+ $Y2=0
cc_166 N_TE_B_c_139_n N_A_340_309#_c_493_n 0.0126872f $X=3.47 $Y=1.47 $X2=0
+ $Y2=0
cc_167 N_TE_B_c_137_n N_A_340_309#_c_494_n 0.0149486f $X=3 $Y=1.47 $X2=0 $Y2=0
cc_168 N_TE_B_c_138_n N_A_340_309#_c_494_n 4.50116e-19 $X=3.38 $Y=1.395 $X2=0
+ $Y2=0
cc_169 N_TE_B_c_139_n N_A_340_309#_c_494_n 0.0174245f $X=3.47 $Y=1.47 $X2=0
+ $Y2=0
cc_170 N_TE_B_c_133_n N_Z_c_545_n 0.0103614f $X=2.06 $Y=1.47 $X2=0 $Y2=0
cc_171 N_TE_B_c_134_n N_Z_c_545_n 0.00508009f $X=2.44 $Y=1.395 $X2=0 $Y2=0
cc_172 N_TE_B_c_135_n N_Z_c_545_n 0.0130132f $X=2.53 $Y=1.47 $X2=0 $Y2=0
cc_173 N_TE_B_c_136_n N_Z_c_545_n 0.00493492f $X=2.91 $Y=1.395 $X2=0 $Y2=0
cc_174 N_TE_B_c_137_n N_Z_c_545_n 0.0130331f $X=3 $Y=1.47 $X2=0 $Y2=0
cc_175 N_TE_B_c_138_n N_Z_c_545_n 0.00755182f $X=3.38 $Y=1.395 $X2=0 $Y2=0
cc_176 N_TE_B_c_139_n N_Z_c_545_n 0.0160447f $X=3.47 $Y=1.47 $X2=0 $Y2=0
cc_177 N_TE_B_c_140_n N_Z_c_545_n 0.00195737f $X=2.06 $Y=1.395 $X2=0 $Y2=0
cc_178 N_TE_B_c_141_n N_Z_c_545_n 0.0017524f $X=2.53 $Y=1.395 $X2=0 $Y2=0
cc_179 N_TE_B_c_142_n N_Z_c_545_n 0.0017524f $X=3 $Y=1.395 $X2=0 $Y2=0
cc_180 N_TE_B_M1009_g N_VGND_c_606_n 0.0153857f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_181 N_TE_B_M1009_g N_VGND_c_611_n 0.00544582f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_182 N_TE_B_M1009_g N_VGND_c_613_n 0.00681521f $X=1.045 $Y=0.56 $X2=0 $Y2=0
cc_183 TE_B N_VGND_c_613_n 0.00771034f $X=1.075 $Y=0.765 $X2=0 $Y2=0
cc_184 N_A_224_47#_c_228_n N_A_27_47#_M1001_g 0.021998f $X=3.97 $Y=1.035 $X2=0
+ $Y2=0
cc_185 N_A_224_47#_c_229_n N_A_27_47#_M1001_g 0.0143433f $X=3.97 $Y=0.96 $X2=0
+ $Y2=0
cc_186 N_A_224_47#_c_226_n N_A_27_47#_c_327_n 3.57817e-19 $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_187 N_A_224_47#_c_223_n N_A_27_47#_c_316_n 0.00627825f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_188 N_A_224_47#_c_225_n N_A_27_47#_c_316_n 0.0140893f $X=1.687 $Y=1.595 $X2=0
+ $Y2=0
cc_189 N_A_224_47#_c_226_n N_A_27_47#_c_316_n 0.0725143f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_190 N_A_224_47#_c_227_n N_A_27_47#_c_316_n 0.0192351f $X=1.687 $Y=1.15 $X2=0
+ $Y2=0
cc_191 N_A_224_47#_c_228_n N_A_27_47#_c_316_n 0.004011f $X=3.97 $Y=1.035 $X2=0
+ $Y2=0
cc_192 N_A_224_47#_c_226_n N_A_27_47#_c_317_n 0.0198098f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_224_47#_c_228_n N_A_27_47#_c_317_n 8.31351e-19 $X=3.97 $Y=1.035 $X2=0
+ $Y2=0
cc_194 N_A_224_47#_c_226_n N_A_27_47#_c_318_n 3.5001e-19 $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_224_47#_c_230_n N_VPWR_c_411_n 0.0173025f $X=1.305 $Y=1.96 $X2=0
+ $Y2=0
cc_196 N_A_224_47#_M1017_d N_VPWR_c_407_n 0.0035638f $X=1.16 $Y=1.485 $X2=0
+ $Y2=0
cc_197 N_A_224_47#_c_230_n N_VPWR_c_407_n 0.00975095f $X=1.305 $Y=1.96 $X2=0
+ $Y2=0
cc_198 N_A_224_47#_c_225_n N_A_340_309#_M1005_d 0.00473819f $X=1.687 $Y=1.595
+ $X2=-0.19 $Y2=-0.24
cc_199 N_A_224_47#_c_230_n N_A_340_309#_c_485_n 0.0247517f $X=1.305 $Y=1.96
+ $X2=0 $Y2=0
cc_200 N_A_224_47#_c_230_n N_A_340_309#_c_486_n 0.0140934f $X=1.305 $Y=1.96
+ $X2=0 $Y2=0
cc_201 N_A_224_47#_c_225_n N_A_340_309#_c_486_n 0.0128275f $X=1.687 $Y=1.595
+ $X2=0 $Y2=0
cc_202 N_A_224_47#_c_226_n N_A_340_309#_c_486_n 0.00290582f $X=3.945 $Y=1.16
+ $X2=0 $Y2=0
cc_203 N_A_224_47#_c_216_n N_Z_c_545_n 9.02704e-19 $X=2.525 $Y=1.035 $X2=0 $Y2=0
cc_204 N_A_224_47#_c_220_n N_Z_c_545_n 0.00103677f $X=3.78 $Y=1.035 $X2=0 $Y2=0
cc_205 N_A_224_47#_c_225_n N_Z_c_545_n 0.023239f $X=1.687 $Y=1.595 $X2=0 $Y2=0
cc_206 N_A_224_47#_c_226_n N_Z_c_545_n 0.141196f $X=3.945 $Y=1.16 $X2=0 $Y2=0
cc_207 N_A_224_47#_c_228_n N_Z_c_545_n 0.00713085f $X=3.97 $Y=1.035 $X2=0 $Y2=0
cc_208 N_A_224_47#_c_223_n N_VGND_c_606_n 0.0232822f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_209 N_A_224_47#_c_214_n N_VGND_c_607_n 0.00877186f $X=2.45 $Y=0.96 $X2=0
+ $Y2=0
cc_210 N_A_224_47#_c_217_n N_VGND_c_607_n 0.00170602f $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_211 N_A_224_47#_c_217_n N_VGND_c_608_n 0.00428022f $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_212 N_A_224_47#_c_219_n N_VGND_c_608_n 0.00199015f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_213 N_A_224_47#_c_217_n N_VGND_c_609_n 6.77692e-19 $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_214 N_A_224_47#_c_219_n N_VGND_c_609_n 0.0100391f $X=3.44 $Y=0.96 $X2=0 $Y2=0
cc_215 N_A_224_47#_c_229_n N_VGND_c_609_n 0.00317372f $X=3.97 $Y=0.96 $X2=0
+ $Y2=0
cc_216 N_A_224_47#_c_214_n N_VGND_c_611_n 0.00341689f $X=2.45 $Y=0.96 $X2=0
+ $Y2=0
cc_217 N_A_224_47#_c_223_n N_VGND_c_611_n 0.0430896f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_218 N_A_224_47#_c_229_n N_VGND_c_612_n 0.00428022f $X=3.97 $Y=0.96 $X2=0
+ $Y2=0
cc_219 N_A_224_47#_M1009_d N_VGND_c_613_n 0.00294208f $X=1.12 $Y=0.235 $X2=0
+ $Y2=0
cc_220 N_A_224_47#_c_214_n N_VGND_c_613_n 0.00540327f $X=2.45 $Y=0.96 $X2=0
+ $Y2=0
cc_221 N_A_224_47#_c_217_n N_VGND_c_613_n 0.00605834f $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_222 N_A_224_47#_c_219_n N_VGND_c_613_n 0.00278819f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_223 N_A_224_47#_c_223_n N_VGND_c_613_n 0.0238257f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_224 N_A_224_47#_c_229_n N_VGND_c_613_n 0.00611632f $X=3.97 $Y=0.96 $X2=0
+ $Y2=0
cc_225 N_A_224_47#_c_223_n N_A_413_47#_c_685_n 0.0298781f $X=1.55 $Y=0.425 $X2=0
+ $Y2=0
cc_226 N_A_224_47#_c_224_n N_A_413_47#_c_685_n 0.00484604f $X=1.687 $Y=1.025
+ $X2=0 $Y2=0
cc_227 N_A_224_47#_c_214_n N_A_413_47#_c_690_n 0.0129432f $X=2.45 $Y=0.96 $X2=0
+ $Y2=0
cc_228 N_A_224_47#_c_215_n N_A_413_47#_c_690_n 0.00393903f $X=2.895 $Y=1.035
+ $X2=0 $Y2=0
cc_229 N_A_224_47#_c_217_n N_A_413_47#_c_690_n 0.0124691f $X=2.97 $Y=0.96 $X2=0
+ $Y2=0
cc_230 N_A_224_47#_c_226_n N_A_413_47#_c_690_n 0.0450705f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_224_47#_c_224_n N_A_413_47#_c_686_n 0.0174646f $X=1.687 $Y=1.025
+ $X2=0 $Y2=0
cc_232 N_A_224_47#_c_226_n N_A_413_47#_c_686_n 0.0256849f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_233 N_A_224_47#_c_219_n N_A_413_47#_c_696_n 0.00408153f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_234 N_A_224_47#_c_218_n N_A_413_47#_c_697_n 2.04719e-19 $X=3.365 $Y=1.035
+ $X2=0 $Y2=0
cc_235 N_A_224_47#_c_219_n N_A_413_47#_c_697_n 0.011362f $X=3.44 $Y=0.96 $X2=0
+ $Y2=0
cc_236 N_A_224_47#_c_220_n N_A_413_47#_c_697_n 0.00290244f $X=3.78 $Y=1.035
+ $X2=0 $Y2=0
cc_237 N_A_224_47#_c_226_n N_A_413_47#_c_697_n 0.0536423f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_238 N_A_224_47#_c_228_n N_A_413_47#_c_697_n 0.00311914f $X=3.97 $Y=1.035
+ $X2=0 $Y2=0
cc_239 N_A_224_47#_c_229_n N_A_413_47#_c_697_n 0.0122701f $X=3.97 $Y=0.96 $X2=0
+ $Y2=0
cc_240 N_A_224_47#_c_218_n N_A_413_47#_c_703_n 0.00279027f $X=3.365 $Y=1.035
+ $X2=0 $Y2=0
cc_241 N_A_224_47#_c_226_n N_A_413_47#_c_703_n 0.012344f $X=3.945 $Y=1.16 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_323_n N_VPWR_c_408_n 0.0484717f $X=0.215 $Y=1.895 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_316_n N_VPWR_c_408_n 0.00679447f $X=4.65 $Y=1.19 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_324_n N_VPWR_c_414_n 0.0182137f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_319_n N_VPWR_c_415_n 0.00429453f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_320_n N_VPWR_c_415_n 0.00429453f $X=4.945 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_27_47#_c_321_n N_VPWR_c_415_n 0.00429453f $X=5.415 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_322_n N_VPWR_c_415_n 0.00429453f $X=5.885 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_M1007_s N_VPWR_c_407_n 0.00425811f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_319_n N_VPWR_c_407_n 0.00743756f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_c_320_n N_VPWR_c_407_n 0.00606499f $X=4.945 $Y=1.41 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_321_n N_VPWR_c_407_n 0.00606499f $X=5.415 $Y=1.41 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_322_n N_VPWR_c_407_n 0.00702766f $X=5.885 $Y=1.41 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_324_n N_VPWR_c_407_n 0.00993674f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_319_n N_A_340_309#_c_487_n 0.0345078f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_320_n N_A_340_309#_c_487_n 0.0206842f $X=4.945 $Y=1.41 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_c_321_n N_A_340_309#_c_487_n 0.0206878f $X=5.415 $Y=1.41 $X2=0
+ $Y2=0
cc_258 N_A_27_47#_c_322_n N_A_340_309#_c_487_n 0.0206878f $X=5.885 $Y=1.41 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1001_g N_Z_c_561_n 0.00331756f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_27_47#_M1003_g N_Z_c_561_n 0.0105863f $X=4.92 $Y=0.56 $X2=0 $Y2=0
cc_261 N_A_27_47#_M1010_g N_Z_c_561_n 0.0106269f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_262 N_A_27_47#_M1019_g N_Z_c_561_n 0.0130285f $X=5.91 $Y=0.56 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_327_n N_Z_c_561_n 0.00193698f $X=4.795 $Y=1.19 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_316_n N_Z_c_561_n 8.60175e-19 $X=4.65 $Y=1.19 $X2=0 $Y2=0
cc_265 N_A_27_47#_c_317_n N_Z_c_561_n 0.0905992f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_318_n N_Z_c_561_n 0.0101976f $X=5.885 $Y=1.217 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_322_n Z 0.00128553f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_27_47#_M1019_g Z 0.0187418f $X=5.91 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_317_n Z 0.0202582f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_319_n N_Z_c_545_n 0.0168017f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_320_n N_Z_c_545_n 0.0135493f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_321_n N_Z_c_545_n 0.0136002f $X=5.415 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_27_47#_c_322_n N_Z_c_545_n 0.0165123f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_27_47#_c_316_n N_Z_c_545_n 0.0775735f $X=4.65 $Y=1.19 $X2=0 $Y2=0
cc_275 N_A_27_47#_c_317_n N_Z_c_545_n 0.113472f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_276 N_A_27_47#_c_318_n N_Z_c_545_n 0.0206381f $X=5.885 $Y=1.217 $X2=0 $Y2=0
cc_277 N_A_27_47#_c_316_n N_VGND_c_606_n 0.00657391f $X=4.65 $Y=1.19 $X2=0 $Y2=0
cc_278 N_A_27_47#_c_313_n N_VGND_c_610_n 0.0154729f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_279 N_A_27_47#_M1001_g N_VGND_c_612_n 0.00357877f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A_27_47#_M1003_g N_VGND_c_612_n 0.00357877f $X=4.92 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_27_47#_M1010_g N_VGND_c_612_n 0.00357877f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_27_47#_M1019_g N_VGND_c_612_n 0.00357877f $X=5.91 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1018_s N_VGND_c_613_n 0.00388065f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_284 N_A_27_47#_M1001_g N_VGND_c_613_n 0.00570108f $X=4.45 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_27_47#_M1003_g N_VGND_c_613_n 0.00548399f $X=4.92 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_27_47#_M1010_g N_VGND_c_613_n 0.00560377f $X=5.39 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_27_47#_M1019_g N_VGND_c_613_n 0.00648381f $X=5.91 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_313_n N_VGND_c_613_n 0.00980171f $X=0.26 $Y=0.445 $X2=0
+ $Y2=0
cc_289 N_A_27_47#_c_316_n N_A_413_47#_c_690_n 0.00417969f $X=4.65 $Y=1.19 $X2=0
+ $Y2=0
cc_290 N_A_27_47#_c_316_n N_A_413_47#_c_686_n 0.00203076f $X=4.65 $Y=1.19 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_316_n N_A_413_47#_c_697_n 0.00958757f $X=4.65 $Y=1.19 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_M1001_g N_A_413_47#_c_687_n 0.011519f $X=4.45 $Y=0.56 $X2=0
+ $Y2=0
cc_293 N_A_27_47#_M1003_g N_A_413_47#_c_687_n 0.00847746f $X=4.92 $Y=0.56 $X2=0
+ $Y2=0
cc_294 N_A_27_47#_M1010_g N_A_413_47#_c_687_n 0.00876725f $X=5.39 $Y=0.56 $X2=0
+ $Y2=0
cc_295 N_A_27_47#_M1019_g N_A_413_47#_c_687_n 0.00876725f $X=5.91 $Y=0.56 $X2=0
+ $Y2=0
cc_296 N_A_27_47#_c_317_n N_A_413_47#_c_687_n 0.00382597f $X=5.77 $Y=1.16 $X2=0
+ $Y2=0
cc_297 N_A_27_47#_c_316_n N_A_413_47#_c_703_n 0.00104304f $X=4.65 $Y=1.19 $X2=0
+ $Y2=0
cc_298 N_VPWR_c_407_n N_A_340_309#_M1005_d 0.00394443f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_299 N_VPWR_c_407_n N_A_340_309#_M1008_d 0.00427219f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_300 N_VPWR_c_407_n N_A_340_309#_M1016_d 0.00690528f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_407_n N_A_340_309#_M1004_d 0.00231289f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_302 N_VPWR_c_407_n N_A_340_309#_M1013_d 0.00233941f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_303 N_VPWR_c_410_n N_A_340_309#_c_485_n 0.0145727f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_411_n N_A_340_309#_c_485_n 0.0168251f $X=2.08 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_407_n N_A_340_309#_c_485_n 0.00929827f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_409_n N_A_340_309#_c_514_n 0.011503f $X=3.235 $Y=2.36 $X2=0
+ $Y2=0
cc_307 N_VPWR_c_410_n N_A_340_309#_c_514_n 0.0116296f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_412_n N_A_340_309#_c_514_n 0.0116627f $X=3.07 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_407_n N_A_340_309#_c_514_n 0.00644035f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_310 N_VPWR_M1005_s N_A_340_309#_c_486_n 0.00350267f $X=2.15 $Y=1.545 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_410_n N_A_340_309#_c_486_n 0.0198898f $X=2.295 $Y=2.36 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_411_n N_A_340_309#_c_486_n 0.00201842f $X=2.08 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_412_n N_A_340_309#_c_486_n 0.00289521f $X=3.07 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_407_n N_A_340_309#_c_486_n 0.00882418f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_409_n N_A_340_309#_c_493_n 0.0127938f $X=3.235 $Y=2.36 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_415_n N_A_340_309#_c_493_n 0.166804f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_317 N_VPWR_c_407_n N_A_340_309#_c_493_n 0.0985906f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_M1012_s N_A_340_309#_c_494_n 0.0035106f $X=3.09 $Y=1.545 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_409_n N_A_340_309#_c_494_n 0.0161796f $X=3.235 $Y=2.36 $X2=0
+ $Y2=0
cc_320 N_VPWR_c_412_n N_A_340_309#_c_494_n 0.00338887f $X=3.07 $Y=2.72 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_415_n N_A_340_309#_c_494_n 0.00338887f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_407_n N_A_340_309#_c_494_n 0.0126775f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_407_n N_Z_M1000_s 0.00232895f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_407_n N_Z_M1011_s 0.00232895f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_325 N_VPWR_M1005_s N_Z_c_545_n 0.00189989f $X=2.15 $Y=1.545 $X2=0 $Y2=0
cc_326 N_VPWR_M1012_s N_Z_c_545_n 0.00190453f $X=3.09 $Y=1.545 $X2=0 $Y2=0
cc_327 N_A_340_309#_c_487_n N_Z_M1000_s 0.0034706f $X=6.12 $Y=2.02 $X2=0 $Y2=0
cc_328 N_A_340_309#_c_487_n N_Z_M1011_s 0.00349548f $X=6.12 $Y=2.02 $X2=0 $Y2=0
cc_329 N_A_340_309#_M1013_d Z 0.0032362f $X=5.975 $Y=1.485 $X2=0 $Y2=0
cc_330 N_A_340_309#_c_487_n Z 0.0160143f $X=6.12 $Y=2.02 $X2=0 $Y2=0
cc_331 N_A_340_309#_M1008_d N_Z_c_545_n 0.0018675f $X=2.62 $Y=1.545 $X2=0 $Y2=0
cc_332 N_A_340_309#_M1016_d N_Z_c_545_n 0.0137539f $X=3.56 $Y=1.545 $X2=0 $Y2=0
cc_333 N_A_340_309#_M1004_d N_Z_c_545_n 0.00190453f $X=5.035 $Y=1.485 $X2=0
+ $Y2=0
cc_334 N_A_340_309#_M1013_d N_Z_c_545_n 7.79125e-19 $X=5.975 $Y=1.485 $X2=0
+ $Y2=0
cc_335 N_A_340_309#_c_486_n N_Z_c_545_n 0.05074f $X=2.85 $Y=2 $X2=0 $Y2=0
cc_336 N_A_340_309#_c_494_n N_Z_c_545_n 0.199569f $X=3.62 $Y=2.18 $X2=0 $Y2=0
cc_337 N_Z_c_542_n N_VGND_c_612_n 0.00105876f $X=6.22 $Y=0.855 $X2=0 $Y2=0
cc_338 N_Z_M1001_d N_VGND_c_613_n 0.00256987f $X=4.525 $Y=0.235 $X2=0 $Y2=0
cc_339 N_Z_M1010_d N_VGND_c_613_n 0.00297142f $X=5.465 $Y=0.235 $X2=0 $Y2=0
cc_340 N_Z_c_542_n N_VGND_c_613_n 0.00200114f $X=6.22 $Y=0.855 $X2=0 $Y2=0
cc_341 N_Z_c_561_n N_A_413_47#_M1003_s 0.00402091f $X=6.105 $Y=0.735 $X2=0 $Y2=0
cc_342 N_Z_c_561_n N_A_413_47#_M1019_s 0.00178753f $X=6.105 $Y=0.735 $X2=0 $Y2=0
cc_343 Z N_A_413_47#_M1019_s 4.99287e-19 $X=6.125 $Y=0.765 $X2=0 $Y2=0
cc_344 N_Z_c_542_n N_A_413_47#_M1019_s 0.00302903f $X=6.22 $Y=0.855 $X2=0 $Y2=0
cc_345 N_Z_c_545_n N_A_413_47#_c_697_n 0.00227192f $X=6.105 $Y=1.585 $X2=0 $Y2=0
cc_346 N_Z_M1001_d N_A_413_47#_c_687_n 0.00400887f $X=4.525 $Y=0.235 $X2=0 $Y2=0
cc_347 N_Z_M1010_d N_A_413_47#_c_687_n 0.00507048f $X=5.465 $Y=0.235 $X2=0 $Y2=0
cc_348 N_Z_c_561_n N_A_413_47#_c_687_n 0.0834719f $X=6.105 $Y=0.735 $X2=0 $Y2=0
cc_349 N_Z_c_542_n N_A_413_47#_c_687_n 0.0139424f $X=6.22 $Y=0.855 $X2=0 $Y2=0
cc_350 N_VGND_c_613_n N_A_413_47#_M1002_d 0.00269999f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_351 N_VGND_c_613_n N_A_413_47#_M1006_d 0.0031681f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_352 N_VGND_c_613_n N_A_413_47#_M1015_d 0.00332861f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_353 N_VGND_c_613_n N_A_413_47#_M1003_s 0.00255381f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_354 N_VGND_c_613_n N_A_413_47#_M1019_s 0.00225742f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_355 N_VGND_c_611_n N_A_413_47#_c_685_n 0.0227423f $X=2.495 $Y=0 $X2=0 $Y2=0
cc_356 N_VGND_c_613_n N_A_413_47#_c_685_n 0.0125906f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_357 N_VGND_M1002_s N_A_413_47#_c_690_n 0.00481305f $X=2.525 $Y=0.235 $X2=0
+ $Y2=0
cc_358 N_VGND_c_607_n N_A_413_47#_c_690_n 0.0219266f $X=2.71 $Y=0.36 $X2=0 $Y2=0
cc_359 N_VGND_c_608_n N_A_413_47#_c_690_n 0.00300242f $X=3.435 $Y=0 $X2=0 $Y2=0
cc_360 N_VGND_c_611_n N_A_413_47#_c_690_n 0.00234306f $X=2.495 $Y=0 $X2=0 $Y2=0
cc_361 N_VGND_c_613_n N_A_413_47#_c_690_n 0.0111856f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_362 N_VGND_c_608_n N_A_413_47#_c_696_n 0.010169f $X=3.435 $Y=0 $X2=0 $Y2=0
cc_363 N_VGND_c_609_n N_A_413_47#_c_696_n 0.0156777f $X=3.65 $Y=0.36 $X2=0 $Y2=0
cc_364 N_VGND_c_613_n N_A_413_47#_c_696_n 0.00637943f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_365 N_VGND_M1014_s N_A_413_47#_c_697_n 0.00388345f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_366 N_VGND_c_608_n N_A_413_47#_c_697_n 0.00233941f $X=3.435 $Y=0 $X2=0 $Y2=0
cc_367 N_VGND_c_609_n N_A_413_47#_c_697_n 0.0216793f $X=3.65 $Y=0.36 $X2=0 $Y2=0
cc_368 N_VGND_c_612_n N_A_413_47#_c_697_n 0.00300242f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_369 N_VGND_c_613_n N_A_413_47#_c_697_n 0.0114174f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_370 N_VGND_c_612_n N_A_413_47#_c_743_n 0.0197284f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_371 N_VGND_c_613_n N_A_413_47#_c_743_n 0.011132f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_372 N_VGND_c_612_n N_A_413_47#_c_687_n 0.11114f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_373 N_VGND_c_613_n N_A_413_47#_c_687_n 0.0702294f $X=6.21 $Y=0 $X2=0 $Y2=0
