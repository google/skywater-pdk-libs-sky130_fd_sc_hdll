* File: sky130_fd_sc_hdll__nor3b_4.pxi.spice
* Created: Wed Sep  2 08:40:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%C_N N_C_N_c_106_n N_C_N_M1001_g N_C_N_c_103_n
+ N_C_N_M1006_g C_N N_C_N_c_105_n C_N PM_SKY130_FD_SC_HDLL__NOR3B_4%C_N
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%A N_A_c_130_n N_A_M1002_g N_A_c_136_n
+ N_A_M1000_g N_A_c_131_n N_A_M1013_g N_A_c_137_n N_A_M1008_g N_A_c_132_n
+ N_A_M1019_g N_A_c_138_n N_A_M1011_g N_A_c_139_n N_A_M1017_g N_A_c_133_n
+ N_A_M1022_g A A A N_A_c_134_n A A A PM_SKY130_FD_SC_HDLL__NOR3B_4%A
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%B N_B_c_201_n N_B_M1004_g N_B_c_207_n
+ N_B_M1003_g N_B_c_202_n N_B_M1014_g N_B_c_208_n N_B_M1010_g N_B_c_203_n
+ N_B_M1021_g N_B_c_209_n N_B_M1015_g N_B_c_210_n N_B_M1020_g N_B_c_204_n
+ N_B_M1024_g B N_B_c_205_n N_B_c_206_n B PM_SKY130_FD_SC_HDLL__NOR3B_4%B
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1001_s
+ N_A_27_47#_c_275_n N_A_27_47#_M1005_g N_A_27_47#_c_287_n N_A_27_47#_M1009_g
+ N_A_27_47#_c_276_n N_A_27_47#_M1007_g N_A_27_47#_c_288_n N_A_27_47#_M1012_g
+ N_A_27_47#_c_277_n N_A_27_47#_M1016_g N_A_27_47#_c_289_n N_A_27_47#_M1018_g
+ N_A_27_47#_c_290_n N_A_27_47#_M1023_g N_A_27_47#_c_278_n N_A_27_47#_M1025_g
+ N_A_27_47#_c_279_n N_A_27_47#_c_291_n N_A_27_47#_c_292_n N_A_27_47#_c_293_n
+ N_A_27_47#_c_280_n N_A_27_47#_c_281_n N_A_27_47#_c_282_n N_A_27_47#_c_295_n
+ N_A_27_47#_c_283_n N_A_27_47#_c_284_n N_A_27_47#_c_285_n N_A_27_47#_c_333_p
+ N_A_27_47#_c_286_n PM_SKY130_FD_SC_HDLL__NOR3B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%VPWR N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1017_d N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n N_VPWR_c_433_n
+ N_VPWR_c_434_n VPWR N_VPWR_c_435_n N_VPWR_c_429_n N_VPWR_c_437_n
+ N_VPWR_c_438_n N_VPWR_c_439_n PM_SKY130_FD_SC_HDLL__NOR3B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%A_215_297# N_A_215_297#_M1000_s
+ N_A_215_297#_M1011_s N_A_215_297#_M1003_s N_A_215_297#_M1015_s
+ N_A_215_297#_c_523_n N_A_215_297#_c_522_n N_A_215_297#_c_527_n
+ N_A_215_297#_c_536_n N_A_215_297#_c_537_n N_A_215_297#_c_538_n
+ N_A_215_297#_c_539_n PM_SKY130_FD_SC_HDLL__NOR3B_4%A_215_297#
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%A_605_297# N_A_605_297#_M1003_d
+ N_A_605_297#_M1010_d N_A_605_297#_M1020_d N_A_605_297#_M1012_d
+ N_A_605_297#_M1023_d N_A_605_297#_c_571_n N_A_605_297#_c_573_n
+ N_A_605_297#_c_579_n N_A_605_297#_c_580_n N_A_605_297#_c_621_p
+ N_A_605_297#_c_570_n N_A_605_297#_c_625_p N_A_605_297#_c_597_n
+ N_A_605_297#_c_600_n N_A_605_297#_c_602_n N_A_605_297#_c_604_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_4%A_605_297#
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%Y N_Y_M1002_d N_Y_M1019_d N_Y_M1004_d
+ N_Y_M1021_d N_Y_M1005_s N_Y_M1016_s N_Y_M1009_s N_Y_M1018_s N_Y_c_646_n
+ N_Y_c_628_n N_Y_c_629_n N_Y_c_658_n N_Y_c_630_n N_Y_c_667_n N_Y_c_631_n
+ N_Y_c_674_n N_Y_c_632_n N_Y_c_677_n N_Y_c_641_n N_Y_c_633_n N_Y_c_703_n
+ N_Y_c_642_n N_Y_c_634_n N_Y_c_635_n N_Y_c_636_n N_Y_c_637_n N_Y_c_638_n
+ N_Y_c_643_n N_Y_c_639_n N_Y_c_644_n Y Y PM_SKY130_FD_SC_HDLL__NOR3B_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR3B_4%VGND N_VGND_M1006_d N_VGND_M1013_s
+ N_VGND_M1022_s N_VGND_M1014_s N_VGND_M1024_s N_VGND_M1007_d N_VGND_M1025_d
+ N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n N_VGND_c_794_n N_VGND_c_795_n
+ N_VGND_c_796_n N_VGND_c_797_n N_VGND_c_798_n N_VGND_c_799_n N_VGND_c_800_n
+ N_VGND_c_801_n N_VGND_c_802_n N_VGND_c_803_n N_VGND_c_804_n N_VGND_c_805_n
+ VGND N_VGND_c_806_n N_VGND_c_807_n N_VGND_c_808_n N_VGND_c_809_n
+ N_VGND_c_810_n N_VGND_c_811_n VGND PM_SKY130_FD_SC_HDLL__NOR3B_4%VGND
cc_1 VNB N_C_N_c_103_n 0.0216587f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=0.995
cc_2 VNB C_N 0.00777182f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_N_c_105_n 0.0422638f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_4 VNB N_A_c_130_n 0.0165954f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_5 VNB N_A_c_131_n 0.0167587f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_c_132_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_7 VNB N_A_c_133_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_c_134_n 0.08147f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A 0.008141f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B_c_201_n 0.021971f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_11 VNB N_B_c_202_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_12 VNB N_B_c_203_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_13 VNB N_B_c_204_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B_c_205_n 0.00314705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B_c_206_n 0.0815017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_275_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_17 VNB N_A_27_47#_c_276_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.54 $Y2=1.202
cc_18 VNB N_A_27_47#_c_277_n 0.0171999f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_278_n 0.0201206f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_279_n 0.0184844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_280_n 9.39746e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_281_n 0.00911773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_282_n 0.00773515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_27_47#_c_283_n 3.4592e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_27_47#_c_284_n 0.00306312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_27_47#_c_285_n 4.00308e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_27_47#_c_286_n 0.0765151f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_429_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_628_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_629_n 0.00335832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_630_n 0.0108431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_631_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_632_n 0.00331095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_633_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_634_n 0.0137904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_635_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_636_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_637_n 0.00277435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_638_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_639_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB Y 0.0227699f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_791_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_792_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_793_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_794_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_795_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_796_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_797_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_798_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_799_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_800_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_801_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_802_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_803_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_804_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_805_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_806_n 0.0128319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_807_n 0.35606f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_808_n 0.0226019f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_809_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_810_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_811_n 0.0208752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VPB N_C_N_c_106_n 0.0204401f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_64 VPB N_C_N_c_105_n 0.0177286f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_65 VPB N_A_c_136_n 0.0160705f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_66 VPB N_A_c_137_n 0.0159553f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_67 VPB N_A_c_138_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_c_139_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_c_134_n 0.0483566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_B_c_207_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=0.995
cc_71 VPB N_B_c_208_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_72 VPB N_B_c_209_n 0.0159557f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_B_c_210_n 0.0160715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B_c_206_n 0.0482824f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_47#_c_287_n 0.0164062f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_76 VPB N_A_27_47#_c_288_n 0.0159548f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_27_47#_c_289_n 0.015956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_27_47#_c_290_n 0.0191692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_27_47#_c_291_n 0.0089398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_27_47#_c_292_n 0.0317613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_27_47#_c_293_n 8.45061e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_27_47#_c_282_n 0.00270512f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_27_47#_c_295_n 0.0289766f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_27_47#_c_283_n 0.00271474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_27_47#_c_286_n 0.0464481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_430_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.18
cc_87 VPB N_VPWR_c_431_n 0.0187819f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_432_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_433_n 0.0180033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_434_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_435_n 0.108918f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_429_n 0.0580545f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_437_n 0.0240584f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_438_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_439_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_215_297#_c_522_n 0.0081428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_605_297#_c_570_n 0.00692367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_641_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_Y_c_642_n 0.0187729f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_Y_c_643_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_Y_c_644_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB Y 0.00874295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 N_C_N_c_103_n N_A_c_130_n 0.0209274f $X=0.54 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_104 N_C_N_c_106_n N_A_c_136_n 0.021612f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_105 N_C_N_c_105_n N_A_c_134_n 0.0209274f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_106 C_N N_A_27_47#_c_291_n 0.0241321f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_107 N_C_N_c_105_n N_A_27_47#_c_291_n 0.00721245f $X=0.515 $Y=1.202 $X2=0
+ $Y2=0
cc_108 N_C_N_c_106_n N_A_27_47#_c_293_n 0.0176372f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_109 C_N N_A_27_47#_c_293_n 0.0027931f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_110 N_C_N_c_105_n N_A_27_47#_c_293_n 8.59828e-19 $X=0.515 $Y=1.202 $X2=0
+ $Y2=0
cc_111 N_C_N_c_103_n N_A_27_47#_c_280_n 0.0118069f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_112 N_C_N_c_105_n N_A_27_47#_c_280_n 6.6226e-19 $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_113 C_N N_A_27_47#_c_281_n 0.0272978f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_114 N_C_N_c_105_n N_A_27_47#_c_281_n 0.0086718f $X=0.515 $Y=1.202 $X2=0 $Y2=0
cc_115 N_C_N_c_106_n N_A_27_47#_c_282_n 0.0010572f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_116 N_C_N_c_103_n N_A_27_47#_c_282_n 0.00911819f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_117 C_N N_A_27_47#_c_282_n 0.0129457f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_118 N_C_N_c_106_n N_VPWR_c_430_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_119 N_C_N_c_106_n N_VPWR_c_429_n 0.0133639f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_120 N_C_N_c_106_n N_VPWR_c_437_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_121 N_C_N_c_103_n N_Y_c_646_n 5.32212e-19 $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_122 N_C_N_c_103_n N_VGND_c_791_n 0.00268723f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_123 N_C_N_c_103_n N_VGND_c_807_n 0.00695342f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_124 N_C_N_c_103_n N_VGND_c_808_n 0.00439206f $X=0.54 $Y=0.995 $X2=0 $Y2=0
cc_125 A N_B_c_205_n 0.00803268f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_126 A N_B_c_206_n 0.00137056f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_127 N_A_c_130_n N_A_27_47#_c_280_n 7.75269e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_130_n N_A_27_47#_c_282_n 0.00970477f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_c_136_n N_A_27_47#_c_282_n 0.0010572f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_130 A N_A_27_47#_c_282_n 0.00914671f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_131 N_A_c_136_n N_A_27_47#_c_295_n 0.0215889f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_137_n N_A_27_47#_c_295_n 0.01191f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_138_n N_A_27_47#_c_295_n 0.01191f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_139_n N_A_27_47#_c_295_n 0.0139099f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_134_n N_A_27_47#_c_295_n 0.0236216f $X=2.395 $Y=1.202 $X2=0 $Y2=0
cc_136 A N_A_27_47#_c_295_n 0.112368f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_137 N_A_c_136_n N_VPWR_c_430_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_136_n N_VPWR_c_431_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_137_n N_VPWR_c_431_n 0.0053025f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_137_n N_VPWR_c_432_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_138_n N_VPWR_c_432_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_138_n N_VPWR_c_433_n 0.0053025f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_139_n N_VPWR_c_433_n 0.0053025f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_139_n N_VPWR_c_434_n 0.00479105f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_136_n N_VPWR_c_429_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_137_n N_VPWR_c_429_n 0.00690493f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_138_n N_VPWR_c_429_n 0.00690493f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_139_n N_VPWR_c_429_n 0.00818727f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_137_n N_A_215_297#_c_523_n 0.0120199f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_138_n N_A_215_297#_c_523_n 0.0120199f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_139_n N_A_215_297#_c_522_n 0.0140197f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_c_130_n N_Y_c_646_n 0.00644736f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_131_n N_Y_c_646_n 0.00686626f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_132_n N_Y_c_646_n 5.45498e-19 $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_131_n N_Y_c_628_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A_c_132_n N_Y_c_628_n 0.00901745f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_c_134_n N_Y_c_628_n 0.00345541f $X=2.395 $Y=1.202 $X2=0 $Y2=0
cc_158 A N_Y_c_628_n 0.0398926f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_159 N_A_c_130_n N_Y_c_629_n 0.00300274f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_c_131_n N_Y_c_629_n 0.00116636f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_c_134_n N_Y_c_629_n 0.00410792f $X=2.395 $Y=1.202 $X2=0 $Y2=0
cc_162 A N_Y_c_629_n 0.0141285f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_163 N_A_c_131_n N_Y_c_658_n 5.24597e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_132_n N_Y_c_658_n 0.00651696f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_c_133_n N_Y_c_630_n 0.01289f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_166 A N_Y_c_630_n 0.0329378f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_167 N_A_c_132_n N_Y_c_635_n 0.00119564f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_c_134_n N_Y_c_635_n 0.00486271f $X=2.395 $Y=1.202 $X2=0 $Y2=0
cc_169 A N_Y_c_635_n 0.030835f $X=2.535 $Y=1.19 $X2=0 $Y2=0
cc_170 N_A_c_130_n N_VGND_c_791_n 0.00268723f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_c_130_n N_VGND_c_792_n 0.00541359f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_131_n N_VGND_c_792_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_131_n N_VGND_c_793_n 0.00379224f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_c_132_n N_VGND_c_793_n 0.00276126f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_130_n N_VGND_c_807_n 0.00965571f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_131_n N_VGND_c_807_n 0.006093f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_132_n N_VGND_c_807_n 0.00608558f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_133_n N_VGND_c_807_n 0.00745263f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_132_n N_VGND_c_810_n 0.00423334f $X=1.9 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_133_n N_VGND_c_810_n 0.00437852f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_133_n N_VGND_c_811_n 0.00481673f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B_c_204_n N_A_27_47#_c_275_n 0.0231917f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_210_n N_A_27_47#_c_287_n 0.0208337f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B_c_207_n N_A_27_47#_c_295_n 0.0139099f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B_c_208_n N_A_27_47#_c_295_n 0.01191f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_209_n N_A_27_47#_c_295_n 0.01191f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_210_n N_A_27_47#_c_295_n 0.0165082f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_205_n N_A_27_47#_c_295_n 0.100766f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_189 N_B_c_206_n N_A_27_47#_c_295_n 0.0229514f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_190 N_B_c_210_n N_A_27_47#_c_283_n 0.00100486f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_206_n N_A_27_47#_c_283_n 0.00290678f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_192 N_B_c_205_n N_A_27_47#_c_284_n 0.0125716f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_193 N_B_c_206_n N_A_27_47#_c_284_n 0.00238026f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_194 N_B_c_206_n N_A_27_47#_c_286_n 0.0231917f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_195 N_B_c_207_n N_VPWR_c_434_n 0.00213395f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_207_n N_VPWR_c_435_n 0.00429453f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_208_n N_VPWR_c_435_n 0.00429453f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B_c_209_n N_VPWR_c_435_n 0.00429453f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_210_n N_VPWR_c_435_n 0.00429453f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_207_n N_VPWR_c_429_n 0.00734734f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_208_n N_VPWR_c_429_n 0.00606499f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_209_n N_VPWR_c_429_n 0.00606499f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_210_n N_VPWR_c_429_n 0.00609021f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_207_n N_A_215_297#_c_522_n 0.0128257f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_c_208_n N_A_215_297#_c_527_n 0.0107828f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_209_n N_A_215_297#_c_527_n 0.0107828f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_207_n N_A_605_297#_c_571_n 0.00991367f $X=3.385 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_208_n N_A_605_297#_c_571_n 0.00991367f $X=3.855 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_209_n N_A_605_297#_c_573_n 0.00995673f $X=4.325 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_210_n N_A_605_297#_c_573_n 0.0115669f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_201_n N_Y_c_630_n 0.0109318f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B_c_205_n N_Y_c_630_n 0.00826974f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_213 N_B_c_201_n N_Y_c_667_n 0.0110728f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_202_n N_Y_c_667_n 0.00686626f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_203_n N_Y_c_667_n 5.45498e-19 $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_216 N_B_c_202_n N_Y_c_631_n 0.00901745f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_217 N_B_c_203_n N_Y_c_631_n 0.00901745f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_218 N_B_c_205_n N_Y_c_631_n 0.0398926f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_219 N_B_c_206_n N_Y_c_631_n 0.00345541f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_220 N_B_c_202_n N_Y_c_674_n 5.24597e-19 $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B_c_203_n N_Y_c_674_n 0.00651696f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B_c_204_n N_Y_c_632_n 0.012453f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B_c_204_n N_Y_c_677_n 5.32212e-19 $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_224 N_B_c_201_n N_Y_c_636_n 0.00116636f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_225 N_B_c_202_n N_Y_c_636_n 0.00116636f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_226 N_B_c_205_n N_Y_c_636_n 0.0307014f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_c_206_n N_Y_c_636_n 0.00358305f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_228 N_B_c_203_n N_Y_c_637_n 0.00119564f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_229 N_B_c_205_n N_Y_c_637_n 0.0287969f $X=4.23 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B_c_206_n N_Y_c_637_n 0.00486271f $X=4.795 $Y=1.202 $X2=0 $Y2=0
cc_231 N_B_c_202_n N_VGND_c_794_n 0.00379224f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B_c_203_n N_VGND_c_794_n 0.00276126f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_204_n N_VGND_c_795_n 0.00268723f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_201_n N_VGND_c_798_n 0.00423334f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B_c_202_n N_VGND_c_798_n 0.00423334f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_203_n N_VGND_c_800_n 0.00423334f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_204_n N_VGND_c_800_n 0.00437852f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_201_n N_VGND_c_807_n 0.00716687f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B_c_202_n N_VGND_c_807_n 0.006093f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B_c_203_n N_VGND_c_807_n 0.00608558f $X=4.3 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B_c_204_n N_VGND_c_807_n 0.00615622f $X=4.82 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B_c_201_n N_VGND_c_811_n 0.00481673f $X=3.36 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_333_p N_VPWR_M1001_d 0.00188126f $X=0.75 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_244 N_A_27_47#_c_295_n N_VPWR_M1008_d 0.00187547f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_245 N_A_27_47#_c_295_n N_VPWR_M1017_d 0.00295153f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_246 N_A_27_47#_c_333_p N_VPWR_c_430_n 0.0153275f $X=0.75 $Y=1.54 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_287_n N_VPWR_c_435_n 0.00429453f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_27_47#_c_288_n N_VPWR_c_435_n 0.00429453f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_27_47#_c_289_n N_VPWR_c_435_n 0.00429453f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_27_47#_c_290_n N_VPWR_c_435_n 0.00429453f $X=6.675 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_27_47#_M1001_s N_VPWR_c_429_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_287_n N_VPWR_c_429_n 0.00609021f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_253 N_A_27_47#_c_288_n N_VPWR_c_429_n 0.00606499f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_c_289_n N_VPWR_c_429_n 0.00606499f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_c_290_n N_VPWR_c_429_n 0.00711127f $X=6.675 $Y=1.41 $X2=0
+ $Y2=0
cc_256 N_A_27_47#_c_292_n N_VPWR_c_429_n 0.0112839f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_292_n N_VPWR_c_437_n 0.0193827f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_295_n N_A_215_297#_M1000_s 0.00187091f $X=4.985 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_259 N_A_27_47#_c_295_n N_A_215_297#_M1011_s 0.00187091f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_260 N_A_27_47#_c_295_n N_A_215_297#_M1003_s 0.00187091f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_261 N_A_27_47#_c_295_n N_A_215_297#_M1015_s 0.00187091f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_262 N_A_27_47#_c_295_n N_A_215_297#_c_523_n 0.0371166f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_295_n N_A_215_297#_c_522_n 0.0756062f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_295_n N_A_215_297#_c_527_n 0.0371166f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_c_295_n N_A_215_297#_c_536_n 0.0143018f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_c_295_n N_A_215_297#_c_537_n 0.0143018f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_295_n N_A_215_297#_c_538_n 0.0135159f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_295_n N_A_215_297#_c_539_n 0.0135159f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_295_n N_A_605_297#_M1003_d 0.00295153f $X=4.985 $Y=1.54
+ $X2=-0.19 $Y2=-0.24
cc_270 N_A_27_47#_c_295_n N_A_605_297#_M1010_d 0.00187547f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_271 N_A_27_47#_c_295_n N_A_605_297#_M1020_d 0.00231948f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_272 N_A_27_47#_c_295_n N_A_605_297#_c_573_n 0.00386609f $X=4.985 $Y=1.54
+ $X2=0 $Y2=0
cc_273 N_A_27_47#_c_295_n N_A_605_297#_c_579_n 0.0152503f $X=4.985 $Y=1.54 $X2=0
+ $Y2=0
cc_274 N_A_27_47#_c_287_n N_A_605_297#_c_580_n 0.0143578f $X=5.265 $Y=1.41 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_c_288_n N_A_605_297#_c_580_n 0.01161f $X=5.735 $Y=1.41 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_c_289_n N_A_605_297#_c_570_n 0.01161f $X=6.205 $Y=1.41 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_c_290_n N_A_605_297#_c_570_n 0.01161f $X=6.675 $Y=1.41 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_280_n N_Y_c_629_n 0.00808484f $X=0.665 $Y=0.82 $X2=0 $Y2=0
cc_279 N_A_27_47#_c_295_n N_Y_c_629_n 0.00717391f $X=4.985 $Y=1.54 $X2=0 $Y2=0
cc_280 N_A_27_47#_c_295_n N_Y_c_630_n 0.0172574f $X=4.985 $Y=1.54 $X2=0 $Y2=0
cc_281 N_A_27_47#_c_275_n N_Y_c_632_n 0.00865686f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_27_47#_c_295_n N_Y_c_632_n 0.0075073f $X=4.985 $Y=1.54 $X2=0 $Y2=0
cc_283 N_A_27_47#_c_284_n N_Y_c_632_n 0.0141654f $X=5.155 $Y=1.18 $X2=0 $Y2=0
cc_284 N_A_27_47#_c_285_n N_Y_c_632_n 0.00899944f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_285 N_A_27_47#_c_275_n N_Y_c_677_n 0.00644736f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_27_47#_c_276_n N_Y_c_677_n 0.00686626f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_27_47#_c_277_n N_Y_c_677_n 5.45498e-19 $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_27_47#_c_288_n N_Y_c_641_n 0.0128188f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_289_n N_Y_c_641_n 0.0128795f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_285_n N_Y_c_641_n 0.0486996f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_27_47#_c_286_n N_Y_c_641_n 0.00864922f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_292 N_A_27_47#_c_276_n N_Y_c_633_n 0.00901745f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_277_n N_Y_c_633_n 0.00901745f $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_27_47#_c_285_n N_Y_c_633_n 0.0398926f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_295 N_A_27_47#_c_286_n N_Y_c_633_n 0.00345541f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_296 N_A_27_47#_c_276_n N_Y_c_703_n 5.24597e-19 $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_27_47#_c_277_n N_Y_c_703_n 0.00651696f $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A_27_47#_c_290_n N_Y_c_642_n 0.0150911f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_299 N_A_27_47#_c_285_n N_Y_c_642_n 0.0107166f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_300 N_A_27_47#_c_286_n N_Y_c_642_n 9.33689e-19 $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_301 N_A_27_47#_c_278_n N_Y_c_634_n 0.0131856f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A_27_47#_c_285_n N_Y_c_634_n 0.00799574f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_27_47#_c_295_n N_Y_c_637_n 8.53266e-19 $X=4.985 $Y=1.54 $X2=0 $Y2=0
cc_304 N_A_27_47#_c_275_n N_Y_c_638_n 0.00116636f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_27_47#_c_276_n N_Y_c_638_n 0.00116636f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_27_47#_c_285_n N_Y_c_638_n 0.0307014f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_307 N_A_27_47#_c_286_n N_Y_c_638_n 0.00358305f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_308 N_A_27_47#_c_287_n N_Y_c_643_n 2.98195e-19 $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_27_47#_c_295_n N_Y_c_643_n 0.00226124f $X=4.985 $Y=1.54 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_285_n N_Y_c_643_n 0.0204252f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_286_n N_Y_c_643_n 0.00655199f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_277_n N_Y_c_639_n 0.00119564f $X=6.18 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_285_n N_Y_c_639_n 0.030835f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_314 N_A_27_47#_c_286_n N_Y_c_639_n 0.00486271f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_315 N_A_27_47#_c_285_n N_Y_c_644_n 0.0204252f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_316 N_A_27_47#_c_286_n N_Y_c_644_n 0.00634604f $X=6.675 $Y=1.202 $X2=0 $Y2=0
cc_317 N_A_27_47#_c_290_n Y 0.00172505f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_318 N_A_27_47#_c_278_n Y 0.0184111f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_27_47#_c_285_n Y 0.0164069f $X=6.5 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_27_47#_c_280_n N_VGND_M1006_d 0.00197558f $X=0.665 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_321 N_A_27_47#_c_280_n N_VGND_c_791_n 0.0128651f $X=0.665 $Y=0.82 $X2=0 $Y2=0
cc_322 N_A_27_47#_c_275_n N_VGND_c_795_n 0.00268723f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_323 N_A_27_47#_c_276_n N_VGND_c_796_n 0.00379224f $X=5.71 $Y=0.995 $X2=0
+ $Y2=0
cc_324 N_A_27_47#_c_277_n N_VGND_c_796_n 0.00276126f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_325 N_A_27_47#_c_278_n N_VGND_c_797_n 0.00438629f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_275_n N_VGND_c_802_n 0.00423334f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_327 N_A_27_47#_c_276_n N_VGND_c_802_n 0.00423334f $X=5.71 $Y=0.995 $X2=0
+ $Y2=0
cc_328 N_A_27_47#_c_277_n N_VGND_c_804_n 0.00423334f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_329 N_A_27_47#_c_278_n N_VGND_c_804_n 0.00437852f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_27_47#_M1006_s N_VGND_c_807_n 0.00275631f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_331 N_A_27_47#_c_275_n N_VGND_c_807_n 0.00587047f $X=5.24 $Y=0.995 $X2=0
+ $Y2=0
cc_332 N_A_27_47#_c_276_n N_VGND_c_807_n 0.006093f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_277_n N_VGND_c_807_n 0.00608558f $X=6.18 $Y=0.995 $X2=0
+ $Y2=0
cc_334 N_A_27_47#_c_278_n N_VGND_c_807_n 0.00722223f $X=6.7 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_279_n N_VGND_c_807_n 0.0128092f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_336 N_A_27_47#_c_280_n N_VGND_c_807_n 0.00563939f $X=0.665 $Y=0.82 $X2=0
+ $Y2=0
cc_337 N_A_27_47#_c_279_n N_VGND_c_808_n 0.0221262f $X=0.28 $Y=0.39 $X2=0 $Y2=0
cc_338 N_A_27_47#_c_280_n N_VGND_c_808_n 0.00248202f $X=0.665 $Y=0.82 $X2=0
+ $Y2=0
cc_339 N_VPWR_c_429_n N_A_215_297#_M1000_s 0.00310186f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_340 N_VPWR_c_429_n N_A_215_297#_M1011_s 0.00250248f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_429_n N_A_215_297#_M1003_s 0.00231289f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_429_n N_A_215_297#_M1015_s 0.00232092f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_M1008_d N_A_215_297#_c_523_n 0.00348263f $X=1.545 $Y=1.485 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_431_n N_A_215_297#_c_523_n 0.00253649f $X=1.565 $Y=2.72 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_432_n N_A_215_297#_c_523_n 0.0138782f $X=1.69 $Y=2.3 $X2=0 $Y2=0
cc_346 N_VPWR_c_433_n N_A_215_297#_c_523_n 0.00253649f $X=2.505 $Y=2.72 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_429_n N_A_215_297#_c_523_n 0.0102844f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_M1017_d N_A_215_297#_c_522_n 0.0053134f $X=2.485 $Y=1.485 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_433_n N_A_215_297#_c_522_n 0.00253649f $X=2.505 $Y=2.72 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_434_n N_A_215_297#_c_522_n 0.016717f $X=2.63 $Y=2.3 $X2=0 $Y2=0
cc_351 N_VPWR_c_435_n N_A_215_297#_c_522_n 0.0039015f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_429_n N_A_215_297#_c_522_n 0.013559f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_353 N_VPWR_c_429_n N_A_215_297#_c_527_n 0.00151263f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_431_n N_A_215_297#_c_536_n 0.0149176f $X=1.565 $Y=2.72 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_429_n N_A_215_297#_c_536_n 0.00954719f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_433_n N_A_215_297#_c_537_n 0.0149176f $X=2.505 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_c_429_n N_A_215_297#_c_537_n 0.00954719f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_429_n N_A_605_297#_M1003_d 0.00215913f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_359 N_VPWR_c_429_n N_A_605_297#_M1010_d 0.00229658f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_429_n N_A_605_297#_M1020_d 0.00231264f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_429_n N_A_605_297#_M1012_d 0.00231264f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_429_n N_A_605_297#_M1023_d 0.00217519f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_VPWR_c_435_n N_A_605_297#_c_571_n 0.0386815f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_364 N_VPWR_c_429_n N_A_605_297#_c_571_n 0.0239184f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_365 N_VPWR_c_435_n N_A_605_297#_c_573_n 0.0386815f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_366 N_VPWR_c_429_n N_A_605_297#_c_573_n 0.0239184f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_367 N_VPWR_c_435_n N_A_605_297#_c_580_n 0.0386815f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_368 N_VPWR_c_429_n N_A_605_297#_c_580_n 0.0239144f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_369 N_VPWR_c_435_n N_A_605_297#_c_570_n 0.0549564f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_370 N_VPWR_c_429_n N_A_605_297#_c_570_n 0.0335386f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_371 N_VPWR_c_434_n N_A_605_297#_c_597_n 0.0180653f $X=2.63 $Y=2.3 $X2=0 $Y2=0
cc_372 N_VPWR_c_435_n N_A_605_297#_c_597_n 0.0154343f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_373 N_VPWR_c_429_n N_A_605_297#_c_597_n 0.00938089f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_374 N_VPWR_c_435_n N_A_605_297#_c_600_n 0.0143076f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_375 N_VPWR_c_429_n N_A_605_297#_c_600_n 0.00938089f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_376 N_VPWR_c_435_n N_A_605_297#_c_602_n 0.0149886f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_377 N_VPWR_c_429_n N_A_605_297#_c_602_n 0.00962421f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_378 N_VPWR_c_435_n N_A_605_297#_c_604_n 0.0149886f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_379 N_VPWR_c_429_n N_A_605_297#_c_604_n 0.00962421f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_429_n N_Y_M1009_s 0.00232895f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_429_n N_Y_M1018_s 0.00232895f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_382 N_A_215_297#_c_522_n N_A_605_297#_M1003_d 0.0053134f $X=3.495 $Y=1.88
+ $X2=-0.19 $Y2=1.305
cc_383 N_A_215_297#_c_527_n N_A_605_297#_M1010_d 0.00348263f $X=4.435 $Y=1.88
+ $X2=0 $Y2=0
cc_384 N_A_215_297#_M1003_s N_A_605_297#_c_571_n 0.00352392f $X=3.475 $Y=1.485
+ $X2=0 $Y2=0
cc_385 N_A_215_297#_c_522_n N_A_605_297#_c_571_n 0.00625304f $X=3.495 $Y=1.88
+ $X2=0 $Y2=0
cc_386 N_A_215_297#_c_527_n N_A_605_297#_c_571_n 0.00625304f $X=4.435 $Y=1.88
+ $X2=0 $Y2=0
cc_387 N_A_215_297#_c_538_n N_A_605_297#_c_571_n 0.0126996f $X=3.62 $Y=1.88
+ $X2=0 $Y2=0
cc_388 N_A_215_297#_M1015_s N_A_605_297#_c_573_n 0.00352392f $X=4.415 $Y=1.485
+ $X2=0 $Y2=0
cc_389 N_A_215_297#_c_527_n N_A_605_297#_c_573_n 0.00625304f $X=4.435 $Y=1.88
+ $X2=0 $Y2=0
cc_390 N_A_215_297#_c_539_n N_A_605_297#_c_573_n 0.0126996f $X=4.56 $Y=1.88
+ $X2=0 $Y2=0
cc_391 N_A_215_297#_c_522_n N_A_605_297#_c_597_n 0.0157703f $X=3.495 $Y=1.88
+ $X2=0 $Y2=0
cc_392 N_A_215_297#_c_527_n N_A_605_297#_c_600_n 0.0130924f $X=4.435 $Y=1.88
+ $X2=0 $Y2=0
cc_393 N_A_605_297#_c_580_n N_Y_M1009_s 0.00352392f $X=5.845 $Y=2.38 $X2=0 $Y2=0
cc_394 N_A_605_297#_c_570_n N_Y_M1018_s 0.00352392f $X=6.785 $Y=2.38 $X2=0 $Y2=0
cc_395 N_A_605_297#_M1012_d N_Y_c_641_n 0.00187091f $X=5.825 $Y=1.485 $X2=0
+ $Y2=0
cc_396 N_A_605_297#_c_580_n N_Y_c_641_n 0.00385532f $X=5.845 $Y=2.38 $X2=0 $Y2=0
cc_397 N_A_605_297#_c_621_p N_Y_c_641_n 0.0143018f $X=5.97 $Y=1.96 $X2=0 $Y2=0
cc_398 N_A_605_297#_c_570_n N_Y_c_641_n 0.00385532f $X=6.785 $Y=2.38 $X2=0 $Y2=0
cc_399 N_A_605_297#_M1023_d N_Y_c_642_n 0.00299663f $X=6.765 $Y=1.485 $X2=0
+ $Y2=0
cc_400 N_A_605_297#_c_570_n N_Y_c_642_n 0.00385532f $X=6.785 $Y=2.38 $X2=0 $Y2=0
cc_401 N_A_605_297#_c_625_p N_Y_c_642_n 0.0183262f $X=6.91 $Y=1.96 $X2=0 $Y2=0
cc_402 N_A_605_297#_c_580_n N_Y_c_643_n 0.013395f $X=5.845 $Y=2.38 $X2=0 $Y2=0
cc_403 N_A_605_297#_c_570_n N_Y_c_644_n 0.013395f $X=6.785 $Y=2.38 $X2=0 $Y2=0
cc_404 N_Y_c_628_n N_VGND_M1013_s 0.00251047f $X=1.945 $Y=0.815 $X2=0 $Y2=0
cc_405 N_Y_c_630_n N_VGND_M1022_s 0.0108248f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_406 N_Y_c_631_n N_VGND_M1014_s 0.00251047f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_407 N_Y_c_632_n N_VGND_M1024_s 0.00162089f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_408 N_Y_c_633_n N_VGND_M1007_d 0.00251047f $X=6.225 $Y=0.815 $X2=0 $Y2=0
cc_409 N_Y_c_634_n N_VGND_M1025_d 0.00322365f $X=6.905 $Y=0.815 $X2=0 $Y2=0
cc_410 N_Y_c_646_n N_VGND_c_792_n 0.0223596f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_411 N_Y_c_628_n N_VGND_c_792_n 0.00266636f $X=1.945 $Y=0.815 $X2=0 $Y2=0
cc_412 N_Y_c_646_n N_VGND_c_793_n 0.0183628f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_413 N_Y_c_628_n N_VGND_c_793_n 0.0127273f $X=1.945 $Y=0.815 $X2=0 $Y2=0
cc_414 N_Y_c_667_n N_VGND_c_794_n 0.0183628f $X=3.62 $Y=0.39 $X2=0 $Y2=0
cc_415 N_Y_c_631_n N_VGND_c_794_n 0.0127273f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_416 N_Y_c_632_n N_VGND_c_795_n 0.0122559f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_417 N_Y_c_677_n N_VGND_c_796_n 0.0183628f $X=5.5 $Y=0.39 $X2=0 $Y2=0
cc_418 N_Y_c_633_n N_VGND_c_796_n 0.0127273f $X=6.225 $Y=0.815 $X2=0 $Y2=0
cc_419 N_Y_c_634_n N_VGND_c_797_n 0.0133978f $X=6.905 $Y=0.815 $X2=0 $Y2=0
cc_420 N_Y_c_630_n N_VGND_c_798_n 0.00198695f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_421 N_Y_c_667_n N_VGND_c_798_n 0.0223596f $X=3.62 $Y=0.39 $X2=0 $Y2=0
cc_422 N_Y_c_631_n N_VGND_c_798_n 0.00266636f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_423 N_Y_c_631_n N_VGND_c_800_n 0.00198695f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_424 N_Y_c_674_n N_VGND_c_800_n 0.0231806f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_425 N_Y_c_632_n N_VGND_c_800_n 0.00254521f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_426 N_Y_c_632_n N_VGND_c_802_n 0.00198695f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_427 N_Y_c_677_n N_VGND_c_802_n 0.0223596f $X=5.5 $Y=0.39 $X2=0 $Y2=0
cc_428 N_Y_c_633_n N_VGND_c_802_n 0.00266636f $X=6.225 $Y=0.815 $X2=0 $Y2=0
cc_429 N_Y_c_633_n N_VGND_c_804_n 0.00198695f $X=6.225 $Y=0.815 $X2=0 $Y2=0
cc_430 N_Y_c_703_n N_VGND_c_804_n 0.0231806f $X=6.44 $Y=0.39 $X2=0 $Y2=0
cc_431 N_Y_c_634_n N_VGND_c_804_n 0.00254521f $X=6.905 $Y=0.815 $X2=0 $Y2=0
cc_432 N_Y_c_634_n N_VGND_c_806_n 0.00420964f $X=6.905 $Y=0.815 $X2=0 $Y2=0
cc_433 N_Y_M1002_d N_VGND_c_807_n 0.0025535f $X=1.035 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Y_M1019_d N_VGND_c_807_n 0.00304143f $X=1.975 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1004_d N_VGND_c_807_n 0.0025535f $X=3.435 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_M1021_d N_VGND_c_807_n 0.00304143f $X=4.375 $Y=0.235 $X2=0 $Y2=0
cc_437 N_Y_M1005_s N_VGND_c_807_n 0.0025535f $X=5.315 $Y=0.235 $X2=0 $Y2=0
cc_438 N_Y_M1016_s N_VGND_c_807_n 0.00304143f $X=6.255 $Y=0.235 $X2=0 $Y2=0
cc_439 N_Y_c_646_n N_VGND_c_807_n 0.0141302f $X=1.22 $Y=0.39 $X2=0 $Y2=0
cc_440 N_Y_c_628_n N_VGND_c_807_n 0.00972452f $X=1.945 $Y=0.815 $X2=0 $Y2=0
cc_441 N_Y_c_658_n N_VGND_c_807_n 0.0143352f $X=2.16 $Y=0.39 $X2=0 $Y2=0
cc_442 N_Y_c_630_n N_VGND_c_807_n 0.0114512f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_443 N_Y_c_667_n N_VGND_c_807_n 0.0141302f $X=3.62 $Y=0.39 $X2=0 $Y2=0
cc_444 N_Y_c_631_n N_VGND_c_807_n 0.00972452f $X=4.345 $Y=0.815 $X2=0 $Y2=0
cc_445 N_Y_c_674_n N_VGND_c_807_n 0.0143352f $X=4.56 $Y=0.39 $X2=0 $Y2=0
cc_446 N_Y_c_632_n N_VGND_c_807_n 0.0094839f $X=5.285 $Y=0.815 $X2=0 $Y2=0
cc_447 N_Y_c_677_n N_VGND_c_807_n 0.0141302f $X=5.5 $Y=0.39 $X2=0 $Y2=0
cc_448 N_Y_c_633_n N_VGND_c_807_n 0.00972452f $X=6.225 $Y=0.815 $X2=0 $Y2=0
cc_449 N_Y_c_703_n N_VGND_c_807_n 0.0143352f $X=6.44 $Y=0.39 $X2=0 $Y2=0
cc_450 N_Y_c_634_n N_VGND_c_807_n 0.0127505f $X=6.905 $Y=0.815 $X2=0 $Y2=0
cc_451 N_Y_c_628_n N_VGND_c_810_n 0.00198695f $X=1.945 $Y=0.815 $X2=0 $Y2=0
cc_452 N_Y_c_658_n N_VGND_c_810_n 0.0231806f $X=2.16 $Y=0.39 $X2=0 $Y2=0
cc_453 N_Y_c_630_n N_VGND_c_810_n 0.00254521f $X=3.405 $Y=0.815 $X2=0 $Y2=0
cc_454 N_Y_c_630_n N_VGND_c_811_n 0.0528344f $X=3.405 $Y=0.815 $X2=0 $Y2=0
