* File: sky130_fd_sc_hdll__or3_1.pex.spice
* Created: Wed Sep  2 08:48:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3_1%C 1 3 6 8 13
r28 13 14 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.505 $Y=1.202
+ $X2=0.53 $Y2=1.202
r29 11 13 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=0.255 $Y=1.202
+ $X2=0.505 $Y2=1.202
r30 8 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r31 4 14 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.53 $Y=0.995
+ $X2=0.53 $Y2=1.202
r32 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.53 $Y=0.995 $X2=0.53
+ $Y2=0.475
r33 1 13 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.202
r34 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.505 $Y=1.41
+ $X2=0.505 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%B 1 2 3 4 6 9 10 11 12 17 22
c42 3 0 1.60095e-19 $X=0.925 $Y=1.41
c43 2 0 8.49032e-20 $X=0.925 $Y=1.31
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.99
+ $Y=2.28 $X2=0.99 $Y2=2.28
r45 12 17 10.1336 $w=2.88e-07 $l=2.55e-07 $layer=LI1_cond $X=0.735 $Y=2.27
+ $X2=0.99 $Y2=2.27
r46 12 22 1.98697 $w=2.88e-07 $l=5e-08 $layer=LI1_cond $X=0.735 $Y=2.27
+ $X2=0.685 $Y2=2.27
r47 11 22 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.225 $Y=2.27
+ $X2=0.685 $Y2=2.27
r48 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.95 $Y=0.475 $X2=0.95
+ $Y2=0.76
r49 4 16 47.4873 $w=2.92e-07 $l=2.7559e-07 $layer=POLY_cond $X=0.925 $Y=2.035
+ $X2=0.99 $Y2=2.28
r50 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.925 $Y=2.035
+ $X2=0.925 $Y2=1.695
r51 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.925 $Y=1.41
+ $X2=0.925 $Y2=1.695
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.925 $Y=1.31 $X2=0.925
+ $Y2=1.41
r53 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.925 $Y=0.86 $X2=0.925
+ $Y2=0.76
r54 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=0.925 $Y=0.86 $X2=0.925
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%A 1 3 6 8 9 10 16 17 23
c50 17 0 1.85985e-19 $X=0.725 $Y=1.325
r51 21 23 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=0.845 $Y=1.16
+ $X2=1.145 $Y2=1.16
r52 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.405
+ $Y=1.16 $X2=1.405 $Y2=1.16
r53 10 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.245 $Y=1.16
+ $X2=1.405 $Y2=1.16
r54 10 23 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.245 $Y=1.16
+ $X2=1.145 $Y2=1.16
r55 9 17 9.84378 $w=2.38e-07 $l=2.05e-07 $layer=LI1_cond $X=0.725 $Y=1.53
+ $X2=0.725 $Y2=1.325
r56 8 17 4.07572 $w=2.4e-07 $l=1.65e-07 $layer=LI1_cond $X=0.725 $Y=1.16
+ $X2=0.725 $Y2=1.325
r57 8 21 2.96416 $w=3.3e-07 $l=1.2e-07 $layer=LI1_cond $X=0.725 $Y=1.16
+ $X2=0.845 $Y2=1.16
r58 4 15 39.1718 $w=2.59e-07 $l=1.93959e-07 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.407 $Y2=1.16
r59 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.475
r60 1 15 51.0578 $w=2.59e-07 $l=2.68328e-07 $layer=POLY_cond $X=1.445 $Y=1.41
+ $X2=1.407 $Y2=1.16
r61 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.445 $Y=1.41
+ $X2=1.445 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%A_29_53# 1 2 3 10 12 13 15 18 20 21 22 26 28
+ 30 35 38 42 43
c91 35 0 1.12758e-19 $X=1.89 $Y=1.16
r92 43 45 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.29 $Y=1.58
+ $X2=1.29 $Y2=1.87
r93 38 40 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=0.267 $Y=1.685
+ $X2=0.267 $Y2=1.87
r94 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.89
+ $Y=1.16 $X2=1.89 $Y2=1.16
r95 33 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.89 $Y=1.495
+ $X2=1.89 $Y2=1.16
r96 32 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.89 $Y=0.825
+ $X2=1.89 $Y2=1.16
r97 31 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.375 $Y=1.58
+ $X2=1.29 $Y2=1.58
r98 30 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.805 $Y=1.58
+ $X2=1.89 $Y2=1.495
r99 30 31 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=1.805 $Y=1.58
+ $X2=1.375 $Y2=1.58
r100 29 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.295 $Y=0.74
+ $X2=1.21 $Y2=0.74
r101 28 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.805 $Y=0.74
+ $X2=1.89 $Y2=0.825
r102 28 29 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=1.805 $Y=0.74
+ $X2=1.295 $Y2=0.74
r103 24 42 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.21 $Y=0.655
+ $X2=1.21 $Y2=0.74
r104 24 26 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.21 $Y=0.655
+ $X2=1.21 $Y2=0.47
r105 23 40 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.43 $Y=1.87
+ $X2=0.267 $Y2=1.87
r106 22 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=1.87
+ $X2=1.29 $Y2=1.87
r107 22 23 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.205 $Y=1.87
+ $X2=0.43 $Y2=1.87
r108 20 42 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.125 $Y=0.74
+ $X2=1.21 $Y2=0.74
r109 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.125 $Y=0.74
+ $X2=0.355 $Y2=0.74
r110 16 21 7.17723 $w=1.7e-07 $l=1.65118e-07 $layer=LI1_cond $X=0.227 $Y=0.655
+ $X2=0.355 $Y2=0.74
r111 16 18 8.36086 $w=2.53e-07 $l=1.85e-07 $layer=LI1_cond $X=0.227 $Y=0.655
+ $X2=0.227 $Y2=0.47
r112 13 36 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=2.01 $Y=0.995
+ $X2=1.92 $Y2=1.16
r113 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.01 $Y=0.995
+ $X2=2.01 $Y2=0.56
r114 10 36 47.6478 $w=3.03e-07 $l=2.80624e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=1.92 $Y2=1.16
r115 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.985 $Y=1.41
+ $X2=1.985 $Y2=1.985
r116 3 38 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.685
r117 2 26 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=1.025
+ $Y=0.265 $X2=1.21 $Y2=0.47
r118 1 18 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=0.145
+ $Y=0.265 $X2=0.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%VPWR 1 6 8 10 17 18 21 26
c24 1 0 1.12758e-19 $X=1.535 $Y=1.485
r25 22 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.23 $Y2=2.72
r26 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r27 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r28 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r29 15 21 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=1.735 $Y2=2.72
r30 15 17 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=1.875 $Y=2.72
+ $X2=2.53 $Y2=2.72
r31 12 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r32 10 21 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=1.595 $Y=2.72
+ $X2=1.735 $Y2=2.72
r33 10 12 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=1.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r34 8 26 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r35 4 21 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.735 $Y=2.635
+ $X2=1.735 $Y2=2.72
r36 4 6 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=1.735 $Y=2.635
+ $X2=1.735 $Y2=2
r37 1 6 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=1.535
+ $Y=1.485 $X2=1.745 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%X 1 2 12 14 15 16
r19 14 16 8.9262 $w=2.73e-07 $l=2.13e-07 $layer=LI1_cond $X=2.477 $Y=1.632
+ $X2=2.477 $Y2=1.845
r20 14 15 7.41084 $w=2.73e-07 $l=1.37e-07 $layer=LI1_cond $X=2.477 $Y=1.632
+ $X2=2.477 $Y2=1.495
r21 10 12 3.50744 $w=3.43e-07 $l=1.05e-07 $layer=LI1_cond $X=2.425 $Y=0.587
+ $X2=2.53 $Y2=0.587
r22 7 12 4.88813 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=2.53 $Y=0.76 $X2=2.53
+ $Y2=0.587
r23 7 15 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.53 $Y=0.76
+ $X2=2.53 $Y2=1.495
r24 2 16 300 $w=1.7e-07 $l=5.05569e-07 $layer=licon1_PDIFF $count=2 $X=2.075
+ $Y=1.485 $X2=2.425 $Y2=1.845
r25 1 10 182 $w=1.7e-07 $l=4.96714e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.425 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3_1%VGND 1 2 9 11 13 18 25 26 29 33 41
r43 33 36 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=1.68 $Y=0 $X2=1.68
+ $Y2=0.4
r44 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r45 30 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r46 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r47 26 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r48 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r49 23 33 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.68
+ $Y2=0
r50 23 25 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.53
+ $Y2=0
r51 22 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r52 22 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r53 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r54 19 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=0.715
+ $Y2=0
r55 19 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=0 $X2=1.15
+ $Y2=0
r56 18 33 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.68
+ $Y2=0
r57 18 21 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.15
+ $Y2=0
r58 15 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r59 13 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.715
+ $Y2=0
r60 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=0 $X2=0.23
+ $Y2=0
r61 11 41 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r62 7 29 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0
r63 7 9 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.715 $Y=0.085
+ $X2=0.715 $Y2=0.4
r64 2 36 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.545
+ $Y=0.265 $X2=1.73 $Y2=0.4
r65 1 9 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=0.605
+ $Y=0.265 $X2=0.74 $Y2=0.4
.ends

