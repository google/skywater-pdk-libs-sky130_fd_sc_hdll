* File: sky130_fd_sc_hdll__o21ai_4.pxi.spice
* Created: Thu Aug 27 19:19:27 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21AI_4%A1 N_A1_c_82_n N_A1_M1003_g N_A1_c_73_n
+ N_A1_M1002_g N_A1_c_83_n N_A1_M1021_g N_A1_c_74_n N_A1_M1007_g N_A1_c_84_n
+ N_A1_M1022_g N_A1_c_75_n N_A1_M1013_g N_A1_c_76_n N_A1_M1023_g N_A1_c_77_n
+ N_A1_M1016_g N_A1_c_92_p N_A1_c_78_n A1 N_A1_c_79_n N_A1_c_80_n A1 N_A1_c_81_n
+ PM_SKY130_FD_SC_HDLL__O21AI_4%A1
x_PM_SKY130_FD_SC_HDLL__O21AI_4%A2 N_A2_c_179_n N_A2_M1001_g N_A2_c_185_n
+ N_A2_M1000_g N_A2_c_180_n N_A2_M1008_g N_A2_c_186_n N_A2_M1004_g N_A2_c_181_n
+ N_A2_M1010_g N_A2_c_187_n N_A2_M1009_g N_A2_c_188_n N_A2_M1015_g N_A2_c_182_n
+ N_A2_M1012_g A2 N_A2_c_183_n N_A2_c_184_n A2 N_A2_X26_noxref_CONDUCTOR
+ PM_SKY130_FD_SC_HDLL__O21AI_4%A2
x_PM_SKY130_FD_SC_HDLL__O21AI_4%B1 N_B1_c_250_n N_B1_M1011_g N_B1_c_256_n
+ N_B1_M1005_g N_B1_c_251_n N_B1_M1017_g N_B1_c_257_n N_B1_M1006_g N_B1_c_252_n
+ N_B1_M1019_g N_B1_c_258_n N_B1_M1014_g N_B1_c_259_n N_B1_M1018_g N_B1_c_253_n
+ N_B1_M1020_g B1 N_B1_c_254_n N_B1_c_255_n B1 PM_SKY130_FD_SC_HDLL__O21AI_4%B1
x_PM_SKY130_FD_SC_HDLL__O21AI_4%VPWR N_VPWR_M1003_d N_VPWR_M1021_d
+ N_VPWR_M1023_d N_VPWR_M1006_d N_VPWR_M1018_d N_VPWR_c_322_n N_VPWR_c_323_n
+ N_VPWR_c_324_n N_VPWR_c_325_n N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_328_n
+ N_VPWR_c_329_n N_VPWR_c_330_n VPWR N_VPWR_c_331_n N_VPWR_c_332_n
+ N_VPWR_c_333_n N_VPWR_c_321_n PM_SKY130_FD_SC_HDLL__O21AI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O21AI_4%A_123_297# N_A_123_297#_M1003_s
+ N_A_123_297#_M1022_s N_A_123_297#_M1004_d N_A_123_297#_M1015_d
+ N_A_123_297#_c_435_n N_A_123_297#_c_418_n N_A_123_297#_c_423_n
+ N_A_123_297#_c_442_n N_A_123_297#_c_425_n
+ PM_SKY130_FD_SC_HDLL__O21AI_4%A_123_297#
x_PM_SKY130_FD_SC_HDLL__O21AI_4%Y N_Y_M1011_d N_Y_M1019_d N_Y_M1000_s
+ N_Y_M1009_s N_Y_M1005_s N_Y_M1014_s N_Y_c_459_n N_Y_c_462_n N_Y_c_503_n
+ N_Y_c_453_n N_Y_c_454_n N_Y_c_512_n N_Y_c_455_n Y N_Y_c_451_n Y
+ PM_SKY130_FD_SC_HDLL__O21AI_4%Y
x_PM_SKY130_FD_SC_HDLL__O21AI_4%A_32_47# N_A_32_47#_M1002_d N_A_32_47#_M1007_d
+ N_A_32_47#_M1001_d N_A_32_47#_M1010_d N_A_32_47#_M1016_d N_A_32_47#_M1017_s
+ N_A_32_47#_M1020_s N_A_32_47#_c_532_n N_A_32_47#_c_569_p N_A_32_47#_c_533_n
+ PM_SKY130_FD_SC_HDLL__O21AI_4%A_32_47#
x_PM_SKY130_FD_SC_HDLL__O21AI_4%VGND N_VGND_M1002_s N_VGND_M1013_s
+ N_VGND_M1008_s N_VGND_M1012_s N_VGND_c_585_n N_VGND_c_586_n VGND
+ N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n
+ N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n
+ PM_SKY130_FD_SC_HDLL__O21AI_4%VGND
cc_1 VNB N_A1_c_73_n 0.0220741f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=0.995
cc_2 VNB N_A1_c_74_n 0.0171564f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=0.995
cc_3 VNB N_A1_c_75_n 0.0163972f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=0.995
cc_4 VNB N_A1_c_76_n 0.0290087f $X=-0.19 $Y=-0.24 $X2=3.885 $Y2=1.41
cc_5 VNB N_A1_c_77_n 0.0172982f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=0.995
cc_6 VNB N_A1_c_78_n 0.00149876f $X=-0.19 $Y=-0.24 $X2=3.88 $Y2=1.16
cc_7 VNB N_A1_c_79_n 0.0117702f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_8 VNB N_A1_c_80_n 0.0792986f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_9 VNB N_A1_c_81_n 0.0029719f $X=-0.19 $Y=-0.24 $X2=1.625 $Y2=1.35
cc_10 VNB N_A2_c_179_n 0.0166765f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.41
cc_11 VNB N_A2_c_180_n 0.0169529f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.41
cc_12 VNB N_A2_c_181_n 0.0173895f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.41
cc_13 VNB N_A2_c_182_n 0.0175233f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=0.995
cc_14 VNB N_A2_c_183_n 0.0026767f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.202
cc_15 VNB N_A2_c_184_n 0.0754023f $X=-0.19 $Y=-0.24 $X2=1.03 $Y2=1.202
cc_16 VNB N_B1_c_250_n 0.0168426f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.41
cc_17 VNB N_B1_c_251_n 0.0170785f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.41
cc_18 VNB N_B1_c_252_n 0.0175833f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.41
cc_19 VNB N_B1_c_253_n 0.0209514f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=0.995
cc_20 VNB N_B1_c_254_n 0.00172607f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.202
cc_21 VNB N_B1_c_255_n 0.0782566f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_22 VNB N_VPWR_c_321_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_Y_c_451_n 0.0114202f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.35
cc_24 VNB Y 0.0208787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_32_47#_c_532_n 0.00946883f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=0.995
cc_26 VNB N_A_32_47#_c_533_n 0.00812227f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_27 VNB N_VGND_c_585_n 0.01367f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.41
cc_28 VNB N_VGND_c_586_n 0.01367f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.985
cc_29 VNB N_VGND_c_587_n 0.0166329f $X=-0.19 $Y=-0.24 $X2=3.885 $Y2=1.41
cc_30 VNB N_VGND_c_588_n 0.0147227f $X=-0.19 $Y=-0.24 $X2=3.95 $Y2=0.56
cc_31 VNB N_VGND_c_589_n 0.0630452f $X=-0.19 $Y=-0.24 $X2=1.165 $Y2=1.445
cc_32 VNB N_VGND_c_590_n 0.317563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_591_n 0.00800334f $X=-0.19 $Y=-0.24 $X2=0.63 $Y2=1.16
cc_34 VNB N_VGND_c_592_n 0.00538475f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_35 VNB N_VGND_c_593_n 0.00538475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_594_n 0.00857211f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_A1_c_82_n 0.0211426f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.41
cc_38 VPB N_A1_c_83_n 0.0153391f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.41
cc_39 VPB N_A1_c_84_n 0.0156704f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.41
cc_40 VPB N_A1_c_76_n 0.0281301f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=1.41
cc_41 VPB N_A1_c_78_n 0.00155178f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.16
cc_42 VPB N_A1_c_79_n 5.70185e-19 $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_43 VPB N_A1_c_80_n 0.0482645f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.202
cc_44 VPB N_A1_c_81_n 0.00286257f $X=-0.19 $Y=1.305 $X2=1.625 $Y2=1.35
cc_45 VPB N_A2_c_185_n 0.0165893f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_46 VPB N_A2_c_186_n 0.0164285f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.995
cc_47 VPB N_A2_c_187_n 0.0164285f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=0.995
cc_48 VPB N_A2_c_188_n 0.016593f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=1.41
cc_49 VPB N_A2_c_183_n 0.00819347f $X=-0.19 $Y=1.305 $X2=1.005 $Y2=1.202
cc_50 VPB N_A2_c_184_n 0.04853f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=1.202
cc_51 VPB N_B1_c_256_n 0.0166831f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=0.995
cc_52 VPB N_B1_c_257_n 0.0156318f $X=-0.19 $Y=1.305 $X2=1.03 $Y2=0.995
cc_53 VPB N_B1_c_258_n 0.0158908f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=0.995
cc_54 VPB N_B1_c_259_n 0.0183865f $X=-0.19 $Y=1.305 $X2=3.885 $Y2=1.41
cc_55 VPB N_B1_c_255_n 0.047238f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_56 VPB N_VPWR_c_322_n 0.0114848f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=0.995
cc_57 VPB N_VPWR_c_323_n 0.0303676f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=0.56
cc_58 VPB N_VPWR_c_324_n 0.0047285f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=0.995
cc_59 VPB N_VPWR_c_325_n 0.0140951f $X=-0.19 $Y=1.305 $X2=3.95 $Y2=0.56
cc_60 VPB N_VPWR_c_326_n 0.0268823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_VPWR_c_327_n 0.0592973f $X=-0.19 $Y=1.305 $X2=3.945 $Y2=1.515
cc_62 VPB N_VPWR_c_328_n 0.00535674f $X=-0.19 $Y=1.305 $X2=3.945 $Y2=1.16
cc_63 VPB N_VPWR_c_329_n 0.00537239f $X=-0.19 $Y=1.305 $X2=3.88 $Y2=1.16
cc_64 VPB N_VPWR_c_330_n 0.0143706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_331_n 0.0158442f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.16
cc_66 VPB N_VPWR_c_332_n 0.0135666f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.35
cc_67 VPB N_VPWR_c_333_n 0.00547531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_321_n 0.0484392f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_Y_c_453_n 0.00245326f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_454_n 0.00147279f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.202
cc_71 VPB N_Y_c_455_n 0.0170968f $X=-0.19 $Y=1.305 $X2=1.41 $Y2=1.16
cc_72 VPB Y 0.0063686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 N_A1_c_75_n N_A2_c_179_n 0.0269803f $X=1.51 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_74 N_A1_c_84_n N_A2_c_185_n 0.0349809f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A1_c_92_p N_A2_c_185_n 0.0190179f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_76 N_A1_c_81_n N_A2_c_185_n 0.00197401f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_77 N_A1_c_92_p N_A2_c_186_n 0.0120284f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_78 N_A1_c_92_p N_A2_c_187_n 0.0120284f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_79 N_A1_c_76_n N_A2_c_188_n 0.0397877f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A1_c_92_p N_A2_c_188_n 0.0119833f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_81 N_A1_c_78_n N_A2_c_188_n 6.5152e-19 $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_82 N_A1_c_77_n N_A2_c_182_n 0.0243143f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A1_c_76_n N_A2_c_183_n 0.0019906f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A1_c_92_p N_A2_c_183_n 0.0944795f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_85 N_A1_c_78_n N_A2_c_183_n 0.0228714f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A1_c_80_n N_A2_c_183_n 2.05897e-19 $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_87 N_A1_c_81_n N_A2_c_183_n 0.0087761f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_88 N_A1_c_76_n N_A2_c_184_n 0.0253694f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A1_c_92_p N_A2_c_184_n 0.00804597f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_90 N_A1_c_78_n N_A2_c_184_n 0.00114258f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A1_c_80_n N_A2_c_184_n 0.0226904f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_92 N_A1_c_81_n N_A2_c_184_n 0.00356041f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_93 N_A1_c_77_n N_B1_c_250_n 0.0231497f $X=3.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_94 N_A1_c_76_n N_B1_c_256_n 0.031848f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A1_c_92_p N_B1_c_256_n 0.00128222f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_96 N_A1_c_78_n N_B1_c_256_n 0.00125971f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A1_c_76_n N_B1_c_254_n 9.20805e-19 $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A1_c_78_n N_B1_c_254_n 0.0172567f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A1_c_76_n N_B1_c_255_n 0.0246319f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A1_c_78_n N_B1_c_255_n 0.00280245f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_81_n N_VPWR_M1021_d 0.00236298f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_102 N_A1_c_92_p N_VPWR_M1023_d 0.00241701f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_103 N_A1_c_78_n N_VPWR_M1023_d 2.88022e-19 $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_104 N_A1_c_82_n N_VPWR_c_323_n 0.0033589f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A1_c_79_n N_VPWR_c_323_n 0.00945755f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A1_c_80_n N_VPWR_c_323_n 0.00514263f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_107 N_A1_c_76_n N_VPWR_c_324_n 0.00291634f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_84_n N_VPWR_c_327_n 0.00467604f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_76_n N_VPWR_c_327_n 0.00512876f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A1_c_82_n N_VPWR_c_331_n 0.00702461f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A1_c_83_n N_VPWR_c_331_n 0.00325906f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A1_c_82_n N_VPWR_c_333_n 5.47792e-19 $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A1_c_83_n N_VPWR_c_333_n 0.00934117f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A1_c_84_n N_VPWR_c_333_n 0.00758326f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A1_c_82_n N_VPWR_c_321_n 0.0133979f $X=0.525 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A1_c_83_n N_VPWR_c_321_n 0.0038791f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A1_c_84_n N_VPWR_c_321_n 0.00532911f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A1_c_76_n N_VPWR_c_321_n 0.006933f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A1_c_81_n N_A_123_297#_M1003_s 0.00293532f $X=1.625 $Y=1.35 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A1_c_92_p N_A_123_297#_M1022_s 0.00935591f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_121 N_A1_c_92_p N_A_123_297#_M1004_d 0.00354953f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_122 N_A1_c_92_p N_A_123_297#_M1015_d 0.00646439f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_123 N_A1_c_83_n N_A_123_297#_c_418_n 0.0131589f $X=1.005 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A1_c_84_n N_A_123_297#_c_418_n 0.0134967f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_92_p N_A_123_297#_c_418_n 0.0118846f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_126 N_A1_c_80_n N_A_123_297#_c_418_n 7.96607e-19 $X=1.485 $Y=1.202 $X2=0
+ $Y2=0
cc_127 N_A1_c_81_n N_A_123_297#_c_418_n 0.0334389f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_128 N_A1_c_80_n N_A_123_297#_c_423_n 7.88489e-19 $X=1.485 $Y=1.202 $X2=0
+ $Y2=0
cc_129 N_A1_c_81_n N_A_123_297#_c_423_n 0.0131161f $X=1.625 $Y=1.35 $X2=0 $Y2=0
cc_130 N_A1_c_76_n N_A_123_297#_c_425_n 0.00251487f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A1_c_92_p N_A_123_297#_c_425_n 0.00280123f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_132 N_A1_c_92_p N_Y_M1000_s 0.00379276f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_133 N_A1_c_92_p N_Y_M1009_s 0.00354953f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_134 N_A1_c_84_n N_Y_c_459_n 3.75967e-19 $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_76_n N_Y_c_459_n 0.0142574f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_92_p N_Y_c_459_n 0.113661f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_137 N_A1_c_77_n N_Y_c_462_n 2.12504e-19 $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A1_c_76_n N_Y_c_454_n 0.00124407f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A1_c_92_p N_Y_c_454_n 0.0113729f $X=3.795 $Y=1.6 $X2=0 $Y2=0
cc_140 N_A1_c_78_n N_Y_c_454_n 0.0044205f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_141 N_A1_c_73_n N_A_32_47#_c_532_n 0.0104839f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_74_n N_A_32_47#_c_532_n 0.0111505f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_75_n N_A_32_47#_c_532_n 0.0100792f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_76_n N_A_32_47#_c_532_n 0.00386458f $X=3.885 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A1_c_77_n N_A_32_47#_c_532_n 0.011962f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A1_c_78_n N_A_32_47#_c_532_n 0.019888f $X=3.88 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A1_c_79_n N_A_32_47#_c_532_n 0.0925128f $X=0.63 $Y=1.16 $X2=0 $Y2=0
cc_148 N_A1_c_80_n N_A_32_47#_c_532_n 0.0147698f $X=1.485 $Y=1.202 $X2=0 $Y2=0
cc_149 N_A1_c_73_n N_VGND_c_587_n 0.00211056f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A1_c_74_n N_VGND_c_588_n 0.00422112f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_75_n N_VGND_c_588_n 0.00211056f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_77_n N_VGND_c_589_n 0.00422112f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_73_n N_VGND_c_590_n 0.00380107f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_74_n N_VGND_c_590_n 0.00590855f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A1_c_75_n N_VGND_c_590_n 0.00289589f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_156 N_A1_c_77_n N_VGND_c_590_n 0.00606048f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A1_c_73_n N_VGND_c_591_n 0.0171546f $X=0.55 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A1_c_74_n N_VGND_c_591_n 0.00165122f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A1_c_74_n N_VGND_c_592_n 0.00118069f $X=1.03 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A1_c_75_n N_VGND_c_592_n 0.0107231f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A1_c_77_n N_VGND_c_594_n 0.0052631f $X=3.95 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A2_c_185_n N_VPWR_c_327_n 0.00429453f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A2_c_186_n N_VPWR_c_327_n 0.00429453f $X=2.445 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A2_c_187_n N_VPWR_c_327_n 0.00429453f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A2_c_188_n N_VPWR_c_327_n 0.00429453f $X=3.405 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A2_c_185_n N_VPWR_c_333_n 9.82843e-19 $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A2_c_185_n N_VPWR_c_321_n 0.00614026f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A2_c_186_n N_VPWR_c_321_n 0.00611674f $X=2.445 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A2_c_187_n N_VPWR_c_321_n 0.00611674f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A2_c_188_n N_VPWR_c_321_n 0.00614026f $X=3.405 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A2_c_185_n N_A_123_297#_c_425_n 0.0112889f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A2_c_186_n N_A_123_297#_c_425_n 0.0101154f $X=2.445 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A2_c_187_n N_A_123_297#_c_425_n 0.0101154f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A2_c_188_n N_A_123_297#_c_425_n 0.0101154f $X=3.405 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A2_c_185_n N_Y_c_459_n 0.00481708f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A2_c_186_n N_Y_c_459_n 0.0103844f $X=2.445 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A2_c_187_n N_Y_c_459_n 0.0103844f $X=2.925 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A2_c_188_n N_Y_c_459_n 0.0103393f $X=3.405 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A2_c_179_n N_A_32_47#_c_532_n 0.0150217f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A2_c_180_n N_A_32_47#_c_532_n 0.0112375f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A2_c_181_n N_A_32_47#_c_532_n 0.0112375f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A2_c_182_n N_A_32_47#_c_532_n 0.0109718f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_183 N_A2_c_183_n N_A_32_47#_c_532_n 0.0687783f $X=3.29 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A2_c_184_n N_A_32_47#_c_532_n 0.0128532f $X=3.405 $Y=1.202 $X2=0 $Y2=0
cc_185 N_A2_c_179_n N_VGND_c_585_n 0.0035176f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A2_c_180_n N_VGND_c_585_n 0.0035176f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A2_c_181_n N_VGND_c_586_n 0.0035176f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A2_c_182_n N_VGND_c_586_n 0.00211056f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A2_c_179_n N_VGND_c_590_n 0.00424616f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A2_c_180_n N_VGND_c_590_n 0.00424616f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A2_c_181_n N_VGND_c_590_n 0.00436366f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A2_c_182_n N_VGND_c_590_n 0.00301339f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A2_c_179_n N_VGND_c_592_n 0.00793528f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A2_c_180_n N_VGND_c_592_n 0.00106058f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A2_c_179_n N_VGND_c_593_n 0.00106058f $X=1.94 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A2_c_180_n N_VGND_c_593_n 0.00819243f $X=2.42 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A2_c_181_n N_VGND_c_593_n 0.00824353f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A2_c_182_n N_VGND_c_593_n 0.00103795f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A2_c_181_n N_VGND_c_594_n 0.0011512f $X=2.9 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A2_c_182_n N_VGND_c_594_n 0.0108692f $X=3.43 $Y=0.995 $X2=0 $Y2=0
cc_201 N_B1_c_256_n N_VPWR_c_324_n 0.00175847f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B1_c_258_n N_VPWR_c_326_n 6.65625e-19 $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B1_c_259_n N_VPWR_c_326_n 0.0153706f $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B1_c_256_n N_VPWR_c_329_n 5.38342e-19 $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B1_c_257_n N_VPWR_c_329_n 0.00928655f $X=4.885 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B1_c_258_n N_VPWR_c_329_n 0.0065955f $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B1_c_259_n N_VPWR_c_329_n 4.82946e-19 $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B1_c_256_n N_VPWR_c_330_n 0.00520311f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B1_c_257_n N_VPWR_c_330_n 0.00325906f $X=4.885 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B1_c_258_n N_VPWR_c_332_n 0.00467604f $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B1_c_259_n N_VPWR_c_332_n 0.00447018f $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B1_c_256_n N_VPWR_c_321_n 0.00685232f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B1_c_257_n N_VPWR_c_321_n 0.0038791f $X=4.885 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B1_c_258_n N_VPWR_c_321_n 0.00530559f $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B1_c_259_n N_VPWR_c_321_n 0.00766229f $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B1_c_256_n N_Y_c_459_n 0.00357251f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B1_c_254_n N_Y_c_459_n 6.28566e-19 $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_218 N_B1_c_250_n N_Y_c_462_n 0.00319406f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B1_c_251_n N_Y_c_462_n 0.0104198f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B1_c_252_n N_Y_c_462_n 0.0104198f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_221 N_B1_c_253_n N_Y_c_462_n 0.00760615f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_222 N_B1_c_254_n N_Y_c_462_n 0.075037f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_223 N_B1_c_255_n N_Y_c_462_n 0.0120647f $X=5.845 $Y=1.202 $X2=0 $Y2=0
cc_224 N_B1_c_257_n N_Y_c_453_n 0.0280082f $X=4.885 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B1_c_258_n N_Y_c_453_n 0.0284027f $X=5.365 $Y=1.41 $X2=0 $Y2=0
cc_226 N_B1_c_254_n N_Y_c_453_n 0.0615666f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B1_c_255_n N_Y_c_453_n 0.0112838f $X=5.845 $Y=1.202 $X2=0 $Y2=0
cc_228 N_B1_c_256_n N_Y_c_454_n 0.0216762f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B1_c_254_n N_Y_c_454_n 0.0326846f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_230 N_B1_c_255_n N_Y_c_454_n 0.00648452f $X=5.845 $Y=1.202 $X2=0 $Y2=0
cc_231 N_B1_c_259_n N_Y_c_455_n 0.0227679f $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B1_c_254_n N_Y_c_455_n 0.00746774f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_233 N_B1_c_255_n N_Y_c_455_n 0.00722359f $X=5.845 $Y=1.202 $X2=0 $Y2=0
cc_234 N_B1_c_253_n N_Y_c_451_n 0.00580029f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B1_c_252_n Y 5.93951e-19 $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B1_c_259_n Y 0.00133231f $X=5.845 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B1_c_253_n Y 0.00615611f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B1_c_254_n Y 0.0125829f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_239 N_B1_c_255_n Y 0.0205506f $X=5.845 $Y=1.202 $X2=0 $Y2=0
cc_240 N_B1_c_250_n N_A_32_47#_c_533_n 0.0110504f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_241 N_B1_c_251_n N_A_32_47#_c_533_n 0.00853857f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_242 N_B1_c_252_n N_A_32_47#_c_533_n 0.00882069f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_243 N_B1_c_253_n N_A_32_47#_c_533_n 0.00881969f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B1_c_254_n N_A_32_47#_c_533_n 0.00324863f $X=5.25 $Y=1.16 $X2=0 $Y2=0
cc_245 N_B1_c_250_n N_VGND_c_589_n 0.00357877f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_246 N_B1_c_251_n N_VGND_c_589_n 0.00357877f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_247 N_B1_c_252_n N_VGND_c_589_n 0.00357877f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_248 N_B1_c_253_n N_VGND_c_589_n 0.00357877f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_249 N_B1_c_250_n N_VGND_c_590_n 0.00547449f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_250 N_B1_c_251_n N_VGND_c_590_n 0.00553284f $X=4.86 $Y=0.995 $X2=0 $Y2=0
cc_251 N_B1_c_252_n N_VGND_c_590_n 0.00565034f $X=5.34 $Y=0.995 $X2=0 $Y2=0
cc_252 N_B1_c_253_n N_VGND_c_590_n 0.00653665f $X=5.87 $Y=0.995 $X2=0 $Y2=0
cc_253 N_VPWR_c_321_n N_A_123_297#_M1003_s 0.00292904f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_254 N_VPWR_c_321_n N_A_123_297#_M1022_s 0.00258996f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_321_n N_A_123_297#_M1004_d 0.00239319f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_321_n N_A_123_297#_M1015_d 0.00239319f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_331_n N_A_123_297#_c_435_n 0.0145465f $X=1.03 $Y=2.72 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_321_n N_A_123_297#_c_435_n 0.008919f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_259 N_VPWR_M1021_d N_A_123_297#_c_418_n 0.00395034f $X=1.095 $Y=1.485 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_327_n N_A_123_297#_c_418_n 0.00323816f $X=4.03 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_331_n N_A_123_297#_c_418_n 0.00241998f $X=1.03 $Y=2.72 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_333_n N_A_123_297#_c_418_n 0.0196796f $X=1.245 $Y=2.34 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_321_n N_A_123_297#_c_418_n 0.011274f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_264 N_VPWR_c_327_n N_A_123_297#_c_442_n 0.0130208f $X=4.03 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_321_n N_A_123_297#_c_442_n 0.00725703f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_327_n N_A_123_297#_c_425_n 0.110952f $X=4.03 $Y=2.72 $X2=0 $Y2=0
cc_267 N_VPWR_c_321_n N_A_123_297#_c_425_n 0.0705948f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_321_n N_Y_M1000_s 0.00240926f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_321_n N_Y_M1009_s 0.00240926f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_270 N_VPWR_c_321_n N_Y_M1005_s 0.00272723f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_271 N_VPWR_c_321_n N_Y_M1014_s 0.00449124f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_272 N_VPWR_M1023_d N_Y_c_459_n 0.00914506f $X=3.975 $Y=1.485 $X2=0 $Y2=0
cc_273 N_VPWR_c_324_n N_Y_c_459_n 0.0175498f $X=4.145 $Y=2.36 $X2=0 $Y2=0
cc_274 N_VPWR_c_327_n N_Y_c_459_n 0.00280993f $X=4.03 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_330_n N_Y_c_459_n 3.13368e-19 $X=4.91 $Y=2.72 $X2=0 $Y2=0
cc_276 N_VPWR_c_321_n N_Y_c_459_n 0.0109801f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_330_n N_Y_c_503_n 0.0138602f $X=4.91 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_321_n N_Y_c_503_n 0.00800522f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_M1006_d N_Y_c_453_n 0.00198123f $X=4.975 $Y=1.485 $X2=0 $Y2=0
cc_280 N_VPWR_c_329_n N_Y_c_453_n 0.0215528f $X=5.125 $Y=2.34 $X2=0 $Y2=0
cc_281 N_VPWR_c_330_n N_Y_c_453_n 0.00259031f $X=4.91 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_332_n N_Y_c_453_n 0.00348255f $X=5.87 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_321_n N_Y_c_453_n 0.0120988f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_284 N_VPWR_c_330_n N_Y_c_454_n 0.00278193f $X=4.91 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_321_n N_Y_c_454_n 0.00471124f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_332_n N_Y_c_512_n 0.0131506f $X=5.87 $Y=2.72 $X2=0 $Y2=0
cc_287 N_VPWR_c_321_n N_Y_c_512_n 0.00722976f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_288 N_VPWR_M1018_d N_Y_c_455_n 0.00354399f $X=5.935 $Y=1.485 $X2=0 $Y2=0
cc_289 N_VPWR_c_326_n N_Y_c_455_n 0.027193f $X=6.085 $Y=1.965 $X2=0 $Y2=0
cc_290 N_A_123_297#_c_425_n N_Y_M1000_s 0.00411534f $X=3.645 $Y=2.36 $X2=0.525
+ $Y2=1.985
cc_291 N_A_123_297#_c_425_n N_Y_M1009_s 0.00411534f $X=3.645 $Y=2.36 $X2=0.55
+ $Y2=0.995
cc_292 N_A_123_297#_M1004_d N_Y_c_459_n 0.00404884f $X=2.535 $Y=1.485 $X2=3.885
+ $Y2=1.41
cc_293 N_A_123_297#_M1015_d N_Y_c_459_n 0.00422785f $X=3.495 $Y=1.485 $X2=3.885
+ $Y2=1.41
cc_294 N_A_123_297#_c_425_n N_Y_c_459_n 0.0654066f $X=3.645 $Y=2.36 $X2=3.885
+ $Y2=1.41
cc_295 N_Y_c_462_n N_A_32_47#_M1017_s 0.00419502f $X=5.92 $Y=0.73 $X2=0 $Y2=0
cc_296 N_Y_c_451_n N_A_32_47#_M1020_s 0.00376009f $X=6.125 $Y=0.845 $X2=0 $Y2=0
cc_297 Y N_A_32_47#_M1020_s 2.26659e-19 $X=6.25 $Y=0.85 $X2=0 $Y2=0
cc_298 N_Y_M1011_d N_A_32_47#_c_533_n 0.0041884f $X=4.455 $Y=0.235 $X2=0 $Y2=0
cc_299 N_Y_M1019_d N_A_32_47#_c_533_n 0.00535007f $X=5.415 $Y=0.235 $X2=0 $Y2=0
cc_300 N_Y_c_462_n N_A_32_47#_c_533_n 0.0789328f $X=5.92 $Y=0.73 $X2=0 $Y2=0
cc_301 N_Y_c_451_n N_A_32_47#_c_533_n 0.0209582f $X=6.125 $Y=0.845 $X2=0 $Y2=0
cc_302 N_Y_c_451_n N_VGND_c_589_n 0.00169401f $X=6.125 $Y=0.845 $X2=0 $Y2=0
cc_303 N_Y_M1011_d N_VGND_c_590_n 0.00265018f $X=4.455 $Y=0.235 $X2=0 $Y2=0
cc_304 N_Y_M1019_d N_VGND_c_590_n 0.00305172f $X=5.415 $Y=0.235 $X2=0 $Y2=0
cc_305 N_Y_c_451_n N_VGND_c_590_n 0.00330181f $X=6.125 $Y=0.845 $X2=0 $Y2=0
cc_306 N_A_32_47#_c_532_n N_VGND_M1002_s 0.00429614f $X=4.03 $Y=0.717 $X2=-0.19
+ $Y2=-0.24
cc_307 N_A_32_47#_c_532_n N_VGND_M1013_s 0.00817986f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_308 N_A_32_47#_c_532_n N_VGND_M1008_s 0.00452812f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_309 N_A_32_47#_c_532_n N_VGND_M1012_s 0.00824222f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_310 N_A_32_47#_c_532_n N_VGND_c_585_n 0.00950223f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_311 N_A_32_47#_c_532_n N_VGND_c_586_n 0.00956125f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_312 N_A_32_47#_c_532_n N_VGND_c_587_n 0.00743655f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_313 N_A_32_47#_c_532_n N_VGND_c_588_n 0.00932634f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_314 N_A_32_47#_c_532_n N_VGND_c_589_n 0.00338335f $X=4.03 $Y=0.717 $X2=0
+ $Y2=0
cc_315 N_A_32_47#_c_569_p N_VGND_c_589_n 0.0137873f $X=4.26 $Y=0.35 $X2=0 $Y2=0
cc_316 N_A_32_47#_c_533_n N_VGND_c_589_n 0.113199f $X=6.085 $Y=0.36 $X2=0 $Y2=0
cc_317 N_A_32_47#_M1002_d N_VGND_c_590_n 0.00363732f $X=0.16 $Y=0.235 $X2=0
+ $Y2=0
cc_318 N_A_32_47#_M1007_d N_VGND_c_590_n 0.00378046f $X=1.105 $Y=0.235 $X2=0
+ $Y2=0
cc_319 N_A_32_47#_M1001_d N_VGND_c_590_n 0.00375928f $X=2.015 $Y=0.235 $X2=0
+ $Y2=0
cc_320 N_A_32_47#_M1010_d N_VGND_c_590_n 0.00435845f $X=2.975 $Y=0.235 $X2=0
+ $Y2=0
cc_321 N_A_32_47#_M1016_d N_VGND_c_590_n 0.00226522f $X=4.025 $Y=0.235 $X2=0
+ $Y2=0
cc_322 N_A_32_47#_M1017_s N_VGND_c_590_n 0.00263412f $X=4.935 $Y=0.235 $X2=0
+ $Y2=0
cc_323 N_A_32_47#_M1020_s N_VGND_c_590_n 0.00229841f $X=5.945 $Y=0.235 $X2=0
+ $Y2=0
cc_324 N_A_32_47#_c_532_n N_VGND_c_590_n 0.0718386f $X=4.03 $Y=0.717 $X2=0 $Y2=0
cc_325 N_A_32_47#_c_569_p N_VGND_c_590_n 0.00881516f $X=4.26 $Y=0.35 $X2=0 $Y2=0
cc_326 N_A_32_47#_c_533_n N_VGND_c_590_n 0.0713494f $X=6.085 $Y=0.36 $X2=0 $Y2=0
cc_327 N_A_32_47#_c_532_n N_VGND_c_591_n 0.0218499f $X=4.03 $Y=0.717 $X2=0 $Y2=0
cc_328 N_A_32_47#_c_532_n N_VGND_c_592_n 0.0196966f $X=4.03 $Y=0.717 $X2=0 $Y2=0
cc_329 N_A_32_47#_c_532_n N_VGND_c_593_n 0.0199417f $X=4.03 $Y=0.717 $X2=0 $Y2=0
cc_330 N_A_32_47#_c_532_n N_VGND_c_594_n 0.0242287f $X=4.03 $Y=0.717 $X2=0 $Y2=0
