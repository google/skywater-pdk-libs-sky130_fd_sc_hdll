* File: sky130_fd_sc_hdll__and2b_2.pxi.spice
* Created: Wed Sep  2 08:21:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND2B_2%A_N N_A_N_c_65_n N_A_N_c_66_n N_A_N_M1001_g
+ N_A_N_M1006_g A_N N_A_N_c_63_n A_N A_N PM_SKY130_FD_SC_HDLL__AND2B_2%A_N
x_PM_SKY130_FD_SC_HDLL__AND2B_2%A_27_413# N_A_27_413#_M1006_d
+ N_A_27_413#_M1001_s N_A_27_413#_c_97_n N_A_27_413#_c_105_n N_A_27_413#_M1008_g
+ N_A_27_413#_M1005_g N_A_27_413#_c_106_n N_A_27_413#_c_107_n
+ N_A_27_413#_c_108_n N_A_27_413#_c_99_n N_A_27_413#_c_100_n N_A_27_413#_c_101_n
+ N_A_27_413#_c_102_n N_A_27_413#_c_103_n
+ PM_SKY130_FD_SC_HDLL__AND2B_2%A_27_413#
x_PM_SKY130_FD_SC_HDLL__AND2B_2%B N_B_c_165_n N_B_M1003_g N_B_M1002_g B
+ PM_SKY130_FD_SC_HDLL__AND2B_2%B
x_PM_SKY130_FD_SC_HDLL__AND2B_2%A_230_413# N_A_230_413#_M1005_s
+ N_A_230_413#_M1008_d N_A_230_413#_c_204_n N_A_230_413#_M1000_g
+ N_A_230_413#_c_196_n N_A_230_413#_M1004_g N_A_230_413#_c_197_n
+ N_A_230_413#_c_198_n N_A_230_413#_c_207_n N_A_230_413#_M1009_g
+ N_A_230_413#_c_199_n N_A_230_413#_M1007_g N_A_230_413#_c_200_n
+ N_A_230_413#_c_209_n N_A_230_413#_c_201_n N_A_230_413#_c_202_n
+ N_A_230_413#_c_203_n N_A_230_413#_c_226_n
+ PM_SKY130_FD_SC_HDLL__AND2B_2%A_230_413#
x_PM_SKY130_FD_SC_HDLL__AND2B_2%VPWR N_VPWR_M1001_d N_VPWR_M1003_d
+ N_VPWR_M1009_d N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n VPWR
+ N_VPWR_c_282_n N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_285_n N_VPWR_c_286_n
+ N_VPWR_c_278_n PM_SKY130_FD_SC_HDLL__AND2B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND2B_2%X N_X_M1004_s N_X_M1000_s N_X_c_325_n X X X
+ N_X_c_322_n PM_SKY130_FD_SC_HDLL__AND2B_2%X
x_PM_SKY130_FD_SC_HDLL__AND2B_2%VGND N_VGND_M1006_s N_VGND_M1002_d
+ N_VGND_M1007_d N_VGND_c_348_n N_VGND_c_349_n N_VGND_c_350_n N_VGND_c_351_n
+ N_VGND_c_352_n N_VGND_c_353_n N_VGND_c_354_n VGND N_VGND_c_355_n
+ N_VGND_c_356_n PM_SKY130_FD_SC_HDLL__AND2B_2%VGND
cc_1 VNB N_A_N_M1006_g 0.0403746f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB N_A_N_c_63_n 0.0357479f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_3 VNB A_N 0.0230148f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0.85
cc_4 VNB N_A_27_413#_c_97_n 0.0112964f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_413#_M1005_g 0.0223654f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_6 VNB N_A_27_413#_c_99_n 0.00425817f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_7 VNB N_A_27_413#_c_100_n 0.00392573f $X=-0.19 $Y=-0.24 $X2=0.297 $Y2=1.53
cc_8 VNB N_A_27_413#_c_101_n 0.00495997f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_413#_c_102_n 0.00816389f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_413#_c_103_n 0.0585635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B_c_165_n 0.0216601f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_12 VNB N_B_M1002_g 0.0396403f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_13 VNB N_A_230_413#_c_196_n 0.0181192f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_14 VNB N_A_230_413#_c_197_n 0.0230077f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_15 VNB N_A_230_413#_c_198_n 0.0195992f $X=-0.19 $Y=-0.24 $X2=0.365 $Y2=1.16
cc_16 VNB N_A_230_413#_c_199_n 0.0227876f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0.85
cc_17 VNB N_A_230_413#_c_200_n 0.0244792f $X=-0.19 $Y=-0.24 $X2=0.297 $Y2=1.16
cc_18 VNB N_A_230_413#_c_201_n 0.00544022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_230_413#_c_202_n 0.0170004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_230_413#_c_203_n 0.00545131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_278_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_X_c_322_n 0.00182827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_348_n 0.0115527f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.445
cc_24 VNB N_VGND_c_349_n 0.0208367f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.16
cc_25 VNB N_VGND_c_350_n 0.00583834f $X=-0.19 $Y=-0.24 $X2=0.397 $Y2=1.325
cc_26 VNB N_VGND_c_351_n 0.0101057f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=0.85
cc_27 VNB N_VGND_c_352_n 0.0256869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_353_n 0.0477866f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_29 VNB N_VGND_c_354_n 0.00709012f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_355_n 0.0232878f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_356_n 0.203283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_N_c_65_n 0.0431934f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_33 VPB N_A_N_c_66_n 0.0267169f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_34 VPB N_A_N_c_63_n 0.00743085f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_35 VPB A_N 0.0149669f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0.85
cc_36 VPB N_A_27_413#_c_97_n 0.0340756f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_37 VPB N_A_27_413#_c_105_n 0.0233346f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_413#_c_106_n 0.00219961f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=0.85
cc_39 VPB N_A_27_413#_c_107_n 0.00909511f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_413#_c_108_n 0.0109634f $X=-0.19 $Y=1.305 $X2=0.297 $Y2=1.16
cc_41 VPB N_A_27_413#_c_100_n 0.00985487f $X=-0.19 $Y=1.305 $X2=0.297 $Y2=1.53
cc_42 VPB N_B_c_165_n 0.101402f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_43 VPB B 0.00752663f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_44 VPB N_A_230_413#_c_204_n 0.0205106f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_45 VPB N_A_230_413#_c_197_n 0.0129686f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_46 VPB N_A_230_413#_c_198_n 0.0117888f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_47 VPB N_A_230_413#_c_207_n 0.0218753f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=0.995
cc_48 VPB N_A_230_413#_c_200_n 0.0098625f $X=-0.19 $Y=1.305 $X2=0.297 $Y2=1.16
cc_49 VPB N_A_230_413#_c_209_n 0.00640752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_230_413#_c_202_n 0.00783822f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_230_413#_c_203_n 0.00249332f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_279_n 0.00287591f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.16
cc_53 VPB N_VPWR_c_280_n 0.0100799f $X=-0.19 $Y=1.305 $X2=0.365 $Y2=1.16
cc_54 VPB N_VPWR_c_281_n 0.0386212f $X=-0.19 $Y=1.305 $X2=0.397 $Y2=1.325
cc_55 VPB N_VPWR_c_282_n 0.015299f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_283_n 0.0255421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_284_n 0.00580026f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_285_n 0.0213675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_VPWR_c_286_n 0.0220531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_278_n 0.044694f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_X_c_322_n 0.00155675f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 N_A_N_c_63_n N_A_27_413#_c_97_n 0.0105067f $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_N_c_65_n N_A_27_413#_c_105_n 0.0105067f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_64 N_A_N_c_66_n N_A_27_413#_c_105_n 0.0119426f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_65 N_A_N_c_66_n N_A_27_413#_c_106_n 0.00550801f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_66 N_A_N_c_65_n N_A_27_413#_c_107_n 0.0125836f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_67 N_A_N_c_66_n N_A_27_413#_c_107_n 0.0100882f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_68 A_N N_A_27_413#_c_107_n 0.00847314f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_69 N_A_N_c_63_n N_A_27_413#_c_108_n 6.06494e-19 $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_70 A_N N_A_27_413#_c_108_n 0.0158932f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_71 N_A_N_M1006_g N_A_27_413#_c_99_n 0.00516557f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_72 A_N N_A_27_413#_c_99_n 0.00250825f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_73 N_A_N_c_63_n N_A_27_413#_c_100_n 0.00893858f $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_74 A_N N_A_27_413#_c_100_n 0.030281f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_75 N_A_N_M1006_g N_A_27_413#_c_102_n 0.00331666f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_76 A_N N_A_27_413#_c_102_n 0.0224269f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_77 N_A_N_M1006_g N_A_27_413#_c_103_n 0.0105067f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_78 A_N N_A_27_413#_c_103_n 3.67811e-19 $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_79 N_A_N_c_65_n N_A_230_413#_c_209_n 2.19769e-19 $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_80 N_A_N_c_66_n N_A_230_413#_c_209_n 5.49995e-19 $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_81 N_A_N_c_66_n N_VPWR_c_279_n 0.0130503f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_82 N_A_N_c_66_n N_VPWR_c_282_n 0.00321743f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_83 N_A_N_c_66_n N_VPWR_c_278_n 0.00482954f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_84 N_A_N_M1006_g N_VGND_c_349_n 0.00511218f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_N_c_63_n N_VGND_c_349_n 9.78244e-19 $X=0.365 $Y=1.16 $X2=0 $Y2=0
cc_86 A_N N_VGND_c_349_n 0.0225521f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_87 N_A_N_M1006_g N_VGND_c_353_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_88 N_A_N_M1006_g N_VGND_c_356_n 0.0128435f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_89 A_N N_VGND_c_356_n 0.00211755f $X=0.23 $Y=0.85 $X2=0 $Y2=0
cc_90 N_A_27_413#_c_97_n N_B_c_165_n 0.02842f $X=1.06 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_91 N_A_27_413#_c_105_n N_B_c_165_n 0.0110119f $X=1.06 $Y=1.99 $X2=-0.19
+ $Y2=-0.24
cc_92 N_A_27_413#_c_103_n N_B_c_165_n 0.00603574f $X=1.14 $Y=0.97 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_27_413#_M1005_g N_B_M1002_g 0.031111f $X=1.56 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_27_413#_c_103_n N_B_M1002_g 0.00233212f $X=1.14 $Y=0.97 $X2=0 $Y2=0
cc_95 N_A_27_413#_c_97_n N_A_230_413#_c_209_n 0.0104126f $X=1.06 $Y=1.89 $X2=0
+ $Y2=0
cc_96 N_A_27_413#_c_105_n N_A_230_413#_c_209_n 0.0114804f $X=1.06 $Y=1.99 $X2=0
+ $Y2=0
cc_97 N_A_27_413#_c_107_n N_A_230_413#_c_209_n 0.0177862f $X=0.67 $Y=1.9 $X2=0
+ $Y2=0
cc_98 N_A_27_413#_c_100_n N_A_230_413#_c_209_n 0.0219212f $X=0.787 $Y=1.785
+ $X2=0 $Y2=0
cc_99 N_A_27_413#_M1005_g N_A_230_413#_c_201_n 0.00605995f $X=1.56 $Y=0.445
+ $X2=0 $Y2=0
cc_100 N_A_27_413#_c_101_n N_A_230_413#_c_201_n 0.00587327f $X=0.73 $Y=0.445
+ $X2=0 $Y2=0
cc_101 N_A_27_413#_c_102_n N_A_230_413#_c_201_n 0.0106411f $X=1.14 $Y=0.97 $X2=0
+ $Y2=0
cc_102 N_A_27_413#_c_103_n N_A_230_413#_c_201_n 0.00587302f $X=1.14 $Y=0.97
+ $X2=0 $Y2=0
cc_103 N_A_27_413#_c_97_n N_A_230_413#_c_202_n 0.00831045f $X=1.06 $Y=1.89 $X2=0
+ $Y2=0
cc_104 N_A_27_413#_c_100_n N_A_230_413#_c_202_n 0.0192972f $X=0.787 $Y=1.785
+ $X2=0 $Y2=0
cc_105 N_A_27_413#_c_102_n N_A_230_413#_c_202_n 0.0315494f $X=1.14 $Y=0.97 $X2=0
+ $Y2=0
cc_106 N_A_27_413#_c_103_n N_A_230_413#_c_202_n 0.0148684f $X=1.14 $Y=0.97 $X2=0
+ $Y2=0
cc_107 N_A_27_413#_M1005_g N_A_230_413#_c_226_n 0.00595503f $X=1.56 $Y=0.445
+ $X2=0 $Y2=0
cc_108 N_A_27_413#_c_101_n N_A_230_413#_c_226_n 0.016358f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_109 N_A_27_413#_c_102_n N_A_230_413#_c_226_n 0.00405807f $X=1.14 $Y=0.97
+ $X2=0 $Y2=0
cc_110 N_A_27_413#_c_103_n N_A_230_413#_c_226_n 0.00734235f $X=1.14 $Y=0.97
+ $X2=0 $Y2=0
cc_111 N_A_27_413#_c_105_n N_VPWR_c_279_n 0.00692624f $X=1.06 $Y=1.99 $X2=0
+ $Y2=0
cc_112 N_A_27_413#_c_106_n N_VPWR_c_279_n 0.0194103f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_113 N_A_27_413#_c_107_n N_VPWR_c_279_n 0.0289845f $X=0.67 $Y=1.9 $X2=0 $Y2=0
cc_114 N_A_27_413#_c_106_n N_VPWR_c_282_n 0.010445f $X=0.26 $Y=2.225 $X2=0 $Y2=0
cc_115 N_A_27_413#_c_107_n N_VPWR_c_282_n 0.00252438f $X=0.67 $Y=1.9 $X2=0 $Y2=0
cc_116 N_A_27_413#_c_105_n N_VPWR_c_285_n 0.00646924f $X=1.06 $Y=1.99 $X2=0
+ $Y2=0
cc_117 N_A_27_413#_M1001_s N_VPWR_c_278_n 0.00388418f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_118 N_A_27_413#_c_105_n N_VPWR_c_278_n 0.0113007f $X=1.06 $Y=1.99 $X2=0 $Y2=0
cc_119 N_A_27_413#_c_106_n N_VPWR_c_278_n 0.00640243f $X=0.26 $Y=2.225 $X2=0
+ $Y2=0
cc_120 N_A_27_413#_c_107_n N_VPWR_c_278_n 0.00600939f $X=0.67 $Y=1.9 $X2=0 $Y2=0
cc_121 N_A_27_413#_M1005_g N_VGND_c_353_n 0.00388886f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_122 N_A_27_413#_c_101_n N_VGND_c_353_n 0.0139933f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_123 N_A_27_413#_M1006_d N_VGND_c_356_n 0.00388065f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_124 N_A_27_413#_M1005_g N_VGND_c_356_n 0.00694043f $X=1.56 $Y=0.445 $X2=0
+ $Y2=0
cc_125 N_A_27_413#_c_101_n N_VGND_c_356_n 0.00898141f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_126 N_A_27_413#_c_102_n N_VGND_c_356_n 0.0116277f $X=1.14 $Y=0.97 $X2=0 $Y2=0
cc_127 N_A_27_413#_c_103_n N_VGND_c_356_n 0.00646506f $X=1.14 $Y=0.97 $X2=0
+ $Y2=0
cc_128 N_B_c_165_n N_A_230_413#_c_204_n 0.0118613f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_129 N_B_M1002_g N_A_230_413#_c_196_n 0.0203093f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_130 N_B_c_165_n N_A_230_413#_c_198_n 0.00283241f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_131 N_B_M1002_g N_A_230_413#_c_198_n 0.0221059f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_132 B N_A_230_413#_c_198_n 0.0017542f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_133 N_B_c_165_n N_A_230_413#_c_209_n 0.0113795f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_134 B N_A_230_413#_c_209_n 0.0212144f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_135 N_B_M1002_g N_A_230_413#_c_201_n 0.00566552f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_136 N_B_c_165_n N_A_230_413#_c_202_n 0.044005f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_137 N_B_M1002_g N_A_230_413#_c_202_n 0.0169217f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_138 B N_A_230_413#_c_202_n 0.0360407f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_139 B N_A_230_413#_c_203_n 0.0151629f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_140 B N_VPWR_M1003_d 0.00847791f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_141 N_B_c_165_n N_VPWR_c_285_n 0.00742462f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_142 N_B_c_165_n N_VPWR_c_286_n 0.0071968f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_143 B N_VPWR_c_286_n 0.0494504f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_144 N_B_c_165_n N_VPWR_c_278_n 0.0144815f $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_145 B N_VPWR_c_278_n 0.00338833f $X=1.985 $Y=1.785 $X2=0 $Y2=0
cc_146 N_B_c_165_n X 5.07933e-19 $X=1.55 $Y=1.99 $X2=0 $Y2=0
cc_147 N_B_M1002_g N_VGND_c_350_n 0.00556028f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_148 N_B_M1002_g N_VGND_c_353_n 0.00583607f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_149 N_B_M1002_g N_VGND_c_356_n 0.0110194f $X=2.03 $Y=0.445 $X2=0 $Y2=0
cc_150 N_A_230_413#_c_209_n N_VPWR_c_279_n 0.0162919f $X=1.305 $Y=2.225 $X2=0
+ $Y2=0
cc_151 N_A_230_413#_c_207_n N_VPWR_c_281_n 0.0116196f $X=3.175 $Y=1.41 $X2=0
+ $Y2=0
cc_152 N_A_230_413#_c_204_n N_VPWR_c_283_n 0.00620778f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_153 N_A_230_413#_c_207_n N_VPWR_c_283_n 0.00696924f $X=3.175 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_230_413#_c_209_n N_VPWR_c_285_n 0.0158266f $X=1.305 $Y=2.225 $X2=0
+ $Y2=0
cc_155 N_A_230_413#_c_204_n N_VPWR_c_286_n 0.015118f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_A_230_413#_M1008_d N_VPWR_c_278_n 0.0033624f $X=1.15 $Y=2.065 $X2=0
+ $Y2=0
cc_157 N_A_230_413#_c_204_n N_VPWR_c_278_n 0.0122048f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_158 N_A_230_413#_c_207_n N_VPWR_c_278_n 0.0138035f $X=3.175 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_230_413#_c_209_n N_VPWR_c_278_n 0.0122726f $X=1.305 $Y=2.225 $X2=0
+ $Y2=0
cc_160 N_A_230_413#_c_197_n N_X_c_325_n 8.20839e-19 $X=3.075 $Y=1.155 $X2=0
+ $Y2=0
cc_161 N_A_230_413#_c_204_n X 0.00835409f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_230_413#_c_197_n X 0.00372899f $X=3.075 $Y=1.155 $X2=0 $Y2=0
cc_163 N_A_230_413#_c_207_n X 0.0106429f $X=3.175 $Y=1.41 $X2=0 $Y2=0
cc_164 N_A_230_413#_c_204_n X 0.0154838f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_230_413#_c_207_n X 0.0151303f $X=3.175 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_230_413#_c_204_n N_X_c_322_n 0.00378092f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_230_413#_c_196_n N_X_c_322_n 0.00506507f $X=2.57 $Y=0.985 $X2=0 $Y2=0
cc_168 N_A_230_413#_c_197_n N_X_c_322_n 0.0302008f $X=3.075 $Y=1.155 $X2=0 $Y2=0
cc_169 N_A_230_413#_c_198_n N_X_c_322_n 0.00126542f $X=2.645 $Y=1.155 $X2=0
+ $Y2=0
cc_170 N_A_230_413#_c_207_n N_X_c_322_n 0.00948517f $X=3.175 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_230_413#_c_199_n N_X_c_322_n 0.00735972f $X=3.2 $Y=0.985 $X2=0 $Y2=0
cc_172 N_A_230_413#_c_200_n N_X_c_322_n 0.0198273f $X=3.175 $Y=1.197 $X2=0 $Y2=0
cc_173 N_A_230_413#_c_202_n N_X_c_322_n 0.00475802f $X=2.105 $Y=1.135 $X2=0
+ $Y2=0
cc_174 N_A_230_413#_c_203_n N_X_c_322_n 0.0246823f $X=2.45 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_230_413#_c_196_n N_VGND_c_350_n 0.00350802f $X=2.57 $Y=0.985 $X2=0
+ $Y2=0
cc_176 N_A_230_413#_c_198_n N_VGND_c_350_n 9.07077e-19 $X=2.645 $Y=1.155 $X2=0
+ $Y2=0
cc_177 N_A_230_413#_c_203_n N_VGND_c_350_n 0.0162705f $X=2.45 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_230_413#_c_199_n N_VGND_c_352_n 0.00681587f $X=3.2 $Y=0.985 $X2=0
+ $Y2=0
cc_179 N_A_230_413#_c_226_n N_VGND_c_353_n 0.0182193f $X=1.3 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_230_413#_c_196_n N_VGND_c_355_n 0.00585385f $X=2.57 $Y=0.985 $X2=0
+ $Y2=0
cc_181 N_A_230_413#_c_199_n N_VGND_c_355_n 0.00585385f $X=3.2 $Y=0.985 $X2=0
+ $Y2=0
cc_182 N_A_230_413#_M1005_s N_VGND_c_356_n 0.00284954f $X=1.175 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_230_413#_c_196_n N_VGND_c_356_n 0.0113965f $X=2.57 $Y=0.985 $X2=0
+ $Y2=0
cc_184 N_A_230_413#_c_199_n N_VGND_c_356_n 0.0121673f $X=3.2 $Y=0.985 $X2=0
+ $Y2=0
cc_185 N_A_230_413#_c_226_n N_VGND_c_356_n 0.0153767f $X=1.3 $Y=0.445 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_278_n N_X_M1000_s 0.00380514f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_c_281_n X 0.0421988f $X=3.41 $Y=1.86 $X2=0 $Y2=0
cc_188 N_VPWR_c_283_n X 0.019433f $X=3.325 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_286_n X 0.0162258f $X=2.395 $Y=2.485 $X2=0 $Y2=0
cc_190 N_VPWR_c_278_n X 0.0183997f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_191 N_X_c_325_n N_VGND_c_355_n 0.0266233f $X=2.78 $Y=0.55 $X2=0 $Y2=0
cc_192 N_X_M1004_s N_VGND_c_356_n 0.00689478f $X=2.645 $Y=0.235 $X2=0 $Y2=0
cc_193 N_X_c_325_n N_VGND_c_356_n 0.0151194f $X=2.78 $Y=0.55 $X2=0 $Y2=0
cc_194 N_VGND_c_356_n A_327_47# 0.0126636f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
