* File: sky130_fd_sc_hdll__o211a_1.pxi.spice
* Created: Wed Sep  2 08:42:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__O211A_1%A_79_21# N_A_79_21#_M1006_d N_A_79_21#_M1005_d
+ N_A_79_21#_M1001_d N_A_79_21#_M1008_g N_A_79_21#_c_62_n N_A_79_21#_M1004_g
+ N_A_79_21#_c_63_n N_A_79_21#_c_64_n N_A_79_21#_c_76_p N_A_79_21#_c_69_n
+ N_A_79_21#_c_77_p N_A_79_21#_c_89_p N_A_79_21#_c_65_n N_A_79_21#_c_71_n
+ N_A_79_21#_c_84_p N_A_79_21#_c_66_n N_A_79_21#_c_72_n
+ PM_SKY130_FD_SC_HDLL__O211A_1%A_79_21#
x_PM_SKY130_FD_SC_HDLL__O211A_1%A1 N_A1_c_143_n N_A1_M1009_g N_A1_c_144_n
+ N_A1_M1007_g A1 A1 PM_SKY130_FD_SC_HDLL__O211A_1%A1
x_PM_SKY130_FD_SC_HDLL__O211A_1%A2 N_A2_c_175_n N_A2_M1000_g N_A2_c_176_n
+ N_A2_M1005_g A2 A2 PM_SKY130_FD_SC_HDLL__O211A_1%A2
x_PM_SKY130_FD_SC_HDLL__O211A_1%B1 N_B1_c_204_n N_B1_M1003_g N_B1_c_205_n
+ N_B1_M1002_g B1 N_B1_c_207_n B1 PM_SKY130_FD_SC_HDLL__O211A_1%B1
x_PM_SKY130_FD_SC_HDLL__O211A_1%C1 N_C1_c_239_n N_C1_M1006_g N_C1_c_243_n
+ N_C1_M1001_g N_C1_c_240_n C1 N_C1_c_242_n C1 PM_SKY130_FD_SC_HDLL__O211A_1%C1
x_PM_SKY130_FD_SC_HDLL__O211A_1%X N_X_M1008_s N_X_M1004_s N_X_c_268_n
+ N_X_c_271_n N_X_c_269_n X X X N_X_c_270_n PM_SKY130_FD_SC_HDLL__O211A_1%X
x_PM_SKY130_FD_SC_HDLL__O211A_1%VPWR N_VPWR_M1004_d N_VPWR_M1007_s
+ N_VPWR_M1002_d N_VPWR_c_290_n N_VPWR_c_291_n N_VPWR_c_292_n N_VPWR_c_293_n
+ VPWR N_VPWR_c_294_n N_VPWR_c_295_n N_VPWR_c_289_n N_VPWR_c_297_n
+ N_VPWR_c_298_n N_VPWR_c_299_n VPWR PM_SKY130_FD_SC_HDLL__O211A_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O211A_1%VGND N_VGND_M1008_d N_VGND_M1009_d
+ N_VGND_c_336_n N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n VGND
+ N_VGND_c_340_n N_VGND_c_341_n N_VGND_c_342_n VGND
+ PM_SKY130_FD_SC_HDLL__O211A_1%VGND
x_PM_SKY130_FD_SC_HDLL__O211A_1%A_225_47# N_A_225_47#_M1009_s
+ N_A_225_47#_M1000_d N_A_225_47#_c_383_n N_A_225_47#_c_384_n
+ N_A_225_47#_c_385_n N_A_225_47#_c_397_n
+ PM_SKY130_FD_SC_HDLL__O211A_1%A_225_47#
cc_1 VNB N_A_79_21#_M1008_g 0.0286055f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_79_21#_c_62_n 0.0413288f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_A_79_21#_c_63_n 0.017371f $X=-0.19 $Y=-0.24 $X2=1.005 $Y2=1.16
cc_4 VNB N_A_79_21#_c_64_n 0.00144235f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.495
cc_5 VNB N_A_79_21#_c_65_n 0.00586187f $X=-0.19 $Y=-0.24 $X2=3.36 $Y2=1.495
cc_6 VNB N_A_79_21#_c_66_n 0.0256142f $X=-0.19 $Y=-0.24 $X2=3.635 $Y2=0.38
cc_7 VNB N_A1_c_143_n 0.0226023f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.235
cc_8 VNB N_A1_c_144_n 0.0263327f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A1 0.00554039f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_10 VNB N_A2_c_175_n 0.018878f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.235
cc_11 VNB N_A2_c_176_n 0.0298171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A2 0.00178553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_B1_c_204_n 0.02028f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.235
cc_14 VNB N_B1_c_205_n 0.028613f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB B1 0.00550411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_B1_c_207_n 0.00167739f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_17 VNB N_C1_c_239_n 0.0216161f $X=-0.19 $Y=-0.24 $X2=3.41 $Y2=0.235
cc_18 VNB N_C1_c_240_n 0.0131496f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB C1 0.0093667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_C1_c_242_n 0.045757f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_21 VNB N_X_c_268_n 0.00778155f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_22 VNB N_X_c_269_n 0.0199656f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_23 VNB N_X_c_270_n 0.0183576f $X=-0.19 $Y=-0.24 $X2=1.09 $Y2=1.245
cc_24 VNB N_VPWR_c_289_n 0.17485f $X=-0.19 $Y=-0.24 $X2=3.635 $Y2=0.38
cc_25 VNB N_VGND_c_336_n 0.0128864f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_26 VNB N_VGND_c_337_n 0.00499625f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_27 VNB N_VGND_c_338_n 0.0194599f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_28 VNB N_VGND_c_339_n 0.00429685f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_29 VNB N_VGND_c_340_n 0.0633238f $X=-0.19 $Y=-0.24 $X2=3.25 $Y2=1.58
cc_30 VNB N_VGND_c_341_n 0.237782f $X=-0.19 $Y=-0.24 $X2=2.465 $Y2=1.58
cc_31 VNB N_VGND_c_342_n 0.0241682f $X=-0.19 $Y=-0.24 $X2=3.635 $Y2=1.665
cc_32 VNB N_A_225_47#_c_383_n 0.00464002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_225_47#_c_384_n 0.00633107f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_34 VNB N_A_225_47#_c_385_n 0.00578617f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_35 VPB N_A_79_21#_c_62_n 0.0317272f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_A_79_21#_c_64_n 0.00518356f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.495
cc_37 VPB N_A_79_21#_c_69_n 0.00555846f $X=-0.19 $Y=1.305 $X2=1.175 $Y2=1.58
cc_38 VPB N_A_79_21#_c_65_n 0.00667971f $X=-0.19 $Y=1.305 $X2=3.36 $Y2=1.495
cc_39 VPB N_A_79_21#_c_71_n 0.0312141f $X=-0.19 $Y=1.305 $X2=3.635 $Y2=2.34
cc_40 VPB N_A_79_21#_c_72_n 0.00740132f $X=-0.19 $Y=1.305 $X2=3.635 $Y2=1.66
cc_41 VPB N_A1_c_144_n 0.0302232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A2_c_176_n 0.0315457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_B1_c_205_n 0.0309112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_C1_c_243_n 0.0208352f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_C1_c_240_n 0.00730163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB C1 0.00143781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_C1_c_242_n 0.0192955f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.56
cc_48 VPB N_X_c_271_n 0.00666696f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_X_c_269_n 0.00910093f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_50 VPB X 0.0316915f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_51 VPB N_VPWR_c_290_n 0.00356354f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_52 VPB N_VPWR_c_291_n 0.0085283f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_53 VPB N_VPWR_c_292_n 0.00956783f $X=-0.19 $Y=1.305 $X2=1.09 $Y2=1.245
cc_54 VPB N_VPWR_c_293_n 0.00562936f $X=-0.19 $Y=1.305 $X2=2.275 $Y2=1.665
cc_55 VPB N_VPWR_c_294_n 0.0416021f $X=-0.19 $Y=1.305 $X2=3.25 $Y2=1.58
cc_56 VPB N_VPWR_c_295_n 0.0324707f $X=-0.19 $Y=1.305 $X2=3.525 $Y2=0.38
cc_57 VPB N_VPWR_c_289_n 0.0636734f $X=-0.19 $Y=1.305 $X2=3.635 $Y2=0.38
cc_58 VPB N_VPWR_c_297_n 0.0226069f $X=-0.19 $Y=1.305 $X2=3.525 $Y2=1.58
cc_59 VPB N_VPWR_c_298_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_299_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_62_n N_A1_c_144_n 0.00476406f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_63_n N_A1_c_144_n 7.43208e-19 $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_64_n N_A1_c_144_n 0.00732921f $X=1.09 $Y=1.495 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_76_p N_A1_c_144_n 0.0220578f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_77_p N_A1_c_144_n 0.00360192f $X=2.3 $Y=2.34 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_62_n A1 3.88392e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_63_n A1 0.0150768f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_64_n A1 0.00228843f $X=1.09 $Y=1.495 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_76_p A1 0.0241967f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_76_p N_A2_c_176_n 0.0154801f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_77_p N_A2_c_176_n 0.0275672f $X=2.3 $Y=2.34 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_84_p N_A2_c_176_n 0.00870654f $X=2.3 $Y=1.66 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_76_p A2 0.00555769f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_84_p A2 0.0166119f $X=2.3 $Y=1.66 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_65_n N_B1_c_204_n 6.99325e-19 $X=3.36 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_79_21#_c_77_p N_B1_c_205_n 0.0119441f $X=2.3 $Y=2.34 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_89_p N_B1_c_205_n 0.022597f $X=3.25 $Y=1.58 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_65_n N_B1_c_205_n 0.00434922f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_89_p B1 0.0179079f $X=3.25 $Y=1.58 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_65_n B1 0.049561f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_89_p N_B1_c_207_n 0.0132911f $X=3.25 $Y=1.58 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_65_n N_C1_c_239_n 0.00524254f $X=3.36 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_79_21#_c_66_n N_C1_c_239_n 0.0279299f $X=3.635 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_79_21#_c_65_n N_C1_c_243_n 0.00350894f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_72_n N_C1_c_243_n 0.0152516f $X=3.635 $Y=1.66 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_65_n N_C1_c_240_n 0.0129503f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_65_n C1 0.0182893f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_66_n C1 0.0109158f $X=3.635 $Y=0.38 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_72_n C1 0.0130317f $X=3.635 $Y=1.66 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_65_n N_C1_c_242_n 0.0075252f $X=3.36 $Y=1.495 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_66_n N_C1_c_242_n 0.0092386f $X=3.635 $Y=0.38 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_72_n N_C1_c_242_n 0.00842771f $X=3.635 $Y=1.66 $X2=0 $Y2=0
cc_93 N_A_79_21#_M1008_g N_X_c_268_n 0.00282668f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_62_n N_X_c_271_n 0.00258239f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_79_21#_M1008_g N_X_c_269_n 0.015656f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_62_n N_X_c_269_n 0.00124306f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_63_n N_X_c_269_n 0.0134533f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_62_n X 0.0100147f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_79_21#_M1008_g N_X_c_270_n 0.00588415f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_76_p N_VPWR_M1007_s 0.00523571f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_69_n N_VPWR_M1007_s 0.00101038f $X=1.175 $Y=1.58 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_89_p N_VPWR_M1002_d 0.0175589f $X=3.25 $Y=1.58 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_62_n N_VPWR_c_290_n 0.0118122f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_63_n N_VPWR_c_290_n 0.00987815f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_69_n N_VPWR_c_290_n 0.0130372f $X=1.175 $Y=1.58 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_76_p N_VPWR_c_292_n 0.0128995f $X=2.085 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_69_n N_VPWR_c_292_n 0.0080326f $X=1.175 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_89_p N_VPWR_c_293_n 0.0237567f $X=3.25 $Y=1.58 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_77_p N_VPWR_c_294_n 0.0245654f $X=2.3 $Y=2.34 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_71_n N_VPWR_c_295_n 0.0218646f $X=3.635 $Y=2.34 $X2=0 $Y2=0
cc_111 N_A_79_21#_M1005_d N_VPWR_c_289_n 0.00704327f $X=2.1 $Y=1.485 $X2=0 $Y2=0
cc_112 N_A_79_21#_M1001_d N_VPWR_c_289_n 0.0031974f $X=3.45 $Y=1.485 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_62_n N_VPWR_c_289_n 0.0140376f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_77_p N_VPWR_c_289_n 0.0144934f $X=2.3 $Y=2.34 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_71_n N_VPWR_c_289_n 0.0126319f $X=3.635 $Y=2.34 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_62_n N_VPWR_c_297_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_76_p A_315_297# 0.0117615f $X=2.085 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_79_21#_M1008_g N_VGND_c_336_n 0.00667329f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_62_n N_VGND_c_336_n 0.00386516f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_63_n N_VGND_c_336_n 0.0183552f $X=1.005 $Y=1.16 $X2=0 $Y2=0
cc_121 N_A_79_21#_c_66_n N_VGND_c_340_n 0.0357845f $X=3.635 $Y=0.38 $X2=0 $Y2=0
cc_122 N_A_79_21#_M1006_d N_VGND_c_341_n 0.00283904f $X=3.41 $Y=0.235 $X2=0
+ $Y2=0
cc_123 N_A_79_21#_M1008_g N_VGND_c_341_n 0.0119046f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_66_n N_VGND_c_341_n 0.0203825f $X=3.635 $Y=0.38 $X2=0 $Y2=0
cc_125 N_A_79_21#_M1008_g N_VGND_c_342_n 0.00541359f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_76_p N_A_225_47#_c_384_n 0.00389298f $X=2.085 $Y=1.58 $X2=0
+ $Y2=0
cc_127 N_A_79_21#_c_84_p N_A_225_47#_c_384_n 0.00148729f $X=2.3 $Y=1.66 $X2=0
+ $Y2=0
cc_128 N_A_79_21#_M1008_g N_A_225_47#_c_385_n 8.16329e-19 $X=0.47 $Y=0.56 $X2=0
+ $Y2=0
cc_129 N_A_79_21#_c_63_n N_A_225_47#_c_385_n 0.00831554f $X=1.005 $Y=1.16 $X2=0
+ $Y2=0
cc_130 N_A_79_21#_c_76_p N_A_225_47#_c_385_n 0.00573213f $X=2.085 $Y=1.58 $X2=0
+ $Y2=0
cc_131 N_A1_c_143_n N_A2_c_175_n 0.0219441f $X=1.46 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_132 N_A1_c_144_n N_A2_c_176_n 0.0696503f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_133 A1 N_A2_c_176_n 0.0013876f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_134 A1 A2 0.016441f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_135 N_A1_c_144_n N_VPWR_c_290_n 0.00524066f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_144_n N_VPWR_c_292_n 0.0182977f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_144_n N_VPWR_c_294_n 0.00702461f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_144_n N_VPWR_c_289_n 0.0140259f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A1_c_143_n N_VGND_c_336_n 0.0022981f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_143_n N_VGND_c_337_n 0.00551294f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_143_n N_VGND_c_338_n 0.00424416f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_143_n N_VGND_c_341_n 0.00750329f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_143_n N_A_225_47#_c_383_n 0.007367f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_143_n N_A_225_47#_c_384_n 0.00901637f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A1_c_144_n N_A_225_47#_c_384_n 0.00425056f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_146 A1 N_A_225_47#_c_384_n 0.0289125f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_147 N_A1_c_143_n N_A_225_47#_c_385_n 0.00126808f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_148 A1 N_A_225_47#_c_385_n 0.00528093f $X=1.635 $Y=1.19 $X2=0 $Y2=0
cc_149 N_A1_c_143_n N_A_225_47#_c_397_n 6.56096e-19 $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A2_c_175_n N_B1_c_204_n 0.0114677f $X=1.985 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_151 N_A2_c_176_n N_B1_c_205_n 0.0521301f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_152 A2 N_B1_c_205_n 6.51034e-19 $X=2.16 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A2_c_176_n B1 3.38293e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A2_c_176_n N_B1_c_207_n 6.58846e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_155 A2 N_B1_c_207_n 0.0174693f $X=2.16 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A2_c_176_n N_VPWR_c_294_n 0.00681208f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A2_c_176_n N_VPWR_c_289_n 0.0127906f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A2_c_175_n N_VGND_c_337_n 0.00291779f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A2_c_175_n N_VGND_c_340_n 0.00424416f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A2_c_175_n N_VGND_c_341_n 0.00647541f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A2_c_175_n N_A_225_47#_c_383_n 6.02202e-19 $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A2_c_175_n N_A_225_47#_c_384_n 0.0111662f $X=1.985 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_176_n N_A_225_47#_c_384_n 0.00735006f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_164 A2 N_A_225_47#_c_384_n 0.0306523f $X=2.16 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A2_c_175_n N_A_225_47#_c_397_n 0.00702357f $X=1.985 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_B1_c_204_n N_C1_c_239_n 0.0139042f $X=2.625 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_167 B1 N_C1_c_239_n 0.0025675f $X=2.62 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_168 N_B1_c_205_n N_C1_c_243_n 0.0165977f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B1_c_205_n N_C1_c_240_n 0.011941f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_170 B1 N_C1_c_240_n 7.91939e-19 $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_171 N_B1_c_205_n N_VPWR_c_293_n 0.00344738f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B1_c_205_n N_VPWR_c_294_n 0.00702461f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B1_c_205_n N_VPWR_c_289_n 0.0133667f $X=2.65 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B1_c_204_n N_VGND_c_340_n 0.00585385f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_175 B1 N_VGND_c_340_n 0.0084617f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_176 N_B1_c_204_n N_VGND_c_341_n 0.0119128f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_177 B1 N_VGND_c_341_n 0.00911787f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_178 N_B1_c_204_n N_A_225_47#_c_384_n 0.0021662f $X=2.625 $Y=0.995 $X2=0 $Y2=0
cc_179 B1 N_A_225_47#_c_384_n 0.00756008f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_180 N_B1_c_204_n N_A_225_47#_c_397_n 0.00843501f $X=2.625 $Y=0.995 $X2=0
+ $Y2=0
cc_181 B1 N_A_225_47#_c_397_n 0.0125864f $X=2.62 $Y=1.105 $X2=0 $Y2=0
cc_182 B1 A_540_47# 0.0184096f $X=2.62 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_183 N_C1_c_243_n N_VPWR_c_293_n 0.00992288f $X=3.36 $Y=1.41 $X2=0 $Y2=0
cc_184 N_C1_c_243_n N_VPWR_c_295_n 0.00702461f $X=3.36 $Y=1.41 $X2=0 $Y2=0
cc_185 N_C1_c_243_n N_VPWR_c_289_n 0.0142837f $X=3.36 $Y=1.41 $X2=0 $Y2=0
cc_186 N_C1_c_239_n N_VGND_c_340_n 0.00357668f $X=3.335 $Y=0.995 $X2=0 $Y2=0
cc_187 N_C1_c_239_n N_VGND_c_341_n 0.00724809f $X=3.335 $Y=0.995 $X2=0 $Y2=0
cc_188 N_X_c_271_n N_VPWR_c_290_n 0.0588307f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_189 N_X_M1004_s N_VPWR_c_289_n 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_190 X N_VPWR_c_289_n 0.0128576f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_191 X N_VPWR_c_297_n 0.0217765f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_192 N_X_c_270_n N_VGND_c_336_n 0.0393237f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_193 N_X_M1008_s N_VGND_c_341_n 0.00209319f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_194 N_X_c_270_n N_VGND_c_341_n 0.0127994f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_195 N_X_c_270_n N_VGND_c_342_n 0.0217139f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_196 N_VPWR_c_289_n A_315_297# 0.0147472f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_197 N_VGND_c_341_n N_A_225_47#_M1009_s 0.00209319f $X=3.91 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_198 N_VGND_c_341_n N_A_225_47#_M1000_d 0.00884338f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_199 N_VGND_c_336_n N_A_225_47#_c_383_n 0.036162f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_200 N_VGND_c_337_n N_A_225_47#_c_383_n 0.0179308f $X=1.75 $Y=0.38 $X2=0 $Y2=0
cc_201 N_VGND_c_338_n N_A_225_47#_c_383_n 0.0209752f $X=1.635 $Y=0 $X2=0 $Y2=0
cc_202 N_VGND_c_341_n N_A_225_47#_c_383_n 0.0124119f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_203 N_VGND_M1009_d N_A_225_47#_c_384_n 0.00331634f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_204 N_VGND_c_337_n N_A_225_47#_c_384_n 0.015465f $X=1.75 $Y=0.38 $X2=0 $Y2=0
cc_205 N_VGND_c_338_n N_A_225_47#_c_384_n 0.00260082f $X=1.635 $Y=0 $X2=0 $Y2=0
cc_206 N_VGND_c_340_n N_A_225_47#_c_384_n 0.00193763f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_207 N_VGND_c_341_n N_A_225_47#_c_384_n 0.00989411f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_208 N_VGND_c_336_n N_A_225_47#_c_385_n 0.0120261f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_209 N_VGND_c_340_n N_A_225_47#_c_397_n 0.0244265f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_210 N_VGND_c_341_n N_A_225_47#_c_397_n 0.0143352f $X=3.91 $Y=0 $X2=0 $Y2=0
cc_211 N_VGND_c_341_n A_540_47# 0.0148121f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
