# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21boi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21boi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 0.995000 3.565000 1.325000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.295000 1.075000 2.675000 1.245000 ;
        RECT 2.300000 1.245000 2.675000 1.495000 ;
        RECT 2.300000 1.495000 4.085000 1.675000 ;
        RECT 3.735000 0.995000 4.085000 1.495000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.120000 0.765000 0.425000 1.805000 ;
    END
  END B1_N
  PIN VGND
    ANTENNADIFFAREA  0.884500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.790000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  0.705500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  0.712500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.525000 0.255000 1.870000 0.615000 ;
        RECT 1.525000 0.615000 3.360000 0.785000 ;
        RECT 1.525000 0.785000 1.865000 2.115000 ;
        RECT 2.980000 0.255000 3.360000 0.615000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.095000  2.080000 0.425000 2.635000 ;
      RECT 0.265000  0.360000 0.825000 0.530000 ;
      RECT 0.645000  0.530000 0.825000 1.070000 ;
      RECT 0.645000  1.070000 1.355000 1.285000 ;
      RECT 0.645000  1.285000 0.825000 2.265000 ;
      RECT 1.085000  0.085000 1.325000 0.885000 ;
      RECT 1.100000  1.795000 1.350000 2.285000 ;
      RECT 1.100000  2.285000 2.415000 2.465000 ;
      RECT 2.035000  1.855000 4.320000 2.025000 ;
      RECT 2.035000  2.025000 2.415000 2.285000 ;
      RECT 2.140000  0.085000 2.470000 0.445000 ;
      RECT 2.635000  2.195000 2.805000 2.635000 ;
      RECT 3.110000  2.025000 4.320000 2.105000 ;
      RECT 3.110000  2.105000 3.280000 2.465000 ;
      RECT 3.460000  2.275000 3.840000 2.635000 ;
      RECT 3.990000  0.085000 4.330000 0.785000 ;
      RECT 4.060000  2.105000 4.320000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21boi_2
END LIBRARY
