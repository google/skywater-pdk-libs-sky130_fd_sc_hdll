# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__clkmux2_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__clkmux2_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.670000 0.255000 3.995000 1.415000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.232200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.160000 0.810000 3.330000 1.615000 ;
        RECT 3.160000 1.615000 4.455000 1.785000 ;
        RECT 4.165000 0.255000 4.455000 1.615000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  0.479400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.995000 2.650000 1.325000 ;
        RECT 2.450000 1.325000 2.650000 2.295000 ;
        RECT 2.450000 2.295000 4.795000 2.465000 ;
        RECT 4.625000 1.440000 5.375000 1.630000 ;
        RECT 4.625000 1.630000 4.795000 2.295000 ;
        RECT 5.185000 1.055000 5.375000 1.440000 ;
    END
  END S
  PIN X
    ANTENNADIFFAREA  0.860800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.565000 1.495000 0.895000 2.465000 ;
        RECT 0.590000 0.255000 0.850000 1.065000 ;
        RECT 0.590000 1.065000 1.745000 1.325000 ;
        RECT 0.590000 1.325000 0.850000 1.495000 ;
        RECT 1.475000 0.255000 1.745000 1.065000 ;
        RECT 1.475000 1.325000 1.745000 1.495000 ;
        RECT 1.475000 1.495000 1.835000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 0.175000  0.085000 0.420000 0.655000 ;
        RECT 1.055000  0.085000 1.305000 0.655000 ;
        RECT 1.915000  0.085000 2.275000 0.485000 ;
        RECT 4.630000  0.085000 5.145000 0.525000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
        RECT 0.135000 1.495000 0.395000 2.635000 ;
        RECT 1.065000 1.495000 1.305000 2.635000 ;
        RECT 2.005000 1.495000 2.280000 2.635000 ;
        RECT 4.965000 1.835000 5.195000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.915000 0.655000 2.990000 0.825000 ;
      RECT 1.915000 0.825000 2.085000 1.325000 ;
      RECT 2.815000 0.255000 3.500000 0.620000 ;
      RECT 2.815000 0.620000 2.990000 0.655000 ;
      RECT 2.820000 0.825000 2.990000 1.955000 ;
      RECT 2.820000 1.955000 4.265000 2.125000 ;
      RECT 4.705000 0.695000 5.765000 0.865000 ;
      RECT 4.705000 0.865000 4.875000 1.185000 ;
      RECT 5.365000 1.835000 5.765000 2.465000 ;
      RECT 5.415000 0.255000 5.660000 0.695000 ;
      RECT 5.595000 0.865000 5.765000 1.835000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__clkmux2_4
