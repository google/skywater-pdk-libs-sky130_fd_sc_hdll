* File: sky130_fd_sc_hdll__or4bb_1.pxi.spice
* Created: Wed Sep  2 08:49:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%C_N N_C_N_c_96_n N_C_N_c_97_n N_C_N_M1011_g
+ N_C_N_M1006_g C_N C_N N_C_N_c_94_n N_C_N_c_95_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_1%C_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%D_N N_D_N_c_126_n N_D_N_M1003_g N_D_N_c_127_n
+ N_D_N_M1012_g D_N D_N PM_SKY130_FD_SC_HDLL__OR4BB_1%D_N
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%A_216_93# N_A_216_93#_M1003_d
+ N_A_216_93#_M1012_d N_A_216_93#_c_167_n N_A_216_93#_c_168_n
+ N_A_216_93#_M1002_g N_A_216_93#_M1010_g N_A_216_93#_c_169_n
+ N_A_216_93#_c_161_n N_A_216_93#_c_162_n N_A_216_93#_c_163_n
+ N_A_216_93#_c_164_n N_A_216_93#_c_165_n N_A_216_93#_c_166_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_1%A_216_93#
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%A_27_410# N_A_27_410#_M1006_s
+ N_A_27_410#_M1011_s N_A_27_410#_M1007_g N_A_27_410#_c_229_n
+ N_A_27_410#_M1013_g N_A_27_410#_c_230_n N_A_27_410#_c_235_n
+ N_A_27_410#_c_236_n N_A_27_410#_c_237_n N_A_27_410#_c_238_n
+ N_A_27_410#_c_239_n N_A_27_410#_c_231_n N_A_27_410#_c_232_n
+ N_A_27_410#_c_241_n PM_SKY130_FD_SC_HDLL__OR4BB_1%A_27_410#
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%B N_B_c_320_n N_B_c_321_n N_B_c_323_n
+ N_B_c_324_n N_B_M1001_g N_B_M1004_g N_B_c_322_n B B
+ PM_SKY130_FD_SC_HDLL__OR4BB_1%B
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%A N_A_c_363_n N_A_M1008_g N_A_M1005_g A
+ N_A_c_365_n A PM_SKY130_FD_SC_HDLL__OR4BB_1%A
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%A_331_413# N_A_331_413#_M1010_d
+ N_A_331_413#_M1004_d N_A_331_413#_M1002_s N_A_331_413#_c_401_n
+ N_A_331_413#_M1000_g N_A_331_413#_c_402_n N_A_331_413#_M1009_g
+ N_A_331_413#_c_410_n N_A_331_413#_c_422_n N_A_331_413#_c_411_n
+ N_A_331_413#_c_403_n N_A_331_413#_c_404_n N_A_331_413#_c_412_n
+ N_A_331_413#_c_419_n N_A_331_413#_c_498_p N_A_331_413#_c_405_n
+ N_A_331_413#_c_457_n N_A_331_413#_c_413_n N_A_331_413#_c_406_n
+ N_A_331_413#_c_414_n N_A_331_413#_c_407_n N_A_331_413#_c_408_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_1%A_331_413#
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%VPWR N_VPWR_M1011_d N_VPWR_M1008_d
+ N_VPWR_c_512_n N_VPWR_c_513_n N_VPWR_c_514_n N_VPWR_c_515_n VPWR
+ N_VPWR_c_516_n N_VPWR_c_517_n N_VPWR_c_511_n N_VPWR_c_519_n
+ PM_SKY130_FD_SC_HDLL__OR4BB_1%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%X N_X_M1009_d N_X_M1000_d N_X_c_569_n
+ N_X_c_571_n N_X_c_570_n X PM_SKY130_FD_SC_HDLL__OR4BB_1%X
x_PM_SKY130_FD_SC_HDLL__OR4BB_1%VGND N_VGND_M1006_d N_VGND_M1010_s
+ N_VGND_M1007_d N_VGND_M1005_d N_VGND_c_587_n N_VGND_c_588_n N_VGND_c_589_n
+ N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n N_VGND_c_593_n N_VGND_c_594_n
+ N_VGND_c_595_n VGND N_VGND_c_596_n N_VGND_c_597_n N_VGND_c_598_n
+ N_VGND_c_599_n PM_SKY130_FD_SC_HDLL__OR4BB_1%VGND
cc_1 VNB C_N 0.00812127f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.105
cc_2 VNB N_C_N_c_94_n 0.024143f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_3 VNB N_C_N_c_95_n 0.0209269f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_4 VNB N_D_N_c_126_n 0.0191088f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_5 VNB N_D_N_c_127_n 0.0273388f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_6 VNB D_N 0.00347298f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.675
cc_7 VNB N_A_216_93#_M1010_g 0.0343207f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_8 VNB N_A_216_93#_c_161_n 0.00648104f $X=-0.19 $Y=-0.24 $X2=0.617 $Y2=1.53
cc_9 VNB N_A_216_93#_c_162_n 0.00126747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_216_93#_c_163_n 0.00792919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_216_93#_c_164_n 0.0257214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_216_93#_c_165_n 0.0127908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_216_93#_c_166_n 0.00204729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_410#_M1007_g 0.0275893f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=1.445
cc_15 VNB N_A_27_410#_c_229_n 0.0252791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_410#_c_230_n 0.0223313f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_17 VNB N_A_27_410#_c_231_n 6.93211e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_410#_c_232_n 0.0186312f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B_c_320_n 0.00670451f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_20 VNB N_B_c_321_n 0.0211181f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.875
cc_21 VNB N_B_c_322_n 0.0158925f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.105
cc_22 VNB N_A_c_363_n 0.0190833f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_23 VNB N_A_M1005_g 0.0293196f $X=-0.19 $Y=-0.24 $X2=0.555 $Y2=0.995
cc_24 VNB N_A_c_365_n 0.00682249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_331_413#_c_401_n 0.0235264f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.105
cc_26 VNB N_A_331_413#_c_402_n 0.0204639f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_27 VNB N_A_331_413#_c_403_n 0.0129372f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_331_413#_c_404_n 0.0047498f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_331_413#_c_405_n 0.00347822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_331_413#_c_406_n 0.0015089f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_331_413#_c_407_n 0.00264294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_331_413#_c_408_n 0.0018431f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VPWR_c_511_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_569_n 0.0150464f $X=-0.19 $Y=-0.24 $X2=0.55 $Y2=1.105
cc_35 VNB N_X_c_570_n 0.0261739f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_36 VNB N_VGND_c_587_n 0.0151265f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_37 VNB N_VGND_c_588_n 0.0200032f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.325
cc_38 VNB N_VGND_c_589_n 0.012349f $X=-0.19 $Y=-0.24 $X2=0.617 $Y2=1.53
cc_39 VNB N_VGND_c_590_n 0.0149555f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_591_n 0.00206109f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_592_n 0.0225599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_593_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_594_n 0.00973217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_595_n 0.0135819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_596_n 0.0224629f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_597_n 0.264989f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_598_n 0.00718038f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_599_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VPB N_C_N_c_96_n 0.0336701f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.875
cc_50 VPB N_C_N_c_97_n 0.0286094f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_51 VPB C_N 0.00247995f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.105
cc_52 VPB N_C_N_c_94_n 0.00328006f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_53 VPB N_D_N_c_127_n 0.0289916f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_54 VPB D_N 0.00146519f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.675
cc_55 VPB N_A_216_93#_c_167_n 0.0386139f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.675
cc_56 VPB N_A_216_93#_c_168_n 0.0307681f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.445
cc_57 VPB N_A_216_93#_c_169_n 0.00838936f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_58 VPB N_A_216_93#_c_162_n 0.0054644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_216_93#_c_164_n 0.00340539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_27_410#_c_229_n 0.0265239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_410#_c_230_n 0.0262129f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_62 VPB N_A_27_410#_c_235_n 0.0164639f $X=-0.19 $Y=1.305 $X2=0.617 $Y2=1.16
cc_63 VPB N_A_27_410#_c_236_n 0.0217044f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_410#_c_237_n 0.00680513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_410#_c_238_n 0.00488674f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_410#_c_239_n 0.00201281f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_410#_c_231_n 9.16142e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_410#_c_241_n 0.0113037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_B_c_323_n 0.00604637f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_70 VPB N_B_c_324_n 0.0514871f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_71 VPB N_B_M1001_g 0.0107583f $X=-0.19 $Y=1.305 $X2=0.555 $Y2=0.995
cc_72 VPB B 0.0144513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_c_363_n 0.0267577f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_74 VPB N_A_c_365_n 0.00378552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_331_413#_c_401_n 0.0318711f $X=-0.19 $Y=1.305 $X2=0.55 $Y2=1.105
cc_76 VPB N_A_331_413#_c_410_n 0.00985638f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_77 VPB N_A_331_413#_c_411_n 0.00256019f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_331_413#_c_412_n 0.00427396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_331_413#_c_413_n 0.00156472f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_331_413#_c_414_n 0.00139492f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_512_n 0.0143673f $X=-0.19 $Y=1.305 $X2=0.525 $Y2=1.445
cc_82 VPB N_VPWR_c_513_n 0.0111765f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_83 VPB N_VPWR_c_514_n 0.0702098f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=0.995
cc_84 VPB N_VPWR_c_515_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.325
cc_85 VPB N_VPWR_c_516_n 0.0145108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_517_n 0.0223347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_511_n 0.0704005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_519_n 0.00593769f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_X_c_571_n 0.00661942f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_90 VPB N_X_c_570_n 0.00946273f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_91 VPB X 0.0336954f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_92 N_C_N_c_95_n N_D_N_c_126_n 0.0103106f $X=0.53 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_C_N_c_96_n N_D_N_c_127_n 0.0219858f $X=0.495 $Y=1.875 $X2=0 $Y2=0
cc_94 N_C_N_c_97_n N_D_N_c_127_n 0.00196932f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_95 C_N N_D_N_c_127_n 0.00906834f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_96 N_C_N_c_94_n N_D_N_c_127_n 0.0149278f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_97 C_N D_N 0.0265444f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_98 N_C_N_c_94_n D_N 3.00501e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_99 C_N N_A_216_93#_c_169_n 0.0110254f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_100 C_N N_A_27_410#_c_230_n 0.0531961f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_101 N_C_N_c_94_n N_A_27_410#_c_230_n 0.0212915f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_102 N_C_N_c_95_n N_A_27_410#_c_230_n 0.00499222f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_103 N_C_N_c_97_n N_A_27_410#_c_235_n 0.00559296f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_104 N_C_N_c_96_n N_A_27_410#_c_236_n 0.00410106f $X=0.495 $Y=1.875 $X2=0
+ $Y2=0
cc_105 N_C_N_c_97_n N_A_27_410#_c_236_n 0.0121812f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_106 C_N N_A_27_410#_c_236_n 0.0305906f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_107 N_C_N_c_94_n N_A_27_410#_c_236_n 2.25066e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_108 N_C_N_c_94_n N_A_27_410#_c_232_n 2.24832e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_109 N_C_N_c_95_n N_A_27_410#_c_232_n 0.00217458f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_110 C_N N_VPWR_M1011_d 0.00399732f $X=0.55 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 N_C_N_c_97_n N_VPWR_c_512_n 0.0127593f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_112 N_C_N_c_97_n N_VPWR_c_516_n 0.00310301f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_113 N_C_N_c_97_n N_VPWR_c_511_n 0.00460685f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_114 C_N N_VGND_c_587_n 0.00948983f $X=0.55 $Y=1.105 $X2=0 $Y2=0
cc_115 N_C_N_c_95_n N_VGND_c_587_n 0.00447907f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C_N_c_95_n N_VGND_c_592_n 0.00510437f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_N_c_95_n N_VGND_c_597_n 0.00512902f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_118 N_D_N_c_127_n N_A_216_93#_c_169_n 0.00640208f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_119 D_N N_A_216_93#_c_169_n 0.0177237f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_120 N_D_N_c_126_n N_A_216_93#_c_161_n 0.00403266f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_121 N_D_N_c_127_n N_A_216_93#_c_161_n 2.26168e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_122 D_N N_A_216_93#_c_161_n 0.00629095f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_123 N_D_N_c_127_n N_A_216_93#_c_162_n 0.00525734f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_124 D_N N_A_216_93#_c_162_n 0.00629095f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_125 N_D_N_c_127_n N_A_216_93#_c_164_n 0.00391977f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_126 D_N N_A_216_93#_c_164_n 5.90824e-19 $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_127 N_D_N_c_126_n N_A_216_93#_c_165_n 0.00207532f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_D_N_c_127_n N_A_216_93#_c_165_n 5.71859e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_129 D_N N_A_216_93#_c_165_n 0.0131611f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_130 N_D_N_c_127_n N_A_216_93#_c_166_n 5.92982e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_131 D_N N_A_216_93#_c_166_n 0.0151326f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_132 N_D_N_c_127_n N_A_27_410#_c_236_n 0.0163179f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_133 D_N N_A_27_410#_c_236_n 0.00166112f $X=1.165 $Y=1.105 $X2=0 $Y2=0
cc_134 N_D_N_c_127_n N_VPWR_c_514_n 0.0031102f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_135 N_D_N_c_127_n N_VPWR_c_511_n 0.00500987f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_136 N_D_N_c_126_n N_VGND_c_587_n 0.0029062f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_137 N_D_N_c_126_n N_VGND_c_588_n 0.00510437f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_138 N_D_N_c_126_n N_VGND_c_589_n 0.0031643f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_139 N_D_N_c_126_n N_VGND_c_597_n 0.00512902f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_216_93#_M1010_g N_A_27_410#_M1007_g 0.0246037f $X=2.04 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_216_93#_c_167_n N_A_27_410#_c_229_n 0.0229713f $X=2.015 $Y=1.89 $X2=0
+ $Y2=0
cc_142 N_A_216_93#_c_168_n N_A_27_410#_c_229_n 0.00116326f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_143 N_A_216_93#_c_163_n N_A_27_410#_c_229_n 0.00114879f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_144 N_A_216_93#_c_164_n N_A_27_410#_c_229_n 0.0209994f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_216_93#_M1012_d N_A_27_410#_c_236_n 0.00269571f $X=1.12 $Y=1.485
+ $X2=0 $Y2=0
cc_146 N_A_216_93#_c_167_n N_A_27_410#_c_236_n 0.00101201f $X=2.015 $Y=1.89
+ $X2=0 $Y2=0
cc_147 N_A_216_93#_c_168_n N_A_27_410#_c_236_n 0.00744737f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_148 N_A_216_93#_c_169_n N_A_27_410#_c_236_n 0.043693f $X=1.505 $Y=1.61 $X2=0
+ $Y2=0
cc_149 N_A_216_93#_c_163_n N_A_27_410#_c_236_n 0.005133f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_150 N_A_216_93#_c_167_n N_A_27_410#_c_237_n 0.0105998f $X=2.015 $Y=1.89 $X2=0
+ $Y2=0
cc_151 N_A_216_93#_c_169_n N_A_27_410#_c_237_n 0.00919945f $X=1.505 $Y=1.61
+ $X2=0 $Y2=0
cc_152 N_A_216_93#_c_167_n N_A_27_410#_c_238_n 0.0079317f $X=2.015 $Y=1.89 $X2=0
+ $Y2=0
cc_153 N_A_216_93#_c_163_n N_A_27_410#_c_238_n 0.00975618f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_154 N_A_216_93#_c_167_n N_A_27_410#_c_239_n 0.00568385f $X=2.015 $Y=1.89
+ $X2=0 $Y2=0
cc_155 N_A_216_93#_c_169_n N_A_27_410#_c_239_n 0.00560512f $X=1.505 $Y=1.61
+ $X2=0 $Y2=0
cc_156 N_A_216_93#_c_162_n N_A_27_410#_c_239_n 0.0092742f $X=1.59 $Y=1.525 $X2=0
+ $Y2=0
cc_157 N_A_216_93#_c_163_n N_A_27_410#_c_239_n 0.0131609f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_216_93#_c_164_n N_A_27_410#_c_239_n 0.00178889f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_159 N_A_216_93#_c_167_n N_A_27_410#_c_231_n 0.00171119f $X=2.015 $Y=1.89
+ $X2=0 $Y2=0
cc_160 N_A_216_93#_c_163_n N_A_27_410#_c_231_n 0.0111379f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_216_93#_c_164_n N_A_27_410#_c_231_n 0.00120304f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_216_93#_c_168_n B 0.00308444f $X=2.015 $Y=1.99 $X2=0 $Y2=0
cc_163 N_A_216_93#_c_168_n N_A_331_413#_c_410_n 0.0121727f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_164 N_A_216_93#_c_168_n N_A_331_413#_c_411_n 0.00679125f $X=2.015 $Y=1.99
+ $X2=0 $Y2=0
cc_165 N_A_216_93#_M1010_g N_A_331_413#_c_404_n 0.00249682f $X=2.04 $Y=0.445
+ $X2=0 $Y2=0
cc_166 N_A_216_93#_c_165_n N_A_331_413#_c_404_n 0.00737188f $X=1.26 $Y=0.66
+ $X2=0 $Y2=0
cc_167 N_A_216_93#_c_167_n N_A_331_413#_c_419_n 0.00151483f $X=2.015 $Y=1.89
+ $X2=0 $Y2=0
cc_168 N_A_216_93#_c_168_n N_VPWR_c_514_n 0.00451183f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_169 N_A_216_93#_c_168_n N_VPWR_c_511_n 0.00874597f $X=2.015 $Y=1.99 $X2=0
+ $Y2=0
cc_170 N_A_216_93#_c_165_n N_VGND_M1010_s 2.1368e-19 $X=1.26 $Y=0.66 $X2=0 $Y2=0
cc_171 N_A_216_93#_c_165_n N_VGND_c_587_n 0.0100868f $X=1.26 $Y=0.66 $X2=0 $Y2=0
cc_172 N_A_216_93#_c_165_n N_VGND_c_588_n 0.00922264f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_173 N_A_216_93#_M1010_g N_VGND_c_589_n 0.00334561f $X=2.04 $Y=0.445 $X2=0
+ $Y2=0
cc_174 N_A_216_93#_c_163_n N_VGND_c_589_n 0.0078586f $X=1.97 $Y=1.16 $X2=0 $Y2=0
cc_175 N_A_216_93#_c_164_n N_VGND_c_589_n 0.00197135f $X=1.97 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A_216_93#_c_165_n N_VGND_c_589_n 0.0113822f $X=1.26 $Y=0.66 $X2=0 $Y2=0
cc_177 N_A_216_93#_M1010_g N_VGND_c_590_n 0.00585385f $X=2.04 $Y=0.445 $X2=0
+ $Y2=0
cc_178 N_A_216_93#_M1010_g N_VGND_c_591_n 6.93631e-19 $X=2.04 $Y=0.445 $X2=0
+ $Y2=0
cc_179 N_A_216_93#_M1010_g N_VGND_c_597_n 0.0120495f $X=2.04 $Y=0.445 $X2=0
+ $Y2=0
cc_180 N_A_216_93#_c_165_n N_VGND_c_597_n 0.0126513f $X=1.26 $Y=0.66 $X2=0 $Y2=0
cc_181 N_A_27_410#_M1007_g N_B_c_320_n 0.0128519f $X=2.525 $Y=0.445 $X2=-0.19
+ $Y2=-0.24
cc_182 N_A_27_410#_c_229_n N_B_c_321_n 0.0259242f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_27_410#_c_231_n N_B_c_321_n 3.37553e-19 $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_27_410#_c_231_n N_B_c_323_n 4.70706e-19 $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_27_410#_c_229_n N_B_M1001_g 0.0359634f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_186 N_A_27_410#_c_238_n N_B_M1001_g 7.32223e-19 $X=2.375 $Y=1.5 $X2=0 $Y2=0
cc_187 N_A_27_410#_M1007_g N_B_c_322_n 0.012133f $X=2.525 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_27_410#_c_229_n N_A_c_365_n 0.00252948f $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_27_410#_c_231_n N_A_c_365_n 0.0187646f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_236_n N_A_331_413#_c_410_n 0.0273036f $X=1.845 $Y=1.95
+ $X2=0 $Y2=0
cc_191 N_A_27_410#_c_238_n N_A_331_413#_c_410_n 0.0049489f $X=2.375 $Y=1.5 $X2=0
+ $Y2=0
cc_192 N_A_27_410#_M1007_g N_A_331_413#_c_422_n 0.00511329f $X=2.525 $Y=0.445
+ $X2=0 $Y2=0
cc_193 N_A_27_410#_c_229_n N_A_331_413#_c_411_n 0.00198717f $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_194 N_A_27_410#_c_236_n N_A_331_413#_c_411_n 0.00508372f $X=1.845 $Y=1.95
+ $X2=0 $Y2=0
cc_195 N_A_27_410#_M1007_g N_A_331_413#_c_403_n 0.0127455f $X=2.525 $Y=0.445
+ $X2=0 $Y2=0
cc_196 N_A_27_410#_c_229_n N_A_331_413#_c_403_n 0.00345912f $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_197 N_A_27_410#_c_238_n N_A_331_413#_c_403_n 0.0012205f $X=2.375 $Y=1.5 $X2=0
+ $Y2=0
cc_198 N_A_27_410#_c_231_n N_A_331_413#_c_403_n 0.012923f $X=2.46 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_27_410#_c_229_n N_A_331_413#_c_404_n 2.86694e-19 $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_200 N_A_27_410#_c_238_n N_A_331_413#_c_404_n 0.00589573f $X=2.375 $Y=1.5
+ $X2=0 $Y2=0
cc_201 N_A_27_410#_c_229_n N_A_331_413#_c_412_n 0.0149855f $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_202 N_A_27_410#_c_238_n N_A_331_413#_c_412_n 0.00590782f $X=2.375 $Y=1.5
+ $X2=0 $Y2=0
cc_203 N_A_27_410#_c_229_n N_A_331_413#_c_419_n 2.30045e-19 $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_204 N_A_27_410#_c_236_n N_A_331_413#_c_419_n 0.00640417f $X=1.845 $Y=1.95
+ $X2=0 $Y2=0
cc_205 N_A_27_410#_c_237_n N_A_331_413#_c_419_n 0.0051505f $X=1.93 $Y=1.865
+ $X2=0 $Y2=0
cc_206 N_A_27_410#_c_238_n N_A_331_413#_c_419_n 0.0117409f $X=2.375 $Y=1.5 $X2=0
+ $Y2=0
cc_207 N_A_27_410#_c_238_n N_A_331_413#_c_414_n 0.00240533f $X=2.375 $Y=1.5
+ $X2=0 $Y2=0
cc_208 N_A_27_410#_c_236_n N_VPWR_M1011_d 0.00620921f $X=1.845 $Y=1.95 $X2=-0.19
+ $Y2=-0.24
cc_209 N_A_27_410#_c_235_n N_VPWR_c_512_n 0.0192602f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_210 N_A_27_410#_c_236_n N_VPWR_c_512_n 0.0265965f $X=1.845 $Y=1.95 $X2=0
+ $Y2=0
cc_211 N_A_27_410#_c_229_n N_VPWR_c_514_n 0.00393512f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_27_410#_c_236_n N_VPWR_c_514_n 0.0114405f $X=1.845 $Y=1.95 $X2=0
+ $Y2=0
cc_213 N_A_27_410#_c_235_n N_VPWR_c_516_n 0.0170546f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_214 N_A_27_410#_c_236_n N_VPWR_c_516_n 0.00257955f $X=1.845 $Y=1.95 $X2=0
+ $Y2=0
cc_215 N_A_27_410#_c_229_n N_VPWR_c_511_n 0.00500987f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_27_410#_c_235_n N_VPWR_c_511_n 0.00987599f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_217 N_A_27_410#_c_236_n N_VPWR_c_511_n 0.0253718f $X=1.845 $Y=1.95 $X2=0
+ $Y2=0
cc_218 N_A_27_410#_c_238_n A_421_413# 0.00275594f $X=2.375 $Y=1.5 $X2=-0.19
+ $Y2=-0.24
cc_219 N_A_27_410#_c_232_n N_VGND_c_587_n 0.0185643f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_220 N_A_27_410#_M1007_g N_VGND_c_590_n 0.00199015f $X=2.525 $Y=0.445 $X2=0
+ $Y2=0
cc_221 N_A_27_410#_M1007_g N_VGND_c_591_n 0.0103553f $X=2.525 $Y=0.445 $X2=0
+ $Y2=0
cc_222 N_A_27_410#_c_232_n N_VGND_c_592_n 0.00957361f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_223 N_A_27_410#_M1007_g N_VGND_c_597_n 0.00284206f $X=2.525 $Y=0.445 $X2=0
+ $Y2=0
cc_224 N_A_27_410#_c_232_n N_VGND_c_597_n 0.0105585f $X=0.295 $Y=0.66 $X2=0
+ $Y2=0
cc_225 N_B_c_321_n N_A_c_363_n 0.0206977f $X=2.955 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_226 N_B_c_323_n N_A_c_363_n 0.00417671f $X=2.955 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_227 N_B_M1001_g N_A_c_363_n 0.0247568f $X=2.955 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_228 B N_A_c_363_n 6.06139e-19 $X=3.155 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_229 N_B_c_322_n N_A_M1005_g 0.0196004f $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_230 N_B_c_321_n N_A_c_365_n 0.0123276f $X=2.955 $Y=1.31 $X2=0 $Y2=0
cc_231 N_B_c_323_n N_A_c_365_n 0.0051106f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B_c_324_n N_A_331_413#_c_410_n 9.05269e-19 $X=2.955 $Y=2.035 $X2=0
+ $Y2=0
cc_233 B N_A_331_413#_c_410_n 0.0113771f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_234 N_B_c_324_n N_A_331_413#_c_411_n 0.00275377f $X=2.955 $Y=2.035 $X2=0
+ $Y2=0
cc_235 B N_A_331_413#_c_411_n 0.00474738f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_236 N_B_c_320_n N_A_331_413#_c_403_n 0.00630115f $X=2.955 $Y=0.86 $X2=0 $Y2=0
cc_237 N_B_c_322_n N_A_331_413#_c_403_n 0.00765134f $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_238 N_B_c_324_n N_A_331_413#_c_412_n 6.90064e-19 $X=2.955 $Y=2.035 $X2=0
+ $Y2=0
cc_239 N_B_M1001_g N_A_331_413#_c_412_n 0.0125693f $X=2.955 $Y=1.695 $X2=0 $Y2=0
cc_240 B N_A_331_413#_c_412_n 0.0385065f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_241 N_B_M1001_g N_A_331_413#_c_414_n 0.00550607f $X=2.955 $Y=1.695 $X2=0
+ $Y2=0
cc_242 B N_A_331_413#_c_414_n 0.0138656f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_243 N_B_c_324_n N_VPWR_c_513_n 0.00478317f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_244 B N_VPWR_c_513_n 0.0239486f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_245 N_B_c_324_n N_VPWR_c_514_n 0.0050964f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_246 B N_VPWR_c_514_n 0.0429955f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_247 N_B_c_324_n N_VPWR_c_511_n 0.00694793f $X=2.955 $Y=2.035 $X2=0 $Y2=0
cc_248 B N_VPWR_c_511_n 0.0247011f $X=3.155 $Y=2.125 $X2=0 $Y2=0
cc_249 N_B_c_322_n N_VGND_c_591_n 0.00167196f $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_250 N_B_c_322_n N_VGND_c_594_n 6.85223e-19 $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_251 N_B_c_322_n N_VGND_c_595_n 0.00428022f $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_252 N_B_c_322_n N_VGND_c_597_n 0.00594333f $X=2.955 $Y=0.76 $X2=0 $Y2=0
cc_253 N_A_c_363_n N_A_331_413#_c_401_n 0.0337925f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_365_n N_A_331_413#_c_401_n 0.0011063f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_255 N_A_M1005_g N_A_331_413#_c_402_n 0.0180817f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_256 N_A_c_365_n N_A_331_413#_c_403_n 0.0225698f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_c_365_n N_A_331_413#_c_412_n 0.0116453f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A_c_363_n N_A_331_413#_c_405_n 0.00240831f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_M1005_g N_A_331_413#_c_405_n 0.0117067f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_c_365_n N_A_331_413#_c_405_n 0.0205685f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_261 N_A_c_363_n N_A_331_413#_c_457_n 0.0141289f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_365_n N_A_331_413#_c_457_n 0.0130503f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_263 N_A_c_363_n N_A_331_413#_c_413_n 0.00173315f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_363_n N_A_331_413#_c_406_n 4.61771e-19 $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_365_n N_A_331_413#_c_406_n 0.0146461f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_c_363_n N_A_331_413#_c_414_n 0.0109312f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_c_365_n N_A_331_413#_c_414_n 0.0112678f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_c_363_n N_A_331_413#_c_407_n 0.00458419f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_365_n N_A_331_413#_c_407_n 0.0287412f $X=3.405 $Y=1.16 $X2=0 $Y2=0
cc_270 N_A_M1005_g N_A_331_413#_c_408_n 0.00177765f $X=3.465 $Y=0.445 $X2=0
+ $Y2=0
cc_271 N_A_c_363_n N_VPWR_c_513_n 0.00330158f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_c_363_n N_VPWR_c_514_n 0.00351015f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_c_363_n N_VPWR_c_511_n 0.00445321f $X=3.44 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_M1005_g N_VGND_c_594_n 0.0105644f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_M1005_g N_VGND_c_595_n 0.00199743f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_276 N_A_M1005_g N_VGND_c_597_n 0.00284206f $X=3.465 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A_331_413#_c_457_n N_VPWR_M1008_d 0.00563715f $X=3.74 $Y=1.58 $X2=0
+ $Y2=0
cc_278 N_A_331_413#_c_401_n N_VPWR_c_513_n 0.00499543f $X=3.98 $Y=1.41 $X2=0
+ $Y2=0
cc_279 N_A_331_413#_c_457_n N_VPWR_c_513_n 0.0204259f $X=3.74 $Y=1.58 $X2=0
+ $Y2=0
cc_280 N_A_331_413#_c_414_n N_VPWR_c_513_n 0.00726621f $X=3.285 $Y=1.58 $X2=0
+ $Y2=0
cc_281 N_A_331_413#_c_410_n N_VPWR_c_514_n 0.0304719f $X=2.235 $Y=2.29 $X2=0
+ $Y2=0
cc_282 N_A_331_413#_c_401_n N_VPWR_c_517_n 0.00702461f $X=3.98 $Y=1.41 $X2=0
+ $Y2=0
cc_283 N_A_331_413#_M1002_s N_VPWR_c_511_n 0.002265f $X=1.655 $Y=2.065 $X2=0
+ $Y2=0
cc_284 N_A_331_413#_c_401_n N_VPWR_c_511_n 0.0148168f $X=3.98 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_331_413#_c_410_n N_VPWR_c_511_n 0.027257f $X=2.235 $Y=2.29 $X2=0
+ $Y2=0
cc_286 N_A_331_413#_c_412_n N_VPWR_c_511_n 0.0102114f $X=3.2 $Y=1.87 $X2=0 $Y2=0
cc_287 N_A_331_413#_c_410_n A_421_413# 0.0046523f $X=2.235 $Y=2.29 $X2=-0.19
+ $Y2=-0.24
cc_288 N_A_331_413#_c_411_n A_421_413# 0.00311349f $X=2.32 $Y=2.205 $X2=-0.19
+ $Y2=-0.24
cc_289 N_A_331_413#_c_419_n A_421_413# 0.00379949f $X=2.405 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_290 N_A_331_413#_c_412_n A_527_297# 0.00442604f $X=3.2 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_291 N_A_331_413#_c_412_n A_609_297# 0.00197899f $X=3.2 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_292 N_A_331_413#_c_414_n A_609_297# 0.00483332f $X=3.285 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_293 N_A_331_413#_c_401_n N_X_c_571_n 0.0122499f $X=3.98 $Y=1.41 $X2=0 $Y2=0
cc_294 N_A_331_413#_c_457_n N_X_c_571_n 0.0112291f $X=3.74 $Y=1.58 $X2=0 $Y2=0
cc_295 N_A_331_413#_c_401_n N_X_c_570_n 7.49618e-19 $X=3.98 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_331_413#_c_402_n N_X_c_570_n 0.0132989f $X=4.005 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_331_413#_c_413_n N_X_c_570_n 0.005373f $X=3.825 $Y=1.495 $X2=0 $Y2=0
cc_298 N_A_331_413#_c_407_n N_X_c_570_n 0.0217737f $X=3.945 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_331_413#_c_408_n N_X_c_570_n 0.00673639f $X=3.885 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A_331_413#_c_405_n N_VGND_M1005_d 0.00652347f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_301 N_A_331_413#_c_408_n N_VGND_M1005_d 6.98847e-19 $X=3.885 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_331_413#_c_422_n N_VGND_c_590_n 0.00861358f $X=2.25 $Y=0.47 $X2=0
+ $Y2=0
cc_303 N_A_331_413#_c_403_n N_VGND_c_590_n 0.00309172f $X=3.12 $Y=0.74 $X2=0
+ $Y2=0
cc_304 N_A_331_413#_c_422_n N_VGND_c_591_n 0.0125877f $X=2.25 $Y=0.47 $X2=0
+ $Y2=0
cc_305 N_A_331_413#_c_403_n N_VGND_c_591_n 0.0242276f $X=3.12 $Y=0.74 $X2=0
+ $Y2=0
cc_306 N_A_331_413#_c_401_n N_VGND_c_594_n 2.73815e-19 $X=3.98 $Y=1.41 $X2=0
+ $Y2=0
cc_307 N_A_331_413#_c_402_n N_VGND_c_594_n 0.00463088f $X=4.005 $Y=0.995 $X2=0
+ $Y2=0
cc_308 N_A_331_413#_c_498_p N_VGND_c_594_n 0.0135697f $X=3.205 $Y=0.47 $X2=0
+ $Y2=0
cc_309 N_A_331_413#_c_405_n N_VGND_c_594_n 0.0298327f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_310 N_A_331_413#_c_403_n N_VGND_c_595_n 0.0035533f $X=3.12 $Y=0.74 $X2=0
+ $Y2=0
cc_311 N_A_331_413#_c_498_p N_VGND_c_595_n 0.00876148f $X=3.205 $Y=0.47 $X2=0
+ $Y2=0
cc_312 N_A_331_413#_c_405_n N_VGND_c_595_n 0.00283814f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_313 N_A_331_413#_c_402_n N_VGND_c_596_n 0.00585385f $X=4.005 $Y=0.995 $X2=0
+ $Y2=0
cc_314 N_A_331_413#_M1010_d N_VGND_c_597_n 0.00494728f $X=2.115 $Y=0.235 $X2=0
+ $Y2=0
cc_315 N_A_331_413#_M1004_d N_VGND_c_597_n 0.00336566f $X=3.055 $Y=0.235 $X2=0
+ $Y2=0
cc_316 N_A_331_413#_c_402_n N_VGND_c_597_n 0.0120637f $X=4.005 $Y=0.995 $X2=0
+ $Y2=0
cc_317 N_A_331_413#_c_422_n N_VGND_c_597_n 0.00625722f $X=2.25 $Y=0.47 $X2=0
+ $Y2=0
cc_318 N_A_331_413#_c_403_n N_VGND_c_597_n 0.0117669f $X=3.12 $Y=0.74 $X2=0
+ $Y2=0
cc_319 N_A_331_413#_c_498_p N_VGND_c_597_n 0.00625722f $X=3.205 $Y=0.47 $X2=0
+ $Y2=0
cc_320 N_A_331_413#_c_405_n N_VGND_c_597_n 0.00690419f $X=3.74 $Y=0.74 $X2=0
+ $Y2=0
cc_321 N_VPWR_c_511_n A_421_413# 0.00222986f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_322 N_VPWR_c_511_n N_X_M1000_d 0.00442383f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_323 N_VPWR_c_517_n X 0.0228497f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_324 N_VPWR_c_511_n X 0.0124393f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_325 N_X_c_569_n N_VGND_c_596_n 0.0109423f $X=4.215 $Y=0.59 $X2=0 $Y2=0
cc_326 N_X_M1009_d N_VGND_c_597_n 0.00419212f $X=4.08 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_c_569_n N_VGND_c_597_n 0.0112582f $X=4.215 $Y=0.59 $X2=0 $Y2=0
