* File: sky130_fd_sc_hdll__einvn_4.pxi.spice
* Created: Thu Aug 27 19:07:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__EINVN_4%TE_B N_TE_B_c_84_n N_TE_B_M1016_g N_TE_B_c_89_n
+ N_TE_B_M1006_g N_TE_B_c_85_n N_TE_B_c_86_n N_TE_B_c_92_n N_TE_B_M1000_g
+ N_TE_B_c_93_n N_TE_B_c_94_n N_TE_B_M1003_g N_TE_B_c_95_n N_TE_B_c_96_n
+ N_TE_B_M1014_g N_TE_B_c_97_n N_TE_B_c_98_n N_TE_B_M1015_g N_TE_B_c_87_n
+ N_TE_B_c_100_n N_TE_B_c_101_n TE_B PM_SKY130_FD_SC_HDLL__EINVN_4%TE_B
x_PM_SKY130_FD_SC_HDLL__EINVN_4%A_27_47# N_A_27_47#_M1016_s N_A_27_47#_M1006_s
+ N_A_27_47#_c_164_n N_A_27_47#_M1004_g N_A_27_47#_c_165_n N_A_27_47#_c_166_n
+ N_A_27_47#_c_167_n N_A_27_47#_M1005_g N_A_27_47#_c_168_n N_A_27_47#_c_169_n
+ N_A_27_47#_M1008_g N_A_27_47#_c_170_n N_A_27_47#_c_171_n N_A_27_47#_M1013_g
+ N_A_27_47#_c_172_n N_A_27_47#_c_173_n N_A_27_47#_c_174_n N_A_27_47#_c_175_n
+ N_A_27_47#_c_179_n N_A_27_47#_c_176_n N_A_27_47#_c_177_n
+ PM_SKY130_FD_SC_HDLL__EINVN_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__EINVN_4%A N_A_c_261_n N_A_M1001_g N_A_c_267_n
+ N_A_M1007_g N_A_c_262_n N_A_M1002_g N_A_c_268_n N_A_M1011_g N_A_c_263_n
+ N_A_M1009_g N_A_c_269_n N_A_M1012_g N_A_c_264_n N_A_M1010_g N_A_c_270_n
+ N_A_M1017_g A A N_A_c_266_n PM_SKY130_FD_SC_HDLL__EINVN_4%A
x_PM_SKY130_FD_SC_HDLL__EINVN_4%VPWR N_VPWR_M1006_d N_VPWR_M1003_d
+ N_VPWR_M1015_d N_VPWR_c_329_n N_VPWR_c_330_n N_VPWR_c_331_n N_VPWR_c_332_n
+ VPWR N_VPWR_c_333_n N_VPWR_c_334_n N_VPWR_c_335_n N_VPWR_c_328_n
+ N_VPWR_c_337_n N_VPWR_c_338_n N_VPWR_c_339_n
+ PM_SKY130_FD_SC_HDLL__EINVN_4%VPWR
x_PM_SKY130_FD_SC_HDLL__EINVN_4%A_222_309# N_A_222_309#_M1000_s
+ N_A_222_309#_M1014_s N_A_222_309#_M1007_d N_A_222_309#_M1011_d
+ N_A_222_309#_M1017_d N_A_222_309#_c_407_n N_A_222_309#_c_402_n
+ N_A_222_309#_c_403_n N_A_222_309#_c_415_n N_A_222_309#_c_404_n
+ N_A_222_309#_c_419_n N_A_222_309#_c_431_n N_A_222_309#_c_405_n
+ N_A_222_309#_c_433_n N_A_222_309#_c_434_n N_A_222_309#_c_436_n
+ N_A_222_309#_c_406_n N_A_222_309#_c_462_n
+ PM_SKY130_FD_SC_HDLL__EINVN_4%A_222_309#
x_PM_SKY130_FD_SC_HDLL__EINVN_4%Z N_Z_M1001_s N_Z_M1009_s N_Z_M1007_s
+ N_Z_M1012_s N_Z_c_474_n N_Z_c_475_n Z Z Z Z N_Z_c_476_n
+ PM_SKY130_FD_SC_HDLL__EINVN_4%Z
x_PM_SKY130_FD_SC_HDLL__EINVN_4%VGND N_VGND_M1016_d N_VGND_M1004_s
+ N_VGND_M1008_s N_VGND_c_518_n N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n
+ N_VGND_c_522_n N_VGND_c_523_n VGND N_VGND_c_524_n N_VGND_c_525_n
+ N_VGND_c_526_n N_VGND_c_527_n N_VGND_c_528_n
+ PM_SKY130_FD_SC_HDLL__EINVN_4%VGND
x_PM_SKY130_FD_SC_HDLL__EINVN_4%A_235_47# N_A_235_47#_M1004_d
+ N_A_235_47#_M1005_d N_A_235_47#_M1013_d N_A_235_47#_M1002_d
+ N_A_235_47#_M1010_d N_A_235_47#_c_592_n N_A_235_47#_c_599_n
+ N_A_235_47#_c_593_n N_A_235_47#_c_605_n N_A_235_47#_c_606_n
+ N_A_235_47#_c_611_n N_A_235_47#_c_612_n N_A_235_47#_c_594_n
+ N_A_235_47#_c_614_n PM_SKY130_FD_SC_HDLL__EINVN_4%A_235_47#
cc_1 VNB N_TE_B_c_84_n 0.0250205f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_TE_B_c_85_n 0.0136496f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_3 VNB N_TE_B_c_86_n 0.0383463f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.25
cc_4 VNB N_TE_B_c_87_n 0.0121778f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.25
cc_5 VNB TE_B 0.0136088f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_6 VNB N_A_27_47#_c_164_n 0.018254f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_7 VNB N_A_27_47#_c_165_n 0.0113615f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=2.015
cc_8 VNB N_A_27_47#_c_166_n 0.00835566f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=2.015
cc_9 VNB N_A_27_47#_c_167_n 0.01485f $X=-0.19 $Y=-0.24 $X2=1.4 $Y2=1.395
cc_10 VNB N_A_27_47#_c_168_n 0.0113601f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_11 VNB N_A_27_47#_c_169_n 0.0150799f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=1.395
cc_12 VNB N_A_27_47#_c_170_n 0.0120821f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=2.015
cc_13 VNB N_A_27_47#_c_171_n 0.0153973f $X=-0.19 $Y=-0.24 $X2=2.34 $Y2=1.395
cc_14 VNB N_A_27_47#_c_172_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_15 VNB N_A_27_47#_c_173_n 0.00391059f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_16 VNB N_A_27_47#_c_174_n 0.0155207f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.25
cc_17 VNB N_A_27_47#_c_175_n 0.0127587f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=1.395
cc_18 VNB N_A_27_47#_c_176_n 0.0149189f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_19 VNB N_A_27_47#_c_177_n 0.0242871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_c_261_n 0.0171736f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_21 VNB N_A_c_262_n 0.0160107f $X=-0.19 $Y=-0.24 $X2=0.92 $Y2=1.25
cc_22 VNB N_A_c_263_n 0.0160107f $X=-0.19 $Y=-0.24 $X2=1.12 $Y2=1.395
cc_23 VNB N_A_c_264_n 0.0191728f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=1.47
cc_24 VNB A 0.0294497f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_25 VNB N_A_c_266_n 0.100357f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_26 VNB N_VPWR_c_328_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_518_n 0.00575291f $X=-0.19 $Y=-0.24 $X2=1.4 $Y2=1.395
cc_28 VNB N_VGND_c_519_n 0.0185905f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=1.47
cc_29 VNB N_VGND_c_520_n 0.00272748f $X=-0.19 $Y=-0.24 $X2=1.58 $Y2=1.395
cc_30 VNB N_VGND_c_521_n 0.00220692f $X=-0.19 $Y=-0.24 $X2=2.34 $Y2=1.395
cc_31 VNB N_VGND_c_522_n 0.0148248f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_32 VNB N_VGND_c_523_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=2.43 $Y2=2.015
cc_33 VNB N_VGND_c_524_n 0.0143218f $X=-0.19 $Y=-0.24 $X2=1.02 $Y2=1.395
cc_34 VNB N_VGND_c_525_n 0.0619423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_526_n 0.284775f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_527_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_528_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_235_47#_c_592_n 0.00646793f $X=-0.19 $Y=-0.24 $X2=1.49 $Y2=2.015
cc_39 VNB N_A_235_47#_c_593_n 0.00271074f $X=-0.19 $Y=-0.24 $X2=1.96 $Y2=2.015
cc_40 VNB N_A_235_47#_c_594_n 0.0124706f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.202
cc_41 VPB N_TE_B_c_89_n 0.0207069f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_TE_B_c_85_n 0.0103502f $X=-0.19 $Y=1.305 $X2=0.92 $Y2=1.25
cc_43 VPB N_TE_B_c_86_n 0.017266f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.25
cc_44 VPB N_TE_B_c_92_n 0.0164357f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.47
cc_45 VPB N_TE_B_c_93_n 0.0146992f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_46 VPB N_TE_B_c_94_n 0.0153558f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.47
cc_47 VPB N_TE_B_c_95_n 0.00980191f $X=-0.19 $Y=1.305 $X2=1.87 $Y2=1.395
cc_48 VPB N_TE_B_c_96_n 0.0156362f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.47
cc_49 VPB N_TE_B_c_97_n 0.0229817f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_50 VPB N_TE_B_c_98_n 0.0187512f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=1.47
cc_51 VPB N_TE_B_c_87_n 0.00718766f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=1.25
cc_52 VPB N_TE_B_c_100_n 0.00533627f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.395
cc_53 VPB N_TE_B_c_101_n 0.0046927f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.395
cc_54 VPB TE_B 0.00311217f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_55 VPB N_A_27_47#_c_175_n 0.00967156f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=1.395
cc_56 VPB N_A_27_47#_c_179_n 0.0307249f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_57 VPB N_A_27_47#_c_176_n 0.00452491f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_58 VPB N_A_27_47#_c_177_n 0.0096023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_c_267_n 0.0206889f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_A_c_268_n 0.0155675f $X=-0.19 $Y=1.305 $X2=1.02 $Y2=2.015
cc_61 VPB N_A_c_269_n 0.0155623f $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_62 VPB N_A_c_270_n 0.0206942f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_63 VPB A 0.013648f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=2.015
cc_64 VPB N_A_c_266_n 0.061513f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_65 VPB N_VPWR_c_329_n 0.00222504f $X=-0.19 $Y=1.305 $X2=1.4 $Y2=1.395
cc_66 VPB N_VPWR_c_330_n 3.28479e-19 $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_67 VPB N_VPWR_c_331_n 0.0140826f $X=-0.19 $Y=1.305 $X2=1.58 $Y2=1.395
cc_68 VPB N_VPWR_c_332_n 0.0114603f $X=-0.19 $Y=1.305 $X2=2.34 $Y2=1.395
cc_69 VPB N_VPWR_c_333_n 0.0150576f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=2.015
cc_70 VPB N_VPWR_c_334_n 0.0157606f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.395
cc_71 VPB N_VPWR_c_335_n 0.0656244f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_328_n 0.0606258f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_337_n 0.00580052f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_338_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_339_n 0.00695794f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_222_309#_c_402_n 0.00278842f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=2.015
cc_77 VPB N_A_222_309#_c_403_n 0.00177529f $X=-0.19 $Y=1.305 $X2=1.96 $Y2=2.015
cc_78 VPB N_A_222_309#_c_404_n 0.0147346f $X=-0.19 $Y=1.305 $X2=2.43 $Y2=2.015
cc_79 VPB N_A_222_309#_c_405_n 0.00141314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_222_309#_c_406_n 0.00106199f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_Z_c_474_n 5.57362e-19 $X=-0.19 $Y=1.305 $X2=1.49 $Y2=2.015
cc_82 VPB N_Z_c_475_n 5.57362e-19 $X=-0.19 $Y=1.305 $X2=1.96 $Y2=1.47
cc_83 VPB N_Z_c_476_n 0.00820234f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 N_TE_B_c_95_n N_A_27_47#_c_165_n 0.0177654f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_85 N_TE_B_c_100_n N_A_27_47#_c_166_n 0.0177654f $X=1.49 $Y=1.395 $X2=0 $Y2=0
cc_86 N_TE_B_c_101_n N_A_27_47#_c_168_n 0.0177654f $X=1.96 $Y=1.395 $X2=0 $Y2=0
cc_87 N_TE_B_c_97_n N_A_27_47#_c_173_n 0.0177654f $X=2.34 $Y=1.395 $X2=0 $Y2=0
cc_88 N_TE_B_c_84_n N_A_27_47#_c_175_n 0.022924f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_89 N_TE_B_c_89_n N_A_27_47#_c_175_n 0.0193828f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_TE_B_c_85_n N_A_27_47#_c_175_n 0.0171587f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_91 N_TE_B_c_86_n N_A_27_47#_c_175_n 0.0220923f $X=0.595 $Y=1.25 $X2=0 $Y2=0
cc_92 N_TE_B_c_92_n N_A_27_47#_c_175_n 0.00196252f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_93 N_TE_B_c_87_n N_A_27_47#_c_175_n 0.00472039f $X=1.02 $Y=1.25 $X2=0 $Y2=0
cc_94 TE_B N_A_27_47#_c_175_n 0.0685238f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_95 N_TE_B_c_89_n N_A_27_47#_c_179_n 0.00783737f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_96 N_TE_B_c_85_n N_A_27_47#_c_176_n 0.00164242f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_97 N_TE_B_c_93_n N_A_27_47#_c_176_n 0.00914812f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_98 N_TE_B_c_95_n N_A_27_47#_c_176_n 0.00618718f $X=1.87 $Y=1.395 $X2=0 $Y2=0
cc_99 N_TE_B_c_97_n N_A_27_47#_c_176_n 0.010621f $X=2.34 $Y=1.395 $X2=0 $Y2=0
cc_100 N_TE_B_c_87_n N_A_27_47#_c_176_n 0.0176781f $X=1.02 $Y=1.25 $X2=0 $Y2=0
cc_101 N_TE_B_c_100_n N_A_27_47#_c_176_n 0.00465183f $X=1.49 $Y=1.395 $X2=0
+ $Y2=0
cc_102 N_TE_B_c_101_n N_A_27_47#_c_176_n 0.00425603f $X=1.96 $Y=1.395 $X2=0
+ $Y2=0
cc_103 N_TE_B_c_97_n N_A_27_47#_c_177_n 3.39336e-19 $X=2.34 $Y=1.395 $X2=0 $Y2=0
cc_104 N_TE_B_c_89_n N_VPWR_c_329_n 0.0170835f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_105 N_TE_B_c_85_n N_VPWR_c_329_n 0.00105584f $X=0.92 $Y=1.25 $X2=0 $Y2=0
cc_106 N_TE_B_c_92_n N_VPWR_c_329_n 0.00524796f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_107 N_TE_B_c_92_n N_VPWR_c_330_n 7.75802e-19 $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_108 N_TE_B_c_94_n N_VPWR_c_330_n 0.0154334f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_109 N_TE_B_c_96_n N_VPWR_c_330_n 0.0117009f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_110 N_TE_B_c_98_n N_VPWR_c_330_n 6.61031e-19 $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_111 N_TE_B_c_96_n N_VPWR_c_331_n 0.00622633f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_112 N_TE_B_c_98_n N_VPWR_c_331_n 0.00427505f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_113 N_TE_B_c_96_n N_VPWR_c_332_n 7.02381e-19 $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_114 N_TE_B_c_98_n N_VPWR_c_332_n 0.0164441f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_115 N_TE_B_c_89_n N_VPWR_c_333_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_116 N_TE_B_c_92_n N_VPWR_c_334_n 0.00635665f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_117 N_TE_B_c_94_n N_VPWR_c_334_n 0.00427505f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_118 N_TE_B_c_89_n N_VPWR_c_328_n 0.00835414f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_119 N_TE_B_c_92_n N_VPWR_c_328_n 0.0111139f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_120 N_TE_B_c_94_n N_VPWR_c_328_n 0.00740765f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_121 N_TE_B_c_96_n N_VPWR_c_328_n 0.010479f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_122 N_TE_B_c_98_n N_VPWR_c_328_n 0.00740765f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_123 N_TE_B_c_89_n N_A_222_309#_c_407_n 7.83445e-19 $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_TE_B_c_92_n N_A_222_309#_c_407_n 0.0127872f $X=1.02 $Y=1.47 $X2=0 $Y2=0
cc_125 N_TE_B_c_94_n N_A_222_309#_c_407_n 0.00614066f $X=1.49 $Y=1.47 $X2=0
+ $Y2=0
cc_126 N_TE_B_c_94_n N_A_222_309#_c_402_n 0.014571f $X=1.49 $Y=1.47 $X2=0 $Y2=0
cc_127 N_TE_B_c_95_n N_A_222_309#_c_402_n 0.00250384f $X=1.87 $Y=1.395 $X2=0
+ $Y2=0
cc_128 N_TE_B_c_96_n N_A_222_309#_c_402_n 0.0160672f $X=1.96 $Y=1.47 $X2=0 $Y2=0
cc_129 N_TE_B_c_92_n N_A_222_309#_c_403_n 0.00430535f $X=1.02 $Y=1.47 $X2=0
+ $Y2=0
cc_130 N_TE_B_c_93_n N_A_222_309#_c_403_n 0.0026331f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_131 N_TE_B_c_96_n N_A_222_309#_c_415_n 0.00600706f $X=1.96 $Y=1.47 $X2=0
+ $Y2=0
cc_132 N_TE_B_c_98_n N_A_222_309#_c_415_n 0.00555086f $X=2.43 $Y=1.47 $X2=0
+ $Y2=0
cc_133 N_TE_B_c_97_n N_A_222_309#_c_404_n 2.27622e-19 $X=2.34 $Y=1.395 $X2=0
+ $Y2=0
cc_134 N_TE_B_c_98_n N_A_222_309#_c_404_n 0.0165379f $X=2.43 $Y=1.47 $X2=0 $Y2=0
cc_135 N_TE_B_c_98_n N_A_222_309#_c_419_n 0.00358253f $X=2.43 $Y=1.47 $X2=0
+ $Y2=0
cc_136 N_TE_B_c_97_n N_A_222_309#_c_406_n 0.0026331f $X=2.34 $Y=1.395 $X2=0
+ $Y2=0
cc_137 N_TE_B_c_84_n N_VGND_c_518_n 0.00977312f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_138 N_TE_B_c_86_n N_VGND_c_518_n 9.2603e-19 $X=0.595 $Y=1.25 $X2=0 $Y2=0
cc_139 N_TE_B_c_84_n N_VGND_c_524_n 0.00341574f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_140 N_TE_B_c_84_n N_VGND_c_526_n 0.00501514f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_141 N_TE_B_c_84_n N_A_235_47#_c_592_n 0.00328724f $X=0.47 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_TE_B_c_84_n N_A_235_47#_c_593_n 6.5289e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_143 N_TE_B_c_93_n N_A_235_47#_c_593_n 0.00101478f $X=1.4 $Y=1.395 $X2=0 $Y2=0
cc_144 N_TE_B_c_87_n N_A_235_47#_c_593_n 2.76908e-19 $X=1.02 $Y=1.25 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_171_n N_A_c_261_n 0.0209158f $X=2.92 $Y=0.96 $X2=-0.19
+ $Y2=-0.24
cc_146 N_A_27_47#_c_176_n N_A_c_266_n 0.00345774f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_177_n N_A_c_266_n 0.0129241f $X=2.9 $Y=1.035 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_175_n N_VPWR_M1006_d 0.00340372f $X=0.215 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_149 N_A_27_47#_c_175_n N_VPWR_c_329_n 0.0266259f $X=0.215 $Y=1.665 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_c_179_n N_VPWR_c_329_n 0.0485357f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_179_n N_VPWR_c_333_n 0.0182101f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_152 N_A_27_47#_M1006_s N_VPWR_c_328_n 0.00430086f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_179_n N_VPWR_c_328_n 0.00993603f $X=0.26 $Y=1.815 $X2=0
+ $Y2=0
cc_154 N_A_27_47#_c_166_n N_A_222_309#_c_402_n 4.62261e-19 $X=1.585 $Y=1.035
+ $X2=0 $Y2=0
cc_155 N_A_27_47#_c_176_n N_A_222_309#_c_402_n 0.0563004f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_27_47#_c_175_n N_A_222_309#_c_403_n 0.00948929f $X=0.215 $Y=1.665
+ $X2=0 $Y2=0
cc_157 N_A_27_47#_c_176_n N_A_222_309#_c_403_n 0.0229519f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_27_47#_c_168_n N_A_222_309#_c_404_n 2.25389e-19 $X=2.375 $Y=1.035
+ $X2=0 $Y2=0
cc_159 N_A_27_47#_c_173_n N_A_222_309#_c_404_n 9.0257e-19 $X=2.45 $Y=1.035 $X2=0
+ $Y2=0
cc_160 N_A_27_47#_c_176_n N_A_222_309#_c_404_n 0.080872f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_161 N_A_27_47#_c_177_n N_A_222_309#_c_404_n 0.00812721f $X=2.9 $Y=1.035 $X2=0
+ $Y2=0
cc_162 N_A_27_47#_c_176_n N_A_222_309#_c_406_n 0.0143361f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_27_47#_c_171_n N_Z_c_476_n 9.60687e-19 $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_176_n N_Z_c_476_n 0.0292385f $X=2.875 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_177_n N_Z_c_476_n 2.33831e-19 $X=2.9 $Y=1.035 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_175_n N_VGND_M1016_d 0.00435803f $X=0.215 $Y=1.665 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_27_47#_c_164_n N_VGND_c_518_n 0.00270009f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_175_n N_VGND_c_518_n 0.0271576f $X=0.215 $Y=1.665 $X2=0
+ $Y2=0
cc_169 N_A_27_47#_c_164_n N_VGND_c_519_n 0.00428022f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_164_n N_VGND_c_520_n 0.00312892f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_167_n N_VGND_c_520_n 0.00733819f $X=1.98 $Y=0.96 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_169_n N_VGND_c_520_n 5.76807e-19 $X=2.45 $Y=0.96 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_169_n N_VGND_c_521_n 0.00167984f $X=2.45 $Y=0.96 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_171_n N_VGND_c_521_n 0.00849499f $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_167_n N_VGND_c_522_n 0.00341689f $X=1.98 $Y=0.96 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_169_n N_VGND_c_522_n 0.00428022f $X=2.45 $Y=0.96 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_174_n N_VGND_c_524_n 0.0177719f $X=0.215 $Y=0.655 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_175_n N_VGND_c_524_n 0.00233078f $X=0.215 $Y=1.665 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_171_n N_VGND_c_525_n 0.00341689f $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_180 N_A_27_47#_M1016_s N_VGND_c_526_n 0.00228937f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_164_n N_VGND_c_526_n 0.00718822f $X=1.51 $Y=0.96 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_167_n N_VGND_c_526_n 0.00415805f $X=1.98 $Y=0.96 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_169_n N_VGND_c_526_n 0.005943f $X=2.45 $Y=0.96 $X2=0 $Y2=0
cc_184 N_A_27_47#_c_171_n N_VGND_c_526_n 0.00429997f $X=2.92 $Y=0.96 $X2=0 $Y2=0
cc_185 N_A_27_47#_c_174_n N_VGND_c_526_n 0.00989054f $X=0.215 $Y=0.655 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_175_n N_VGND_c_526_n 0.00599845f $X=0.215 $Y=1.665 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_164_n N_A_235_47#_c_599_n 0.0115119f $X=1.51 $Y=0.96 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_165_n N_A_235_47#_c_599_n 0.00278658f $X=1.905 $Y=1.035
+ $X2=0 $Y2=0
cc_189 N_A_27_47#_c_167_n N_A_235_47#_c_599_n 0.0106628f $X=1.98 $Y=0.96 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_176_n N_A_235_47#_c_599_n 0.0481586f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_175_n N_A_235_47#_c_593_n 0.0159284f $X=0.215 $Y=1.665 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_176_n N_A_235_47#_c_593_n 0.0272529f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_167_n N_A_235_47#_c_605_n 0.00437226f $X=1.98 $Y=0.96 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_169_n N_A_235_47#_c_606_n 0.0109748f $X=2.45 $Y=0.96 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_170_n N_A_235_47#_c_606_n 0.00282823f $X=2.74 $Y=1.035 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_171_n N_A_235_47#_c_606_n 0.0119624f $X=2.92 $Y=0.96 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_176_n N_A_235_47#_c_606_n 0.0649758f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_177_n N_A_235_47#_c_606_n 0.00133229f $X=2.9 $Y=1.035 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_171_n N_A_235_47#_c_611_n 0.00413107f $X=2.92 $Y=0.96 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_171_n N_A_235_47#_c_612_n 0.00182697f $X=2.92 $Y=0.96 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_176_n N_A_235_47#_c_594_n 7.29254e-19 $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_168_n N_A_235_47#_c_614_n 0.00268716f $X=2.375 $Y=1.035
+ $X2=0 $Y2=0
cc_203 N_A_27_47#_c_176_n N_A_235_47#_c_614_n 0.0135367f $X=2.875 $Y=1.16 $X2=0
+ $Y2=0
cc_204 N_A_c_267_n N_VPWR_c_332_n 0.00326066f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_267_n N_VPWR_c_335_n 0.00429453f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_268_n N_VPWR_c_335_n 0.00429453f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_c_269_n N_VPWR_c_335_n 0.00429453f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_270_n N_VPWR_c_335_n 0.00429453f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_c_267_n N_VPWR_c_328_n 0.00743756f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_268_n N_VPWR_c_328_n 0.00610589f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_c_269_n N_VPWR_c_328_n 0.00610589f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_c_270_n N_VPWR_c_328_n 0.00716615f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_c_267_n N_A_222_309#_c_404_n 0.00313438f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_c_267_n N_A_222_309#_c_431_n 0.0145999f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_268_n N_A_222_309#_c_431_n 0.0152369f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_266_n N_A_222_309#_c_433_n 9.17414e-19 $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A_c_269_n N_A_222_309#_c_434_n 0.0137645f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_270_n N_A_222_309#_c_434_n 0.0159498f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_219 A N_A_222_309#_c_436_n 0.0089194f $X=5.195 $Y=0.765 $X2=0 $Y2=0
cc_220 N_A_c_266_n N_A_222_309#_c_436_n 0.00122612f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_221 N_A_c_267_n N_Z_c_474_n 0.010453f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_268_n N_Z_c_474_n 0.00844867f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_269_n N_Z_c_474_n 5.60154e-19 $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_266_n N_Z_c_474_n 0.00153779f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_225 N_A_c_268_n N_Z_c_475_n 5.90635e-19 $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_269_n N_Z_c_475_n 0.0109729f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_c_270_n N_Z_c_475_n 0.0130795f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_266_n N_Z_c_475_n 0.00153779f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_229 N_A_c_261_n N_Z_c_476_n 0.00779807f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_230 N_A_c_267_n N_Z_c_476_n 0.00453579f $X=3.47 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_c_262_n N_Z_c_476_n 0.013797f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_268_n N_Z_c_476_n 0.0112444f $X=3.94 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_c_263_n N_Z_c_476_n 0.013797f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_c_269_n N_Z_c_476_n 0.0088063f $X=4.41 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_264_n N_Z_c_476_n 0.00598378f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_c_270_n N_Z_c_476_n 0.00410424f $X=4.88 $Y=1.41 $X2=0 $Y2=0
cc_237 A N_Z_c_476_n 0.0473397f $X=5.195 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A_c_266_n N_Z_c_476_n 0.0900036f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A_c_261_n N_VGND_c_521_n 0.00111107f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_c_261_n N_VGND_c_525_n 0.00357877f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_c_262_n N_VGND_c_525_n 0.00357877f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_c_263_n N_VGND_c_525_n 0.00357877f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A_c_264_n N_VGND_c_525_n 0.00357877f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_c_261_n N_VGND_c_526_n 0.00566968f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_c_262_n N_VGND_c_526_n 0.00548399f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_c_263_n N_VGND_c_526_n 0.00548399f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_c_264_n N_VGND_c_526_n 0.0064529f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_248 A N_A_235_47#_M1010_d 0.00576272f $X=5.195 $Y=0.765 $X2=0 $Y2=0
cc_249 N_A_c_261_n N_A_235_47#_c_606_n 0.00107493f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_261_n N_A_235_47#_c_594_n 0.0135958f $X=3.445 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_262_n N_A_235_47#_c_594_n 0.00855322f $X=3.915 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_263_n N_A_235_47#_c_594_n 0.00861661f $X=4.385 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_c_264_n N_A_235_47#_c_594_n 0.0123256f $X=4.855 $Y=0.995 $X2=0 $Y2=0
cc_254 A N_A_235_47#_c_594_n 0.0335786f $X=5.195 $Y=0.765 $X2=0 $Y2=0
cc_255 N_A_c_266_n N_A_235_47#_c_594_n 0.00232829f $X=4.88 $Y=1.202 $X2=0 $Y2=0
cc_256 N_VPWR_c_328_n N_A_222_309#_M1000_s 0.00444633f $X=5.29 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_257 N_VPWR_c_328_n N_A_222_309#_M1014_s 0.00656398f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_328_n N_A_222_309#_M1007_d 0.00218326f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_328_n N_A_222_309#_M1011_d 0.00232878f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_260 N_VPWR_c_328_n N_A_222_309#_M1017_d 0.00357188f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_261 N_VPWR_c_330_n N_A_222_309#_c_407_n 0.0487409f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_334_n N_A_222_309#_c_407_n 0.0171175f $X=1.51 $Y=2.72 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_328_n N_A_222_309#_c_407_n 0.0103125f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_264 N_VPWR_M1003_d N_A_222_309#_c_402_n 0.00187091f $X=1.58 $Y=1.545 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_330_n N_A_222_309#_c_402_n 0.0209383f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_330_n N_A_222_309#_c_415_n 0.0385613f $X=1.725 $Y=2.02 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_331_n N_A_222_309#_c_415_n 0.0118139f $X=2.45 $Y=2.72 $X2=0
+ $Y2=0
cc_268 N_VPWR_c_332_n N_A_222_309#_c_415_n 0.0475804f $X=2.665 $Y=2 $X2=0 $Y2=0
cc_269 N_VPWR_c_328_n N_A_222_309#_c_415_n 0.00646998f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_270 N_VPWR_M1015_d N_A_222_309#_c_404_n 0.00285703f $X=2.52 $Y=1.545 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_332_n N_A_222_309#_c_404_n 0.0309049f $X=2.665 $Y=2 $X2=0 $Y2=0
cc_272 N_VPWR_c_332_n N_A_222_309#_c_419_n 0.0309218f $X=2.665 $Y=2 $X2=0 $Y2=0
cc_273 N_VPWR_c_335_n N_A_222_309#_c_431_n 0.0415557f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_328_n N_A_222_309#_c_431_n 0.027018f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_332_n N_A_222_309#_c_405_n 0.0124912f $X=2.665 $Y=2 $X2=0 $Y2=0
cc_276 N_VPWR_c_335_n N_A_222_309#_c_405_n 0.0147673f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_328_n N_A_222_309#_c_405_n 0.00808747f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_335_n N_A_222_309#_c_434_n 0.0535102f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_328_n N_A_222_309#_c_434_n 0.033565f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_335_n N_A_222_309#_c_462_n 0.0119545f $X=5.29 $Y=2.72 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_328_n N_A_222_309#_c_462_n 0.006547f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_c_328_n N_Z_M1007_s 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_328_n N_Z_M1012_s 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_284 N_A_222_309#_c_431_n N_Z_M1007_s 0.00374708f $X=4.09 $Y=2.38 $X2=0 $Y2=0
cc_285 N_A_222_309#_c_434_n N_Z_M1012_s 0.00374708f $X=5.03 $Y=2.38 $X2=0 $Y2=0
cc_286 N_A_222_309#_c_404_n N_Z_c_474_n 0.0141783f $X=3.11 $Y=1.58 $X2=0 $Y2=0
cc_287 N_A_222_309#_c_419_n N_Z_c_474_n 0.0310503f $X=3.235 $Y=1.815 $X2=0 $Y2=0
cc_288 N_A_222_309#_c_431_n N_Z_c_474_n 0.0154815f $X=4.09 $Y=2.38 $X2=0 $Y2=0
cc_289 N_A_222_309#_c_433_n N_Z_c_474_n 0.0260136f $X=4.175 $Y=1.815 $X2=0 $Y2=0
cc_290 N_A_222_309#_c_433_n N_Z_c_475_n 0.0317284f $X=4.175 $Y=1.815 $X2=0 $Y2=0
cc_291 N_A_222_309#_c_434_n N_Z_c_475_n 0.0154815f $X=5.03 $Y=2.38 $X2=0 $Y2=0
cc_292 N_A_222_309#_c_436_n N_Z_c_475_n 0.0260136f $X=5.115 $Y=1.815 $X2=0 $Y2=0
cc_293 N_A_222_309#_c_433_n N_Z_c_476_n 0.0153778f $X=4.175 $Y=1.815 $X2=0 $Y2=0
cc_294 N_Z_M1001_s N_VGND_c_526_n 0.00256987f $X=3.52 $Y=0.235 $X2=0 $Y2=0
cc_295 N_Z_M1009_s N_VGND_c_526_n 0.00256987f $X=4.46 $Y=0.235 $X2=0 $Y2=0
cc_296 N_Z_c_476_n N_A_235_47#_M1002_d 0.00219732f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_297 N_Z_c_476_n N_A_235_47#_c_606_n 0.0133517f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_298 N_Z_c_476_n N_A_235_47#_c_611_n 0.0023689f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_299 N_Z_M1001_s N_A_235_47#_c_594_n 0.00399896f $X=3.52 $Y=0.235 $X2=0 $Y2=0
cc_300 N_Z_M1009_s N_A_235_47#_c_594_n 0.00399896f $X=4.46 $Y=0.235 $X2=0 $Y2=0
cc_301 N_Z_c_476_n N_A_235_47#_c_594_n 0.0732838f $X=4.645 $Y=0.74 $X2=0 $Y2=0
cc_302 N_VGND_c_526_n N_A_235_47#_M1004_d 0.00229009f $X=5.29 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_303 N_VGND_c_526_n N_A_235_47#_M1005_d 0.00314422f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_304 N_VGND_c_526_n N_A_235_47#_M1013_d 0.00352323f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_305 N_VGND_c_526_n N_A_235_47#_M1002_d 0.00255381f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_306 N_VGND_c_526_n N_A_235_47#_M1010_d 0.00266737f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_307 N_VGND_c_518_n N_A_235_47#_c_592_n 0.0193139f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_308 N_VGND_c_519_n N_A_235_47#_c_592_n 0.0220167f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_309 N_VGND_c_526_n N_A_235_47#_c_592_n 0.0121907f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_310 N_VGND_M1004_s N_A_235_47#_c_599_n 0.0038973f $X=1.585 $Y=0.235 $X2=0
+ $Y2=0
cc_311 N_VGND_c_519_n N_A_235_47#_c_599_n 0.0029785f $X=1.605 $Y=0 $X2=0 $Y2=0
cc_312 N_VGND_c_520_n N_A_235_47#_c_599_n 0.0178569f $X=1.77 $Y=0.36 $X2=0 $Y2=0
cc_313 N_VGND_c_522_n N_A_235_47#_c_599_n 0.00310196f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_314 N_VGND_c_526_n N_A_235_47#_c_599_n 0.0122777f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_315 N_VGND_c_520_n N_A_235_47#_c_605_n 0.0139248f $X=1.77 $Y=0.36 $X2=0 $Y2=0
cc_316 N_VGND_c_522_n N_A_235_47#_c_605_n 0.011459f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_317 N_VGND_c_526_n N_A_235_47#_c_605_n 0.00644035f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_318 N_VGND_M1008_s N_A_235_47#_c_606_n 0.00397655f $X=2.525 $Y=0.235 $X2=0
+ $Y2=0
cc_319 N_VGND_c_521_n N_A_235_47#_c_606_n 0.0178569f $X=2.71 $Y=0.36 $X2=0 $Y2=0
cc_320 N_VGND_c_522_n N_A_235_47#_c_606_n 0.0029785f $X=2.545 $Y=0 $X2=0 $Y2=0
cc_321 N_VGND_c_525_n N_A_235_47#_c_606_n 0.00361096f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_322 N_VGND_c_526_n N_A_235_47#_c_606_n 0.0131245f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_323 N_VGND_c_521_n N_A_235_47#_c_611_n 0.00189407f $X=2.71 $Y=0.36 $X2=0
+ $Y2=0
cc_324 N_VGND_c_521_n N_A_235_47#_c_612_n 0.0119692f $X=2.71 $Y=0.36 $X2=0 $Y2=0
cc_325 N_VGND_c_525_n N_A_235_47#_c_612_n 0.0118015f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_326 N_VGND_c_526_n N_A_235_47#_c_612_n 0.00651702f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_327 N_VGND_c_525_n N_A_235_47#_c_594_n 0.122757f $X=5.29 $Y=0 $X2=0 $Y2=0
cc_328 N_VGND_c_526_n N_A_235_47#_c_594_n 0.0769936f $X=5.29 $Y=0 $X2=0 $Y2=0
