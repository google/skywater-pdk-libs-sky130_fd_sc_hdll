* File: sky130_fd_sc_hdll__dlygate4sd3_1.pex.spice
* Created: Thu Aug 27 19:06:47 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A 3 7 9 10 18
c32 18 0 9.35701e-20 $X=0.51 $Y=1.16
r33 17 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.51 $Y2=1.16
r34 14 17 32.3493 $w=3.3e-07 $l=1.85e-07 $layer=POLY_cond $X=0.31 $Y=1.16
+ $X2=0.495 $Y2=1.16
r35 9 10 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.345 $Y=1.16
+ $X2=0.345 $Y2=1.53
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.16 $X2=0.31 $Y2=1.16
r37 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.51 $Y=0.995
+ $X2=0.51 $Y2=1.16
r38 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.51 $Y=0.995 $X2=0.51
+ $Y2=0.445
r39 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r40 1 3 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 28 31 32 34
c70 34 0 1.21278e-19 $X=0.86 $Y=0.8
c71 32 0 7.01046e-20 $X=1.27 $Y=1.16
c72 25 0 9.35701e-20 $X=0.775 $Y=1.895
r73 32 39 16.3701 $w=6.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=1.325
r74 32 38 16.3701 $w=6.1e-07 $l=1.65e-07 $layer=POLY_cond $X=1.1 $Y=1.16 $X2=1.1
+ $Y2=0.995
r75 31 32 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r76 29 34 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.86 $Y=1.16
+ $X2=0.86 $Y2=0.8
r77 29 31 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.945 $Y=1.16
+ $X2=1.27 $Y2=1.16
r78 27 29 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=0.86 $Y=1.325
+ $X2=0.86 $Y2=1.16
r79 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.86 $Y=1.325
+ $X2=0.86 $Y2=1.785
r80 25 28 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.775 $Y=1.895
+ $X2=0.86 $Y2=1.785
r81 25 26 20.6916 $w=2.18e-07 $l=3.95e-07 $layer=LI1_cond $X=0.775 $Y=1.895
+ $X2=0.38 $Y2=1.895
r82 23 34 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=0.8
+ $X2=0.86 $Y2=0.8
r83 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.775 $Y=0.8
+ $X2=0.38 $Y2=0.8
r84 19 24 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.38 $Y2=0.8
r85 19 21 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.237 $Y2=0.51
r86 15 26 7.00622 $w=2.2e-07 $l=1.95407e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.38 $Y2=1.895
r87 15 17 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.232 $Y2=2.21
r88 13 39 101.656 $w=5e-07 $l=9.5e-07 $layer=POLY_cond $X=1.115 $Y=2.275
+ $X2=1.115 $Y2=1.325
r89 9 38 58.8532 $w=5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.115 $Y=0.445
+ $X2=1.115 $Y2=0.995
r90 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.21
r91 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_273_47# 1 2 7 9 12 14 16 19 25 30
+ 32
c57 19 0 1.76659e-19 $X=2.31 $Y=1.16
c58 7 0 1.2273e-19 $X=2.405 $Y=0.995
r59 28 30 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.5 $Y=2.32
+ $X2=1.655 $Y2=2.32
r60 23 25 6.15961 $w=2.88e-07 $l=1.55e-07 $layer=LI1_cond $X=1.5 $Y=0.4
+ $X2=1.655 $Y2=0.4
r61 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.31
+ $Y=1.16 $X2=2.31 $Y2=1.16
r62 17 32 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.74 $Y=1.175
+ $X2=1.655 $Y2=1.175
r63 17 19 31.6091 $w=1.98e-07 $l=5.7e-07 $layer=LI1_cond $X=1.74 $Y=1.175
+ $X2=2.31 $Y2=1.175
r64 16 30 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.655 $Y=2.175
+ $X2=1.655 $Y2=2.32
r65 15 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.655 $Y=1.275
+ $X2=1.655 $Y2=1.175
r66 15 16 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.655 $Y=1.275
+ $X2=1.655 $Y2=2.175
r67 14 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.655 $Y=1.075
+ $X2=1.655 $Y2=1.175
r68 13 25 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.655 $Y=0.545
+ $X2=1.655 $Y2=0.4
r69 13 14 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.655 $Y=0.545
+ $X2=1.655 $Y2=1.075
r70 7 20 16.6118 $w=3.3e-07 $l=9.5e-08 $layer=POLY_cond $X=2.405 $Y=1.16
+ $X2=2.31 $Y2=1.16
r71 7 12 56.876 $w=5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.405 $Y=1.325 $X2=2.405
+ $Y2=1.915
r72 7 9 30.848 $w=5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.405 $Y=0.995 $X2=2.405
+ $Y2=0.675
r73 2 28 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.365
+ $Y=2.065 $X2=1.5 $Y2=2.34
r74 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.365
+ $Y=0.235 $X2=1.5 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_379_93# 1 2 9 13 16 18 19 20 22 23
+ 25 32 34
c57 32 0 1.76659e-19 $X=3.03 $Y=1.16
r58 32 35 40.7387 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.037 $Y=1.16
+ $X2=3.037 $Y2=1.325
r59 32 34 46.3655 $w=3.45e-07 $l=1.65e-07 $layer=POLY_cond $X=3.037 $Y=1.16
+ $X2=3.037 $Y2=0.995
r60 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.03
+ $Y=1.16 $X2=3.03 $Y2=1.16
r61 29 31 14.5544 $w=2.85e-07 $l=3.4e-07 $layer=LI1_cond $X=2.982 $Y=0.82
+ $X2=2.982 $Y2=1.16
r62 25 27 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=2.025 $Y=0.675
+ $X2=2.025 $Y2=0.82
r63 22 31 7.93228 $w=2.85e-07 $l=1.95653e-07 $layer=LI1_cond $X=2.915 $Y=1.325
+ $X2=2.982 $Y2=1.16
r64 22 23 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=2.915 $Y=1.325
+ $X2=2.915 $Y2=1.575
r65 21 27 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.14 $Y=0.82
+ $X2=2.025 $Y2=0.82
r66 20 29 3.76007 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=2.81 $Y=0.82
+ $X2=2.982 $Y2=0.82
r67 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.81 $Y=0.82
+ $X2=2.14 $Y2=0.82
r68 18 23 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.81 $Y=1.66
+ $X2=2.915 $Y2=1.575
r69 18 19 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.81 $Y=1.66
+ $X2=2.13 $Y2=1.66
r70 14 19 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.02 $Y=1.745
+ $X2=2.13 $Y2=1.66
r71 14 16 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=2.02 $Y=1.745
+ $X2=2.02 $Y2=1.915
r72 13 34 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.135 $Y=0.56
+ $X2=3.135 $Y2=0.995
r73 9 35 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=3.12 $Y=1.985
+ $X2=3.12 $Y2=1.325
r74 2 16 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=1.895
+ $Y=1.705 $X2=2.02 $Y2=1.915
r75 1 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.465 $X2=2.02 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VPWR 1 2 9 13 18 19 20 22 35 36 39
+ 44
r40 40 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r41 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r42 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r43 33 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r44 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r45 30 33 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r46 30 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 29 32 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.53 $Y2=2.72
r48 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 27 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=0.73 $Y2=2.72
r50 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.855 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 24 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 22 39 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.73 $Y2=2.72
r53 22 24 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 20 44 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 18 32 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=2.72
+ $X2=2.855 $Y2=2.72
r57 17 35 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=2.72
+ $X2=2.855 $Y2=2.72
r59 13 16 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=2.855 $Y=2 $X2=2.855
+ $Y2=2.34
r60 11 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=2.635
+ $X2=2.855 $Y2=2.72
r61 11 16 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.855 $Y=2.635
+ $X2=2.855 $Y2=2.34
r62 7 39 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r63 7 9 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.34
r64 2 16 600 $w=1.7e-07 $l=7.28166e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=1.705 $X2=2.855 $Y2=2.34
r65 2 13 600 $w=1.7e-07 $l=3.82132e-07 $layer=licon1_PDIFF $count=1 $X=2.655
+ $Y=1.705 $X2=2.855 $Y2=2
r66 1 9 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%X 1 2 7 8 9 10 11 12 24 38 45
c19 45 0 1.2273e-19 $X=3.45 $Y=1.53
r20 45 46 2.27943 $w=4.03e-07 $l=3.5e-08 $layer=LI1_cond $X=3.392 $Y=1.53
+ $X2=3.392 $Y2=1.495
r21 29 49 1.05285 $w=4.03e-07 $l=3.7e-08 $layer=LI1_cond $X=3.392 $Y=1.697
+ $X2=3.392 $Y2=1.66
r22 24 43 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.46 $Y=0.85
+ $X2=3.46 $Y2=0.825
r23 12 35 3.6992 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=3.392 $Y=2.21
+ $X2=3.392 $Y2=2.34
r24 11 12 9.67483 $w=4.03e-07 $l=3.4e-07 $layer=LI1_cond $X=3.392 $Y=1.87
+ $X2=3.392 $Y2=2.21
r25 11 29 4.92278 $w=4.03e-07 $l=1.73e-07 $layer=LI1_cond $X=3.392 $Y=1.87
+ $X2=3.392 $Y2=1.697
r26 10 49 2.98782 $w=4.03e-07 $l=1.05e-07 $layer=LI1_cond $X=3.392 $Y=1.555
+ $X2=3.392 $Y2=1.66
r27 10 45 0.711385 $w=4.03e-07 $l=2.5e-08 $layer=LI1_cond $X=3.392 $Y=1.555
+ $X2=3.392 $Y2=1.53
r28 10 46 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.46 $Y=1.47
+ $X2=3.46 $Y2=1.495
r29 9 10 11.9513 $w=2.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.46 $Y=1.19 $X2=3.46
+ $Y2=1.47
r30 8 43 2.13715 $w=4.03e-07 $l=3e-08 $layer=LI1_cond $X=3.392 $Y=0.795
+ $X2=3.392 $Y2=0.825
r31 8 9 13.2318 $w=2.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.46 $Y=0.88 $X2=3.46
+ $Y2=1.19
r32 8 24 1.28049 $w=2.68e-07 $l=3e-08 $layer=LI1_cond $X=3.46 $Y=0.88 $X2=3.46
+ $Y2=0.85
r33 7 8 8.10978 $w=4.03e-07 $l=2.85e-07 $layer=LI1_cond $X=3.392 $Y=0.51
+ $X2=3.392 $Y2=0.795
r34 7 38 3.6992 $w=4.03e-07 $l=1.3e-07 $layer=LI1_cond $X=3.392 $Y=0.51
+ $X2=3.392 $Y2=0.38
r35 2 49 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.485 $X2=3.355 $Y2=1.66
r36 2 35 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.21
+ $Y=1.485 $X2=3.355 $Y2=2.34
r37 1 38 91 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=2 $X=3.21
+ $Y=0.235 $X2=3.355 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VGND 1 2 9 13 16 17 18 20 33 34 37
+ 42
c45 9 0 7.01046e-20 $X=0.73 $Y=0.38
r46 38 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r47 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r48 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r50 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r51 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r52 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r53 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r54 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r55 25 37 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.707
+ $Y2=0
r56 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r57 22 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r58 20 37 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.707
+ $Y2=0
r59 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.23
+ $Y2=0
r60 18 42 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r61 16 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.53
+ $Y2=0
r62 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.69 $Y=0 $X2=2.855
+ $Y2=0
r63 15 33 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=3.45
+ $Y2=0
r64 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.02 $Y=0 $X2=2.855
+ $Y2=0
r65 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0
r66 11 13 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.855 $Y=0.085
+ $X2=2.855 $Y2=0.44
r67 7 37 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0
r68 7 9 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0.38
r69 2 13 182 $w=1.7e-07 $l=2.12132e-07 $layer=licon1_NDIFF $count=1 $X=2.655
+ $Y=0.465 $X2=2.855 $Y2=0.44
r70 1 9 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=0.585
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

