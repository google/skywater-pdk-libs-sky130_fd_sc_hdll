# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a2bb2oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a2bb2oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.545000 1.075000 8.070000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.440000 1.075000 9.965000 1.275000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.075000 1.705000 1.285000 ;
        RECT 1.535000 1.285000 1.705000 1.445000 ;
        RECT 1.535000 1.445000 3.975000 1.615000 ;
        RECT 3.595000 1.075000 3.975000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.875000 1.075000 3.425000 1.275000 ;
    END
  END B2
  PIN Y
    ANTENNADIFFAREA  1.477000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.645000 3.295000 0.725000 ;
        RECT 1.925000 0.725000 5.595000 0.905000 ;
        RECT 4.145000 0.905000 4.365000 1.415000 ;
        RECT 4.145000 1.415000 5.515000 1.615000 ;
        RECT 4.275000 0.275000 4.655000 0.725000 ;
        RECT 4.365000 1.615000 4.615000 2.125000 ;
        RECT 5.215000 0.275000 5.595000 0.725000 ;
        RECT 5.245000 1.615000 5.515000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.085000  1.455000  1.315000 1.625000 ;
      RECT  0.085000  1.625000  0.425000 2.465000 ;
      RECT  0.175000  0.085000  0.345000 0.895000 ;
      RECT  0.515000  0.255000  0.895000 0.725000 ;
      RECT  0.515000  0.725000  1.755000 0.905000 ;
      RECT  0.645000  1.795000  0.855000 2.635000 ;
      RECT  1.075000  1.625000  1.315000 1.795000 ;
      RECT  1.075000  1.795000  4.145000 1.965000 ;
      RECT  1.075000  1.965000  1.315000 2.465000 ;
      RECT  1.115000  0.085000  1.285000 0.555000 ;
      RECT  1.455000  0.255000  3.715000 0.475000 ;
      RECT  1.455000  0.475000  1.755000 0.725000 ;
      RECT  1.545000  2.135000  1.795000 2.635000 ;
      RECT  2.015000  1.965000  2.265000 2.465000 ;
      RECT  2.485000  2.135000  2.735000 2.635000 ;
      RECT  2.955000  1.965000  3.205000 2.465000 ;
      RECT  3.425000  2.135000  3.675000 2.635000 ;
      RECT  3.895000  1.965000  4.145000 2.295000 ;
      RECT  3.895000  2.295000  6.065000 2.465000 ;
      RECT  3.935000  0.085000  4.105000 0.555000 ;
      RECT  4.535000  1.075000  6.325000 1.245000 ;
      RECT  4.835000  1.795000  5.075000 2.295000 ;
      RECT  4.875000  0.085000  5.045000 0.555000 ;
      RECT  5.685000  1.455000  6.065000 2.295000 ;
      RECT  5.815000  0.085000  6.505000 0.555000 ;
      RECT  6.155000  0.735000 10.460000 0.905000 ;
      RECT  6.155000  0.905000  6.325000 1.075000 ;
      RECT  6.255000  1.455000  8.425000 1.625000 ;
      RECT  6.255000  1.625000  6.585000 2.465000 ;
      RECT  6.675000  0.255000  7.055000 0.725000 ;
      RECT  6.675000  0.725000  9.875000 0.735000 ;
      RECT  6.805000  1.795000  7.015000 2.635000 ;
      RECT  7.240000  1.625000  7.480000 2.465000 ;
      RECT  7.275000  0.085000  7.445000 0.555000 ;
      RECT  7.615000  0.255000  7.995000 0.725000 ;
      RECT  7.705000  1.795000  7.955000 2.635000 ;
      RECT  8.175000  1.625000  8.425000 2.295000 ;
      RECT  8.175000  2.295000 10.310000 2.465000 ;
      RECT  8.215000  0.085000  8.385000 0.555000 ;
      RECT  8.555000  0.255000  8.935000 0.725000 ;
      RECT  8.645000  1.455000 10.460000 1.625000 ;
      RECT  8.645000  1.625000  8.895000 2.125000 ;
      RECT  9.115000  1.795000  9.365000 2.295000 ;
      RECT  9.155000  0.085000  9.325000 0.555000 ;
      RECT  9.495000  0.255000  9.875000 0.725000 ;
      RECT  9.585000  1.625000  9.835000 2.125000 ;
      RECT 10.060000  1.795000 10.310000 2.295000 ;
      RECT 10.095000  0.085000 10.265000 0.555000 ;
      RECT 10.135000  0.905000 10.460000 1.455000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a2bb2oi_4
END LIBRARY
