* File: sky130_fd_sc_hdll__or4_2.spice
* Created: Thu Aug 27 19:24:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4_2.pex.spice"
.subckt sky130_fd_sc_hdll__or4_2  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 N_A_27_297#_M1000_d N_D_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.1302 PD=0.8 PS=1.46 NRD=7.14 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.9 A=0.063 P=1.14 MULT=1
MM1006 N_VGND_M1006_d N_C_M1006_g N_A_27_297#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0798 PD=0.74 PS=0.8 NRD=0 NRS=21.42 M=1 R=2.8 SA=75000.8
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1005 N_A_27_297#_M1005_d N_B_M1005_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0672 PD=0.74 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.2
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_A_27_297#_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0799766 AS=0.0672 PD=0.777196 PS=0.74 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_X_M1002_d N_A_27_297#_M1002_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.173875 AS=0.123773 PD=1.185 PS=1.2028 NRD=38.76 NRS=2.76 M=1 R=4.33333
+ SA=75001.5 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1002_d N_A_27_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.173875 AS=0.19825 PD=1.185 PS=1.91 NRD=8.304 NRS=3.684 M=1 R=4.33333
+ SA=75002.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_117_297# N_D_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0735 AS=0.1134 PD=0.77 PS=1.38 NRD=56.2829 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.9 A=0.0756 P=1.2 MULT=1
MM1010 A_223_297# N_C_M1010_g A_117_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0483
+ AS=0.0735 PD=0.65 PS=0.77 NRD=28.1316 NRS=56.2829 M=1 R=2.33333 SA=90000.7
+ SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1011 A_305_297# N_B_M1011_g A_223_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0735
+ AS=0.0483 PD=0.77 PS=0.65 NRD=56.2829 NRS=28.1316 M=1 R=2.33333 SA=90001.1
+ SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_305_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0735 PD=0.804507 PS=0.77 NRD=76.83 NRS=56.2829 M=1 R=2.33333
+ SA=90001.6 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1004_d N_A_27_297#_M1007_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.218803 AS=0.2275 PD=1.91549 PS=1.455 NRD=1.9503 NRS=33.4703 M=1 R=5.55556
+ SA=90001 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_27_297#_M1009_g N_X_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.315 AS=0.2275 PD=2.63 PS=1.455 NRD=5.91 NRS=0.9653 M=1 R=5.55556
+ SA=90001.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX13_noxref noxref_14 A A PROBETYPE=1
c_66 VPB 0 8.49032e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or4_2.pxi.spice"
*
.ends
*
*
