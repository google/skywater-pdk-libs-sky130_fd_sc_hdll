# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sedfxbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sedfxbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  16.56000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.795000 0.765000 2.155000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.325000 0.765000 2.765000 1.185000 ;
        RECT 2.325000 1.185000 2.525000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.530500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.320000 0.255000 15.700000 2.420000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.935000 1.065000 13.430000 1.300000 ;
        RECT 12.935000 1.300000 13.315000 2.465000 ;
        RECT 13.100000 0.255000 13.430000 1.065000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.445000 1.105000 6.950000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.605000 1.105000 5.885000 1.615000 ;
    END
  END SCE
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 16.560000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  2.385000  0.085000  2.765000 0.515000 ;
        RECT  3.385000  0.085000  3.765000 0.610000 ;
        RECT  6.445000  0.085000  6.695000 0.905000 ;
        RECT  9.180000  0.085000  9.575000 0.560000 ;
        RECT 10.450000  0.085000 10.725000 0.615000 ;
        RECT 12.630000  0.085000 12.880000 0.900000 ;
        RECT 13.650000  0.085000 13.900000 0.900000 ;
        RECT 14.915000  0.085000 15.150000 0.900000 ;
        RECT 15.920000  0.085000 16.180000 0.900000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
        RECT 14.865000 -0.085000 15.035000 0.085000 ;
        RECT 15.325000 -0.085000 15.495000 0.085000 ;
        RECT 15.785000 -0.085000 15.955000 0.085000 ;
        RECT 16.245000 -0.085000 16.415000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 16.560000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 16.560000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  2.385000 1.890000  2.765000 2.635000 ;
        RECT  3.515000 1.825000  3.710000 2.635000 ;
        RECT  6.350000 2.175000  6.695000 2.635000 ;
        RECT  9.360000 1.835000  9.595000 2.635000 ;
        RECT 10.355000 2.105000 10.645000 2.635000 ;
        RECT 12.595000 1.495000 12.765000 2.635000 ;
        RECT 13.535000 1.465000 13.785000 2.635000 ;
        RECT 14.915000 1.465000 15.150000 2.635000 ;
        RECT 15.920000 1.465000 16.180000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
        RECT 14.405000 2.635000 14.575000 2.805000 ;
        RECT 14.865000 2.635000 15.035000 2.805000 ;
        RECT 15.325000 2.635000 15.495000 2.805000 ;
        RECT 15.785000 2.635000 15.955000 2.805000 ;
        RECT 16.245000 2.635000 16.415000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 16.560000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.175000 0.345000  0.345000 0.635000 ;
      RECT  0.175000 0.635000  0.895000 0.805000 ;
      RECT  0.175000 1.795000  0.895000 1.965000 ;
      RECT  0.175000 1.965000  0.345000 2.465000 ;
      RECT  0.665000 0.805000  0.895000 1.795000 ;
      RECT  1.115000 0.345000  1.285000 2.465000 ;
      RECT  1.455000 0.255000  1.885000 0.515000 ;
      RECT  1.455000 0.515000  1.625000 1.890000 ;
      RECT  1.455000 1.890000  1.885000 2.465000 ;
      RECT  2.695000 1.355000  3.285000 1.720000 ;
      RECT  2.955000 1.720000  3.285000 2.425000 ;
      RECT  2.980000 0.255000  3.205000 0.845000 ;
      RECT  2.980000 0.845000  3.885000 1.175000 ;
      RECT  2.980000 1.175000  3.285000 1.355000 ;
      RECT  4.105000 0.685000  4.275000 1.320000 ;
      RECT  4.105000 1.320000  4.525000 1.650000 ;
      RECT  4.425000 1.820000  4.865000 2.020000 ;
      RECT  4.425000 2.020000  4.805000 2.465000 ;
      RECT  4.445000 0.255000  4.765000 0.980000 ;
      RECT  4.445000 0.980000  4.865000 1.150000 ;
      RECT  4.695000 1.150000  4.865000 1.820000 ;
      RECT  4.995000 0.255000  5.195000 0.645000 ;
      RECT  4.995000 0.645000  5.255000 0.825000 ;
      RECT  5.035000 2.210000  5.365000 2.465000 ;
      RECT  5.085000 0.825000  5.255000 1.785000 ;
      RECT  5.085000 1.785000  5.365000 2.210000 ;
      RECT  5.365000 0.255000  6.225000 0.515000 ;
      RECT  5.790000 1.835000  7.370000 2.005000 ;
      RECT  5.790000 2.005000  6.130000 2.465000 ;
      RECT  5.895000 0.515000  6.225000 0.935000 ;
      RECT  6.055000 0.935000  6.225000 1.835000 ;
      RECT  7.120000 1.355000  7.370000 1.835000 ;
      RECT  7.300000 0.255000  7.920000 0.565000 ;
      RECT  7.300000 0.565000  7.710000 1.185000 ;
      RECT  7.460000 2.150000  7.790000 2.465000 ;
      RECT  7.540000 1.185000  7.710000 1.865000 ;
      RECT  7.540000 1.865000  7.790000 2.150000 ;
      RECT  7.880000 1.125000  8.115000 1.720000 ;
      RECT  7.900000 0.735000  8.455000 0.955000 ;
      RECT  8.000000 2.175000  9.190000 2.375000 ;
      RECT  8.140000 0.255000  8.865000 0.565000 ;
      RECT  8.285000 0.955000  8.455000 1.655000 ;
      RECT  8.285000 1.655000  8.800000 2.005000 ;
      RECT  8.695000 0.565000  8.865000 1.315000 ;
      RECT  8.695000 1.315000  9.595000 1.485000 ;
      RECT  8.970000 1.485000  9.595000 1.575000 ;
      RECT  8.970000 1.575000  9.190000 2.175000 ;
      RECT  9.055000 0.765000 10.220000 1.045000 ;
      RECT  9.055000 1.045000 10.730000 1.065000 ;
      RECT  9.055000 1.065000  9.305000 1.095000 ;
      RECT  9.425000 1.245000  9.595000 1.315000 ;
      RECT  9.765000 0.255000 10.220000 0.765000 ;
      RECT  9.765000 1.065000 10.730000 1.375000 ;
      RECT  9.765000 1.375000 10.145000 2.465000 ;
      RECT 11.125000 1.245000 11.365000 1.965000 ;
      RECT 11.260000 2.165000 12.375000 2.355000 ;
      RECT 11.390000 0.705000 11.905000 1.035000 ;
      RECT 11.410000 0.330000 12.375000 0.535000 ;
      RECT 11.535000 1.035000 11.905000 1.995000 ;
      RECT 12.125000 0.535000 12.375000 2.165000 ;
      RECT 13.955000 1.575000 14.185000 2.010000 ;
      RECT 14.070000 0.890000 14.695000 1.220000 ;
      RECT 14.355000 0.255000 14.695000 0.890000 ;
      RECT 14.355000 1.220000 14.695000 2.465000 ;
    LAYER mcon ;
      RECT  0.685000 1.785000  0.855000 1.955000 ;
      RECT  1.115000 1.445000  1.285000 1.615000 ;
      RECT  1.455000 0.425000  1.625000 0.595000 ;
      RECT  4.105000 0.765000  4.275000 0.935000 ;
      RECT  4.535000 0.425000  4.705000 0.595000 ;
      RECT  5.015000 0.425000  5.185000 0.595000 ;
      RECT  7.315000 0.425000  7.485000 0.595000 ;
      RECT  7.910000 1.445000  8.080000 1.615000 ;
      RECT  8.345000 1.785000  8.515000 1.955000 ;
      RECT 11.160000 1.785000 11.330000 1.955000 ;
      RECT 11.630000 1.445000 11.800000 1.615000 ;
      RECT 12.165000 1.785000 12.335000 1.955000 ;
      RECT 13.985000 1.785000 14.155000 1.955000 ;
      RECT 14.445000 0.765000 14.615000 0.935000 ;
    LAYER met1 ;
      RECT  0.625000 1.755000  0.915000 1.800000 ;
      RECT  0.625000 1.800000 11.415000 1.940000 ;
      RECT  0.625000 1.940000  0.915000 1.985000 ;
      RECT  1.005000 1.415000  1.345000 1.460000 ;
      RECT  1.005000 1.460000 11.885000 1.600000 ;
      RECT  1.005000 1.600000  1.345000 1.645000 ;
      RECT  1.395000 0.395000  4.765000 0.580000 ;
      RECT  1.395000 0.580000  1.685000 0.625000 ;
      RECT  4.045000 0.735000  4.335000 0.780000 ;
      RECT  4.045000 0.780000 14.675000 0.920000 ;
      RECT  4.045000 0.920000  4.335000 0.965000 ;
      RECT  4.425000 0.580000  4.765000 0.625000 ;
      RECT  4.905000 0.395000  7.545000 0.580000 ;
      RECT  4.905000 0.580000  5.245000 0.625000 ;
      RECT  7.205000 0.580000  7.545000 0.625000 ;
      RECT  7.825000 1.415000  8.165000 1.460000 ;
      RECT  7.825000 1.600000  8.165000 1.645000 ;
      RECT  8.285000 1.755000  8.625000 1.800000 ;
      RECT  8.285000 1.940000  8.625000 1.985000 ;
      RECT 11.075000 1.755000 11.415000 1.800000 ;
      RECT 11.075000 1.940000 11.415000 1.985000 ;
      RECT 11.545000 1.415000 11.885000 1.460000 ;
      RECT 11.545000 1.600000 11.885000 1.645000 ;
      RECT 12.105000 1.755000 12.395000 1.800000 ;
      RECT 12.105000 1.800000 14.215000 1.940000 ;
      RECT 12.105000 1.940000 12.395000 1.985000 ;
      RECT 13.925000 1.755000 14.215000 1.800000 ;
      RECT 13.925000 1.940000 14.215000 1.985000 ;
      RECT 14.385000 0.735000 14.675000 0.780000 ;
      RECT 14.385000 0.920000 14.675000 0.965000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sedfxbp_2
