# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nor4bb_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nor4bb_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.465000 1.075000 6.330000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.400000 1.075000 5.295000 1.275000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.000000 0.995000 1.270000 1.325000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.830000 1.695000 ;
    END
  END D_N
  PIN VGND
    ANTENNADIFFAREA  1.295950 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 6.440000 0.085000 ;
        RECT 0.685000  0.085000 0.855000 0.825000 ;
        RECT 1.595000  0.085000 1.925000 0.480000 ;
        RECT 2.695000  0.085000 2.865000 0.555000 ;
        RECT 3.635000  0.085000 4.345000 0.555000 ;
        RECT 5.115000  0.085000 5.285000 0.555000 ;
        RECT 6.055000  0.085000 6.330000 0.905000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.543625 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 6.440000 2.805000 ;
        RECT 0.515000 2.240000 0.895000 2.635000 ;
        RECT 5.545000 1.795000 5.755000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.219500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.095000 0.255000 2.475000 0.725000 ;
        RECT 2.095000 0.725000 5.835000 0.905000 ;
        RECT 3.035000 0.255000 3.415000 0.725000 ;
        RECT 3.035000 1.445000 4.230000 1.705000 ;
        RECT 3.810000 0.905000 4.230000 1.445000 ;
        RECT 4.515000 0.255000 4.895000 0.725000 ;
        RECT 5.455000 0.255000 5.835000 0.725000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.085000 0.450000 0.465000 0.825000 ;
      RECT 0.085000 0.825000 0.255000 1.885000 ;
      RECT 0.085000 1.885000 1.950000 2.055000 ;
      RECT 0.085000 2.055000 0.345000 2.455000 ;
      RECT 1.045000 1.525000 1.610000 1.715000 ;
      RECT 1.155000 0.450000 1.350000 0.655000 ;
      RECT 1.155000 0.655000 1.610000 0.825000 ;
      RECT 1.440000 0.825000 1.610000 1.075000 ;
      RECT 1.440000 1.075000 2.475000 1.245000 ;
      RECT 1.440000 1.245000 1.610000 1.525000 ;
      RECT 1.675000 2.225000 3.885000 2.465000 ;
      RECT 1.780000 1.415000 2.865000 1.585000 ;
      RECT 1.780000 1.585000 1.950000 1.885000 ;
      RECT 2.145000 1.875000 4.895000 2.045000 ;
      RECT 2.695000 1.075000 3.640000 1.275000 ;
      RECT 2.695000 1.275000 2.865000 1.415000 ;
      RECT 4.095000 2.215000 5.325000 2.465000 ;
      RECT 4.605000 1.455000 4.895000 1.875000 ;
      RECT 5.115000 1.455000 6.305000 1.625000 ;
      RECT 5.115000 1.625000 5.325000 2.215000 ;
      RECT 5.925000 1.625000 6.305000 2.465000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nor4bb_2
