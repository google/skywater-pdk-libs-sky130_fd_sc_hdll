* File: sky130_fd_sc_hdll__isobufsrc_4.pxi.spice
* Created: Thu Aug 27 19:10:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%SLEEP N_SLEEP_c_86_n N_SLEEP_M1002_g
+ N_SLEEP_c_92_n N_SLEEP_M1001_g N_SLEEP_c_87_n N_SLEEP_M1007_g N_SLEEP_c_93_n
+ N_SLEEP_M1003_g N_SLEEP_c_88_n N_SLEEP_M1008_g N_SLEEP_c_94_n N_SLEEP_M1006_g
+ N_SLEEP_c_95_n N_SLEEP_M1012_g N_SLEEP_c_89_n N_SLEEP_M1015_g SLEEP
+ N_SLEEP_c_90_n N_SLEEP_c_91_n SLEEP PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%SLEEP
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A_459_21# N_A_459_21#_M1011_s
+ N_A_459_21#_M1010_s N_A_459_21#_c_164_n N_A_459_21#_M1004_g
+ N_A_459_21#_c_174_n N_A_459_21#_M1000_g N_A_459_21#_c_165_n
+ N_A_459_21#_M1005_g N_A_459_21#_c_175_n N_A_459_21#_M1009_g
+ N_A_459_21#_c_166_n N_A_459_21#_M1013_g N_A_459_21#_c_176_n
+ N_A_459_21#_M1014_g N_A_459_21#_c_177_n N_A_459_21#_M1017_g
+ N_A_459_21#_c_167_n N_A_459_21#_M1016_g N_A_459_21#_c_210_p
+ N_A_459_21#_c_168_n N_A_459_21#_c_169_n N_A_459_21#_c_170_n
+ N_A_459_21#_c_179_n N_A_459_21#_c_171_n N_A_459_21#_c_172_n
+ N_A_459_21#_c_180_n N_A_459_21#_c_181_n N_A_459_21#_c_173_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A_459_21#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A N_A_c_280_n N_A_M1011_g N_A_c_283_n
+ N_A_M1010_g A N_A_c_282_n A PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A_27_297# N_A_27_297#_M1001_s
+ N_A_27_297#_M1003_s N_A_27_297#_M1012_s N_A_27_297#_M1009_s
+ N_A_27_297#_M1017_s N_A_27_297#_c_308_n N_A_27_297#_c_309_n
+ N_A_27_297#_c_310_n N_A_27_297#_c_355_p N_A_27_297#_c_311_n
+ N_A_27_297#_c_312_n N_A_27_297#_c_328_n N_A_27_297#_c_336_n
+ N_A_27_297#_c_338_n N_A_27_297#_c_313_n N_A_27_297#_c_314_n
+ N_A_27_297#_c_315_n N_A_27_297#_c_347_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%VPWR N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1010_d N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n
+ VPWR N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n
+ N_VPWR_c_405_n N_VPWR_c_396_n PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%VPWR
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%X N_X_M1002_s N_X_M1008_s N_X_M1004_d
+ N_X_M1013_d N_X_M1000_d N_X_M1014_d N_X_c_479_n N_X_c_468_n N_X_c_469_n
+ N_X_c_490_n N_X_c_470_n N_X_c_494_n N_X_c_471_n N_X_c_533_n N_X_c_472_n
+ N_X_c_516_n N_X_c_476_n N_X_c_537_n N_X_c_473_n N_X_c_474_n N_X_c_477_n
+ N_X_c_478_n X PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%X
x_PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%VGND N_VGND_M1002_d N_VGND_M1007_d
+ N_VGND_M1015_d N_VGND_M1005_s N_VGND_M1016_s N_VGND_M1011_d N_VGND_c_582_n
+ N_VGND_c_583_n N_VGND_c_584_n N_VGND_c_585_n N_VGND_c_586_n N_VGND_c_587_n
+ N_VGND_c_588_n N_VGND_c_589_n N_VGND_c_590_n N_VGND_c_591_n N_VGND_c_592_n
+ N_VGND_c_593_n N_VGND_c_594_n N_VGND_c_595_n N_VGND_c_596_n VGND
+ N_VGND_c_597_n N_VGND_c_598_n N_VGND_c_599_n
+ PM_SKY130_FD_SC_HDLL__ISOBUFSRC_4%VGND
cc_1 VNB N_SLEEP_c_86_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_SLEEP_c_87_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_SLEEP_c_88_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_SLEEP_c_89_n 0.0169164f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_SLEEP_c_90_n 0.0105081f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_6 VNB N_SLEEP_c_91_n 0.081832f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_A_459_21#_c_164_n 0.0164599f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_8 VNB N_A_459_21#_c_165_n 0.0163741f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_9 VNB N_A_459_21#_c_166_n 0.0171716f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_10 VNB N_A_459_21#_c_167_n 0.0207384f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_11 VNB N_A_459_21#_c_168_n 0.0442418f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_12 VNB N_A_459_21#_c_169_n 0.00335056f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_13 VNB N_A_459_21#_c_170_n 0.00363351f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_14 VNB N_A_459_21#_c_171_n 0.00134522f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_459_21#_c_172_n 0.00117446f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_459_21#_c_173_n 0.0706411f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_c_280_n 0.024631f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_18 VNB A 0.0154621f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_19 VNB N_A_c_282_n 0.0436188f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_20 VNB N_VPWR_c_396_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_468_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_22 VNB N_X_c_469_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_23 VNB N_X_c_470_n 0.0042799f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.202
cc_24 VNB N_X_c_471_n 8.90776e-19 $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.202
cc_25 VNB N_X_c_472_n 0.00582316f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_26 VNB N_X_c_473_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_474_n 0.00375367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_582_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_29 VNB N_VGND_c_583_n 0.0354575f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_30 VNB N_VGND_c_584_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_31 VNB N_VGND_c_585_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_32 VNB N_VGND_c_586_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_33 VNB N_VGND_c_587_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_34 VNB N_VGND_c_588_n 0.0142632f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_35 VNB N_VGND_c_589_n 0.0159132f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_36 VNB N_VGND_c_590_n 0.0336476f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_37 VNB N_VGND_c_591_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.175
cc_38 VNB N_VGND_c_592_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_593_n 0.019174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_594_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_595_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_596_n 0.00557808f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_597_n 0.0199516f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_598_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_599_n 0.289053f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VPB N_SLEEP_c_92_n 0.0198936f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_47 VPB N_SLEEP_c_93_n 0.0158033f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_48 VPB N_SLEEP_c_94_n 0.015524f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_49 VPB N_SLEEP_c_95_n 0.0160989f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_50 VPB N_SLEEP_c_91_n 0.0483884f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_51 VPB N_A_459_21#_c_174_n 0.0162273f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_52 VPB N_A_459_21#_c_175_n 0.0157312f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_53 VPB N_A_459_21#_c_176_n 0.0158699f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_54 VPB N_A_459_21#_c_177_n 0.0196978f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_55 VPB N_A_459_21#_c_168_n 0.021667f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_56 VPB N_A_459_21#_c_179_n 0.00630951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_459_21#_c_180_n 0.00139033f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_459_21#_c_181_n 0.00516618f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_459_21#_c_173_n 0.0497241f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_c_283_n 0.023968f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_61 VPB A 0.00365733f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=0.995
cc_62 VPB N_A_c_282_n 0.0193015f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_63 VPB N_A_27_297#_c_308_n 0.0133505f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_64 VPB N_A_27_297#_c_309_n 0.0309889f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_65 VPB N_A_27_297#_c_310_n 0.00262139f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_66 VPB N_A_27_297#_c_311_n 0.00210179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_297#_c_312_n 0.00441003f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_68 VPB N_A_27_297#_c_313_n 0.00218233f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=1.202
cc_69 VPB N_A_27_297#_c_314_n 0.00755385f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_70 VPB N_A_27_297#_c_315_n 0.00104475f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.175
cc_71 VPB N_VPWR_c_397_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_72 VPB N_VPWR_c_398_n 0.00229677f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_73 VPB N_VPWR_c_399_n 0.014431f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_74 VPB N_VPWR_c_400_n 0.0516989f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_75 VPB N_VPWR_c_401_n 0.0155059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_402_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_77 VPB N_VPWR_c_403_n 0.0760872f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_78 VPB N_VPWR_c_404_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.175
cc_79 VPB N_VPWR_c_405_n 0.00426137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_396_n 0.0537008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_X_c_471_n 0.00117186f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_82 VPB N_X_c_476_n 0.00148925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_X_c_477_n 3.0028e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_X_c_478_n 0.00233651f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 N_SLEEP_c_89_n N_A_459_21#_c_164_n 0.0243795f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_86 N_SLEEP_c_95_n N_A_459_21#_c_174_n 0.00965962f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_87 N_SLEEP_c_90_n N_A_459_21#_c_173_n 8.57065e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_88 N_SLEEP_c_91_n N_A_459_21#_c_173_n 0.0243795f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_89 N_SLEEP_c_90_n N_A_27_297#_c_308_n 4.10066e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_90 N_SLEEP_c_92_n N_A_27_297#_c_310_n 0.0151455f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_91 N_SLEEP_c_93_n N_A_27_297#_c_310_n 0.0164876f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_92 N_SLEEP_c_90_n N_A_27_297#_c_310_n 0.0530179f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_93 N_SLEEP_c_91_n N_A_27_297#_c_310_n 0.00953178f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_94 N_SLEEP_c_94_n N_A_27_297#_c_311_n 0.01491f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_95 N_SLEEP_c_95_n N_A_27_297#_c_311_n 0.0111858f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_96 N_SLEEP_c_90_n N_A_27_297#_c_311_n 0.0439319f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_97 N_SLEEP_c_91_n N_A_27_297#_c_311_n 0.00905881f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_98 N_SLEEP_c_95_n N_A_27_297#_c_312_n 0.00359583f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_99 N_SLEEP_c_90_n N_A_27_297#_c_312_n 3.67829e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_100 N_SLEEP_c_91_n N_A_27_297#_c_312_n 3.8543e-19 $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_101 N_SLEEP_c_94_n N_A_27_297#_c_328_n 4.84481e-19 $X=1.455 $Y=1.41 $X2=0
+ $Y2=0
cc_102 N_SLEEP_c_95_n N_A_27_297#_c_328_n 0.0132763f $X=1.925 $Y=1.41 $X2=0
+ $Y2=0
cc_103 N_SLEEP_c_90_n N_A_27_297#_c_315_n 0.0132791f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_104 N_SLEEP_c_91_n N_A_27_297#_c_315_n 0.00435155f $X=1.925 $Y=1.202 $X2=0
+ $Y2=0
cc_105 N_SLEEP_c_92_n N_VPWR_c_397_n 0.0171285f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_106 N_SLEEP_c_93_n N_VPWR_c_397_n 0.0117009f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_107 N_SLEEP_c_94_n N_VPWR_c_397_n 6.2189e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_108 N_SLEEP_c_93_n N_VPWR_c_398_n 6.52114e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_109 N_SLEEP_c_94_n N_VPWR_c_398_n 0.014932f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_110 N_SLEEP_c_95_n N_VPWR_c_398_n 0.00519421f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_111 N_SLEEP_c_92_n N_VPWR_c_401_n 0.00427505f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_112 N_SLEEP_c_93_n N_VPWR_c_402_n 0.00622633f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_113 N_SLEEP_c_94_n N_VPWR_c_402_n 0.00427505f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_114 N_SLEEP_c_95_n N_VPWR_c_403_n 0.00596194f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_115 N_SLEEP_c_92_n N_VPWR_c_396_n 0.00825932f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_116 N_SLEEP_c_93_n N_VPWR_c_396_n 0.0104011f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_117 N_SLEEP_c_94_n N_VPWR_c_396_n 0.00732977f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_118 N_SLEEP_c_95_n N_VPWR_c_396_n 0.0099828f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_119 N_SLEEP_c_86_n N_X_c_479_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_120 N_SLEEP_c_87_n N_X_c_479_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_121 N_SLEEP_c_88_n N_X_c_479_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_122 N_SLEEP_c_87_n N_X_c_468_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_123 N_SLEEP_c_88_n N_X_c_468_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_124 N_SLEEP_c_90_n N_X_c_468_n 0.0397461f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_125 N_SLEEP_c_91_n N_X_c_468_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_126 N_SLEEP_c_86_n N_X_c_469_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_127 N_SLEEP_c_87_n N_X_c_469_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_128 N_SLEEP_c_90_n N_X_c_469_n 0.0306016f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_129 N_SLEEP_c_91_n N_X_c_469_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_130 N_SLEEP_c_87_n N_X_c_490_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_131 N_SLEEP_c_88_n N_X_c_490_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_132 N_SLEEP_c_89_n N_X_c_470_n 0.01152f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_133 N_SLEEP_c_90_n N_X_c_470_n 0.00658691f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_134 N_SLEEP_c_89_n N_X_c_494_n 5.32212e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_135 N_SLEEP_c_90_n N_X_c_471_n 0.0055903f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_136 N_SLEEP_c_91_n N_X_c_471_n 0.0012283f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_137 N_SLEEP_c_88_n N_X_c_473_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_138 N_SLEEP_c_90_n N_X_c_473_n 0.0307352f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_139 N_SLEEP_c_91_n N_X_c_473_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_140 N_SLEEP_c_86_n N_VGND_c_583_n 0.00497314f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_141 N_SLEEP_c_86_n N_VGND_c_584_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_142 N_SLEEP_c_87_n N_VGND_c_584_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_143 N_SLEEP_c_87_n N_VGND_c_585_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_144 N_SLEEP_c_88_n N_VGND_c_585_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_145 N_SLEEP_c_89_n N_VGND_c_586_n 0.00268723f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_146 N_SLEEP_c_88_n N_VGND_c_591_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_147 N_SLEEP_c_89_n N_VGND_c_591_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_148 N_SLEEP_c_86_n N_VGND_c_599_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_149 N_SLEEP_c_87_n N_VGND_c_599_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_150 N_SLEEP_c_88_n N_VGND_c_599_n 0.00608558f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_151 N_SLEEP_c_89_n N_VGND_c_599_n 0.00615622f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_459_21#_c_169_n N_A_c_280_n 0.00508485f $X=4.59 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_153 N_A_459_21#_c_170_n N_A_c_280_n 0.00619296f $X=4.55 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_459_21#_c_171_n N_A_c_280_n 0.00342967f $X=4.59 $Y=0.815 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_459_21#_c_179_n N_A_c_283_n 0.00908916f $X=4.59 $Y=2.34 $X2=0 $Y2=0
cc_156 N_A_459_21#_c_180_n N_A_c_283_n 0.00297076f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_157 N_A_459_21#_c_181_n N_A_c_283_n 0.00367998f $X=4.59 $Y=1.575 $X2=0 $Y2=0
cc_158 N_A_459_21#_c_172_n A 0.0175378f $X=4.55 $Y=1.175 $X2=0 $Y2=0
cc_159 N_A_459_21#_c_181_n A 0.00353171f $X=4.59 $Y=1.575 $X2=0 $Y2=0
cc_160 N_A_459_21#_c_168_n N_A_c_282_n 0.0210908f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_459_21#_c_172_n N_A_c_282_n 0.00166662f $X=4.55 $Y=1.175 $X2=0 $Y2=0
cc_162 N_A_459_21#_c_181_n N_A_c_282_n 0.00406149f $X=4.59 $Y=1.575 $X2=0 $Y2=0
cc_163 N_A_459_21#_c_174_n N_A_27_297#_c_312_n 0.00336534f $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_164 N_A_459_21#_c_173_n N_A_27_297#_c_312_n 3.8543e-19 $X=3.905 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_459_21#_c_174_n N_A_27_297#_c_328_n 0.00892871f $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_166 N_A_459_21#_c_175_n N_A_27_297#_c_328_n 5.45102e-19 $X=2.865 $Y=1.41
+ $X2=0 $Y2=0
cc_167 N_A_459_21#_c_174_n N_A_27_297#_c_336_n 0.0129846f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_459_21#_c_175_n N_A_27_297#_c_336_n 0.0080971f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_169 N_A_459_21#_c_176_n N_A_27_297#_c_338_n 0.010646f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_170 N_A_459_21#_c_177_n N_A_27_297#_c_338_n 0.00955151f $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_171 N_A_459_21#_c_177_n N_A_27_297#_c_313_n 0.00169565f $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_172 N_A_459_21#_c_179_n N_A_27_297#_c_313_n 0.0150382f $X=4.59 $Y=2.34 $X2=0
+ $Y2=0
cc_173 N_A_459_21#_c_176_n N_A_27_297#_c_314_n 5.7646e-19 $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_174 N_A_459_21#_c_177_n N_A_27_297#_c_314_n 0.0127031f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_459_21#_c_210_p N_A_27_297#_c_314_n 0.0202987f $X=4.425 $Y=1.175
+ $X2=0 $Y2=0
cc_176 N_A_459_21#_c_168_n N_A_27_297#_c_314_n 0.00778953f $X=4.38 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_459_21#_c_180_n N_A_27_297#_c_314_n 0.0610922f $X=4.59 $Y=1.66 $X2=0
+ $Y2=0
cc_178 N_A_459_21#_c_174_n N_A_27_297#_c_347_n 6.08324e-19 $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_179 N_A_459_21#_c_175_n N_A_27_297#_c_347_n 0.00957505f $X=2.865 $Y=1.41
+ $X2=0 $Y2=0
cc_180 N_A_459_21#_c_176_n N_A_27_297#_c_347_n 0.00657656f $X=3.335 $Y=1.41
+ $X2=0 $Y2=0
cc_181 N_A_459_21#_c_177_n N_A_27_297#_c_347_n 5.59969e-19 $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_182 N_A_459_21#_c_180_n N_VPWR_c_400_n 0.0575527f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_183 N_A_459_21#_c_181_n N_VPWR_c_400_n 0.00417777f $X=4.59 $Y=1.575 $X2=0
+ $Y2=0
cc_184 N_A_459_21#_c_174_n N_VPWR_c_403_n 0.00429425f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_459_21#_c_175_n N_VPWR_c_403_n 0.00430873f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_459_21#_c_176_n N_VPWR_c_403_n 0.00430943f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_459_21#_c_177_n N_VPWR_c_403_n 0.00429355f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_459_21#_c_179_n N_VPWR_c_403_n 0.0210458f $X=4.59 $Y=2.34 $X2=0 $Y2=0
cc_189 N_A_459_21#_M1010_s N_VPWR_c_396_n 0.00225715f $X=4.455 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_459_21#_c_174_n N_VPWR_c_396_n 0.00609019f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_459_21#_c_175_n N_VPWR_c_396_n 0.00605584f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_459_21#_c_176_n N_VPWR_c_396_n 0.0060559f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_459_21#_c_177_n N_VPWR_c_396_n 0.00734727f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_459_21#_c_179_n N_VPWR_c_396_n 0.0124725f $X=4.59 $Y=2.34 $X2=0 $Y2=0
cc_195 N_A_459_21#_c_164_n N_X_c_470_n 0.0117455f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_459_21#_c_164_n N_X_c_494_n 0.00644736f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_459_21#_c_165_n N_X_c_494_n 0.00686626f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_459_21#_c_166_n N_X_c_494_n 5.45498e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_199 N_A_459_21#_c_164_n N_X_c_471_n 0.00232392f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_459_21#_c_174_n N_X_c_471_n 9.2652e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_459_21#_c_165_n N_X_c_471_n 0.00309297f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_459_21#_c_175_n N_X_c_471_n 0.00112479f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_459_21#_c_166_n N_X_c_471_n 4.96717e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_459_21#_c_210_p N_X_c_471_n 0.0128469f $X=4.425 $Y=1.175 $X2=0 $Y2=0
cc_205 N_A_459_21#_c_173_n N_X_c_471_n 0.0402787f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_459_21#_c_165_n N_X_c_472_n 0.00499466f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_459_21#_c_166_n N_X_c_472_n 0.010179f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_459_21#_c_167_n N_X_c_472_n 2.15189e-19 $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_209 N_A_459_21#_c_210_p N_X_c_472_n 0.0491542f $X=4.425 $Y=1.175 $X2=0 $Y2=0
cc_210 N_A_459_21#_c_173_n N_X_c_472_n 0.00872135f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_459_21#_c_165_n N_X_c_516_n 5.24597e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_459_21#_c_166_n N_X_c_516_n 0.00651696f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_459_21#_c_177_n N_X_c_476_n 0.00437462f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_459_21#_c_210_p N_X_c_476_n 0.0138618f $X=4.425 $Y=1.175 $X2=0 $Y2=0
cc_215 N_A_459_21#_c_173_n N_X_c_476_n 0.00419992f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_459_21#_c_164_n N_X_c_474_n 0.00224457f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_217 N_A_459_21#_c_165_n N_X_c_474_n 0.00412844f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_459_21#_c_173_n N_X_c_474_n 4.78733e-19 $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_459_21#_c_174_n N_X_c_477_n 0.00184921f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_459_21#_c_175_n N_X_c_477_n 0.00588782f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_459_21#_c_175_n N_X_c_478_n 0.00905398f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_459_21#_c_176_n N_X_c_478_n 0.0160369f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_459_21#_c_210_p N_X_c_478_n 0.0287801f $X=4.425 $Y=1.175 $X2=0 $Y2=0
cc_224 N_A_459_21#_c_173_n N_X_c_478_n 0.0100381f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_225 N_A_459_21#_c_164_n N_VGND_c_586_n 0.00268723f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_459_21#_c_165_n N_VGND_c_587_n 0.00379224f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_459_21#_c_166_n N_VGND_c_587_n 0.00276126f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_228 N_A_459_21#_c_167_n N_VGND_c_588_n 0.00499982f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_229 N_A_459_21#_c_210_p N_VGND_c_588_n 0.0234825f $X=4.425 $Y=1.175 $X2=0
+ $Y2=0
cc_230 N_A_459_21#_c_168_n N_VGND_c_588_n 0.00739466f $X=4.38 $Y=1.16 $X2=0
+ $Y2=0
cc_231 N_A_459_21#_c_169_n N_VGND_c_588_n 0.0512575f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_232 N_A_459_21#_c_169_n N_VGND_c_590_n 0.0352721f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_233 N_A_459_21#_c_170_n N_VGND_c_590_n 0.00287218f $X=4.55 $Y=1.075 $X2=0
+ $Y2=0
cc_234 N_A_459_21#_c_164_n N_VGND_c_593_n 0.00423334f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_235 N_A_459_21#_c_165_n N_VGND_c_593_n 0.00423261f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_236 N_A_459_21#_c_166_n N_VGND_c_595_n 0.00423334f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_237 N_A_459_21#_c_167_n N_VGND_c_595_n 0.00585385f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_238 N_A_459_21#_c_169_n N_VGND_c_597_n 0.020984f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_239 N_A_459_21#_M1011_s N_VGND_c_599_n 0.00225715f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_240 N_A_459_21#_c_164_n N_VGND_c_599_n 0.00587047f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_459_21#_c_165_n N_VGND_c_599_n 0.00609168f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_242 N_A_459_21#_c_166_n N_VGND_c_599_n 0.00608558f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_459_21#_c_167_n N_VGND_c_599_n 0.0121055f $X=3.83 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_459_21#_c_169_n N_VGND_c_599_n 0.0124119f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_245 N_A_c_283_n N_VPWR_c_400_n 0.00923983f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_246 A N_VPWR_c_400_n 0.032799f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_247 N_A_c_282_n N_VPWR_c_400_n 0.0058213f $X=4.825 $Y=1.202 $X2=0 $Y2=0
cc_248 N_A_c_283_n N_VPWR_c_403_n 0.00673617f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A_c_283_n N_VPWR_c_396_n 0.0141776f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_c_280_n N_VGND_c_588_n 0.0023653f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_c_280_n N_VGND_c_590_n 0.00734095f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_252 A N_VGND_c_590_n 0.0239559f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_253 N_A_c_282_n N_VGND_c_590_n 0.0063933f $X=4.825 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_c_280_n N_VGND_c_597_n 0.00541359f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_c_280_n N_VGND_c_599_n 0.0120732f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_27_297#_c_310_n N_VPWR_M1001_d 0.00188315f $X=1.135 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_257 N_A_27_297#_c_311_n N_VPWR_M1006_d 0.00184035f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_258 N_A_27_297#_c_309_n N_VPWR_c_397_n 0.0488071f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_259 N_A_27_297#_c_310_n N_VPWR_c_397_n 0.0212439f $X=1.135 $Y=1.56 $X2=0
+ $Y2=0
cc_260 N_A_27_297#_c_355_p N_VPWR_c_397_n 0.0385613f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_261 N_A_27_297#_c_355_p N_VPWR_c_398_n 0.0461742f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_262 N_A_27_297#_c_311_n N_VPWR_c_398_n 0.0194872f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_c_328_n N_VPWR_c_398_n 0.0496968f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_c_309_n N_VPWR_c_401_n 0.0196165f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_265 N_A_27_297#_c_355_p N_VPWR_c_402_n 0.0118139f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_328_n N_VPWR_c_403_n 0.0224921f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_267 N_A_27_297#_c_336_n N_VPWR_c_403_n 0.0317606f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_c_338_n N_VPWR_c_403_n 0.0317606f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_c_313_n N_VPWR_c_403_n 0.0281657f $X=4.04 $Y=2.295 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_c_347_n N_VPWR_c_403_n 0.0220286f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_271 N_A_27_297#_M1001_s N_VPWR_c_396_n 0.00442207f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_272 N_A_27_297#_M1003_s N_VPWR_c_396_n 0.00647849f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_273 N_A_27_297#_M1012_s N_VPWR_c_396_n 0.00231261f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_274 N_A_27_297#_M1009_s N_VPWR_c_396_n 0.00231261f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_M1017_s N_VPWR_c_396_n 0.00233913f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_309_n N_VPWR_c_396_n 0.0107063f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_277 N_A_27_297#_c_355_p N_VPWR_c_396_n 0.00646998f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_328_n N_VPWR_c_396_n 0.014078f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_279 N_A_27_297#_c_336_n N_VPWR_c_396_n 0.0196262f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_338_n N_VPWR_c_396_n 0.0196262f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_c_313_n N_VPWR_c_396_n 0.0161675f $X=4.04 $Y=2.295 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_347_n N_VPWR_c_396_n 0.0139179f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_283 N_A_27_297#_c_336_n N_X_M1000_d 0.0034107f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_338_n N_X_M1014_d 0.0034107f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_285 N_A_27_297#_c_312_n N_X_c_470_n 0.0132538f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_286 N_A_27_297#_c_328_n N_X_c_533_n 0.0232292f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_287 N_A_27_297#_c_336_n N_X_c_533_n 0.0128008f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_347_n N_X_c_533_n 0.0141845f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_289 N_A_27_297#_c_314_n N_X_c_476_n 0.0143033f $X=4.04 $Y=1.66 $X2=0 $Y2=0
cc_290 N_A_27_297#_c_338_n N_X_c_537_n 0.0128008f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_291 N_A_27_297#_c_314_n N_X_c_537_n 0.0286107f $X=4.04 $Y=1.66 $X2=0 $Y2=0
cc_292 N_A_27_297#_c_347_n N_X_c_537_n 0.0116296f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_293 N_A_27_297#_c_312_n N_X_c_477_n 0.0150774f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_294 N_A_27_297#_c_328_n N_X_c_477_n 0.00543755f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_295 N_A_27_297#_c_336_n N_X_c_477_n 0.00296569f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_296 N_A_27_297#_M1009_s N_X_c_478_n 0.00199621f $X=2.955 $Y=1.485 $X2=0 $Y2=0
cc_297 N_A_27_297#_c_336_n N_X_c_478_n 2.56171e-19 $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_298 N_A_27_297#_c_338_n N_X_c_478_n 0.00435577f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_299 N_A_27_297#_c_347_n N_X_c_478_n 0.0196167f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_300 N_A_27_297#_c_308_n N_VGND_c_583_n 0.0113923f $X=0.225 $Y=1.665 $X2=0
+ $Y2=0
cc_301 N_VPWR_c_396_n N_X_M1000_d 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_396_n N_X_M1014_d 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_303 N_X_c_468_n N_VGND_M1007_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_304 N_X_c_470_n N_VGND_M1015_d 0.00162089f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_305 N_X_c_472_n N_VGND_M1005_s 0.00251047f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_306 N_X_c_469_n N_VGND_c_583_n 0.00835667f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_307 N_X_c_479_n N_VGND_c_584_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_308 N_X_c_468_n N_VGND_c_584_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_309 N_X_c_479_n N_VGND_c_585_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_310 N_X_c_468_n N_VGND_c_585_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_311 N_X_c_470_n N_VGND_c_586_n 0.0122559f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_312 N_X_c_494_n N_VGND_c_587_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_313 N_X_c_472_n N_VGND_c_587_n 0.0127273f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_314 N_X_c_472_n N_VGND_c_588_n 0.00138734f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_315 N_X_c_468_n N_VGND_c_591_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_316 N_X_c_490_n N_VGND_c_591_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_317 N_X_c_470_n N_VGND_c_591_n 0.00254521f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_318 N_X_c_470_n N_VGND_c_593_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_319 N_X_c_494_n N_VGND_c_593_n 0.0224037f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_320 N_X_c_472_n N_VGND_c_593_n 0.00159127f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_321 N_X_c_474_n N_VGND_c_593_n 0.00118043f $X=2.645 $Y=0.815 $X2=0 $Y2=0
cc_322 N_X_c_472_n N_VGND_c_595_n 0.00198695f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_323 N_X_c_516_n N_VGND_c_595_n 0.0231806f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_324 N_X_M1002_s N_VGND_c_599_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_325 N_X_M1008_s N_VGND_c_599_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_326 N_X_M1004_d N_VGND_c_599_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_327 N_X_M1013_d N_VGND_c_599_n 0.00364931f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_328 N_X_c_479_n N_VGND_c_599_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_329 N_X_c_468_n N_VGND_c_599_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_330 N_X_c_490_n N_VGND_c_599_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_331 N_X_c_470_n N_VGND_c_599_n 0.0094839f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_332 N_X_c_494_n N_VGND_c_599_n 0.0141415f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_333 N_X_c_472_n N_VGND_c_599_n 0.00800459f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_334 N_X_c_516_n N_VGND_c_599_n 0.0143352f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_335 N_X_c_474_n N_VGND_c_599_n 0.001841f $X=2.645 $Y=0.815 $X2=0 $Y2=0
