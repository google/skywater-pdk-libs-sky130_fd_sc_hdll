# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__and4b_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__and4b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.135000 0.740000 0.335000 1.630000 ;
    END
  END A_N
  PIN B
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.895000 0.420000 2.155000 1.745000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.375000 0.420000 2.615000 1.615000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 0.645000 3.115000 1.615000 ;
    END
  END D
  PIN VGND
    ANTENNADIFFAREA  0.539650 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.095000  0.085000 0.425000 0.465000 ;
        RECT 3.010000  0.085000 3.390000 0.465000 ;
        RECT 4.065000  0.085000 4.450000 0.465000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.856300 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.515000 2.195000 0.895000 2.635000 ;
        RECT 1.705000 2.255000 2.425000 2.635000 ;
        RECT 3.140000 2.195000 3.470000 2.635000 ;
        RECT 4.195000 1.835000 4.450000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.555750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.560000 0.255000 3.895000 0.640000 ;
        RECT 3.560000 0.640000 4.455000 0.825000 ;
        RECT 3.690000 1.535000 4.455000 1.665000 ;
        RECT 3.690000 1.665000 3.995000 2.465000 ;
        RECT 3.775000 0.825000 4.455000 1.535000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.175000 1.830000 0.855000 2.000000 ;
      RECT 0.175000 2.000000 0.345000 2.465000 ;
      RECT 0.645000 0.255000 0.855000 0.585000 ;
      RECT 0.685000 0.585000 0.855000 0.995000 ;
      RECT 0.685000 0.995000 1.075000 1.325000 ;
      RECT 0.685000 1.325000 0.855000 1.830000 ;
      RECT 1.115000 1.660000 1.415000 1.915000 ;
      RECT 1.115000 1.915000 3.465000 1.965000 ;
      RECT 1.115000 1.965000 2.860000 2.085000 ;
      RECT 1.115000 2.085000 1.285000 2.465000 ;
      RECT 1.195000 0.255000 1.415000 0.585000 ;
      RECT 1.245000 0.585000 1.415000 1.660000 ;
      RECT 2.670000 2.085000 2.860000 2.465000 ;
      RECT 2.690000 1.795000 3.465000 1.915000 ;
      RECT 3.295000 0.995000 3.555000 1.325000 ;
      RECT 3.295000 1.325000 3.465000 1.795000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__and4b_2
