* File: sky130_fd_sc_hdll__ebufn_4.spice
* Created: Thu Aug 27 19:07:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__ebufn_4.pex.spice"
.subckt sky130_fd_sc_hdll__ebufn_4  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_27_47#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.138125 AS=0.169 PD=1.075 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1009 N_A_224_47#_M1009_d N_TE_B_M1009_g N_VGND_M1018_d VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.138125 PD=1.92 PS=1.075 NRD=8.304 NRS=18.456 M=1
+ R=4.33333 SA=75000.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_413_47#_M1002_d N_A_224_47#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.12025 PD=1.92 PS=1.02 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_413_47#_M1006_d N_A_224_47#_M1006_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.8 SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1014 N_A_413_47#_M1006_d N_A_224_47#_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75002.7 A=0.0975 P=1.6 MULT=1
MM1015 N_A_413_47#_M1015_d N_A_224_47#_M1015_g N_VGND_M1014_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12675 AS=0.104 PD=1.04 PS=0.97 NRD=10.152 NRS=8.304 M=1 R=4.33333
+ SA=75001.7 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1001 N_Z_M1001_d N_A_27_47#_M1001_g N_A_413_47#_M1015_d VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.12675 PD=0.97 PS=1.04 NRD=8.304 NRS=10.152 M=1 R=4.33333
+ SA=75002.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1003 N_Z_M1001_d N_A_27_47#_M1003_g N_A_413_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75002.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1010 N_Z_M1010_d N_A_27_47#_M1010_g N_A_413_47#_M1003_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_Z_M1010_d N_A_27_47#_M1019_g N_A_413_47#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.182 PD=1.02 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_A_27_47#_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1975 AS=0.27 PD=1.395 PS=2.54 NRD=8.8453 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1017 N_A_224_47#_M1017_d N_TE_B_M1017_g N_VPWR_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.1975 PD=2.54 PS=1.395 NRD=0.9653 NRS=13.7703 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_340_309#_M1005_d N_TE_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.2538 AS=0.1363 PD=2.42 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.2 SB=90004 A=0.1692 P=2.24 MULT=1
MM1008 N_A_340_309#_M1008_d N_TE_B_M1008_g N_VPWR_M1005_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90000.6 SB=90003.6 A=0.1692 P=2.24 MULT=1
MM1012 N_A_340_309#_M1008_d N_TE_B_M1012_g N_VPWR_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.1363 AS=0.1363 PD=1.23 PS=1.23 NRD=1.0441 NRS=1.0441 M=1 R=5.22222
+ SA=90001.1 SB=90003.1 A=0.1692 P=2.24 MULT=1
MM1016 N_A_340_309#_M1016_d N_TE_B_M1016_g N_VPWR_M1012_s VPB PHIGHVT L=0.18
+ W=0.94 AD=0.397271 AS=0.1363 PD=1.76856 PS=1.23 NRD=19.897 NRS=1.0441 M=1
+ R=5.22222 SA=90001.6 SB=90002.6 A=0.1692 P=2.24 MULT=1
MM1000 N_A_340_309#_M1016_d N_A_27_47#_M1000_g N_Z_M1000_s VPB PHIGHVT L=0.18
+ W=1 AD=0.422629 AS=0.145 PD=1.88144 PS=1.29 NRD=11.8003 NRS=0.9653 M=1
+ R=5.55556 SA=90002.5 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1004 N_A_340_309#_M1004_d N_A_27_47#_M1004_g N_Z_M1000_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.9 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 N_A_340_309#_M1004_d N_A_27_47#_M1011_g N_Z_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.4 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1013 N_A_340_309#_M1013_d N_A_27_47#_M1013_g N_Z_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
*
.include "sky130_fd_sc_hdll__ebufn_4.pxi.spice"
*
.ends
*
*
