* File: sky130_fd_sc_hdll__and3b_2.pex.spice
* Created: Thu Aug 27 18:58:25 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%A_N 1 3 6 8 9
r24 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r25 8 9 13.4814 $w=2.63e-07 $l=3.1e-07 $layer=LI1_cond $X=0.277 $Y=0.85
+ $X2=0.277 $Y2=1.16
r26 4 13 39.4323 $w=3.92e-07 $l=2.38642e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.35 $Y2=1.16
r27 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r28 1 13 53.5809 $w=3.92e-07 $l=3.85746e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.35 $Y2=1.16
r29 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.48
+ $X2=0.495 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%A_117_311# 1 2 7 9 12 16 20 24 27
r41 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.27
+ $Y=1.16 $X2=1.27 $Y2=1.16
r42 22 27 1.99325 $w=2.3e-07 $l=1.38e-07 $layer=LI1_cond $X=0.905 $Y=1.13
+ $X2=0.767 $Y2=1.13
r43 22 24 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.905 $Y=1.13
+ $X2=1.27 $Y2=1.13
r44 18 27 4.44123 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=0.767 $Y=1.245
+ $X2=0.767 $Y2=1.13
r45 18 20 20.744 $w=2.73e-07 $l=4.95e-07 $layer=LI1_cond $X=0.767 $Y=1.245
+ $X2=0.767 $Y2=1.74
r46 14 27 4.44123 $w=2.75e-07 $l=1.15e-07 $layer=LI1_cond $X=0.767 $Y=1.015
+ $X2=0.767 $Y2=1.13
r47 14 16 22.8393 $w=2.73e-07 $l=5.45e-07 $layer=LI1_cond $X=0.767 $Y=1.015
+ $X2=0.767 $Y2=0.47
r48 10 25 39.0558 $w=3.7e-07 $l=2.2798e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.36 $Y2=1.16
r49 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.475
r50 7 25 54.4254 $w=3.7e-07 $l=3.77359e-07 $layer=POLY_cond $X=1.485 $Y=1.48
+ $X2=1.36 $Y2=1.16
r51 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.48
+ $X2=1.485 $Y2=1.765
r52 2 20 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.555 $X2=0.73 $Y2=1.74
r53 1 16 182 $w=1.7e-07 $l=2.71662e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=0.75 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%B 1 2 4 7 10 19
c40 2 0 1.704e-19 $X=1.955 $Y=2.105
r41 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=2.3
+ $X2=2 $Y2=2.3
r42 10 19 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=2.09 $Y=2.295
+ $X2=2.095 $Y2=2.295
r43 10 14 3.05058 $w=3.38e-07 $l=9e-08 $layer=LI1_cond $X=2.09 $Y=2.295 $X2=2
+ $Y2=2.295
r44 7 9 371.755 $w=1.5e-07 $l=7.25e-07 $layer=POLY_cond $X=1.98 $Y=0.475
+ $X2=1.98 $Y2=1.2
r45 2 13 38.5229 $w=3.2e-07 $l=2.25167e-07 $layer=POLY_cond $X=1.955 $Y=2.105
+ $X2=2.02 $Y2=2.3
r46 2 4 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.955 $Y=2.105
+ $X2=1.955 $Y2=1.765
r47 1 9 110.989 $w=1.8e-07 $l=2.8e-07 $layer=POLY_cond $X=1.955 $Y=1.48
+ $X2=1.955 $Y2=1.2
r48 1 4 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.955 $Y=1.48
+ $X2=1.955 $Y2=1.765
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%C 3 5 7 8 9 15 21
r45 15 24 5.55678 $w=4.78e-07 $l=2.23e-07 $layer=LI1_cond $X=2.4 $Y=1.005
+ $X2=2.177 $Y2=1.005
r46 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.16 $X2=2.4 $Y2=1.16
r47 8 24 1.91871 $w=4.78e-07 $l=7.7e-08 $layer=LI1_cond $X=2.1 $Y=1.005
+ $X2=2.177 $Y2=1.005
r48 8 24 2.04398 $w=3.85e-07 $l=2.4e-07 $layer=LI1_cond $X=2.177 $Y=0.765
+ $X2=2.177 $Y2=1.005
r49 8 21 0.124591 $w=4.78e-07 $l=5e-09 $layer=LI1_cond $X=2.1 $Y=1.005 $X2=2.095
+ $Y2=1.005
r50 8 9 6.62929 $w=5.53e-07 $l=2.55e-07 $layer=LI1_cond $X=2.177 $Y=0.765
+ $X2=2.177 $Y2=0.51
r51 5 14 48.3784 $w=2.91e-07 $l=2.77489e-07 $layer=POLY_cond $X=2.48 $Y=1.41
+ $X2=2.422 $Y2=1.16
r52 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.48 $Y=1.41 $X2=2.48
+ $Y2=1.695
r53 1 14 38.6072 $w=2.91e-07 $l=2.01879e-07 $layer=POLY_cond $X=2.34 $Y=0.995
+ $X2=2.422 $Y2=1.16
r54 1 3 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.34 $Y=0.995 $X2=2.34
+ $Y2=0.475
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%A_225_311# 1 2 3 10 12 13 15 16 18 19 21
+ 24 26 30 31 33 34 38 40 44 47 48 52
c106 38 0 1.704e-19 $X=2.245 $Y=1.725
c107 30 0 1.27873e-19 $X=1.645 $Y=1.51
r108 52 53 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.485 $Y=1.202
+ $X2=3.51 $Y2=1.202
r109 51 52 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=3.04 $Y=1.202
+ $X2=3.485 $Y2=1.202
r110 50 51 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.015 $Y=1.202
+ $X2=3.04 $Y2=1.202
r111 45 50 10.3378 $w=3.73e-07 $l=8e-08 $layer=POLY_cond $X=2.935 $Y=1.202
+ $X2=3.015 $Y2=1.202
r112 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.935
+ $Y=1.16 $X2=2.935 $Y2=1.16
r113 42 44 13.2781 $w=2.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.905 $Y=1.425
+ $X2=2.905 $Y2=1.16
r114 41 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.35 $Y=1.51
+ $X2=2.255 $Y2=1.51
r115 40 42 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=2.79 $Y=1.51
+ $X2=2.905 $Y2=1.425
r116 40 41 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=2.79 $Y=1.51
+ $X2=2.35 $Y2=1.51
r117 36 48 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=1.595
+ $X2=2.255 $Y2=1.51
r118 36 38 7.58852 $w=1.88e-07 $l=1.3e-07 $layer=LI1_cond $X=2.255 $Y=1.595
+ $X2=2.255 $Y2=1.725
r119 35 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=1.51
+ $X2=1.73 $Y2=1.51
r120 34 48 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.16 $Y=1.51
+ $X2=2.255 $Y2=1.51
r121 34 35 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.16 $Y=1.51
+ $X2=1.815 $Y2=1.51
r122 33 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=1.425
+ $X2=1.73 $Y2=1.51
r123 32 33 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.73 $Y=0.57
+ $X2=1.73 $Y2=1.425
r124 30 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.51
+ $X2=1.73 $Y2=1.51
r125 30 31 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.645 $Y=1.51
+ $X2=1.335 $Y2=1.51
r126 26 32 7.24806 $w=2.65e-07 $l=1.70276e-07 $layer=LI1_cond $X=1.645 $Y=0.437
+ $X2=1.73 $Y2=0.57
r127 26 28 16.3082 $w=2.63e-07 $l=3.75e-07 $layer=LI1_cond $X=1.645 $Y=0.437
+ $X2=1.27 $Y2=0.437
r128 22 31 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=1.217 $Y=1.595
+ $X2=1.335 $Y2=1.51
r129 22 24 8.09162 $w=2.33e-07 $l=1.65e-07 $layer=LI1_cond $X=1.217 $Y=1.595
+ $X2=1.217 $Y2=1.76
r130 19 53 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=1.202
r131 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r132 16 52 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.202
r133 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.985
r134 13 51 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.04 $Y=0.995
+ $X2=3.04 $Y2=1.202
r135 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.04 $Y=0.995
+ $X2=3.04 $Y2=0.56
r136 10 50 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.202
r137 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.015 $Y=1.41
+ $X2=3.015 $Y2=1.985
r138 3 38 600 $w=1.7e-07 $l=2.72029e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.555 $X2=2.245 $Y2=1.725
r139 2 24 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.555 $X2=1.25 $Y2=1.76
r140 1 28 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=1.145
+ $Y=0.265 $X2=1.27 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%VPWR 1 2 3 4 13 15 17 23 25 27 32 35 36 37
+ 43 51 59
c58 2 0 1.27873e-19 $X=1.575 $Y=1.555
r59 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 53 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 46 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r62 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 43 58 4.13553 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.76 $Y=2.72 $X2=3.95
+ $Y2=2.72
r64 43 45 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=2.72
+ $X2=3.45 $Y2=2.72
r65 42 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r66 42 55 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r68 39 41 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=1.745 $Y=2.72
+ $X2=2.53 $Y2=2.72
r69 37 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r70 37 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 35 41 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=2.66 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 35 36 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.66 $Y=2.72
+ $X2=2.767 $Y2=2.72
r73 34 45 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=3.45 $Y2=2.72
r74 34 36 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=2.875 $Y=2.72
+ $X2=2.767 $Y2=2.72
r75 25 58 3.11253 $w=2.65e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.95 $Y2=2.72
r76 25 27 29.3547 $w=2.63e-07 $l=6.75e-07 $layer=LI1_cond $X=3.892 $Y=2.635
+ $X2=3.892 $Y2=1.96
r77 21 36 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.767 $Y=2.635
+ $X2=2.767 $Y2=2.72
r78 21 23 36.4494 $w=2.13e-07 $l=6.8e-07 $layer=LI1_cond $X=2.767 $Y=2.635
+ $X2=2.767 $Y2=1.955
r79 19 32 5.54545 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=1.625 $Y=1.86
+ $X2=1.72 $Y2=1.86
r80 19 51 8.40323 $w=2.38e-07 $l=1.75e-07 $layer=LI1_cond $X=1.625 $Y=1.955
+ $X2=1.625 $Y2=2.13
r81 18 48 4.67309 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r82 17 39 8.98481 $w=1.7e-07 $l=3.33e-07 $layer=LI1_cond $X=1.412 $Y=2.72
+ $X2=1.745 $Y2=2.72
r83 17 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r84 17 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r85 17 51 15.7657 $w=6.63e-07 $l=5.9e-07 $layer=LI1_cond $X=1.412 $Y=2.72
+ $X2=1.412 $Y2=2.13
r86 17 18 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.08 $Y=2.72 $X2=0.4
+ $Y2=2.72
r87 13 48 2.96741 $w=3.15e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.2 $Y2=2.72
r88 13 15 32.744 $w=3.13e-07 $l=8.95e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.74
r89 4 27 300 $w=1.7e-07 $l=5.96867e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.485 $X2=3.85 $Y2=1.96
r90 3 23 300 $w=1.7e-07 $l=5.65332e-07 $layer=licon1_PDIFF $count=2 $X=2.57
+ $Y=1.485 $X2=2.78 $Y2=1.955
r91 2 32 600 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.555 $X2=1.72 $Y2=1.85
r92 1 15 600 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.555 $X2=0.26 $Y2=1.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%X 1 2 8 11 12 13 24 25 33
r33 31 33 7.36048 $w=5.18e-07 $l=3.2e-07 $layer=LI1_cond $X=3.415 $Y=1.185
+ $X2=3.735 $Y2=1.185
r34 29 31 0.230015 $w=5.18e-07 $l=1e-08 $layer=LI1_cond $X=3.405 $Y=1.185
+ $X2=3.415 $Y2=1.185
r35 24 25 5.00312 $w=4.63e-07 $l=1.65e-07 $layer=LI1_cond $X=3.357 $Y=1.96
+ $X2=3.357 $Y2=1.795
r36 21 22 5.69342 $w=4.03e-07 $l=1.85e-07 $layer=LI1_cond $X=3.367 $Y=0.53
+ $X2=3.367 $Y2=0.715
r37 13 33 3.91026 $w=5.18e-07 $l=1.7e-07 $layer=LI1_cond $X=3.905 $Y=1.185
+ $X2=3.735 $Y2=1.185
r38 12 24 6.43053 $w=4.63e-07 $l=2.5e-07 $layer=LI1_cond $X=3.357 $Y=2.21
+ $X2=3.357 $Y2=1.96
r39 11 21 0.569108 $w=4.03e-07 $l=2e-08 $layer=LI1_cond $X=3.367 $Y=0.51
+ $X2=3.367 $Y2=0.53
r40 9 31 3.05479 $w=3.5e-07 $l=2.6e-07 $layer=LI1_cond $X=3.415 $Y=1.445
+ $X2=3.415 $Y2=1.185
r41 9 25 11.5244 $w=3.48e-07 $l=3.5e-07 $layer=LI1_cond $X=3.415 $Y=1.445
+ $X2=3.415 $Y2=1.795
r42 8 29 3.39791 $w=3.3e-07 $l=2.6e-07 $layer=LI1_cond $X=3.405 $Y=0.925
+ $X2=3.405 $Y2=1.185
r43 8 22 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=3.405 $Y=0.925
+ $X2=3.405 $Y2=0.715
r44 2 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.105
+ $Y=1.485 $X2=3.25 $Y2=1.96
r45 1 21 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=3.115
+ $Y=0.235 $X2=3.25 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND3B_2%VGND 1 2 3 10 12 16 18 20 23 24 25 34 43
r46 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r47 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r48 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r49 34 42 4.13553 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.95
+ $Y2=0
r50 34 36 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=3.76 $Y=0 $X2=3.45
+ $Y2=0
r51 33 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r52 32 33 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r53 30 33 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r54 29 32 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r55 29 30 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 27 39 4.2375 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.177
+ $Y2=0
r57 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.69
+ $Y2=0
r58 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r59 25 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r60 23 32 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=2.61 $Y=0 $X2=2.53
+ $Y2=0
r61 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.61 $Y=0 $X2=2.775
+ $Y2=0
r62 22 36 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=3.45
+ $Y2=0
r63 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.775
+ $Y2=0
r64 18 42 3.11253 $w=2.65e-07 $l=1.1025e-07 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.95 $Y2=0
r65 18 20 18.7 $w=2.63e-07 $l=4.3e-07 $layer=LI1_cond $X=3.892 $Y=0.085
+ $X2=3.892 $Y2=0.515
r66 14 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.775 $Y=0.085
+ $X2=2.775 $Y2=0
r67 14 16 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.775 $Y=0.085
+ $X2=2.775 $Y2=0.495
r68 10 39 3.04719 $w=2.7e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.177 $Y2=0
r69 10 12 13.872 $w=2.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.22 $Y=0.085
+ $X2=0.22 $Y2=0.41
r70 3 20 182 $w=1.7e-07 $l=3.90641e-07 $layer=licon1_NDIFF $count=1 $X=3.585
+ $Y=0.235 $X2=3.85 $Y2=0.515
r71 2 16 182 $w=1.7e-07 $l=4.60869e-07 $layer=licon1_NDIFF $count=1 $X=2.415
+ $Y=0.265 $X2=2.775 $Y2=0.495
r72 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.41
.ends

