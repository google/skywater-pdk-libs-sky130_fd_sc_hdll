* File: sky130_fd_sc_hdll__nor4bb_1.pxi.spice
* Created: Thu Aug 27 19:17:49 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%C_N N_C_N_c_75_n N_C_N_c_76_n N_C_N_M1008_g
+ N_C_N_M1000_g C_N C_N N_C_N_c_72_n N_C_N_c_73_n N_C_N_c_74_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_1%C_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%D_N N_D_N_c_106_n N_D_N_M1002_g N_D_N_c_107_n
+ N_D_N_M1009_g D_N D_N PM_SKY130_FD_SC_HDLL__NOR4BB_1%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_216_93# N_A_216_93#_M1002_d
+ N_A_216_93#_M1009_d N_A_216_93#_c_142_n N_A_216_93#_M1005_g
+ N_A_216_93#_c_136_n N_A_216_93#_M1003_g N_A_216_93#_c_137_n
+ N_A_216_93#_c_138_n N_A_216_93#_c_145_n N_A_216_93#_c_139_n
+ N_A_216_93#_c_140_n N_A_216_93#_c_141_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_216_93#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_27_410# N_A_27_410#_M1000_s
+ N_A_27_410#_M1008_s N_A_27_410#_c_196_n N_A_27_410#_M1011_g
+ N_A_27_410#_c_197_n N_A_27_410#_M1006_g N_A_27_410#_c_198_n
+ N_A_27_410#_c_203_n N_A_27_410#_c_204_n N_A_27_410#_c_205_n
+ N_A_27_410#_c_206_n N_A_27_410#_c_207_n N_A_27_410#_c_199_n
+ N_A_27_410#_c_200_n N_A_27_410#_c_209_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_1%A_27_410#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%B N_B_c_273_n N_B_M1010_g N_B_c_274_n
+ N_B_M1001_g B N_B_c_275_n PM_SKY130_FD_SC_HDLL__NOR4BB_1%B
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%A N_A_c_301_n N_A_M1004_g N_A_c_302_n
+ N_A_M1007_g A PM_SKY130_FD_SC_HDLL__NOR4BB_1%A
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%VPWR N_VPWR_M1008_d N_VPWR_M1007_d
+ N_VPWR_c_322_n N_VPWR_c_323_n N_VPWR_c_324_n VPWR N_VPWR_c_325_n
+ N_VPWR_c_326_n N_VPWR_c_327_n N_VPWR_c_321_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%Y N_Y_M1003_d N_Y_M1001_d N_Y_M1005_s
+ N_Y_c_367_n N_Y_c_366_n N_Y_c_401_p N_Y_c_390_n N_Y_c_380_n Y
+ PM_SKY130_FD_SC_HDLL__NOR4BB_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR4BB_1%VGND N_VGND_M1000_d N_VGND_M1003_s
+ N_VGND_M1006_d N_VGND_M1004_d N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n
+ N_VGND_c_424_n N_VGND_c_425_n N_VGND_c_426_n N_VGND_c_427_n N_VGND_c_428_n
+ N_VGND_c_429_n N_VGND_c_430_n N_VGND_c_431_n VGND N_VGND_c_432_n
+ N_VGND_c_433_n VGND PM_SKY130_FD_SC_HDLL__NOR4BB_1%VGND
cc_1 VNB N_C_N_c_72_n 0.0241133f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_2 VNB N_C_N_c_73_n 0.00809375f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_3 VNB N_C_N_c_74_n 0.0208834f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=0.995
cc_4 VNB N_D_N_c_106_n 0.0194283f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_5 VNB N_D_N_c_107_n 0.0263977f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_6 VNB D_N 0.00339436f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_7 VNB N_A_216_93#_c_136_n 0.0200732f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_8 VNB N_A_216_93#_c_137_n 0.0283765f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_9 VNB N_A_216_93#_c_138_n 0.0116018f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_10 VNB N_A_216_93#_c_139_n 0.0118762f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_216_93#_c_140_n 0.0029106f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_216_93#_c_141_n 0.00201956f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_410#_c_196_n 0.0209242f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_14 VNB N_A_27_410#_c_197_n 0.0177203f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_15 VNB N_A_27_410#_c_198_n 0.0224941f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_16 VNB N_A_27_410#_c_199_n 0.00282949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_410#_c_200_n 0.0187907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B_c_273_n 0.0200131f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_19 VNB N_B_c_274_n 0.0173702f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_20 VNB N_B_c_275_n 0.00568771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_c_301_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_22 VNB N_A_c_302_n 0.024698f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_23 VNB A 0.0148243f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=0.675
cc_24 VNB N_VPWR_c_321_n 0.17485f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_Y_c_366_n 0.0040131f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_26 VNB N_VGND_c_421_n 0.0151242f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_27 VNB N_VGND_c_422_n 0.0112341f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_423_n 0.0022216f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_424_n 0.0149757f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_425_n 0.0351548f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_426_n 0.0225278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_427_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_428_n 0.0213827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_429_n 0.00631534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_430_n 0.0156907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_431_n 0.00519124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_432_n 0.0150439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_433_n 0.245086f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_C_N_c_75_n 0.0336761f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.875
cc_40 VPB N_C_N_c_76_n 0.0283674f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_41 VPB N_C_N_c_72_n 0.00327867f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_42 VPB N_C_N_c_73_n 0.00249829f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_43 VPB N_D_N_c_107_n 0.0285733f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_44 VPB D_N 0.00132037f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_45 VPB N_A_216_93#_c_142_n 0.0189871f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_46 VPB N_A_216_93#_c_137_n 0.0115294f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_47 VPB N_A_216_93#_c_138_n 0.00608661f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_48 VPB N_A_216_93#_c_145_n 0.0124103f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_49 VPB N_A_216_93#_c_140_n 0.00351783f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_A_27_410#_c_196_n 0.0252331f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_51 VPB N_A_27_410#_c_198_n 0.0273499f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_52 VPB N_A_27_410#_c_203_n 0.0149581f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.325
cc_53 VPB N_A_27_410#_c_204_n 0.00747461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_410#_c_205_n 0.00612227f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.53
cc_55 VPB N_A_27_410#_c_206_n 0.0097009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_410#_c_207_n 0.00373498f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_410#_c_199_n 0.00223652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_410#_c_209_n 0.0117133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B_c_273_n 0.023903f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_60 VPB N_B_c_275_n 0.00244362f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_c_302_n 0.0275299f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_62 VPB A 0.00788878f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=0.675
cc_63 VPB N_VPWR_c_322_n 0.00684542f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_64 VPB N_VPWR_c_323_n 0.0147131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_324_n 0.035898f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_66 VPB N_VPWR_c_325_n 0.0144618f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.325
cc_67 VPB N_VPWR_c_326_n 0.0642391f $X=-0.19 $Y=1.305 $X2=0.63 $Y2=1.53
cc_68 VPB N_VPWR_c_327_n 0.00593536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_321_n 0.0550457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_Y_c_367_n 0.00358877f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.445
cc_71 VPB N_Y_c_366_n 0.00109751f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_72 N_C_N_c_74_n N_D_N_c_106_n 0.0105153f $X=0.53 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_73 N_C_N_c_75_n N_D_N_c_107_n 0.0219527f $X=0.495 $Y=1.875 $X2=0 $Y2=0
cc_74 N_C_N_c_76_n N_D_N_c_107_n 0.00196013f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_75 N_C_N_c_72_n N_D_N_c_107_n 0.0149638f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_76 N_C_N_c_73_n N_D_N_c_107_n 0.00951774f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_77 N_C_N_c_72_n D_N 2.83086e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_N_c_73_n D_N 0.0265431f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_79 N_C_N_c_75_n N_A_216_93#_c_145_n 2.14279e-19 $X=0.495 $Y=1.875 $X2=0 $Y2=0
cc_80 N_C_N_c_73_n N_A_216_93#_c_145_n 0.00989496f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_81 N_C_N_c_72_n N_A_27_410#_c_198_n 0.0221654f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_82 N_C_N_c_73_n N_A_27_410#_c_198_n 0.0534696f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_83 N_C_N_c_74_n N_A_27_410#_c_198_n 0.00501087f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_84 N_C_N_c_76_n N_A_27_410#_c_203_n 0.00479178f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_85 N_C_N_c_76_n N_A_27_410#_c_204_n 0.0176421f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_86 N_C_N_c_72_n N_A_27_410#_c_204_n 2.27401e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_87 N_C_N_c_73_n N_A_27_410#_c_204_n 0.0294214f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_88 N_C_N_c_76_n N_A_27_410#_c_205_n 0.00268221f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_89 N_C_N_c_72_n N_A_27_410#_c_200_n 4.49664e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_90 N_C_N_c_74_n N_A_27_410#_c_200_n 0.00215399f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_91 N_C_N_c_73_n N_VPWR_M1008_d 0.00464392f $X=0.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_92 N_C_N_c_76_n N_VPWR_c_322_n 0.0122493f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_93 N_C_N_c_76_n N_VPWR_c_325_n 0.00306699f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_94 N_C_N_c_76_n N_VPWR_c_321_n 0.00454334f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_95 N_C_N_c_73_n N_VGND_c_421_n 0.0113325f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_96 N_C_N_c_74_n N_VGND_c_421_n 0.00448195f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_97 N_C_N_c_74_n N_VGND_c_426_n 0.00510437f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_98 N_C_N_c_74_n N_VGND_c_433_n 0.00512902f $X=0.53 $Y=0.995 $X2=0 $Y2=0
cc_99 N_D_N_c_107_n N_A_216_93#_c_137_n 0.0110158f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_100 D_N N_A_216_93#_c_137_n 0.00278531f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_101 N_D_N_c_107_n N_A_216_93#_c_145_n 0.00501309f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_102 D_N N_A_216_93#_c_145_n 0.0143223f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_103 N_D_N_c_106_n N_A_216_93#_c_140_n 0.00358705f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_104 N_D_N_c_107_n N_A_216_93#_c_140_n 0.00480292f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_105 D_N N_A_216_93#_c_140_n 0.0172045f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_106 N_D_N_c_106_n N_A_216_93#_c_141_n 0.00187001f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_D_N_c_107_n N_A_216_93#_c_141_n 0.00100647f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_108 D_N N_A_216_93#_c_141_n 0.0134146f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_109 N_D_N_c_107_n N_A_27_410#_c_204_n 0.0155252f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_110 D_N N_A_27_410#_c_204_n 0.00269637f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_111 N_D_N_c_107_n N_VPWR_c_326_n 6.50559e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_112 N_D_N_c_107_n N_Y_c_367_n 4.09148e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_113 N_D_N_c_106_n N_VGND_c_421_n 0.00289791f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_114 N_D_N_c_106_n N_VGND_c_422_n 0.00295956f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_115 N_D_N_c_106_n N_VGND_c_428_n 0.00510437f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_116 N_D_N_c_106_n N_VGND_c_433_n 0.00512902f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_216_93#_c_142_n N_A_27_410#_c_196_n 0.0500918f $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_216_93#_c_138_n N_A_27_410#_c_196_n 0.0240929f $X=2.02 $Y=1.202 $X2=0
+ $Y2=0
cc_119 N_A_216_93#_c_136_n N_A_27_410#_c_197_n 0.0181699f $X=2.045 $Y=0.995
+ $X2=0 $Y2=0
cc_120 N_A_216_93#_M1009_d N_A_27_410#_c_204_n 0.00174577f $X=1.12 $Y=1.485
+ $X2=0 $Y2=0
cc_121 N_A_216_93#_c_145_n N_A_27_410#_c_204_n 0.0117002f $X=1.62 $Y=1.62 $X2=0
+ $Y2=0
cc_122 N_A_216_93#_c_142_n N_A_27_410#_c_205_n 0.00250018f $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_123 N_A_216_93#_c_142_n N_A_27_410#_c_206_n 0.0129905f $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_124 N_A_216_93#_c_145_n N_A_27_410#_c_206_n 0.00859714f $X=1.62 $Y=1.62 $X2=0
+ $Y2=0
cc_125 N_A_216_93#_c_142_n N_A_27_410#_c_199_n 6.57659e-19 $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_126 N_A_216_93#_c_138_n N_A_27_410#_c_199_n 5.44754e-19 $X=2.02 $Y=1.202
+ $X2=0 $Y2=0
cc_127 N_A_216_93#_c_142_n N_VPWR_c_326_n 0.00429453f $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A_216_93#_c_142_n N_VPWR_c_321_n 0.00748834f $X=2.02 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A_216_93#_c_145_n N_Y_M1005_s 0.00456525f $X=1.62 $Y=1.62 $X2=0 $Y2=0
cc_130 N_A_216_93#_c_140_n N_Y_M1005_s 4.5056e-19 $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_216_93#_c_142_n N_Y_c_367_n 0.00770296f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_216_93#_c_137_n N_Y_c_367_n 0.00313319f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_216_93#_c_145_n N_Y_c_367_n 0.0134649f $X=1.62 $Y=1.62 $X2=0 $Y2=0
cc_134 N_A_216_93#_c_142_n N_Y_c_366_n 0.0206668f $X=2.02 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_216_93#_c_136_n N_Y_c_366_n 0.00587656f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_216_93#_c_138_n N_Y_c_366_n 0.0135423f $X=2.02 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_216_93#_c_145_n N_Y_c_366_n 0.0154101f $X=1.62 $Y=1.62 $X2=0 $Y2=0
cc_138 N_A_216_93#_c_140_n N_Y_c_366_n 0.0482774f $X=1.705 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_216_93#_c_136_n N_Y_c_380_n 0.0100657f $X=2.045 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_216_93#_c_139_n N_VGND_M1003_s 0.00400305f $X=1.62 $Y=0.74 $X2=0
+ $Y2=0
cc_141 N_A_216_93#_c_140_n N_VGND_M1003_s 4.95468e-19 $X=1.705 $Y=1.16 $X2=0
+ $Y2=0
cc_142 N_A_216_93#_c_141_n N_VGND_c_421_n 0.00934005f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_143 N_A_216_93#_c_136_n N_VGND_c_422_n 0.00341589f $X=2.045 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A_216_93#_c_137_n N_VGND_c_422_n 0.00490246f $X=1.92 $Y=1.16 $X2=0
+ $Y2=0
cc_145 N_A_216_93#_c_139_n N_VGND_c_422_n 0.0140929f $X=1.62 $Y=0.74 $X2=0 $Y2=0
cc_146 N_A_216_93#_c_141_n N_VGND_c_422_n 0.00168088f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_147 N_A_216_93#_c_136_n N_VGND_c_423_n 6.74955e-19 $X=2.045 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_216_93#_c_139_n N_VGND_c_428_n 0.00477097f $X=1.62 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_216_93#_c_141_n N_VGND_c_428_n 0.00512277f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_150 N_A_216_93#_c_136_n N_VGND_c_430_n 0.00427876f $X=2.045 $Y=0.995 $X2=0
+ $Y2=0
cc_151 N_A_216_93#_c_136_n N_VGND_c_433_n 0.00718208f $X=2.045 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_216_93#_c_139_n N_VGND_c_433_n 0.00849895f $X=1.62 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_216_93#_c_141_n N_VGND_c_433_n 0.00563626f $X=1.26 $Y=0.66 $X2=0
+ $Y2=0
cc_154 N_A_27_410#_c_196_n N_B_c_273_n 0.0633358f $X=2.5 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_27_410#_c_199_n N_B_c_273_n 0.00205316f $X=2.465 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_27_410#_c_197_n N_B_c_274_n 0.0229401f $X=2.525 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_27_410#_c_196_n N_B_c_275_n 0.00501752f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_27_410#_c_199_n N_B_c_275_n 0.0626832f $X=2.465 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_27_410#_c_204_n N_VPWR_M1008_d 0.00604817f $X=1.135 $Y=1.977
+ $X2=-0.19 $Y2=-0.24
cc_160 N_A_27_410#_c_203_n N_VPWR_c_322_n 0.0165638f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_161 N_A_27_410#_c_204_n N_VPWR_c_322_n 0.0244739f $X=1.135 $Y=1.977 $X2=0
+ $Y2=0
cc_162 N_A_27_410#_c_205_n N_VPWR_c_322_n 0.00343759f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_163 N_A_27_410#_c_207_n N_VPWR_c_322_n 0.0119283f $X=1.305 $Y=2.38 $X2=0
+ $Y2=0
cc_164 N_A_27_410#_c_203_n N_VPWR_c_325_n 0.0170443f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_165 N_A_27_410#_c_204_n N_VPWR_c_325_n 0.00230305f $X=1.135 $Y=1.977 $X2=0
+ $Y2=0
cc_166 N_A_27_410#_c_196_n N_VPWR_c_326_n 0.00429201f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_27_410#_c_204_n N_VPWR_c_326_n 0.00425784f $X=1.135 $Y=1.977 $X2=0
+ $Y2=0
cc_168 N_A_27_410#_c_206_n N_VPWR_c_326_n 0.0784054f $X=2.38 $Y=2.38 $X2=0 $Y2=0
cc_169 N_A_27_410#_c_207_n N_VPWR_c_326_n 0.0120427f $X=1.305 $Y=2.38 $X2=0
+ $Y2=0
cc_170 N_A_27_410#_c_196_n N_VPWR_c_321_n 0.00630133f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_27_410#_c_203_n N_VPWR_c_321_n 0.00987378f $X=0.26 $Y=2.29 $X2=0
+ $Y2=0
cc_172 N_A_27_410#_c_204_n N_VPWR_c_321_n 0.0126415f $X=1.135 $Y=1.977 $X2=0
+ $Y2=0
cc_173 N_A_27_410#_c_206_n N_VPWR_c_321_n 0.047429f $X=2.38 $Y=2.38 $X2=0 $Y2=0
cc_174 N_A_27_410#_c_207_n N_VPWR_c_321_n 0.00651993f $X=1.305 $Y=2.38 $X2=0
+ $Y2=0
cc_175 N_A_27_410#_c_206_n N_Y_M1005_s 0.00509651f $X=2.38 $Y=2.38 $X2=0 $Y2=0
cc_176 N_A_27_410#_c_196_n N_Y_c_367_n 6.31334e-19 $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_27_410#_c_204_n N_Y_c_367_n 0.00767905f $X=1.135 $Y=1.977 $X2=0 $Y2=0
cc_178 N_A_27_410#_c_205_n N_Y_c_367_n 0.00325524f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_179 N_A_27_410#_c_206_n N_Y_c_367_n 0.0363558f $X=2.38 $Y=2.38 $X2=0 $Y2=0
cc_180 N_A_27_410#_c_196_n N_Y_c_366_n 0.00394949f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_27_410#_c_197_n N_Y_c_366_n 0.00354194f $X=2.525 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_27_410#_c_204_n N_Y_c_366_n 0.00203753f $X=1.135 $Y=1.977 $X2=0 $Y2=0
cc_183 N_A_27_410#_c_199_n N_Y_c_366_n 0.0556376f $X=2.465 $Y=1.16 $X2=0 $Y2=0
cc_184 N_A_27_410#_c_196_n N_Y_c_390_n 7.53888e-19 $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A_27_410#_c_197_n N_Y_c_390_n 0.0120196f $X=2.525 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_27_410#_c_199_n N_Y_c_390_n 0.0154237f $X=2.465 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_410#_c_196_n N_Y_c_380_n 0.00171206f $X=2.5 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_410#_c_206_n A_422_297# 0.00764964f $X=2.38 $Y=2.38 $X2=-0.19
+ $Y2=-0.24
cc_189 N_A_27_410#_c_200_n N_VGND_c_421_n 0.0188143f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_190 N_A_27_410#_c_197_n N_VGND_c_423_n 0.00675938f $X=2.525 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_27_410#_c_200_n N_VGND_c_426_n 0.00972557f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_192 N_A_27_410#_c_197_n N_VGND_c_430_n 0.00398759f $X=2.525 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_27_410#_c_197_n N_VGND_c_433_n 0.00477752f $X=2.525 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_27_410#_c_200_n N_VGND_c_433_n 0.0107261f $X=0.3 $Y=0.66 $X2=0 $Y2=0
cc_195 N_B_c_274_n N_A_c_301_n 0.0219255f $X=3.045 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_196 N_B_c_273_n N_A_c_302_n 0.0725978f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_275_n N_A_c_302_n 0.00183289f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_198 N_B_c_273_n A 0.00192033f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_275_n A 0.0326486f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_200 N_B_c_273_n N_VPWR_c_324_n 0.00201585f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_273_n N_VPWR_c_326_n 0.00442707f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_275_n N_VPWR_c_326_n 0.0137325f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_203 N_B_c_273_n N_VPWR_c_321_n 0.00630585f $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_275_n N_VPWR_c_321_n 0.0106827f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_205 N_B_c_273_n N_Y_c_390_n 7.17521e-19 $X=3.02 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_274_n N_Y_c_390_n 0.0115184f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_207 N_B_c_275_n N_Y_c_390_n 0.0216097f $X=2.985 $Y=1.16 $X2=0 $Y2=0
cc_208 N_B_c_275_n A_518_297# 0.00923928f $X=2.985 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_209 N_B_c_274_n N_VGND_c_423_n 0.00294569f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_210 N_B_c_274_n N_VGND_c_425_n 8.85097e-19 $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_211 N_B_c_274_n N_VGND_c_432_n 0.00428022f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B_c_274_n N_VGND_c_433_n 0.00609388f $X=3.045 $Y=0.995 $X2=0 $Y2=0
cc_213 A N_VPWR_M1007_d 0.00928569f $X=3.44 $Y=1.105 $X2=0 $Y2=0
cc_214 N_A_c_302_n N_VPWR_c_324_n 0.0202129f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_215 A N_VPWR_c_324_n 0.00830984f $X=3.44 $Y=1.105 $X2=0 $Y2=0
cc_216 N_A_c_302_n N_VPWR_c_326_n 0.00427505f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_302_n N_VPWR_c_321_n 0.00743383f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_301_n N_VGND_c_425_n 0.0123719f $X=3.465 $Y=0.995 $X2=0 $Y2=0
cc_219 N_A_c_302_n N_VGND_c_425_n 0.00279043f $X=3.49 $Y=1.41 $X2=0 $Y2=0
cc_220 A N_VGND_c_425_n 0.0107812f $X=3.44 $Y=1.105 $X2=0 $Y2=0
cc_221 N_A_c_301_n N_VGND_c_432_n 0.0046653f $X=3.465 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_c_301_n N_VGND_c_433_n 0.00799591f $X=3.465 $Y=0.995 $X2=0 $Y2=0
cc_223 N_VPWR_c_321_n N_Y_M1005_s 0.00218346f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_224 N_VPWR_c_321_n A_422_297# 0.00240923f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_225 N_VPWR_c_321_n A_518_297# 0.0098973f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_226 N_VPWR_c_321_n A_622_297# 0.0117394f $X=3.91 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_227 N_Y_c_367_n A_422_297# 0.0019205f $X=1.96 $Y=2.04 $X2=-0.19 $Y2=-0.24
cc_228 N_Y_c_366_n A_422_297# 0.00401421f $X=2.085 $Y=1.955 $X2=-0.19 $Y2=-0.24
cc_229 N_Y_c_390_n N_VGND_M1006_d 0.00980742f $X=3.14 $Y=0.74 $X2=0 $Y2=0
cc_230 N_Y_c_401_p N_VGND_c_423_n 0.0113373f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_231 N_Y_c_390_n N_VGND_c_423_n 0.0202581f $X=3.14 $Y=0.74 $X2=0 $Y2=0
cc_232 N_Y_c_401_p N_VGND_c_430_n 0.0104733f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_233 N_Y_c_390_n N_VGND_c_430_n 0.00307941f $X=3.14 $Y=0.74 $X2=0 $Y2=0
cc_234 N_Y_c_380_n N_VGND_c_430_n 0.00312613f $X=2.165 $Y=0.74 $X2=0 $Y2=0
cc_235 N_Y_c_390_n N_VGND_c_432_n 0.0029785f $X=3.14 $Y=0.74 $X2=0 $Y2=0
cc_236 Y N_VGND_c_432_n 0.00906533f $X=3.16 $Y=0.425 $X2=0 $Y2=0
cc_237 N_Y_M1003_d N_VGND_c_433_n 0.00316568f $X=2.12 $Y=0.235 $X2=0 $Y2=0
cc_238 N_Y_M1001_d N_VGND_c_433_n 0.00403782f $X=3.12 $Y=0.235 $X2=0 $Y2=0
cc_239 N_Y_c_401_p N_VGND_c_433_n 0.0074087f $X=2.255 $Y=0.495 $X2=0 $Y2=0
cc_240 N_Y_c_390_n N_VGND_c_433_n 0.012226f $X=3.14 $Y=0.74 $X2=0 $Y2=0
cc_241 N_Y_c_380_n N_VGND_c_433_n 0.00540169f $X=2.165 $Y=0.74 $X2=0 $Y2=0
cc_242 Y N_VGND_c_433_n 0.00735151f $X=3.16 $Y=0.425 $X2=0 $Y2=0
