* File: sky130_fd_sc_hdll__or4_2.pxi.spice
* Created: Wed Sep  2 08:49:19 2020
* 
x_PM_SKY130_FD_SC_HDLL__OR4_2%D N_D_c_70_n N_D_M1003_g N_D_M1000_g D D
+ N_D_c_69_n PM_SKY130_FD_SC_HDLL__OR4_2%D
x_PM_SKY130_FD_SC_HDLL__OR4_2%C N_C_c_95_n N_C_M1010_g N_C_M1006_g C C C C C C
+ PM_SKY130_FD_SC_HDLL__OR4_2%C
x_PM_SKY130_FD_SC_HDLL__OR4_2%B N_B_c_130_n N_B_c_133_n N_B_c_134_n N_B_M1011_g
+ N_B_M1005_g N_B_c_131_n N_B_c_132_n B B B B B B PM_SKY130_FD_SC_HDLL__OR4_2%B
x_PM_SKY130_FD_SC_HDLL__OR4_2%A N_A_c_174_n N_A_M1004_g N_A_M1001_g A
+ N_A_c_176_n A PM_SKY130_FD_SC_HDLL__OR4_2%A
x_PM_SKY130_FD_SC_HDLL__OR4_2%A_27_297# N_A_27_297#_M1000_d N_A_27_297#_M1005_d
+ N_A_27_297#_M1003_s N_A_27_297#_c_215_n N_A_27_297#_M1002_g
+ N_A_27_297#_c_226_n N_A_27_297#_M1007_g N_A_27_297#_c_227_n
+ N_A_27_297#_M1009_g N_A_27_297#_c_216_n N_A_27_297#_M1008_g
+ N_A_27_297#_c_217_n N_A_27_297#_c_218_n N_A_27_297#_c_219_n
+ N_A_27_297#_c_231_n N_A_27_297#_c_245_n N_A_27_297#_c_220_n
+ N_A_27_297#_c_221_n N_A_27_297#_c_322_p N_A_27_297#_c_222_n
+ N_A_27_297#_c_257_n N_A_27_297#_c_223_n N_A_27_297#_c_232_n
+ N_A_27_297#_c_233_n N_A_27_297#_c_224_n N_A_27_297#_c_234_n
+ N_A_27_297#_c_225_n PM_SKY130_FD_SC_HDLL__OR4_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__OR4_2%VPWR N_VPWR_M1004_d N_VPWR_M1009_d N_VPWR_c_344_n
+ N_VPWR_c_345_n N_VPWR_c_346_n N_VPWR_c_347_n N_VPWR_c_348_n VPWR
+ N_VPWR_c_349_n N_VPWR_c_343_n PM_SKY130_FD_SC_HDLL__OR4_2%VPWR
x_PM_SKY130_FD_SC_HDLL__OR4_2%X N_X_M1002_d N_X_M1007_s N_X_c_376_n N_X_c_380_n
+ N_X_c_374_n X PM_SKY130_FD_SC_HDLL__OR4_2%X
x_PM_SKY130_FD_SC_HDLL__OR4_2%VGND N_VGND_M1000_s N_VGND_M1006_d N_VGND_M1001_d
+ N_VGND_M1008_s N_VGND_c_405_n N_VGND_c_406_n N_VGND_c_407_n N_VGND_c_408_n
+ N_VGND_c_409_n VGND N_VGND_c_410_n N_VGND_c_411_n N_VGND_c_412_n
+ N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n PM_SKY130_FD_SC_HDLL__OR4_2%VGND
cc_1 VNB N_D_M1000_g 0.033863f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB D 0.0266761f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_D_c_69_n 0.0389134f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_C_c_95_n 0.0210104f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_C_M1006_g 0.026662f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_6 VNB C 0.00949415f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_B_c_130_n 0.0205225f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_8 VNB N_B_c_131_n 0.0147582f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_c_132_n 0.0135779f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_c_174_n 0.0246492f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_A_M1001_g 0.0272047f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_12 VNB N_A_c_176_n 0.00216296f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_13 VNB N_A_27_297#_c_215_n 0.0185579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_297#_c_216_n 0.020717f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_297#_c_217_n 0.0108766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_218_n 0.0280807f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_219_n 0.0235634f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_220_n 0.00390934f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_221_n 0.00325027f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_297#_c_222_n 0.00135955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_297#_c_223_n 0.00147549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_297#_c_224_n 0.00149272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_297#_c_225_n 0.00226413f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_343_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_374_n 0.00103657f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_26 VNB N_VGND_c_405_n 0.0114891f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_27 VNB N_VGND_c_406_n 0.0195472f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_28 VNB N_VGND_c_407_n 0.00270623f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_408_n 0.0110579f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_409_n 0.0138237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_410_n 0.0164929f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_411_n 0.0138146f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_412_n 0.0253862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_413_n 0.00602632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_414_n 0.00664852f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_415_n 0.210194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VPB N_D_c_70_n 0.0213198f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_38 VPB D 0.00363797f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_39 VPB N_D_c_69_n 0.0178473f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_40 VPB N_C_c_95_n 0.0238977f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB C 0.00371969f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B_c_133_n 0.0062896f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.695
cc_43 VPB N_B_c_134_n 0.0498712f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_44 VPB N_B_M1011_g 0.0111652f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_45 VPB B 0.0507627f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_46 VPB N_A_c_174_n 0.0289584f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_47 VPB N_A_c_176_n 0.00295988f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.202
cc_48 VPB N_A_27_297#_c_226_n 0.0198853f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_49 VPB N_A_27_297#_c_227_n 0.0211129f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_50 VPB N_A_27_297#_c_217_n 0.00660177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_27_297#_c_218_n 0.0179529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_27_297#_c_219_n 0.00987427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_297#_c_231_n 0.00581573f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_297#_c_232_n 0.0019714f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_297#_c_233_n 0.0213018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_297#_c_234_n 0.00205005f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_297#_c_225_n 5.11682e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_344_n 0.0129735f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_59 VPB N_VPWR_c_345_n 0.011032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_346_n 0.00961147f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_61 VPB N_VPWR_c_347_n 0.0540305f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_348_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_349_n 0.0262176f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_343_n 0.0652749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_X_c_374_n 0.00146684f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_66 N_D_c_70_n N_C_c_95_n 0.0216164f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_67 D N_C_c_95_n 2.25554e-19 $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_68 N_D_c_69_n N_C_c_95_n 0.0236421f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_69 N_D_M1000_g N_C_M1006_g 0.0191389f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_70 N_D_c_70_n C 0.00325995f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_71 D C 0.0279202f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_72 N_D_c_69_n C 0.00584047f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_73 N_D_c_70_n B 0.00528936f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_D_c_70_n N_A_27_297#_c_231_n 0.0141565f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 D N_A_27_297#_c_231_n 8.01096e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_76 N_D_M1000_g N_A_27_297#_c_221_n 0.00385395f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_77 D N_A_27_297#_c_221_n 0.00487517f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_78 N_D_c_70_n N_A_27_297#_c_233_n 0.00647329f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_79 D N_A_27_297#_c_233_n 0.0248263f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_80 N_D_c_69_n N_A_27_297#_c_233_n 0.00192889f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_81 N_D_M1000_g N_VGND_c_406_n 0.00427003f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_82 D N_VGND_c_406_n 0.0276393f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_83 N_D_c_69_n N_VGND_c_406_n 0.00130319f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_84 N_D_M1000_g N_VGND_c_407_n 5.72193e-19 $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_85 N_D_M1000_g N_VGND_c_410_n 0.00555245f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_86 N_D_M1000_g N_VGND_c_415_n 0.0113233f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_87 D N_VGND_c_415_n 0.00184222f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_88 N_C_c_95_n N_B_c_130_n 0.0201924f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_89 C N_B_c_130_n 0.00524431f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_90 N_C_c_95_n N_B_M1011_g 0.0355231f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_91 C N_B_M1011_g 0.00282307f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_92 N_C_M1006_g N_B_c_131_n 0.0112508f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_93 N_C_M1006_g N_B_c_132_n 0.0201924f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_94 N_C_c_95_n B 0.00527095f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_95 N_C_c_95_n N_A_c_176_n 2.36343e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_96 C N_A_c_176_n 0.0290697f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_97 N_C_c_95_n N_A_27_297#_c_231_n 0.0109955f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_98 C N_A_27_297#_c_231_n 0.0418289f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_99 N_C_M1006_g N_A_27_297#_c_245_n 0.00520782f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_100 N_C_c_95_n N_A_27_297#_c_220_n 0.00308093f $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_101 N_C_M1006_g N_A_27_297#_c_220_n 0.01115f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_102 C N_A_27_297#_c_220_n 0.0365281f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_103 N_C_c_95_n N_A_27_297#_c_221_n 9.23324e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_104 C N_A_27_297#_c_221_n 0.0152593f $X=1.105 $Y=1.445 $X2=0 $Y2=0
cc_105 N_C_c_95_n N_A_27_297#_c_233_n 9.0777e-19 $X=1.025 $Y=1.41 $X2=0 $Y2=0
cc_106 C A_117_297# 0.0032015f $X=1.105 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_107 C A_223_297# 0.00128624f $X=1.105 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_108 N_C_M1006_g N_VGND_c_407_n 0.0101294f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_109 N_C_M1006_g N_VGND_c_410_n 0.00187556f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_110 N_C_M1006_g N_VGND_c_415_n 0.00271727f $X=1.05 $Y=0.475 $X2=0 $Y2=0
cc_111 N_B_c_130_n N_A_c_174_n 0.0167852f $X=1.435 $Y=1.31 $X2=-0.19 $Y2=-0.24
cc_112 N_B_c_133_n N_A_c_174_n 0.0034991f $X=1.435 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_113 N_B_M1011_g N_A_c_174_n 0.0195328f $X=1.435 $Y=1.695 $X2=-0.19 $Y2=-0.24
cc_114 B N_A_c_174_n 6.66635e-19 $X=1.515 $Y=2.125 $X2=-0.19 $Y2=-0.24
cc_115 N_B_c_130_n N_A_M1001_g 0.00330916f $X=1.435 $Y=1.31 $X2=0 $Y2=0
cc_116 N_B_c_131_n N_A_M1001_g 0.0154918f $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_117 N_B_c_130_n N_A_c_176_n 0.00849267f $X=1.435 $Y=1.31 $X2=0 $Y2=0
cc_118 N_B_c_133_n N_A_c_176_n 0.00171029f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B_c_132_n N_A_c_176_n 0.00177283f $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_120 N_B_c_134_n N_A_27_297#_c_231_n 0.00108081f $X=1.435 $Y=2.035 $X2=0 $Y2=0
cc_121 N_B_M1011_g N_A_27_297#_c_231_n 0.0153201f $X=1.435 $Y=1.695 $X2=0 $Y2=0
cc_122 B N_A_27_297#_c_231_n 0.0923567f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_123 N_B_c_131_n N_A_27_297#_c_220_n 0.00747646f $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_124 N_B_c_132_n N_A_27_297#_c_220_n 0.0122051f $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_125 B N_A_27_297#_c_257_n 0.00163296f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_126 B N_A_27_297#_c_233_n 0.0265285f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_127 N_B_M1011_g N_A_27_297#_c_234_n 0.0051945f $X=1.435 $Y=1.695 $X2=0 $Y2=0
cc_128 B N_A_27_297#_c_234_n 0.0138062f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_129 N_B_c_134_n N_VPWR_c_344_n 0.00350357f $X=1.435 $Y=2.035 $X2=0 $Y2=0
cc_130 B N_VPWR_c_344_n 0.0210031f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_131 N_B_c_134_n N_VPWR_c_347_n 0.00793506f $X=1.435 $Y=2.035 $X2=0 $Y2=0
cc_132 B N_VPWR_c_347_n 0.0911538f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_133 N_B_c_134_n N_VPWR_c_343_n 0.0113914f $X=1.435 $Y=2.035 $X2=0 $Y2=0
cc_134 B N_VPWR_c_343_n 0.0660152f $X=1.515 $Y=2.125 $X2=0 $Y2=0
cc_135 N_B_c_131_n N_VGND_c_407_n 0.00166902f $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_136 N_B_c_132_n N_VGND_c_407_n 4.40092e-19 $X=1.465 $Y=0.91 $X2=0 $Y2=0
cc_137 N_B_c_131_n N_VGND_c_411_n 0.00403348f $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_138 N_B_c_131_n N_VGND_c_414_n 5.85623e-19 $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_139 N_B_c_131_n N_VGND_c_415_n 0.00564418f $X=1.465 $Y=0.76 $X2=0 $Y2=0
cc_140 N_A_M1001_g N_A_27_297#_c_215_n 0.0175538f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_141 N_A_c_174_n N_A_27_297#_c_226_n 0.0162601f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_174_n N_A_27_297#_c_217_n 0.015987f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_176_n N_A_27_297#_c_217_n 3.16637e-19 $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A_c_176_n N_A_27_297#_c_231_n 0.00573381f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_c_176_n N_A_27_297#_c_220_n 0.0127413f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_146 N_A_c_174_n N_A_27_297#_c_222_n 0.0034911f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_M1001_g N_A_27_297#_c_222_n 0.0114522f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_148 N_A_c_176_n N_A_27_297#_c_222_n 0.0204446f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_c_174_n N_A_27_297#_c_257_n 0.0156215f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_176_n N_A_27_297#_c_257_n 0.0160437f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_M1001_g N_A_27_297#_c_223_n 0.00346969f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_152 N_A_c_174_n N_A_27_297#_c_232_n 0.00349984f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_c_174_n N_A_27_297#_c_224_n 5.77159e-19 $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_c_176_n N_A_27_297#_c_224_n 0.0146254f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_c_174_n N_A_27_297#_c_234_n 0.00266894f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_c_176_n N_A_27_297#_c_234_n 0.0135132f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_157 N_A_c_174_n N_A_27_297#_c_225_n 0.00232056f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_176_n N_A_27_297#_c_225_n 0.0280505f $X=1.925 $Y=1.16 $X2=0 $Y2=0
cc_159 N_A_c_174_n N_VPWR_c_344_n 0.00342204f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_174_n N_VPWR_c_347_n 0.00351268f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A_c_174_n N_VPWR_c_343_n 0.00445321f $X=1.965 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_M1001_g N_VGND_c_411_n 0.00188229f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_163 N_A_M1001_g N_VGND_c_414_n 0.0101041f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_164 N_A_M1001_g N_VGND_c_415_n 0.00261357f $X=1.99 $Y=0.475 $X2=0 $Y2=0
cc_165 N_A_27_297#_c_231_n A_117_297# 0.00241926f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_166 N_A_27_297#_c_231_n A_223_297# 0.00123611f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_167 N_A_27_297#_c_231_n A_305_297# 0.00163933f $X=1.66 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_27_297#_c_234_n A_305_297# 0.00577191f $X=1.745 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_169 N_A_27_297#_c_257_n N_VPWR_M1004_d 0.00561585f $X=2.265 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_27_297#_c_226_n N_VPWR_c_344_n 0.00482583f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_27_297#_c_257_n N_VPWR_c_344_n 0.0200207f $X=2.265 $Y=1.58 $X2=0
+ $Y2=0
cc_172 N_A_27_297#_c_234_n N_VPWR_c_344_n 0.00457307f $X=1.745 $Y=1.58 $X2=0
+ $Y2=0
cc_173 N_A_27_297#_c_227_n N_VPWR_c_346_n 0.00826499f $X=3.14 $Y=1.41 $X2=0
+ $Y2=0
cc_174 N_A_27_297#_c_226_n N_VPWR_c_349_n 0.00702461f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_27_297#_c_227_n N_VPWR_c_349_n 0.00590121f $X=3.14 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_27_297#_c_226_n N_VPWR_c_343_n 0.0141458f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_27_297#_c_227_n N_VPWR_c_343_n 0.0112403f $X=3.14 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_27_297#_c_215_n N_X_c_376_n 0.00550306f $X=2.48 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_27_297#_c_216_n N_X_c_376_n 0.00459562f $X=3.165 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_27_297#_c_218_n N_X_c_376_n 0.00261904f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_181 N_A_27_297#_c_222_n N_X_c_376_n 0.00456953f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_182 N_A_27_297#_c_226_n N_X_c_380_n 0.0118214f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_27_297#_c_227_n N_X_c_380_n 0.00426092f $X=3.14 $Y=1.41 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_218_n N_X_c_380_n 0.00306645f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_185 N_A_27_297#_c_257_n N_X_c_380_n 0.00731128f $X=2.265 $Y=1.58 $X2=0 $Y2=0
cc_186 N_A_27_297#_c_215_n N_X_c_374_n 0.00198383f $X=2.48 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_226_n N_X_c_374_n 7.29791e-19 $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_27_297#_c_227_n N_X_c_374_n 0.00355795f $X=3.14 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_27_297#_c_216_n N_X_c_374_n 0.00553389f $X=3.165 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_27_297#_c_217_n N_X_c_374_n 7.46749e-19 $X=2.505 $Y=1.202 $X2=0 $Y2=0
cc_191 N_A_27_297#_c_218_n N_X_c_374_n 0.0155949f $X=3.04 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_297#_c_219_n N_X_c_374_n 0.0206423f $X=3.14 $Y=1.202 $X2=0 $Y2=0
cc_193 N_A_27_297#_c_222_n N_X_c_374_n 0.00240973f $X=2.265 $Y=0.74 $X2=0 $Y2=0
cc_194 N_A_27_297#_c_223_n N_X_c_374_n 0.00586618f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_27_297#_c_232_n N_X_c_374_n 0.00592343f $X=2.35 $Y=1.495 $X2=0 $Y2=0
cc_196 N_A_27_297#_c_225_n N_X_c_374_n 0.0225345f $X=2.615 $Y=1.16 $X2=0 $Y2=0
cc_197 N_A_27_297#_c_227_n X 0.0142571f $X=3.14 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_27_297#_c_220_n N_VGND_M1006_d 0.00211434f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_199 N_A_27_297#_c_222_n N_VGND_M1001_d 0.00479994f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_200 N_A_27_297#_c_223_n N_VGND_M1001_d 6.98847e-19 $X=2.35 $Y=0.995 $X2=0
+ $Y2=0
cc_201 N_A_27_297#_c_245_n N_VGND_c_407_n 0.0118543f $X=0.76 $Y=0.47 $X2=0 $Y2=0
cc_202 N_A_27_297#_c_220_n N_VGND_c_407_n 0.0214496f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_203 N_A_27_297#_c_216_n N_VGND_c_409_n 0.0118948f $X=3.165 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A_27_297#_c_245_n N_VGND_c_410_n 0.00876148f $X=0.76 $Y=0.47 $X2=0
+ $Y2=0
cc_205 N_A_27_297#_c_220_n N_VGND_c_410_n 0.00282959f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_206 N_A_27_297#_c_220_n N_VGND_c_411_n 0.0029785f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_207 N_A_27_297#_c_322_p N_VGND_c_411_n 0.00861358f $X=1.73 $Y=0.47 $X2=0
+ $Y2=0
cc_208 N_A_27_297#_c_222_n N_VGND_c_411_n 0.00232988f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_209 N_A_27_297#_c_215_n N_VGND_c_412_n 0.00525358f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_210 N_A_27_297#_c_216_n N_VGND_c_412_n 0.00540845f $X=3.165 $Y=0.995 $X2=0
+ $Y2=0
cc_211 N_A_27_297#_c_222_n N_VGND_c_412_n 3.28435e-19 $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_212 N_A_27_297#_c_215_n N_VGND_c_414_n 0.00986338f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_213 N_A_27_297#_c_216_n N_VGND_c_414_n 0.00140294f $X=3.165 $Y=0.995 $X2=0
+ $Y2=0
cc_214 N_A_27_297#_c_322_p N_VGND_c_414_n 0.0135697f $X=1.73 $Y=0.47 $X2=0 $Y2=0
cc_215 N_A_27_297#_c_222_n N_VGND_c_414_n 0.0239317f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_216 N_A_27_297#_c_215_n N_VGND_c_415_n 0.00908624f $X=2.48 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_27_297#_c_216_n N_VGND_c_415_n 0.011021f $X=3.165 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_27_297#_c_245_n N_VGND_c_415_n 0.00625722f $X=0.76 $Y=0.47 $X2=0
+ $Y2=0
cc_219 N_A_27_297#_c_220_n N_VGND_c_415_n 0.0122608f $X=1.645 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_27_297#_c_322_p N_VGND_c_415_n 0.00625722f $X=1.73 $Y=0.47 $X2=0
+ $Y2=0
cc_221 N_A_27_297#_c_222_n N_VGND_c_415_n 0.00676015f $X=2.265 $Y=0.74 $X2=0
+ $Y2=0
cc_222 N_VPWR_c_343_n N_X_M1007_s 0.0115153f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_346_n N_X_c_374_n 0.0692746f $X=3.4 $Y=1.66 $X2=0 $Y2=0
cc_224 N_VPWR_c_349_n X 0.0191629f $X=3.315 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_343_n X 0.0113307f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_226 N_VPWR_c_346_n N_VGND_c_409_n 0.0102904f $X=3.4 $Y=1.66 $X2=0 $Y2=0
cc_227 N_X_c_376_n N_VGND_c_409_n 0.0399486f $X=2.905 $Y=0.59 $X2=0 $Y2=0
cc_228 N_X_c_376_n N_VGND_c_412_n 0.00930659f $X=2.905 $Y=0.59 $X2=0 $Y2=0
cc_229 N_X_c_376_n N_VGND_c_414_n 0.0028217f $X=2.905 $Y=0.59 $X2=0 $Y2=0
cc_230 N_X_M1002_d N_VGND_c_415_n 0.0137969f $X=2.555 $Y=0.235 $X2=0 $Y2=0
cc_231 N_X_c_376_n N_VGND_c_415_n 0.0104048f $X=2.905 $Y=0.59 $X2=0 $Y2=0
