* File: sky130_fd_sc_hdll__a32oi_4.pex.spice
* Created: Wed Sep  2 08:21:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%B2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 29 30 37 51 53 61 68
c84 22 0 1.16491e-19 $X=1.93 $Y=0.995
r85 59 61 18.2888 $w=2.28e-07 $l=3.65e-07 $layer=LI1_cond $X=0.33 $Y=1.19
+ $X2=0.695 $Y2=1.19
r86 51 52 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r87 50 51 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=1.46 $Y=1.202
+ $X2=1.905 $Y2=1.202
r88 49 50 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r89 47 49 5.19677 $w=3.71e-07 $l=4e-08 $layer=POLY_cond $X=1.395 $Y=1.202
+ $X2=1.435 $Y2=1.202
r90 47 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.395
+ $Y=1.16 $X2=1.395 $Y2=1.16
r91 45 47 52.6173 $w=3.71e-07 $l=4.05e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.395 $Y2=1.202
r92 44 45 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r93 43 44 57.814 $w=3.71e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r94 42 43 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r95 37 42 16.004 $w=3.71e-07 $l=1.17047e-07 $layer=POLY_cond $X=0.395 $Y=1.165
+ $X2=0.495 $Y2=1.202
r96 37 39 25.7087 $w=2.8e-07 $l=1.2e-07 $layer=POLY_cond $X=0.395 $Y=1.165
+ $X2=0.275 $Y2=1.165
r97 30 68 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=1.19
+ $X2=1.615 $Y2=1.19
r98 30 48 10.7728 $w=2.28e-07 $l=2.15e-07 $layer=LI1_cond $X=1.61 $Y=1.19
+ $X2=1.395 $Y2=1.19
r99 29 48 12.0255 $w=2.28e-07 $l=2.4e-07 $layer=LI1_cond $X=1.155 $Y=1.19
+ $X2=1.395 $Y2=1.19
r100 28 29 22.7983 $w=2.28e-07 $l=4.55e-07 $layer=LI1_cond $X=0.7 $Y=1.19
+ $X2=1.155 $Y2=1.19
r101 28 61 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=0.7 $Y=1.19
+ $X2=0.695 $Y2=1.19
r102 26 27 17.8105 $w=2.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.22 $Y=1.53
+ $X2=0.22 $Y2=1.87
r103 26 53 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=0.22 $Y=1.53
+ $X2=0.22 $Y2=1.305
r104 25 53 3.48622 $w=2.2e-07 $l=1.15e-07 $layer=LI1_cond $X=0.22 $Y=1.19
+ $X2=0.22 $Y2=1.305
r105 25 59 3.33465 $w=2.3e-07 $l=1.1e-07 $layer=LI1_cond $X=0.22 $Y=1.19
+ $X2=0.33 $Y2=1.19
r106 25 39 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r107 22 52 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r108 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r109 19 51 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r110 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r111 16 50 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r112 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r113 13 49 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r114 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r115 10 45 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r116 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r117 7 44 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r118 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r119 4 43 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r120 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=0.56
r121 1 42 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r122 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 40 41 46 49
r78 41 42 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r79 40 49 8.55602 $w=3.28e-07 $l=2.45e-07 $layer=LI1_cond $X=3.7 $Y=1.16
+ $X2=3.455 $Y2=1.16
r80 39 41 11.0134 $w=3.72e-07 $l=8.5e-08 $layer=POLY_cond $X=3.7 $Y=1.202
+ $X2=3.785 $Y2=1.202
r81 39 40 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.7
+ $Y=1.16 $X2=3.7 $Y2=1.16
r82 37 39 49.8844 $w=3.72e-07 $l=3.85e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.7 $Y2=1.202
r83 36 37 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r84 34 36 47.9409 $w=3.72e-07 $l=3.7e-07 $layer=POLY_cond $X=2.92 $Y=1.202
+ $X2=3.29 $Y2=1.202
r85 32 34 9.71774 $w=3.72e-07 $l=7.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.92 $Y2=1.202
r86 31 32 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r87 30 31 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r88 29 30 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r89 26 49 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=3.455 $Y2=1.16
r90 26 46 15.8897 $w=3.28e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.16
+ $X2=2.995 $Y2=1.16
r91 25 46 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=2.92 $Y=1.16
+ $X2=2.995 $Y2=1.16
r92 25 34 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.92
+ $Y=1.16 $X2=2.92 $Y2=1.16
r93 22 42 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r94 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r95 19 41 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r96 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r97 16 37 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r98 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r99 13 36 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r100 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r101 10 32 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r102 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r103 7 31 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r104 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r105 4 30 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r106 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r107 1 29 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r108 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 50 53 56
c69 28 0 1.71753e-19 $X=5.855 $Y=1.19
r70 45 46 15.6748 $w=3.69e-07 $l=1.2e-07 $layer=POLY_cond $X=6.14 $Y=1.202
+ $X2=6.26 $Y2=1.202
r71 43 45 37.8808 $w=3.69e-07 $l=2.9e-07 $layer=POLY_cond $X=5.85 $Y=1.202
+ $X2=6.14 $Y2=1.202
r72 41 43 7.8374 $w=3.69e-07 $l=6e-08 $layer=POLY_cond $X=5.79 $Y=1.202 $X2=5.85
+ $Y2=1.202
r73 40 41 61.393 $w=3.69e-07 $l=4.7e-07 $layer=POLY_cond $X=5.32 $Y=1.202
+ $X2=5.79 $Y2=1.202
r74 39 40 13.7154 $w=3.69e-07 $l=1.05e-07 $layer=POLY_cond $X=5.215 $Y=1.202
+ $X2=5.32 $Y2=1.202
r75 38 39 47.6775 $w=3.69e-07 $l=3.65e-07 $layer=POLY_cond $X=4.85 $Y=1.202
+ $X2=5.215 $Y2=1.202
r76 37 38 13.7154 $w=3.69e-07 $l=1.05e-07 $layer=POLY_cond $X=4.745 $Y=1.202
+ $X2=4.85 $Y2=1.202
r77 35 37 52.9024 $w=3.69e-07 $l=4.05e-07 $layer=POLY_cond $X=4.34 $Y=1.202
+ $X2=4.745 $Y2=1.202
r78 33 35 8.49051 $w=3.69e-07 $l=6.5e-08 $layer=POLY_cond $X=4.275 $Y=1.202
+ $X2=4.34 $Y2=1.202
r79 28 56 24.2944 $w=2.08e-07 $l=4.6e-07 $layer=LI1_cond $X=5.775 $Y=1.18
+ $X2=5.315 $Y2=1.18
r80 28 43 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.85
+ $Y=1.16 $X2=5.85 $Y2=1.16
r81 27 56 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=5.29 $Y=1.18
+ $X2=5.315 $Y2=1.18
r82 27 53 22.974 $w=2.08e-07 $l=4.35e-07 $layer=LI1_cond $X=5.29 $Y=1.18
+ $X2=4.855 $Y2=1.18
r83 26 53 1.84848 $w=2.08e-07 $l=3.5e-08 $layer=LI1_cond $X=4.82 $Y=1.18
+ $X2=4.855 $Y2=1.18
r84 26 50 22.4459 $w=2.08e-07 $l=4.25e-07 $layer=LI1_cond $X=4.82 $Y=1.18
+ $X2=4.395 $Y2=1.18
r85 25 50 2.90476 $w=2.08e-07 $l=5.5e-08 $layer=LI1_cond $X=4.34 $Y=1.18
+ $X2=4.395 $Y2=1.18
r86 25 35 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.34
+ $Y=1.16 $X2=4.34 $Y2=1.16
r87 22 46 23.9013 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.26 $Y=1.01
+ $X2=6.26 $Y2=1.202
r88 22 24 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=6.26 $Y=1.01 $X2=6.26
+ $Y2=0.56
r89 19 45 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.14 $Y=1.41 $X2=6.14
+ $Y2=1.202
r90 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.14 $Y=1.41
+ $X2=6.14 $Y2=1.985
r91 16 41 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=1.202
r92 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.79 $Y=0.995
+ $X2=5.79 $Y2=0.56
r93 13 40 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=1.202
r94 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.32 $Y=0.995
+ $X2=5.32 $Y2=0.56
r95 10 39 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.202
r96 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.215 $Y=1.41
+ $X2=5.215 $Y2=1.985
r97 7 38 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.85 $Y=0.995
+ $X2=4.85 $Y2=1.202
r98 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.85 $Y=0.995 $X2=4.85
+ $Y2=0.56
r99 4 37 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.202
r100 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.745 $Y=1.41
+ $X2=4.745 $Y2=1.985
r101 1 33 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.202
r102 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.275 $Y=1.41
+ $X2=4.275 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 45 50 58
c67 45 0 1.71753e-19 $X=8.255 $Y=1.202
r68 45 46 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=8.255 $Y=1.202
+ $X2=8.28 $Y2=1.202
r69 43 45 22.374 $w=3.77e-07 $l=1.75e-07 $layer=POLY_cond $X=8.08 $Y=1.202
+ $X2=8.255 $Y2=1.202
r70 41 43 37.7162 $w=3.77e-07 $l=2.95e-07 $layer=POLY_cond $X=7.785 $Y=1.202
+ $X2=8.08 $Y2=1.202
r71 40 41 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=7.76 $Y=1.202
+ $X2=7.785 $Y2=1.202
r72 39 40 56.8939 $w=3.77e-07 $l=4.45e-07 $layer=POLY_cond $X=7.315 $Y=1.202
+ $X2=7.76 $Y2=1.202
r73 38 39 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=7.29 $Y=1.202
+ $X2=7.315 $Y2=1.202
r74 37 50 10.5 $w=2.23e-07 $l=2.05e-07 $layer=LI1_cond $X=6.91 $Y=1.187
+ $X2=7.115 $Y2=1.187
r75 36 38 48.5836 $w=3.77e-07 $l=3.8e-07 $layer=POLY_cond $X=6.91 $Y=1.202
+ $X2=7.29 $Y2=1.202
r76 36 37 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.91
+ $Y=1.16 $X2=6.91 $Y2=1.16
r77 34 36 8.31034 $w=3.77e-07 $l=6.5e-08 $layer=POLY_cond $X=6.845 $Y=1.202
+ $X2=6.91 $Y2=1.202
r78 33 34 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=6.82 $Y=1.202
+ $X2=6.845 $Y2=1.202
r79 28 58 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=8.45 $Y=1.187
+ $X2=8.455 $Y2=1.187
r80 27 28 19.7196 $w=2.23e-07 $l=3.85e-07 $layer=LI1_cond $X=8.065 $Y=1.187
+ $X2=8.45 $Y2=1.187
r81 27 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=8.08
+ $Y=1.16 $X2=8.08 $Y2=1.16
r82 26 27 25.0976 $w=2.23e-07 $l=4.9e-07 $layer=LI1_cond $X=7.575 $Y=1.187
+ $X2=8.065 $Y2=1.187
r83 25 26 23.305 $w=2.23e-07 $l=4.55e-07 $layer=LI1_cond $X=7.12 $Y=1.187
+ $X2=7.575 $Y2=1.187
r84 25 50 0.256098 $w=2.23e-07 $l=5e-09 $layer=LI1_cond $X=7.12 $Y=1.187
+ $X2=7.115 $Y2=1.187
r85 22 46 24.4204 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.28 $Y=1.01
+ $X2=8.28 $Y2=1.202
r86 22 24 144.6 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=8.28 $Y=1.01 $X2=8.28
+ $Y2=0.56
r87 19 45 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.255 $Y=1.41
+ $X2=8.255 $Y2=1.202
r88 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.255 $Y=1.41
+ $X2=8.255 $Y2=1.985
r89 16 41 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.785 $Y=1.41
+ $X2=7.785 $Y2=1.202
r90 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.785 $Y=1.41
+ $X2=7.785 $Y2=1.985
r91 13 40 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.76 $Y=0.995
+ $X2=7.76 $Y2=1.202
r92 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.76 $Y=0.995
+ $X2=7.76 $Y2=0.56
r93 10 39 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.315 $Y=1.41
+ $X2=7.315 $Y2=1.202
r94 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.315 $Y=1.41
+ $X2=7.315 $Y2=1.985
r95 7 38 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.29 $Y=0.995
+ $X2=7.29 $Y2=1.202
r96 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.29 $Y=0.995 $X2=7.29
+ $Y2=0.56
r97 4 34 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.845 $Y=1.41
+ $X2=6.845 $Y2=1.202
r98 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.845 $Y=1.41
+ $X2=6.845 $Y2=1.985
r99 1 33 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.82 $Y=0.995
+ $X2=6.82 $Y2=1.202
r100 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.82 $Y=0.995
+ $X2=6.82 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A3 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 27 28 29 49 53 58 60 65
r78 58 60 24.8869 $w=2.03e-07 $l=4.6e-07 $layer=LI1_cond $X=9.435 $Y=1.177
+ $X2=9.895 $Y2=1.177
r79 49 51 25.4389 $w=3.6e-07 $l=1.9e-07 $layer=POLY_cond $X=10.68 $Y=1.202
+ $X2=10.87 $Y2=1.202
r80 48 49 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=10.655 $Y=1.202
+ $X2=10.68 $Y2=1.202
r81 46 48 23.4306 $w=3.6e-07 $l=1.75e-07 $layer=POLY_cond $X=10.48 $Y=1.202
+ $X2=10.655 $Y2=1.202
r82 46 47 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.48
+ $Y=1.16 $X2=10.48 $Y2=1.16
r83 44 46 39.4972 $w=3.6e-07 $l=2.95e-07 $layer=POLY_cond $X=10.185 $Y=1.202
+ $X2=10.48 $Y2=1.202
r84 43 44 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=10.16 $Y=1.202
+ $X2=10.185 $Y2=1.202
r85 42 43 59.5806 $w=3.6e-07 $l=4.45e-07 $layer=POLY_cond $X=9.715 $Y=1.202
+ $X2=10.16 $Y2=1.202
r86 41 42 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=9.69 $Y=1.202
+ $X2=9.715 $Y2=1.202
r87 39 41 50.8778 $w=3.6e-07 $l=3.8e-07 $layer=POLY_cond $X=9.31 $Y=1.202
+ $X2=9.69 $Y2=1.202
r88 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.31
+ $Y=1.16 $X2=9.31 $Y2=1.16
r89 37 39 8.70278 $w=3.6e-07 $l=6.5e-08 $layer=POLY_cond $X=9.245 $Y=1.202
+ $X2=9.31 $Y2=1.202
r90 36 37 3.34722 $w=3.6e-07 $l=2.5e-08 $layer=POLY_cond $X=9.22 $Y=1.202
+ $X2=9.245 $Y2=1.202
r91 29 65 9.2607 $w=2.78e-07 $l=2.25e-07 $layer=LI1_cond $X=10.895 $Y=0.85
+ $X2=10.895 $Y2=1.075
r92 28 65 2.96334 $w=2.8e-07 $l=1.02e-07 $layer=LI1_cond $X=10.895 $Y=1.177
+ $X2=10.895 $Y2=1.075
r93 28 53 4.06733 $w=2.05e-07 $l=1.4e-07 $layer=LI1_cond $X=10.895 $Y=1.177
+ $X2=10.755 $Y2=1.177
r94 28 53 0.703326 $w=2.03e-07 $l=1.3e-08 $layer=LI1_cond $X=10.742 $Y=1.177
+ $X2=10.755 $Y2=1.177
r95 28 47 14.1747 $w=2.03e-07 $l=2.62e-07 $layer=LI1_cond $X=10.742 $Y=1.177
+ $X2=10.48 $Y2=1.177
r96 28 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.87
+ $Y=1.16 $X2=10.87 $Y2=1.16
r97 27 47 6.22173 $w=2.03e-07 $l=1.15e-07 $layer=LI1_cond $X=10.365 $Y=1.177
+ $X2=10.48 $Y2=1.177
r98 26 27 23.8049 $w=2.03e-07 $l=4.4e-07 $layer=LI1_cond $X=9.925 $Y=1.177
+ $X2=10.365 $Y2=1.177
r99 26 60 1.62306 $w=2.03e-07 $l=3e-08 $layer=LI1_cond $X=9.925 $Y=1.177
+ $X2=9.895 $Y2=1.177
r100 25 58 0.27051 $w=2.03e-07 $l=5e-09 $layer=LI1_cond $X=9.43 $Y=1.177
+ $X2=9.435 $Y2=1.177
r101 25 40 6.49224 $w=2.03e-07 $l=1.2e-07 $layer=LI1_cond $X=9.43 $Y=1.177
+ $X2=9.31 $Y2=1.177
r102 22 49 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.68 $Y=0.995
+ $X2=10.68 $Y2=1.202
r103 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.68 $Y=0.995
+ $X2=10.68 $Y2=0.56
r104 19 48 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.655 $Y=1.41
+ $X2=10.655 $Y2=1.202
r105 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.655 $Y=1.41
+ $X2=10.655 $Y2=1.985
r106 16 44 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.185 $Y=1.41
+ $X2=10.185 $Y2=1.202
r107 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.185 $Y=1.41
+ $X2=10.185 $Y2=1.985
r108 13 43 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.16 $Y=0.995
+ $X2=10.16 $Y2=1.202
r109 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.16 $Y=0.995
+ $X2=10.16 $Y2=0.56
r110 10 42 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.715 $Y=1.41
+ $X2=9.715 $Y2=1.202
r111 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.715 $Y=1.41
+ $X2=9.715 $Y2=1.985
r112 7 41 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.69 $Y=0.995
+ $X2=9.69 $Y2=1.202
r113 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.69 $Y=0.995
+ $X2=9.69 $Y2=0.56
r114 4 37 18.9685 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.245 $Y=1.41
+ $X2=9.245 $Y2=1.202
r115 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.245 $Y=1.41
+ $X2=9.245 $Y2=1.985
r116 1 36 23.3057 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.22 $Y=0.995
+ $X2=9.22 $Y2=1.202
r117 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.22 $Y=0.995
+ $X2=9.22 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_297# 1 2 3 4 5 6 7 8 9 10 11 34 45 46
+ 47 50 52 56 58 62 64 68 70 74 76 80 84 85 86 87 88
r125 78 80 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.89 $Y=1.745
+ $X2=10.89 $Y2=1.96
r126 77 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.035 $Y=1.66
+ $X2=9.95 $Y2=1.66
r127 76 78 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.805 $Y=1.66
+ $X2=10.89 $Y2=1.745
r128 76 77 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=10.805 $Y=1.66
+ $X2=10.035 $Y2=1.66
r129 72 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.95 $Y=1.745
+ $X2=9.95 $Y2=1.66
r130 72 74 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.95 $Y=1.745
+ $X2=9.95 $Y2=1.96
r131 71 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.575 $Y=1.66
+ $X2=8.49 $Y2=1.66
r132 70 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.865 $Y=1.66
+ $X2=9.95 $Y2=1.66
r133 70 71 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.865 $Y=1.66
+ $X2=8.575 $Y2=1.66
r134 66 87 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.49 $Y=1.745
+ $X2=8.49 $Y2=1.66
r135 66 68 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=8.49 $Y=1.745
+ $X2=8.49 $Y2=1.96
r136 65 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.635 $Y=1.66
+ $X2=7.55 $Y2=1.66
r137 64 87 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=1.66
+ $X2=8.49 $Y2=1.66
r138 64 65 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=8.405 $Y=1.66
+ $X2=7.635 $Y2=1.66
r139 60 86 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.55 $Y=1.745
+ $X2=7.55 $Y2=1.66
r140 60 62 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.55 $Y=1.745
+ $X2=7.55 $Y2=1.96
r141 59 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.46 $Y=1.66
+ $X2=6.375 $Y2=1.66
r142 58 86 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.465 $Y=1.66
+ $X2=7.55 $Y2=1.66
r143 58 59 65.5668 $w=1.68e-07 $l=1.005e-06 $layer=LI1_cond $X=7.465 $Y=1.66
+ $X2=6.46 $Y2=1.66
r144 54 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.375 $Y=1.745
+ $X2=6.375 $Y2=1.66
r145 54 56 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=6.375 $Y=1.745
+ $X2=6.375 $Y2=1.96
r146 53 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.065 $Y=1.66
+ $X2=4.98 $Y2=1.66
r147 52 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.29 $Y=1.66
+ $X2=6.375 $Y2=1.66
r148 52 53 79.9198 $w=1.68e-07 $l=1.225e-06 $layer=LI1_cond $X=6.29 $Y=1.66
+ $X2=5.065 $Y2=1.66
r149 48 84 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.98 $Y=1.745
+ $X2=4.98 $Y2=1.66
r150 48 50 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.98 $Y=1.745
+ $X2=4.98 $Y2=1.96
r151 46 84 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.895 $Y=1.66
+ $X2=4.98 $Y2=1.66
r152 46 47 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=4.895 $Y=1.66
+ $X2=4.105 $Y2=1.66
r153 45 83 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.255
+ $X2=4.02 $Y2=2.34
r154 44 47 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.02 $Y=1.745
+ $X2=4.105 $Y2=1.66
r155 44 45 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=4.02 $Y=1.745
+ $X2=4.02 $Y2=2.255
r156 41 43 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.14 $Y=2.34
+ $X2=3.08 $Y2=2.34
r157 39 41 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=2.34
+ $X2=2.14 $Y2=2.34
r158 36 39 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=1.2 $Y2=2.34
r159 34 83 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=2.34
+ $X2=4.02 $Y2=2.34
r160 34 43 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=3.935 $Y=2.34
+ $X2=3.08 $Y2=2.34
r161 11 80 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=10.745
+ $Y=1.485 $X2=10.89 $Y2=1.96
r162 10 74 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.805
+ $Y=1.485 $X2=9.95 $Y2=1.96
r163 9 68 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.345
+ $Y=1.485 $X2=8.49 $Y2=1.96
r164 8 62 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.405
+ $Y=1.485 $X2=7.55 $Y2=1.96
r165 7 56 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.23
+ $Y=1.485 $X2=6.375 $Y2=1.96
r166 6 50 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.835
+ $Y=1.485 $X2=4.98 $Y2=1.96
r167 5 83 600 $w=1.7e-07 $l=8.44393e-07 $layer=licon1_PDIFF $count=1 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2.26
r168 4 43 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2.34
r169 3 41 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.34
r170 2 39 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r171 1 36 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%Y 1 2 3 4 5 6 7 8 25 27 29 37 39 42 47 53
+ 55 56 57 68 71 73
c102 29 0 1.16491e-19 $X=2.505 $Y=0.805
r103 68 76 1.17863 $w=4.38e-07 $l=4.5e-08 $layer=LI1_cond $X=2.395 $Y=1.53
+ $X2=2.395 $Y2=1.575
r104 63 73 0.523838 $w=4.38e-07 $l=2e-08 $layer=LI1_cond $X=2.395 $Y=1.21
+ $X2=2.395 $Y2=1.19
r105 57 78 4.18627 $w=5.98e-07 $l=2.1e-07 $layer=LI1_cond $X=2.475 $Y=1.87
+ $X2=2.475 $Y2=1.66
r106 56 78 1.29575 $w=5.98e-07 $l=6.5e-08 $layer=LI1_cond $X=2.475 $Y=1.595
+ $X2=2.475 $Y2=1.66
r107 56 76 1.27213 $w=5.98e-07 $l=2e-08 $layer=LI1_cond $X=2.475 $Y=1.595
+ $X2=2.475 $Y2=1.575
r108 56 68 0.523838 $w=4.38e-07 $l=2e-08 $layer=LI1_cond $X=2.395 $Y=1.51
+ $X2=2.395 $Y2=1.53
r109 55 73 0.864332 $w=4.38e-07 $l=3.3e-08 $layer=LI1_cond $X=2.395 $Y=1.157
+ $X2=2.395 $Y2=1.19
r110 55 71 7.25322 $w=4.38e-07 $l=1.67e-07 $layer=LI1_cond $X=2.395 $Y=1.157
+ $X2=2.395 $Y2=0.99
r111 55 56 7.01943 $w=4.38e-07 $l=2.68e-07 $layer=LI1_cond $X=2.395 $Y=1.242
+ $X2=2.395 $Y2=1.51
r112 55 63 0.83814 $w=4.38e-07 $l=3.2e-08 $layer=LI1_cond $X=2.395 $Y=1.242
+ $X2=2.395 $Y2=1.21
r113 40 78 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=2.775 $Y=1.66
+ $X2=2.475 $Y2=1.66
r114 39 53 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.335 $Y=1.66
+ $X2=3.525 $Y2=1.66
r115 39 40 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.335 $Y=1.66
+ $X2=2.775 $Y2=1.66
r116 35 37 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.06 $Y=0.72 $X2=6
+ $Y2=0.72
r117 33 35 98.5134 $w=1.68e-07 $l=1.51e-06 $layer=LI1_cond $X=3.55 $Y=0.72
+ $X2=5.06 $Y2=0.72
r118 31 50 3.92798 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=2.615 $Y=0.72
+ $X2=2.505 $Y2=0.72
r119 31 33 61 $w=1.68e-07 $l=9.35e-07 $layer=LI1_cond $X=2.615 $Y=0.72 $X2=3.55
+ $Y2=0.72
r120 29 50 3.03526 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=2.505 $Y=0.805
+ $X2=2.505 $Y2=0.72
r121 29 71 9.691 $w=2.18e-07 $l=1.85e-07 $layer=LI1_cond $X=2.505 $Y=0.805
+ $X2=2.505 $Y2=0.99
r122 28 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.66
+ $X2=1.645 $Y2=1.66
r123 27 78 8.31678 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=2.175 $Y=1.66
+ $X2=2.475 $Y2=1.66
r124 27 28 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.175 $Y=1.66
+ $X2=1.835 $Y2=1.66
r125 26 42 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.66
+ $X2=0.705 $Y2=1.66
r126 25 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.66
+ $X2=1.645 $Y2=1.66
r127 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.66
+ $X2=0.895 $Y2=1.66
r128 8 53 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r129 7 78 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r130 6 47 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r131 5 42 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r132 4 37 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.865
+ $Y=0.235 $X2=6 $Y2=0.72
r133 3 35 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.925
+ $Y=0.235 $X2=5.06 $Y2=0.72
r134 2 33 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.72
r135 1 50 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%VPWR 1 2 3 4 5 6 21 25 29 33 37 39 41 46
+ 51 56 61 66 71 74 76 79 86 89 92 95
r131 95 96 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r132 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r133 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r134 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r135 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r136 79 82 11.9608 $w=7.18e-07 $l=7.2e-07 $layer=LI1_cond $X=5.68 $Y=2 $X2=5.68
+ $Y2=2.72
r137 76 77 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 74 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=10.35 $Y2=2.72
r139 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r140 71 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.585 $Y=2.72
+ $X2=10.395 $Y2=2.72
r141 71 73 16.1471 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=10.585 $Y=2.72
+ $X2=10.81 $Y2=2.72
r142 70 96 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r143 70 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r144 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r145 67 92 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.645 $Y=2.72
+ $X2=9.455 $Y2=2.72
r146 67 69 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=9.645 $Y=2.72
+ $X2=9.89 $Y2=2.72
r147 66 95 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.205 $Y=2.72
+ $X2=10.395 $Y2=2.72
r148 66 69 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.205 $Y=2.72
+ $X2=9.89 $Y2=2.72
r149 65 93 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r150 65 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.05 $Y2=2.72
r151 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r152 62 89 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.185 $Y=2.72
+ $X2=7.995 $Y2=2.72
r153 62 64 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=8.185 $Y=2.72
+ $X2=8.97 $Y2=2.72
r154 61 92 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=9.455 $Y2=2.72
r155 61 64 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.265 $Y=2.72
+ $X2=8.97 $Y2=2.72
r156 60 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r157 60 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r158 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r159 57 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.245 $Y=2.72
+ $X2=7.055 $Y2=2.72
r160 57 59 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=7.245 $Y=2.72
+ $X2=7.59 $Y2=2.72
r161 56 89 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.805 $Y=2.72
+ $X2=7.995 $Y2=2.72
r162 56 59 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.805 $Y=2.72
+ $X2=7.59 $Y2=2.72
r163 55 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r164 55 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=5.75 $Y2=2.72
r165 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r166 52 82 9.50744 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=6.04 $Y=2.72
+ $X2=5.68 $Y2=2.72
r167 52 54 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.04 $Y=2.72
+ $X2=6.67 $Y2=2.72
r168 51 86 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.865 $Y=2.72
+ $X2=7.055 $Y2=2.72
r169 51 54 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.865 $Y=2.72
+ $X2=6.67 $Y2=2.72
r170 50 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r171 50 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r172 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r173 47 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=4.485 $Y2=2.72
r174 47 49 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=4.675 $Y=2.72
+ $X2=5.29 $Y2=2.72
r175 46 82 9.50744 $w=1.7e-07 $l=3.6e-07 $layer=LI1_cond $X=5.32 $Y=2.72
+ $X2=5.68 $Y2=2.72
r176 46 49 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.32 $Y=2.72 $X2=5.29
+ $Y2=2.72
r177 41 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=4.485 $Y2=2.72
r178 41 43 265.203 $w=1.68e-07 $l=4.065e-06 $layer=LI1_cond $X=4.295 $Y=2.72
+ $X2=0.23 $Y2=2.72
r179 39 77 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=4.37 $Y2=2.72
r180 39 43 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r181 35 95 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.395 $Y=2.635
+ $X2=10.395 $Y2=2.72
r182 35 37 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=10.395 $Y=2.635
+ $X2=10.395 $Y2=2
r183 31 92 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.455 $Y=2.635
+ $X2=9.455 $Y2=2.72
r184 31 33 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=9.455 $Y=2.635
+ $X2=9.455 $Y2=2
r185 27 89 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.995 $Y=2.635
+ $X2=7.995 $Y2=2.72
r186 27 29 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=7.995 $Y=2.635
+ $X2=7.995 $Y2=2.34
r187 23 86 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.055 $Y=2.635
+ $X2=7.055 $Y2=2.72
r188 23 25 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=7.055 $Y=2.635
+ $X2=7.055 $Y2=2
r189 19 76 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.485 $Y=2.635
+ $X2=4.485 $Y2=2.72
r190 19 21 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=4.485 $Y=2.635
+ $X2=4.485 $Y2=2
r191 6 37 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.275
+ $Y=1.485 $X2=10.42 $Y2=2
r192 5 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.335
+ $Y=1.485 $X2=9.48 $Y2=2
r193 4 29 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.875
+ $Y=1.485 $X2=8.02 $Y2=2.34
r194 3 25 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.935
+ $Y=1.485 $X2=7.08 $Y2=2
r195 2 79 150 $w=1.7e-07 $l=7.33621e-07 $layer=licon1_PDIFF $count=4 $X=5.305
+ $Y=1.485 $X2=5.825 $Y2=2
r196 1 21 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.365
+ $Y=1.485 $X2=4.51 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A_27_47# 1 2 3 4 5 18 20 21 24 26 28 34 36
r56 32 34 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.08 $Y=0.38
+ $X2=4.02 $Y2=0.38
r57 30 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.38
+ $X2=2.14 $Y2=0.38
r58 30 32 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.38
+ $X2=3.08 $Y2=0.38
r59 28 38 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.465
+ $X2=2.14 $Y2=0.38
r60 28 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.14 $Y=0.465
+ $X2=2.14 $Y2=0.635
r61 27 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.72 $X2=1.2
+ $Y2=0.72
r62 26 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=2.14 $Y2=0.635
r63 26 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0.72
+ $X2=1.285 $Y2=0.72
r64 22 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.635 $X2=1.2
+ $Y2=0.72
r65 22 24 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.2 $Y=0.635
+ $X2=1.2 $Y2=0.42
r66 20 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0.72 $X2=1.2
+ $Y2=0.72
r67 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0.72
+ $X2=0.345 $Y2=0.72
r68 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r69 16 18 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.42
r70 5 34 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.38
r71 4 32 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.38
r72 3 38 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.46
r73 2 24 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.42
r74 1 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%VGND 1 2 3 4 5 18 22 24 29 34 42 47 54 61
+ 67 71 78 79
r131 78 81 11.2289 $w=3.88e-07 $l=3.8e-07 $layer=LI1_cond $X=10.88 $Y=0
+ $X2=10.88 $Y2=0.38
r132 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r133 71 74 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=9.925 $Y=0
+ $X2=9.925 $Y2=0.38
r134 71 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r135 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r136 61 64 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.645 $Y=0
+ $X2=1.645 $Y2=0.38
r137 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r138 54 57 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r139 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r140 51 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r141 51 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=9.89 $Y2=0
r142 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r143 48 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=9.925 $Y2=0
r144 48 50 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=10.115 $Y=0
+ $X2=10.35 $Y2=0
r145 47 78 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=10.685 $Y=0
+ $X2=10.88 $Y2=0
r146 47 50 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=10.685 $Y=0
+ $X2=10.35 $Y2=0
r147 46 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=9.89
+ $Y2=0
r148 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.97
+ $Y2=0
r149 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r150 43 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.175 $Y=0 $X2=9.01
+ $Y2=0
r151 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=9.175 $Y=0
+ $X2=9.43 $Y2=0
r152 42 71 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.735 $Y=0 $X2=9.925
+ $Y2=0
r153 42 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.735 $Y=0
+ $X2=9.43 $Y2=0
r154 41 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0 $X2=8.97
+ $Y2=0
r155 40 41 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r156 38 41 1.83245 $w=4.8e-07 $l=6.44e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=8.51
+ $Y2=0
r157 38 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r158 37 40 420.15 $w=1.68e-07 $l=6.44e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=8.51
+ $Y2=0
r159 37 38 1.24 $w=1.7e-07 $l=1.275e-06 $layer=mcon $count=7 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r160 35 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.645
+ $Y2=0
r161 35 37 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=1.835 $Y=0
+ $X2=2.07 $Y2=0
r162 34 67 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.845 $Y=0 $X2=9.01
+ $Y2=0
r163 34 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=8.845 $Y=0
+ $X2=8.51 $Y2=0
r164 33 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r165 33 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r166 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r167 30 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r168 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r169 29 61 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0 $X2=1.645
+ $Y2=0
r170 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=0
+ $X2=1.15 $Y2=0
r171 24 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r172 24 26 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r173 22 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r174 22 26 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r175 16 67 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0
r176 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=9.01 $Y=0.085
+ $X2=9.01 $Y2=0.38
r177 5 81 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=10.755
+ $Y=0.235 $X2=10.9 $Y2=0.38
r178 4 74 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=9.765
+ $Y=0.235 $X2=9.95 $Y2=0.38
r179 3 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=8.885
+ $Y=0.235 $X2=9.01 $Y2=0.38
r180 2 64 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r181 1 57 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A_893_47# 1 2 3 4 5 26
r29 24 26 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.55 $Y=0.38
+ $X2=8.49 $Y2=0.38
r30 22 24 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=6.47 $Y=0.38
+ $X2=7.55 $Y2=0.38
r31 20 22 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=5.53 $Y=0.38
+ $X2=6.47 $Y2=0.38
r32 17 20 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=4.59 $Y=0.38
+ $X2=5.53 $Y2=0.38
r33 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.355
+ $Y=0.235 $X2=8.49 $Y2=0.38
r34 4 24 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.365
+ $Y=0.235 $X2=7.55 $Y2=0.38
r35 3 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.47 $Y2=0.38
r36 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.395
+ $Y=0.235 $X2=5.53 $Y2=0.38
r37 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.465
+ $Y=0.235 $X2=4.59 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_4%A_1379_47# 1 2 3 4 13 21 23 27 29
r47 25 27 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=10.42 $Y=0.635
+ $X2=10.42 $Y2=0.42
r48 24 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.565 $Y=0.72
+ $X2=9.48 $Y2=0.72
r49 23 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.335 $Y=0.72
+ $X2=10.42 $Y2=0.635
r50 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=10.335 $Y=0.72
+ $X2=9.565 $Y2=0.72
r51 19 29 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.48 $Y=0.635
+ $X2=9.48 $Y2=0.72
r52 19 21 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=9.48 $Y=0.635
+ $X2=9.48 $Y2=0.42
r53 15 18 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=7.08 $Y=0.72
+ $X2=8.02 $Y2=0.72
r54 13 29 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.395 $Y=0.72
+ $X2=9.48 $Y2=0.72
r55 13 18 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=9.395 $Y=0.72
+ $X2=8.02 $Y2=0.72
r56 4 27 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=10.235
+ $Y=0.235 $X2=10.42 $Y2=0.42
r57 3 21 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.235 $X2=9.48 $Y2=0.42
r58 2 18 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=7.835
+ $Y=0.235 $X2=8.02 $Y2=0.72
r59 1 15 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=6.895
+ $Y=0.235 $X2=7.08 $Y2=0.72
.ends

