* File: sky130_fd_sc_hdll__o31ai_4.pex.spice
* Created: Wed Sep  2 08:46:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A1 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 54 61 66 70
c88 70 0 1.155e-20 $X=1.78 $Y=1.19
c89 22 0 1.07883e-19 $X=1.925 $Y=1.41
r90 54 55 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.217
+ $X2=1.95 $Y2=1.217
r91 52 54 23.5841 $w=3.27e-07 $l=1.6e-07 $layer=POLY_cond $X=1.765 $Y=1.217
+ $X2=1.925 $Y2=1.217
r92 50 52 45.6942 $w=3.27e-07 $l=3.1e-07 $layer=POLY_cond $X=1.455 $Y=1.217
+ $X2=1.765 $Y2=1.217
r93 49 50 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.217
+ $X2=1.455 $Y2=1.217
r94 48 66 3.42618 $w=3.68e-07 $l=1.1e-07 $layer=LI1_cond $X=1.375 $Y=1.24
+ $X2=1.265 $Y2=1.24
r95 47 49 8.10703 $w=3.27e-07 $l=5.5e-08 $layer=POLY_cond $X=1.375 $Y=1.217
+ $X2=1.43 $Y2=1.217
r96 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.375
+ $Y=1.16 $X2=1.375 $Y2=1.16
r97 44 47 57.4862 $w=3.27e-07 $l=3.9e-07 $layer=POLY_cond $X=0.985 $Y=1.217
+ $X2=1.375 $Y2=1.217
r98 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.985
+ $Y=1.16 $X2=0.985 $Y2=1.16
r99 42 44 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.217
+ $X2=0.985 $Y2=1.217
r100 41 61 3.11471 $w=3.68e-07 $l=1e-07 $layer=LI1_cond $X=0.595 $Y=1.24
+ $X2=0.695 $Y2=1.24
r101 40 42 53.8012 $w=3.27e-07 $l=3.65e-07 $layer=POLY_cond $X=0.595 $Y=1.217
+ $X2=0.96 $Y2=1.217
r102 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r103 38 40 11.792 $w=3.27e-07 $l=8e-08 $layer=POLY_cond $X=0.515 $Y=1.217
+ $X2=0.595 $Y2=1.217
r104 37 38 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.217
+ $X2=0.515 $Y2=1.217
r105 32 70 0.467207 $w=3.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.765 $Y=1.24
+ $X2=1.78 $Y2=1.24
r106 32 48 12.1474 $w=3.68e-07 $l=3.9e-07 $layer=LI1_cond $X=1.765 $Y=1.24
+ $X2=1.375 $Y2=1.24
r107 32 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.765
+ $Y=1.16 $X2=1.765 $Y2=1.16
r108 31 66 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=1.255 $Y=1.24
+ $X2=1.265 $Y2=1.24
r109 31 45 8.40972 $w=3.68e-07 $l=2.7e-07 $layer=LI1_cond $X=1.255 $Y=1.24
+ $X2=0.985 $Y2=1.24
r110 30 45 7.47531 $w=3.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.745 $Y=1.24
+ $X2=0.985 $Y2=1.24
r111 30 61 1.55736 $w=3.68e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.24
+ $X2=0.695 $Y2=1.24
r112 29 41 11.213 $w=3.68e-07 $l=3.6e-07 $layer=LI1_cond $X=0.235 $Y=1.24
+ $X2=0.595 $Y2=1.24
r113 25 55 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.95 $Y=1.025
+ $X2=1.95 $Y2=1.217
r114 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.95 $Y=1.025
+ $X2=1.95 $Y2=0.56
r115 22 54 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.217
r116 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r117 19 50 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.217
r118 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r119 15 49 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.43 $Y=1.025
+ $X2=1.43 $Y2=1.217
r120 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.43 $Y=1.025
+ $X2=1.43 $Y2=0.56
r121 12 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.217
r122 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r123 8 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.96 $Y=1.025
+ $X2=0.96 $Y2=1.217
r124 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.96 $Y=1.025
+ $X2=0.96 $Y2=0.56
r125 5 38 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.217
r126 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r127 1 37 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=1.217
r128 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.49 $Y=1.025
+ $X2=0.49 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A2 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 55 58 64 66 70
c92 32 0 1.07883e-19 $X=3.72 $Y=1.105
c93 5 0 1.155e-20 $X=2.395 $Y=1.41
r94 64 66 13.8605 $w=3.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.795 $Y=1.24
+ $X2=3.24 $Y2=1.24
r95 55 56 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.805 $Y=1.217
+ $X2=3.83 $Y2=1.217
r96 54 70 3.73765 $w=3.68e-07 $l=1.2e-07 $layer=LI1_cond $X=3.63 $Y=1.24
+ $X2=3.75 $Y2=1.24
r97 53 55 25.7951 $w=3.27e-07 $l=1.75e-07 $layer=POLY_cond $X=3.63 $Y=1.217
+ $X2=3.805 $Y2=1.217
r98 53 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.63
+ $Y=1.16 $X2=3.63 $Y2=1.16
r99 51 53 43.4832 $w=3.27e-07 $l=2.95e-07 $layer=POLY_cond $X=3.335 $Y=1.217
+ $X2=3.63 $Y2=1.217
r100 50 51 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.31 $Y=1.217
+ $X2=3.335 $Y2=1.217
r101 48 50 10.318 $w=3.27e-07 $l=7e-08 $layer=POLY_cond $X=3.24 $Y=1.217
+ $X2=3.31 $Y2=1.217
r102 48 66 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.24
+ $Y=1.16 $X2=3.24 $Y2=1.16
r103 46 48 55.2752 $w=3.27e-07 $l=3.75e-07 $layer=POLY_cond $X=2.865 $Y=1.217
+ $X2=3.24 $Y2=1.217
r104 44 46 2.21101 $w=3.27e-07 $l=1.5e-08 $layer=POLY_cond $X=2.85 $Y=1.217
+ $X2=2.865 $Y2=1.217
r105 44 64 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.85
+ $Y=1.16 $X2=2.85 $Y2=1.16
r106 42 44 1.47401 $w=3.27e-07 $l=1e-08 $layer=POLY_cond $X=2.84 $Y=1.217
+ $X2=2.85 $Y2=1.217
r107 40 42 56.0122 $w=3.27e-07 $l=3.8e-07 $layer=POLY_cond $X=2.46 $Y=1.217
+ $X2=2.84 $Y2=1.217
r108 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.46
+ $Y=1.16 $X2=2.46 $Y2=1.16
r109 38 40 9.58104 $w=3.27e-07 $l=6.5e-08 $layer=POLY_cond $X=2.395 $Y=1.217
+ $X2=2.46 $Y2=1.217
r110 37 38 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.37 $Y=1.217
+ $X2=2.395 $Y2=1.217
r111 32 70 1.71309 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.805 $Y=1.24
+ $X2=3.75 $Y2=1.24
r112 31 54 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.295 $Y=1.24
+ $X2=3.63 $Y2=1.24
r113 31 66 1.71309 $w=3.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.295 $Y=1.24
+ $X2=3.24 $Y2=1.24
r114 30 64 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=2.785 $Y=1.24
+ $X2=2.795 $Y2=1.24
r115 30 41 10.1228 $w=3.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.785 $Y=1.24
+ $X2=2.46 $Y2=1.24
r116 29 41 5.76222 $w=3.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.275 $Y=1.24
+ $X2=2.46 $Y2=1.24
r117 29 58 0.311471 $w=3.68e-07 $l=1e-08 $layer=LI1_cond $X=2.275 $Y=1.24
+ $X2=2.265 $Y2=1.24
r118 25 56 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=1.217
r119 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.83 $Y=1.025
+ $X2=3.83 $Y2=0.56
r120 22 55 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.217
r121 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.805 $Y=1.41
+ $X2=3.805 $Y2=1.985
r122 19 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.217
r123 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.335 $Y=1.41
+ $X2=3.335 $Y2=1.985
r124 15 50 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.31 $Y=1.025
+ $X2=3.31 $Y2=1.217
r125 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.31 $Y=1.025
+ $X2=3.31 $Y2=0.56
r126 12 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.217
r127 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.865 $Y=1.41
+ $X2=2.865 $Y2=1.985
r128 8 42 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.84 $Y=1.025
+ $X2=2.84 $Y2=1.217
r129 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.84 $Y=1.025
+ $X2=2.84 $Y2=0.56
r130 5 38 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.217
r131 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.395 $Y=1.41
+ $X2=2.395 $Y2=1.985
r132 1 37 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.37 $Y=1.025
+ $X2=2.37 $Y2=1.217
r133 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.37 $Y=1.025
+ $X2=2.37 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A3 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 32 33 34 40 52 57 60 62 65 69
c73 27 0 1.07318e-19 $X=6.295 $Y=0.56
c74 22 0 1.73812e-19 $X=6.27 $Y=1.41
r75 60 62 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=4.83 $Y=1.165
+ $X2=5.29 $Y2=1.165
r76 52 53 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.27 $Y=1.217
+ $X2=6.295 $Y2=1.217
r77 50 52 54.5382 $w=3.27e-07 $l=3.7e-07 $layer=POLY_cond $X=5.9 $Y=1.217
+ $X2=6.27 $Y2=1.217
r78 48 50 14.7401 $w=3.27e-07 $l=1e-07 $layer=POLY_cond $X=5.8 $Y=1.217 $X2=5.9
+ $Y2=1.217
r79 47 48 21.3731 $w=3.27e-07 $l=1.45e-07 $layer=POLY_cond $X=5.655 $Y=1.217
+ $X2=5.8 $Y2=1.217
r80 46 47 47.9052 $w=3.27e-07 $l=3.25e-07 $layer=POLY_cond $X=5.33 $Y=1.217
+ $X2=5.655 $Y2=1.217
r81 45 46 21.3731 $w=3.27e-07 $l=1.45e-07 $layer=POLY_cond $X=5.185 $Y=1.217
+ $X2=5.33 $Y2=1.217
r82 44 45 47.9052 $w=3.27e-07 $l=3.25e-07 $layer=POLY_cond $X=4.86 $Y=1.217
+ $X2=5.185 $Y2=1.217
r83 40 44 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=4.76 $Y=1.16
+ $X2=4.86 $Y2=1.217
r84 40 42 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=4.76 $Y=1.16 $X2=4.34
+ $Y2=1.16
r85 34 69 0.261919 $w=2.18e-07 $l=5e-09 $layer=LI1_cond $X=6.35 $Y=1.165
+ $X2=6.355 $Y2=1.165
r86 33 34 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=5.89 $Y=1.165
+ $X2=6.35 $Y2=1.165
r87 33 65 0.785757 $w=2.18e-07 $l=1.5e-08 $layer=LI1_cond $X=5.89 $Y=1.165
+ $X2=5.875 $Y2=1.165
r88 33 50 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=5.9
+ $Y=1.16 $X2=5.9 $Y2=1.16
r89 32 65 28.5492 $w=2.18e-07 $l=5.45e-07 $layer=LI1_cond $X=5.33 $Y=1.165
+ $X2=5.875 $Y2=1.165
r90 32 62 2.09535 $w=2.18e-07 $l=4e-08 $layer=LI1_cond $X=5.33 $Y=1.165 $X2=5.29
+ $Y2=1.165
r91 31 60 0.523838 $w=2.18e-07 $l=1e-08 $layer=LI1_cond $X=4.82 $Y=1.165
+ $X2=4.83 $Y2=1.165
r92 31 57 23.5727 $w=2.18e-07 $l=4.5e-07 $layer=LI1_cond $X=4.82 $Y=1.165
+ $X2=4.37 $Y2=1.165
r93 30 57 1.57151 $w=2.18e-07 $l=3e-08 $layer=LI1_cond $X=4.34 $Y=1.165 $X2=4.37
+ $Y2=1.165
r94 30 42 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=4.34
+ $Y=1.16 $X2=4.34 $Y2=1.16
r95 29 42 3.33261 $w=2.7e-07 $l=1.5e-08 $layer=POLY_cond $X=4.325 $Y=1.16
+ $X2=4.34 $Y2=1.16
r96 25 53 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.295 $Y=1.025
+ $X2=6.295 $Y2=1.217
r97 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.295 $Y=1.025
+ $X2=6.295 $Y2=0.56
r98 22 52 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.27 $Y=1.41
+ $X2=6.27 $Y2=1.217
r99 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.27 $Y=1.41
+ $X2=6.27 $Y2=1.985
r100 19 48 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.8 $Y=1.41
+ $X2=5.8 $Y2=1.217
r101 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.8 $Y=1.41
+ $X2=5.8 $Y2=1.985
r102 15 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.655 $Y=1.025
+ $X2=5.655 $Y2=1.217
r103 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.655 $Y=1.025
+ $X2=5.655 $Y2=0.56
r104 12 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.33 $Y=1.41
+ $X2=5.33 $Y2=1.217
r105 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.33 $Y=1.41
+ $X2=5.33 $Y2=1.985
r106 8 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.185 $Y=1.025
+ $X2=5.185 $Y2=1.217
r107 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.185 $Y=1.025
+ $X2=5.185 $Y2=0.56
r108 5 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.217
r109 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.86 $Y=1.41
+ $X2=4.86 $Y2=1.985
r110 1 29 29.8935 $w=2.7e-07 $l=1.68375e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.325 $Y2=1.16
r111 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.25 $Y=1.025
+ $X2=4.25 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%B1 3 5 7 10 12 14 17 19 21 24 26 28 29 30
+ 31 47 51 55
r71 47 48 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=8.125 $Y=1.217
+ $X2=8.15 $Y2=1.217
r72 46 55 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=8.11 $Y=1.165
+ $X2=7.94 $Y2=1.165
r73 45 47 2.23148 $w=3.24e-07 $l=1.5e-08 $layer=POLY_cond $X=8.11 $Y=1.217
+ $X2=8.125 $Y2=1.217
r74 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=8.11
+ $Y=1.16 $X2=8.11 $Y2=1.16
r75 43 45 63.9691 $w=3.24e-07 $l=4.3e-07 $layer=POLY_cond $X=7.68 $Y=1.217
+ $X2=8.11 $Y2=1.217
r76 42 43 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=7.655 $Y=1.217
+ $X2=7.68 $Y2=1.217
r77 40 42 48.3488 $w=3.24e-07 $l=3.25e-07 $layer=POLY_cond $X=7.33 $Y=1.217
+ $X2=7.655 $Y2=1.217
r78 40 51 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.33
+ $Y=1.16 $X2=7.33 $Y2=1.16
r79 38 40 17.8519 $w=3.24e-07 $l=1.2e-07 $layer=POLY_cond $X=7.21 $Y=1.217
+ $X2=7.33 $Y2=1.217
r80 37 38 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=7.185 $Y=1.217
+ $X2=7.21 $Y2=1.217
r81 36 37 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=6.74 $Y=1.217
+ $X2=7.185 $Y2=1.217
r82 35 36 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=6.715 $Y=1.217
+ $X2=6.74 $Y2=1.217
r83 31 46 17.2866 $w=2.18e-07 $l=3.3e-07 $layer=LI1_cond $X=8.44 $Y=1.165
+ $X2=8.11 $Y2=1.165
r84 30 55 0.523838 $w=2.18e-07 $l=1e-08 $layer=LI1_cond $X=7.93 $Y=1.165
+ $X2=7.94 $Y2=1.165
r85 29 30 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=7.42 $Y=1.165
+ $X2=7.93 $Y2=1.165
r86 29 51 4.71454 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=7.42 $Y=1.165 $X2=7.33
+ $Y2=1.165
r87 26 48 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.217
r88 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.15 $Y=1.41
+ $X2=8.15 $Y2=1.985
r89 22 47 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.125 $Y=1.025
+ $X2=8.125 $Y2=1.217
r90 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.125 $Y=1.025
+ $X2=8.125 $Y2=0.56
r91 19 43 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.68 $Y=1.41
+ $X2=7.68 $Y2=1.217
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.68 $Y=1.41
+ $X2=7.68 $Y2=1.985
r93 15 42 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.655 $Y=1.025
+ $X2=7.655 $Y2=1.217
r94 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.655 $Y=1.025
+ $X2=7.655 $Y2=0.56
r95 12 38 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.21 $Y=1.41
+ $X2=7.21 $Y2=1.217
r96 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.21 $Y=1.41
+ $X2=7.21 $Y2=1.985
r97 8 37 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.185 $Y=1.025
+ $X2=7.185 $Y2=1.217
r98 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.185 $Y=1.025
+ $X2=7.185 $Y2=0.56
r99 5 36 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.74 $Y=1.41
+ $X2=6.74 $Y2=1.217
r100 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.74 $Y=1.41
+ $X2=6.74 $Y2=1.985
r101 1 35 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.715 $Y=1.025
+ $X2=6.715 $Y2=1.217
r102 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.715 $Y=1.025
+ $X2=6.715 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 28 29
+ 30 34 39 45
r82 45 47 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=3.075 $Y=2.02
+ $X2=3.075 $Y2=2.335
r83 32 47 2.9592 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=3.265 $Y=2.335
+ $X2=3.075 $Y2=2.335
r84 32 34 34.3517 $w=2.58e-07 $l=7.75e-07 $layer=LI1_cond $X=3.265 $Y=2.335
+ $X2=4.04 $Y2=2.335
r85 31 43 4.23515 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=2.335
+ $X2=2.135 $Y2=2.335
r86 30 47 2.9592 $w=2.6e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=2.335
+ $X2=3.075 $Y2=2.335
r87 30 31 24.8218 $w=2.58e-07 $l=5.6e-07 $layer=LI1_cond $X=2.885 $Y=2.335
+ $X2=2.325 $Y2=2.335
r88 29 43 2.89773 $w=3.8e-07 $l=1.3e-07 $layer=LI1_cond $X=2.135 $Y=2.205
+ $X2=2.135 $Y2=2.335
r89 28 41 3.06173 $w=3.8e-07 $l=1.5e-07 $layer=LI1_cond $X=2.135 $Y=1.895
+ $X2=2.135 $Y2=1.745
r90 28 29 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=2.135 $Y=1.895
+ $X2=2.135 $Y2=2.205
r91 27 39 6.25931 $w=3e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=1.745
+ $X2=1.195 $Y2=1.745
r92 26 41 3.87819 $w=3e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=1.745
+ $X2=2.135 $Y2=1.745
r93 26 27 21.5123 $w=2.98e-07 $l=5.6e-07 $layer=LI1_cond $X=1.945 $Y=1.745
+ $X2=1.385 $Y2=1.745
r94 22 39 0.506867 $w=3.8e-07 $l=1.5e-07 $layer=LI1_cond $X=1.195 $Y=1.895
+ $X2=1.195 $Y2=1.745
r95 22 24 14.1023 $w=3.78e-07 $l=4.65e-07 $layer=LI1_cond $X=1.195 $Y=1.895
+ $X2=1.195 $Y2=2.36
r96 21 37 3.73322 $w=3e-07 $l=1.78e-07 $layer=LI1_cond $X=0.445 $Y=1.745
+ $X2=0.267 $Y2=1.745
r97 20 39 6.25931 $w=3e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=1.745
+ $X2=1.195 $Y2=1.745
r98 20 21 21.5123 $w=2.98e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=1.745
+ $X2=0.445 $Y2=1.745
r99 16 37 3.14597 $w=3.55e-07 $l=1.5e-07 $layer=LI1_cond $X=0.267 $Y=1.895
+ $X2=0.267 $Y2=1.745
r100 16 18 15.0954 $w=3.53e-07 $l=4.65e-07 $layer=LI1_cond $X=0.267 $Y=1.895
+ $X2=0.267 $Y2=2.36
r101 5 34 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.895
+ $Y=1.485 $X2=4.04 $Y2=2.36
r102 4 45 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=2.955
+ $Y=1.485 $X2=3.1 $Y2=2.02
r103 3 43 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=2.36
r104 3 41 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.68
r105 2 39 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.68
r106 2 24 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.36
r107 1 37 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.68
r108 1 18 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%VPWR 1 2 3 4 17 19 23 27 31 34 35 37 38 39
+ 52 53 56 59
r112 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r113 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r116 50 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r117 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r118 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r119 46 47 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r120 44 47 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=6.67 $Y2=2.72
r121 44 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r122 43 46 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=6.67 $Y2=2.72
r123 43 44 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 41 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=1.69 $Y2=2.72
r125 41 43 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.775 $Y=2.72
+ $X2=2.07 $Y2=2.72
r126 39 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r127 37 49 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=7.7 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 37 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.7 $Y=2.72 $X2=7.89
+ $Y2=2.72
r129 36 52 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.08 $Y=2.72
+ $X2=8.51 $Y2=2.72
r130 36 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.08 $Y=2.72
+ $X2=7.89 $Y2=2.72
r131 34 46 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.76 $Y=2.72 $X2=6.67
+ $Y2=2.72
r132 34 35 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.76 $Y=2.72
+ $X2=6.95 $Y2=2.72
r133 33 49 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=7.14 $Y=2.72
+ $X2=7.59 $Y2=2.72
r134 33 35 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.14 $Y=2.72
+ $X2=6.95 $Y2=2.72
r135 29 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.89 $Y=2.635
+ $X2=7.89 $Y2=2.72
r136 29 31 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=7.89 $Y=2.635
+ $X2=7.89 $Y2=2.02
r137 25 35 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.95 $Y=2.635
+ $X2=6.95 $Y2=2.72
r138 25 27 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=6.95 $Y=2.635
+ $X2=6.95 $Y2=2.02
r139 21 59 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.72
r140 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.69 $Y=2.635
+ $X2=1.69 $Y2=2.34
r141 20 56 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.75 $Y2=2.72
r142 19 59 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=1.69 $Y2=2.72
r143 19 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.605 $Y=2.72
+ $X2=0.835 $Y2=2.72
r144 15 56 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r145 15 17 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.34
r146 4 31 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=7.77
+ $Y=1.485 $X2=7.915 $Y2=2.02
r147 3 27 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=6.83
+ $Y=1.485 $X2=6.975 $Y2=2.02
r148 2 23 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2.34
r149 1 17 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A_497_297# 1 2 3 4 17 19 23 27 28 31
r48 30 31 18.1299 $w=5.98e-07 $l=5.65e-07 $layer=LI1_cond $X=5.095 $Y=2.165
+ $X2=4.53 $Y2=2.165
r49 28 31 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=4.005 $Y=1.95
+ $X2=4.53 $Y2=1.95
r50 26 28 15.9071 $w=4.38e-07 $l=4.35e-07 $layer=LI1_cond $X=3.57 $Y=1.815
+ $X2=4.005 $Y2=1.815
r51 26 27 6.73996 $w=4.38e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=1.815
+ $X2=3.485 $Y2=1.815
r52 17 30 0.697712 $w=5.98e-07 $l=3.5e-08 $layer=LI1_cond $X=5.13 $Y=2.165
+ $X2=5.095 $Y2=2.165
r53 17 19 18.0408 $w=5.98e-07 $l=9.05e-07 $layer=LI1_cond $X=5.13 $Y=2.165
+ $X2=6.035 $Y2=2.165
r54 14 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=1.68
+ $X2=2.63 $Y2=1.68
r55 14 27 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.715 $Y=1.68
+ $X2=3.485 $Y2=1.68
r56 4 19 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=5.89
+ $Y=1.485 $X2=6.035 $Y2=1.95
r57 3 30 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=4.95
+ $Y=1.485 $X2=5.095 $Y2=1.95
r58 2 26 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=3.425
+ $Y=1.485 $X2=3.57 $Y2=1.76
r59 1 23 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=2.485
+ $Y=1.485 $X2=2.63 $Y2=1.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%Y 1 2 3 4 5 6 7 24 28 32 34 37 38 39 40 41
+ 42 43 44 45 46 47 62 66 71 73 78 82 83 84 86 90 91 103
c83 42 0 1.73812e-19 $X=6.81 $Y=1.445
c84 34 0 1.07318e-19 $X=6.877 $Y=0.885
r85 101 103 0.368782 $w=2.48e-07 $l=8e-09 $layer=LI1_cond $X=6.877 $Y=1.57
+ $X2=6.885 $Y2=1.57
r86 86 90 16.3647 $w=2.48e-07 $l=3.55e-07 $layer=LI1_cond $X=8.3 $Y=1.57
+ $X2=7.945 $Y2=1.57
r87 76 78 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=5.565 $Y=1.57
+ $X2=5.88 $Y2=1.57
r88 71 73 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=4.83 $Y=1.57 $X2=5.29
+ $Y2=1.57
r89 66 68 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.37 $Y=1.57
+ $X2=4.625 $Y2=1.57
r90 62 82 2.53537 $w=2.48e-07 $l=5.5e-08 $layer=LI1_cond $X=6.42 $Y=1.57
+ $X2=6.365 $Y2=1.57
r91 46 47 12.0563 $w=3.23e-07 $l=3.4e-07 $layer=LI1_cond $X=8.462 $Y=1.87
+ $X2=8.462 $Y2=2.21
r92 46 91 6.20546 $w=3.23e-07 $l=1.75e-07 $layer=LI1_cond $X=8.462 $Y=1.87
+ $X2=8.462 $Y2=1.695
r93 45 91 3.03503 $w=3.25e-07 $l=1.25e-07 $layer=LI1_cond $X=8.462 $Y=1.57
+ $X2=8.462 $Y2=1.695
r94 45 86 3.93339 $w=2.5e-07 $l=1.62e-07 $layer=LI1_cond $X=8.462 $Y=1.57
+ $X2=8.3 $Y2=1.57
r95 44 90 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=7.93 $Y=1.57
+ $X2=7.945 $Y2=1.57
r96 44 87 18.4391 $w=2.48e-07 $l=4e-07 $layer=LI1_cond $X=7.93 $Y=1.57 $X2=7.53
+ $Y2=1.57
r97 43 83 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=1.57
+ $X2=7.36 $Y2=1.57
r98 43 87 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=1.57
+ $X2=7.53 $Y2=1.57
r99 43 83 0.59927 $w=2.48e-07 $l=1.3e-08 $layer=LI1_cond $X=7.347 $Y=1.57
+ $X2=7.36 $Y2=1.57
r100 43 84 16.2264 $w=2.48e-07 $l=3.52e-07 $layer=LI1_cond $X=7.347 $Y=1.57
+ $X2=6.995 $Y2=1.57
r101 42 84 4.60977 $w=2.48e-07 $l=1e-07 $layer=LI1_cond $X=6.895 $Y=1.57
+ $X2=6.995 $Y2=1.57
r102 42 103 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.895 $Y=1.57
+ $X2=6.885 $Y2=1.57
r103 42 101 1.11538 $w=2.35e-07 $l=1.25e-07 $layer=LI1_cond $X=6.877 $Y=1.445
+ $X2=6.877 $Y2=1.57
r104 41 101 20.1447 $w=2.48e-07 $l=4.37e-07 $layer=LI1_cond $X=6.44 $Y=1.57
+ $X2=6.877 $Y2=1.57
r105 41 62 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=6.44 $Y=1.57
+ $X2=6.42 $Y2=1.57
r106 41 82 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=6.355 $Y=1.57
+ $X2=6.365 $Y2=1.57
r107 40 41 21.4354 $w=2.48e-07 $l=4.65e-07 $layer=LI1_cond $X=5.89 $Y=1.57
+ $X2=6.355 $Y2=1.57
r108 40 78 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=5.89 $Y=1.57
+ $X2=5.88 $Y2=1.57
r109 39 76 11.2939 $w=2.48e-07 $l=2.45e-07 $layer=LI1_cond $X=5.32 $Y=1.57
+ $X2=5.565 $Y2=1.57
r110 39 73 1.38293 $w=2.48e-07 $l=3e-08 $layer=LI1_cond $X=5.32 $Y=1.57 $X2=5.29
+ $Y2=1.57
r111 38 71 0.460977 $w=2.48e-07 $l=1e-08 $layer=LI1_cond $X=4.82 $Y=1.57
+ $X2=4.83 $Y2=1.57
r112 38 68 8.98906 $w=2.48e-07 $l=1.95e-07 $layer=LI1_cond $X=4.82 $Y=1.57
+ $X2=4.625 $Y2=1.57
r113 37 66 0.921954 $w=2.48e-07 $l=2e-08 $layer=LI1_cond $X=4.35 $Y=1.57
+ $X2=4.37 $Y2=1.57
r114 34 42 17.061 $w=4.03e-07 $l=5.6e-07 $layer=LI1_cond $X=6.877 $Y=0.885
+ $X2=6.877 $Y2=1.445
r115 34 36 3.43738 $w=2.35e-07 $l=1.2e-07 $layer=LI1_cond $X=6.877 $Y=0.885
+ $X2=6.877 $Y2=0.765
r116 30 43 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.445 $Y=1.695
+ $X2=7.445 $Y2=1.57
r117 30 32 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.445 $Y=1.695
+ $X2=7.445 $Y2=1.95
r118 26 36 3.38009 $w=2.4e-07 $l=1.18e-07 $layer=LI1_cond $X=6.995 $Y=0.765
+ $X2=6.877 $Y2=0.765
r119 26 28 44.177 $w=2.38e-07 $l=9.2e-07 $layer=LI1_cond $X=6.995 $Y=0.765
+ $X2=7.915 $Y2=0.765
r120 22 41 2.99516 $w=1.7e-07 $l=1.5411e-07 $layer=LI1_cond $X=6.505 $Y=1.695
+ $X2=6.44 $Y2=1.57
r121 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.505 $Y=1.695
+ $X2=6.505 $Y2=1.95
r122 7 45 300 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=2 $X=8.24
+ $Y=1.485 $X2=8.385 $Y2=1.69
r123 6 43 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.3
+ $Y=1.485 $X2=7.445 $Y2=1.61
r124 6 32 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=7.3
+ $Y=1.485 $X2=7.445 $Y2=1.95
r125 5 41 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=6.36
+ $Y=1.485 $X2=6.505 $Y2=1.61
r126 5 24 300 $w=1.7e-07 $l=5.32588e-07 $layer=licon1_PDIFF $count=2 $X=6.36
+ $Y=1.485 $X2=6.505 $Y2=1.95
r127 4 76 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.42
+ $Y=1.485 $X2=5.565 $Y2=1.61
r128 3 68 600 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=1 $X=4.475
+ $Y=1.485 $X2=4.625 $Y2=1.61
r129 2 28 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=7.73
+ $Y=0.235 $X2=7.915 $Y2=0.76
r130 1 36 182 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_NDIFF $count=1 $X=6.79
+ $Y=0.235 $X2=6.975 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%A_31_47# 1 2 3 4 5 6 7 8 9 30 32 33 36 38
+ 42 44 48 50 54 56 60 62 68 69 72 74 76 77 78 79 80
r150 72 82 3.04002 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=8.442 $Y=0.475
+ $X2=8.442 $Y2=0.365
r151 72 74 9.90697 $w=2.83e-07 $l=2.45e-07 $layer=LI1_cond $X=8.442 $Y=0.475
+ $X2=8.442 $Y2=0.72
r152 69 71 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=6.59 $Y=0.365
+ $X2=7.445 $Y2=0.365
r153 68 82 3.92439 $w=2.2e-07 $l=1.42e-07 $layer=LI1_cond $X=8.3 $Y=0.365
+ $X2=8.442 $Y2=0.365
r154 68 71 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=8.3 $Y=0.365
+ $X2=7.445 $Y2=0.365
r155 65 67 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=6.505 $Y=0.715
+ $X2=6.505 $Y2=0.56
r156 64 69 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.505 $Y=0.475
+ $X2=6.59 $Y2=0.365
r157 64 67 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0.475
+ $X2=6.505 $Y2=0.56
r158 63 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.53 $Y=0.8
+ $X2=5.445 $Y2=0.8
r159 62 65 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.42 $Y=0.8
+ $X2=6.505 $Y2=0.715
r160 62 63 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=6.42 $Y=0.8
+ $X2=5.53 $Y2=0.8
r161 58 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.445 $Y=0.715
+ $X2=5.445 $Y2=0.8
r162 58 60 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.445 $Y=0.715
+ $X2=5.445 $Y2=0.56
r163 57 79 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.205 $Y=0.8
+ $X2=4.015 $Y2=0.8
r164 56 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.36 $Y=0.8
+ $X2=5.445 $Y2=0.8
r165 56 57 75.3529 $w=1.68e-07 $l=1.155e-06 $layer=LI1_cond $X=5.36 $Y=0.8
+ $X2=4.205 $Y2=0.8
r166 52 79 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.015 $Y=0.715
+ $X2=4.015 $Y2=0.8
r167 52 54 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=4.015 $Y=0.715
+ $X2=4.015 $Y2=0.36
r168 51 78 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.265 $Y=0.8
+ $X2=3.075 $Y2=0.8
r169 50 79 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.825 $Y=0.8
+ $X2=4.015 $Y2=0.8
r170 50 51 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.825 $Y=0.8
+ $X2=3.265 $Y2=0.8
r171 46 78 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.715
+ $X2=3.075 $Y2=0.8
r172 46 48 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=3.075 $Y=0.715
+ $X2=3.075 $Y2=0.36
r173 45 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=0.8
+ $X2=2.135 $Y2=0.8
r174 44 78 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=0.8
+ $X2=3.075 $Y2=0.8
r175 44 45 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.885 $Y=0.8
+ $X2=2.325 $Y2=0.8
r176 40 77 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.135 $Y=0.715
+ $X2=2.135 $Y2=0.8
r177 40 42 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=2.135 $Y=0.715
+ $X2=2.135 $Y2=0.36
r178 39 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=0.8
+ $X2=1.195 $Y2=0.8
r179 38 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.945 $Y=0.8
+ $X2=2.135 $Y2=0.8
r180 38 39 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.945 $Y=0.8
+ $X2=1.385 $Y2=0.8
r181 34 76 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.715
+ $X2=1.195 $Y2=0.8
r182 34 36 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.195 $Y=0.715
+ $X2=1.195 $Y2=0.36
r183 32 76 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0.8
+ $X2=1.195 $Y2=0.8
r184 32 33 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=0.8
+ $X2=0.445 $Y2=0.8
r185 28 33 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.445 $Y2=0.8
r186 28 30 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.267 $Y2=0.38
r187 9 82 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=8.2
+ $Y=0.235 $X2=8.385 $Y2=0.38
r188 9 74 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=8.2
+ $Y=0.235 $X2=8.385 $Y2=0.72
r189 8 71 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=7.26
+ $Y=0.235 $X2=7.445 $Y2=0.36
r190 7 67 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=6.37
+ $Y=0.235 $X2=6.505 $Y2=0.56
r191 6 60 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=5.26
+ $Y=0.235 $X2=5.445 $Y2=0.56
r192 5 54 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.905
+ $Y=0.235 $X2=4.04 $Y2=0.36
r193 4 48 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=2.915
+ $Y=0.235 $X2=3.1 $Y2=0.36
r194 3 42 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.36
r195 2 36 91 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=2 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.36
r196 1 30 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.155
+ $Y=0.235 $X2=0.28 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_4%VGND 1 2 3 4 5 6 23 25 29 33 37 41 44 45
+ 47 48 50 51 52 73 74 77 80 85 88
r130 87 88 11.301 $w=6.28e-07 $l=2.15e-07 $layer=LI1_cond $X=4.925 $Y=0.23
+ $X2=5.14 $Y2=0.23
r131 83 87 1.80361 $w=6.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.83 $Y=0.23
+ $X2=4.925 $Y2=0.23
r132 83 85 14.5285 $w=6.28e-07 $l=3.85e-07 $layer=LI1_cond $X=4.83 $Y=0.23
+ $X2=4.445 $Y2=0.23
r133 83 84 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r134 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r135 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r136 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r137 73 74 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r138 71 74 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=6.21 $Y=0 $X2=8.51
+ $Y2=0
r139 70 73 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=6.21 $Y=0 $X2=8.51
+ $Y2=0
r140 70 71 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r141 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r142 68 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=4.83
+ $Y2=0
r143 67 88 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=5.14
+ $Y2=0
r144 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r145 64 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r146 63 85 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.445
+ $Y2=0
r147 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r148 60 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r149 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r150 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r151 57 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r152 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r153 54 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.775 $Y=0 $X2=1.69
+ $Y2=0
r154 54 56 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=1.775 $Y=0
+ $X2=2.53 $Y2=0
r155 52 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r156 50 67 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=5.79 $Y=0 $X2=5.75
+ $Y2=0
r157 50 51 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=5.79 $Y=0 $X2=5.975
+ $Y2=0
r158 49 70 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=6.16 $Y=0 $X2=6.21
+ $Y2=0
r159 49 51 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.16 $Y=0 $X2=5.975
+ $Y2=0
r160 47 59 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.45
+ $Y2=0
r161 47 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.485 $Y=0 $X2=3.57
+ $Y2=0
r162 46 63 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=3.655 $Y=0
+ $X2=4.37 $Y2=0
r163 46 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.655 $Y=0 $X2=3.57
+ $Y2=0
r164 44 56 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r165 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.63
+ $Y2=0
r166 43 59 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.715 $Y=0
+ $X2=3.45 $Y2=0
r167 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.63
+ $Y2=0
r168 39 51 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0
r169 39 41 8.56545 $w=3.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.975 $Y=0.085
+ $X2=5.975 $Y2=0.36
r170 35 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0
r171 35 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.57 $Y=0.085
+ $X2=3.57 $Y2=0.38
r172 31 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0
r173 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.63 $Y=0.085
+ $X2=2.63 $Y2=0.38
r174 27 80 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0
r175 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.69 $Y=0.085
+ $X2=1.69 $Y2=0.38
r176 26 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.75
+ $Y2=0
r177 25 80 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.69
+ $Y2=0
r178 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.835 $Y2=0
r179 21 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r180 21 23 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r181 6 41 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=5.73
+ $Y=0.235 $X2=5.975 $Y2=0.36
r182 5 87 91 $w=1.7e-07 $l=6.59545e-07 $layer=licon1_NDIFF $count=2 $X=4.325
+ $Y=0.235 $X2=4.925 $Y2=0.36
r183 4 37 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.385
+ $Y=0.235 $X2=3.57 $Y2=0.38
r184 3 33 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.445
+ $Y=0.235 $X2=2.63 $Y2=0.38
r185 2 29 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.38
r186 1 23 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.38
.ends

