* NGSPICE file created from sky130_fd_sc_hdll__clkmux2_4.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkmux2_4 A0 A1 S VGND VNB VPB VPWR X
M1000 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=1.3588e+12p pd=1.066e+07u as=5.8e+11p ps=5.16e+06u
M1001 VGND a_925_21# a_754_47# VNB nshort w=420000u l=150000u
+  ad=8.016e+11p pd=7.42e+06u as=3.591e+11p ps=2.55e+06u
M1002 a_925_21# S VGND VNB nshort w=520000u l=150000u
+  ad=1.352e+11p pd=1.56e+06u as=0p ps=0u
M1003 X a_79_199# VGND VNB nshort w=520000u l=150000u
+  ad=2.808e+11p pd=3.16e+06u as=0p ps=0u
M1004 X a_79_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_79_199# A1 a_525_47# VNB nshort w=420000u l=150000u
+  ad=2.121e+11p pd=1.85e+06u as=1.428e+11p ps=1.52e+06u
M1006 a_925_21# S VPWR VPB phighvt w=940000u l=180000u
+  ad=2.726e+11p pd=2.46e+06u as=0p ps=0u
M1007 a_875_309# A1 a_79_199# VPB phighvt w=940000u l=180000u
+  ad=2.444e+11p pd=2.4e+06u as=9.447e+11p ps=3.89e+06u
M1008 X a_79_199# VGND VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_754_47# A0 a_79_199# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND a_79_199# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_523_309# S VPWR VPB phighvt w=940000u l=180000u
+  ad=3.713e+11p pd=2.67e+06u as=0p ps=0u
M1013 a_79_199# A0 a_523_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 VGND a_79_199# X VNB nshort w=520000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_79_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_525_47# S VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_925_21# a_875_309# VPB phighvt w=940000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

