* File: sky130_fd_sc_hdll__a32o_2.spice
* Created: Wed Sep  2 08:20:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a32o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a32o_2  VNB VPB B2 B1 A1 A2 A3 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A3	A3
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* VPB	VPB
* VNB	VNB
MM1001 N_VGND_M1001_d N_A_21_199#_M1001_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75003.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A_21_199#_M1009_g N_X_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.225875 AS=0.104 PD=1.345 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75003.2 A=0.0975 P=1.6 MULT=1
MM1012 A_382_47# N_B2_M1012_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.225875 PD=1.005 PS=1.345 NRD=22.608 NRS=8.304 M=1 R=4.33333
+ SA=75001.5 SB=75002.4 A=0.0975 P=1.6 MULT=1
MM1004 N_A_21_199#_M1004_d N_B1_M1004_g A_382_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.115375 PD=1.03 PS=1.005 NRD=11.988 NRS=22.608 M=1 R=4.33333
+ SA=75002.1 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1007 A_589_47# N_A1_M1007_g N_A_21_199#_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.1235 PD=1.18 PS=1.03 NRD=38.76 NRS=6.456 M=1 R=4.33333
+ SA=75002.6 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1010 A_725_47# N_A2_M1010_g A_589_47# VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.17225 PD=0.92 PS=1.18 NRD=14.76 NRS=38.76 M=1 R=4.33333 SA=75003.3
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1013 N_VGND_M1013_d N_A3_M1013_g A_725_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333 SA=75003.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_X_M1000_d N_A_21_199#_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_X_M1003_d N_A_21_199#_M1003_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1008 N_A_21_199#_M1008_d N_B2_M1008_g N_A_319_297#_M1008_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_319_297#_M1005_d N_B1_M1005_g N_A_21_199#_M1008_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_319_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.225 AS=0.145 PD=1.45 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1011 N_A_319_297#_M1011_d N_A2_M1011_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.225 PD=1.29 PS=1.45 NRD=0.9653 NRS=32.4853 M=1 R=5.55556
+ SA=90001.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_A3_M1006_g N_A_319_297#_M1011_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
pX15_noxref noxref_16 A2 A2 PROBETYPE=1
pX16_noxref noxref_17 A2 A2 PROBETYPE=1
pX17_noxref noxref_18 A2 A2 PROBETYPE=1
pX18_noxref noxref_19 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__a32o_2.pxi.spice"
*
.ends
*
*
