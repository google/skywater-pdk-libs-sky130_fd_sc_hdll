* NGSPICE file created from sky130_fd_sc_hdll__and4_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and4_2 A B C D VGND VNB VPB VPWR X
M1000 VGND a_27_47# X VNB nshort w=650000u l=150000u
+  ad=5.1575e+11p pd=4.24e+06u as=2.795e+11p ps=2.16e+06u
M1001 VGND D a_301_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.386e+11p ps=1.5e+06u
M1002 a_27_47# A VPWR VPB phighvt w=420000u l=180000u
+  ad=2.478e+11p pd=2.86e+06u as=9.943e+11p ps=8.44e+06u
M1003 a_27_47# C VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.5e+11p pd=2.7e+06u as=0p ps=0u
M1005 X a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_203_47# B a_119_47# VNB nshort w=420000u l=150000u
+  ad=1.428e+11p pd=1.52e+06u as=1.134e+11p ps=1.38e+06u
M1007 a_119_47# A a_27_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1008 VPWR B a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_301_47# C a_203_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VPWR D a_27_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

