* NGSPICE file created from sky130_fd_sc_hdll__or2_8.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__or2_8 A B VGND VNB VPB VPWR X
M1000 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=1.71e+12p pd=1.542e+07u as=8.5e+11p ps=7.7e+06u
M1001 VGND A a_123_47# VNB nshort w=650000u l=150000u
+  ad=1.963e+12p pd=1.514e+07u as=3.51e+11p ps=3.68e+06u
M1002 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=1.16e+12p pd=1.032e+07u as=0p ps=0u
M1003 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=7.02e+11p ps=7.36e+06u
M1004 a_123_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_27_297# B a_123_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_123_47# B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_123_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VGND B a_123_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR a_123_47# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 X a_123_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 VGND a_123_47# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_123_47# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

