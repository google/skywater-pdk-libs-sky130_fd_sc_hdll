* File: sky130_fd_sc_hdll__o21ai_4.pex.spice
* Created: Thu Aug 27 19:19:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%A1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 27 31 34 40 46 52 56
c106 31 0 2.07545e-19 $X=3.88 $Y=1.16
r107 46 47 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r108 45 56 11.5043 $w=6.68e-07 $l=2.15e-07 $layer=LI1_cond $X=1.41 $Y=1.35
+ $X2=1.625 $Y2=1.35
r109 44 46 9.93132 $w=3.64e-07 $l=7.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.485 $Y2=1.202
r110 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.41
+ $Y=1.16 $X2=1.41 $Y2=1.16
r111 42 44 50.3187 $w=3.64e-07 $l=3.8e-07 $layer=POLY_cond $X=1.03 $Y=1.202
+ $X2=1.41 $Y2=1.202
r112 41 42 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=1.005 $Y=1.202
+ $X2=1.03 $Y2=1.202
r113 40 52 9.283 $w=6.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.63 $Y=1.35 $X2=1.15
+ $Y2=1.35
r114 39 41 49.6566 $w=3.64e-07 $l=3.75e-07 $layer=POLY_cond $X=0.63 $Y=1.202
+ $X2=1.005 $Y2=1.202
r115 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.63
+ $Y=1.16 $X2=0.63 $Y2=1.16
r116 37 39 10.5934 $w=3.64e-07 $l=8e-08 $layer=POLY_cond $X=0.55 $Y=1.202
+ $X2=0.63 $Y2=1.202
r117 36 37 3.31044 $w=3.64e-07 $l=2.5e-08 $layer=POLY_cond $X=0.525 $Y=1.202
+ $X2=0.55 $Y2=1.202
r118 34 45 2.85631 $w=6.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.25 $Y=1.35
+ $X2=1.41 $Y2=1.35
r119 34 52 1.78519 $w=6.68e-07 $l=1e-07 $layer=LI1_cond $X=1.25 $Y=1.35 $X2=1.15
+ $Y2=1.35
r120 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r121 29 31 13.6372 $w=2.98e-07 $l=3.55e-07 $layer=LI1_cond $X=3.945 $Y=1.515
+ $X2=3.945 $Y2=1.16
r122 27 29 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.795 $Y=1.6
+ $X2=3.945 $Y2=1.515
r123 27 56 141.572 $w=1.68e-07 $l=2.17e-06 $layer=LI1_cond $X=3.795 $Y=1.6
+ $X2=1.625 $Y2=1.6
r124 22 32 38.7084 $w=3.43e-07 $l=1.86145e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.905 $Y2=1.16
r125 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.95 $Y=0.995
+ $X2=3.95 $Y2=0.56
r126 19 32 45.964 $w=3.43e-07 $l=2.59808e-07 $layer=POLY_cond $X=3.885 $Y=1.41
+ $X2=3.905 $Y2=1.16
r127 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.885 $Y=1.41
+ $X2=3.885 $Y2=1.985
r128 16 47 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=1.202
r129 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.56
r130 13 46 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r131 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r132 10 42 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.03 $Y=0.995
+ $X2=1.03 $Y2=1.202
r133 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.03 $Y=0.995
+ $X2=1.03 $Y2=0.56
r134 7 41 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.005 $Y=1.41
+ $X2=1.005 $Y2=1.202
r135 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.005 $Y=1.41
+ $X2=1.005 $Y2=1.985
r136 4 37 23.572 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.55 $Y2=1.202
r137 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.55 $Y=0.995
+ $X2=0.55 $Y2=0.56
r138 1 36 19.2285 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.525 $Y=1.41
+ $X2=0.525 $Y2=1.202
r139 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.525 $Y=1.41
+ $X2=0.525 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%A2 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 41 42 47 49
c71 22 0 1.00539e-19 $X=3.43 $Y=0.995
r72 47 49 0.041907 $w=2.73e-07 $l=1e-09 $layer=LI1_cond $X=2.36 $Y=1.207
+ $X2=2.361 $Y2=1.207
r73 42 43 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=3.405 $Y=1.202
+ $X2=3.43 $Y2=1.202
r74 40 42 14.9407 $w=3.71e-07 $l=1.15e-07 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.405 $Y2=1.202
r75 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.29
+ $Y=1.16 $X2=3.29 $Y2=1.16
r76 38 40 47.4205 $w=3.71e-07 $l=3.65e-07 $layer=POLY_cond $X=2.925 $Y=1.202
+ $X2=3.29 $Y2=1.202
r77 37 38 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.9 $Y=1.202
+ $X2=2.925 $Y2=1.202
r78 36 41 18.8582 $w=2.73e-07 $l=4.5e-07 $layer=LI1_cond $X=2.84 $Y=1.207
+ $X2=3.29 $Y2=1.207
r79 36 49 20.0735 $w=2.73e-07 $l=4.79e-07 $layer=LI1_cond $X=2.84 $Y=1.207
+ $X2=2.361 $Y2=1.207
r80 35 37 7.79515 $w=3.71e-07 $l=6e-08 $layer=POLY_cond $X=2.84 $Y=1.202 $X2=2.9
+ $Y2=1.202
r81 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.84
+ $Y=1.16 $X2=2.84 $Y2=1.16
r82 33 35 51.3181 $w=3.71e-07 $l=3.95e-07 $layer=POLY_cond $X=2.445 $Y=1.202
+ $X2=2.84 $Y2=1.202
r83 32 33 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=2.42 $Y=1.202
+ $X2=2.445 $Y2=1.202
r84 30 32 7.79515 $w=3.71e-07 $l=6e-08 $layer=POLY_cond $X=2.36 $Y=1.202
+ $X2=2.42 $Y2=1.202
r85 30 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.36
+ $Y=1.16 $X2=2.36 $Y2=1.16
r86 28 30 51.3181 $w=3.71e-07 $l=3.95e-07 $layer=POLY_cond $X=1.965 $Y=1.202
+ $X2=2.36 $Y2=1.202
r87 27 28 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=1.94 $Y=1.202
+ $X2=1.965 $Y2=1.202
r88 25 47 3.77163 $w=2.73e-07 $l=9e-08 $layer=LI1_cond $X=2.27 $Y=1.207 $X2=2.36
+ $Y2=1.207
r89 22 43 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=1.202
r90 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.43 $Y=0.995
+ $X2=3.43 $Y2=0.56
r91 19 42 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.405 $Y=1.41
+ $X2=3.405 $Y2=1.202
r92 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.405 $Y=1.41
+ $X2=3.405 $Y2=1.985
r93 16 38 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.202
r94 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.925 $Y=1.41
+ $X2=2.925 $Y2=1.985
r95 13 37 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.9 $Y=0.995 $X2=2.9
+ $Y2=1.202
r96 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.9 $Y=0.995 $X2=2.9
+ $Y2=0.56
r97 10 33 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.445 $Y=1.41
+ $X2=2.445 $Y2=1.202
r98 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.445 $Y=1.41
+ $X2=2.445 $Y2=1.985
r99 7 32 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=1.202
r100 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.42 $Y=0.995
+ $X2=2.42 $Y2=0.56
r101 4 28 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.202
r102 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.985
r103 1 27 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.94 $Y=0.995
+ $X2=1.94 $Y2=1.202
r104 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.94 $Y=0.995
+ $X2=1.94 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%B1 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 36 39 45
c71 16 0 1.53101e-19 $X=5.365 $Y=1.41
c72 1 0 1.07005e-19 $X=4.38 $Y=0.995
r73 39 40 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=5.845 $Y=1.202
+ $X2=5.87 $Y2=1.202
r74 38 39 62.3612 $w=3.71e-07 $l=4.8e-07 $layer=POLY_cond $X=5.365 $Y=1.202
+ $X2=5.845 $Y2=1.202
r75 37 38 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=5.34 $Y=1.202
+ $X2=5.365 $Y2=1.202
r76 36 45 18.6164 $w=2.58e-07 $l=4.2e-07 $layer=LI1_cond $X=5.25 $Y=1.145
+ $X2=4.83 $Y2=1.145
r77 35 37 11.6927 $w=3.71e-07 $l=9e-08 $layer=POLY_cond $X=5.25 $Y=1.202
+ $X2=5.34 $Y2=1.202
r78 35 36 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r79 33 35 47.4205 $w=3.71e-07 $l=3.65e-07 $layer=POLY_cond $X=4.885 $Y=1.202
+ $X2=5.25 $Y2=1.202
r80 32 33 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.86 $Y=1.202
+ $X2=4.885 $Y2=1.202
r81 30 32 50.6685 $w=3.71e-07 $l=3.9e-07 $layer=POLY_cond $X=4.47 $Y=1.202
+ $X2=4.86 $Y2=1.202
r82 30 31 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=4.47
+ $Y=1.16 $X2=4.47 $Y2=1.16
r83 28 30 8.44474 $w=3.71e-07 $l=6.5e-08 $layer=POLY_cond $X=4.405 $Y=1.202
+ $X2=4.47 $Y2=1.202
r84 27 28 3.24798 $w=3.71e-07 $l=2.5e-08 $layer=POLY_cond $X=4.38 $Y=1.202
+ $X2=4.405 $Y2=1.202
r85 25 45 0.443247 $w=2.58e-07 $l=1e-08 $layer=LI1_cond $X=4.82 $Y=1.145
+ $X2=4.83 $Y2=1.145
r86 25 31 15.5137 $w=2.58e-07 $l=3.5e-07 $layer=LI1_cond $X=4.82 $Y=1.145
+ $X2=4.47 $Y2=1.145
r87 22 40 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.87 $Y=0.995
+ $X2=5.87 $Y2=1.202
r88 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.87 $Y=0.995
+ $X2=5.87 $Y2=0.56
r89 19 39 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.845 $Y=1.41
+ $X2=5.845 $Y2=1.202
r90 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.845 $Y=1.41
+ $X2=5.845 $Y2=1.985
r91 16 38 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.202
r92 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.365 $Y=1.41
+ $X2=5.365 $Y2=1.985
r93 13 37 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=1.202
r94 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.34 $Y=0.995
+ $X2=5.34 $Y2=0.56
r95 10 33 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.885 $Y=1.41
+ $X2=4.885 $Y2=1.202
r96 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.885 $Y=1.41
+ $X2=4.885 $Y2=1.985
r97 7 32 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.86 $Y=0.995
+ $X2=4.86 $Y2=1.202
r98 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.86 $Y=0.995 $X2=4.86
+ $Y2=0.56
r99 4 28 19.6776 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.202
r100 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.405 $Y=1.41
+ $X2=4.405 $Y2=1.985
r101 1 27 24.032 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=1.202
r102 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.38 $Y=0.995
+ $X2=4.38 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%VPWR 1 2 3 4 5 16 18 22 24 26 29 30 32 35
+ 38 40 55 63 71
r93 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r94 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r95 63 66 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.22 $Y=2.34
+ $X2=1.22 $Y2=2.72
r96 58 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r97 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r98 55 70 5.02378 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=5.87 $Y=2.72
+ $X2=6.155 $Y2=2.72
r99 55 57 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=5.87 $Y=2.72
+ $X2=5.75 $Y2=2.72
r100 54 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r101 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 50 51 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 48 51 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 48 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r106 47 50 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r107 47 48 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r108 45 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.22 $Y2=2.72
r109 45 47 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=1.41 $Y=2.72 $X2=1.61
+ $Y2=2.72
r110 44 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r111 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r112 41 60 4.31589 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.202 $Y2=2.72
r113 41 43 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.405 $Y=2.72
+ $X2=0.69 $Y2=2.72
r114 40 66 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.03 $Y=2.72
+ $X2=1.22 $Y2=2.72
r115 40 43 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=1.03 $Y=2.72
+ $X2=0.69 $Y2=2.72
r116 38 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r117 38 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r118 36 57 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r119 35 53 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.91 $Y=2.72 $X2=4.83
+ $Y2=2.72
r120 34 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=2.72 $X2=5.29
+ $Y2=2.72
r121 34 35 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.1 $Y=2.72 $X2=4.91
+ $Y2=2.72
r122 32 34 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=5.1 $Y=2.34 $X2=5.1
+ $Y2=2.72
r123 29 50 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=4.03 $Y=2.72
+ $X2=3.91 $Y2=2.72
r124 29 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.03 $Y=2.72 $X2=4.17
+ $Y2=2.72
r125 28 53 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=4.31 $Y=2.72
+ $X2=4.83 $Y2=2.72
r126 28 30 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=4.31 $Y=2.72 $X2=4.17
+ $Y2=2.72
r127 24 70 3.17291 $w=3.8e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.06 $Y=2.635
+ $X2=6.155 $Y2=2.72
r128 24 26 20.3194 $w=3.78e-07 $l=6.7e-07 $layer=LI1_cond $X=6.06 $Y=2.635
+ $X2=6.06 $Y2=1.965
r129 20 30 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2.72
r130 20 22 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=4.17 $Y=2.635
+ $X2=4.17 $Y2=2.36
r131 16 60 3.08278 $w=2.85e-07 $l=1.11018e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.202 $Y2=2.72
r132 16 18 25.6772 $w=2.83e-07 $l=6.35e-07 $layer=LI1_cond $X=0.262 $Y=2.635
+ $X2=0.262 $Y2=2
r133 5 26 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=5.935
+ $Y=1.485 $X2=6.085 $Y2=1.965
r134 4 32 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.975
+ $Y=1.485 $X2=5.125 $Y2=2.34
r135 3 22 600 $w=1.7e-07 $l=9.5623e-07 $layer=licon1_PDIFF $count=1 $X=3.975
+ $Y=1.485 $X2=4.145 $Y2=2.36
r136 2 63 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=1.095
+ $Y=1.485 $X2=1.245 $Y2=2.34
r137 1 18 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.16
+ $Y=1.485 $X2=0.285 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%A_123_297# 1 2 3 4 15 17 18 20 25
r37 23 25 56.0383 $w=1.88e-07 $l=9.6e-07 $layer=LI1_cond $X=2.685 $Y=2.37
+ $X2=3.645 $Y2=2.37
r38 21 28 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.82 $Y=2.37
+ $X2=1.725 $Y2=2.37
r39 21 23 50.4928 $w=1.88e-07 $l=8.65e-07 $layer=LI1_cond $X=1.82 $Y=2.37
+ $X2=2.685 $Y2=2.37
r40 20 28 3.40825 $w=1.9e-07 $l=9.5e-08 $layer=LI1_cond $X=1.725 $Y=2.275
+ $X2=1.725 $Y2=2.37
r41 19 20 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=1.725 $Y=2.085
+ $X2=1.725 $Y2=2.275
r42 17 19 6.84389 $w=1.7e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.63 $Y=2
+ $X2=1.725 $Y2=2.085
r43 17 18 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.63 $Y=2 $X2=0.86
+ $Y2=2
r44 13 18 7.04737 $w=1.7e-07 $l=1.54771e-07 $layer=LI1_cond $X=0.742 $Y=2.085
+ $X2=0.86 $Y2=2
r45 13 15 10.5436 $w=2.33e-07 $l=2.15e-07 $layer=LI1_cond $X=0.742 $Y=2.085
+ $X2=0.742 $Y2=2.3
r46 4 25 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=3.495
+ $Y=1.485 $X2=3.645 $Y2=2.36
r47 3 23 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=1.485 $X2=2.685 $Y2=2.36
r48 2 28 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.725 $Y2=2.3
r49 1 15 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=0.615
+ $Y=1.485 $X2=0.765 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%Y 1 2 3 4 5 6 19 25 33 35 36 39 45 48 51
+ 53
c81 53 0 1.53101e-19 $X=6.25 $Y=0.85
r82 51 53 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=6.125 $Y=0.845
+ $X2=6.125 $Y2=0.85
r83 48 51 2.71052 $w=4.1e-07 $l=1.15e-07 $layer=LI1_cond $X=6.125 $Y=0.73
+ $X2=6.125 $Y2=0.845
r84 48 53 1.12433 $w=4.08e-07 $l=4e-08 $layer=LI1_cond $X=6.125 $Y=0.89
+ $X2=6.125 $Y2=0.85
r85 47 48 15.6001 $w=4.08e-07 $l=5.55e-07 $layer=LI1_cond $X=6.125 $Y=1.445
+ $X2=6.125 $Y2=0.89
r86 45 47 18.4419 $w=3.44e-07 $l=5.2e-07 $layer=LI1_cond $X=5.605 $Y=1.7
+ $X2=6.125 $Y2=1.7
r87 41 43 0.199673 $w=6.11e-07 $l=1e-08 $layer=LI1_cond $X=4.635 $Y=1.765
+ $X2=4.645 $Y2=1.765
r88 37 45 4.21186 $w=1.9e-07 $l=3.85e-07 $layer=LI1_cond $X=5.605 $Y=2.085
+ $X2=5.605 $Y2=1.7
r89 37 39 12.5502 $w=1.88e-07 $l=2.15e-07 $layer=LI1_cond $X=5.605 $Y=2.085
+ $X2=5.605 $Y2=2.3
r90 36 43 1.81094 $w=6.4e-07 $l=9.5e-08 $layer=LI1_cond $X=4.74 $Y=1.765
+ $X2=4.645 $Y2=1.765
r91 35 45 4.40409 $w=6.4e-07 $l=1.23288e-07 $layer=LI1_cond $X=5.51 $Y=1.765
+ $X2=5.605 $Y2=1.7
r92 35 36 14.3903 $w=6.38e-07 $l=7.7e-07 $layer=LI1_cond $X=5.51 $Y=1.765
+ $X2=4.74 $Y2=1.765
r93 31 41 7.0888 $w=2.1e-07 $l=3.2e-07 $layer=LI1_cond $X=4.635 $Y=2.085
+ $X2=4.635 $Y2=1.765
r94 31 33 11.355 $w=2.08e-07 $l=2.15e-07 $layer=LI1_cond $X=4.635 $Y=2.085
+ $X2=4.635 $Y2=2.3
r95 27 30 48.102 $w=2.28e-07 $l=9.6e-07 $layer=LI1_cond $X=4.645 $Y=0.73
+ $X2=5.605 $Y2=0.73
r96 25 48 4.8318 $w=2.3e-07 $l=2.05e-07 $layer=LI1_cond $X=5.92 $Y=0.73
+ $X2=6.125 $Y2=0.73
r97 25 30 15.7835 $w=2.28e-07 $l=3.15e-07 $layer=LI1_cond $X=5.92 $Y=0.73
+ $X2=5.605 $Y2=0.73
r98 21 24 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=2.205 $Y=1.94
+ $X2=3.165 $Y2=1.94
r99 19 41 13.1279 $w=6.11e-07 $l=3.77492e-07 $layer=LI1_cond $X=4.335 $Y=1.94
+ $X2=4.635 $Y2=1.765
r100 19 24 76.3316 $w=1.68e-07 $l=1.17e-06 $layer=LI1_cond $X=4.335 $Y=1.94
+ $X2=3.165 $Y2=1.94
r101 6 45 600 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=1.485 $X2=5.605 $Y2=1.825
r102 6 39 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=5.455
+ $Y=1.485 $X2=5.605 $Y2=2.3
r103 5 43 600 $w=1.7e-07 $l=4.08167e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.485 $X2=4.645 $Y2=1.825
r104 5 33 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=4.495
+ $Y=1.485 $X2=4.645 $Y2=2.3
r105 4 24 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=3.015
+ $Y=1.485 $X2=3.165 $Y2=1.94
r106 3 21 600 $w=1.7e-07 $l=5.24667e-07 $layer=licon1_PDIFF $count=1 $X=2.055
+ $Y=1.485 $X2=2.205 $Y2=1.94
r107 2 30 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.605 $Y2=0.7
r108 1 27 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=4.455
+ $Y=0.235 $X2=4.645 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%A_32_47# 1 2 3 4 5 6 7 22 36 40
r53 38 40 56.0383 $w=1.88e-07 $l=9.6e-07 $layer=LI1_cond $X=5.125 $Y=0.35
+ $X2=6.085 $Y2=0.35
r54 36 38 50.4928 $w=1.88e-07 $l=8.65e-07 $layer=LI1_cond $X=4.26 $Y=0.35
+ $X2=5.125 $Y2=0.35
r55 33 35 3.75797 $w=2.28e-07 $l=7.5e-08 $layer=LI1_cond $X=4.145 $Y=0.615
+ $X2=4.145 $Y2=0.54
r56 32 36 6.89722 $w=1.9e-07 $l=1.55403e-07 $layer=LI1_cond $X=4.145 $Y=0.445
+ $X2=4.26 $Y2=0.35
r57 32 35 4.76009 $w=2.28e-07 $l=9.5e-08 $layer=LI1_cond $X=4.145 $Y=0.445
+ $X2=4.145 $Y2=0.54
r58 29 31 51.9379 $w=2.03e-07 $l=9.6e-07 $layer=LI1_cond $X=2.205 $Y=0.717
+ $X2=3.165 $Y2=0.717
r59 27 29 51.9379 $w=2.03e-07 $l=9.6e-07 $layer=LI1_cond $X=1.245 $Y=0.717
+ $X2=2.205 $Y2=0.717
r60 24 27 51.9379 $w=2.03e-07 $l=9.6e-07 $layer=LI1_cond $X=0.285 $Y=0.717
+ $X2=1.245 $Y2=0.717
r61 22 33 6.84582 $w=2.05e-07 $l=1.57972e-07 $layer=LI1_cond $X=4.03 $Y=0.717
+ $X2=4.145 $Y2=0.615
r62 22 31 46.7982 $w=2.03e-07 $l=8.65e-07 $layer=LI1_cond $X=4.03 $Y=0.717
+ $X2=3.165 $Y2=0.717
r63 7 40 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=5.945
+ $Y=0.235 $X2=6.085 $Y2=0.36
r64 6 38 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=4.935
+ $Y=0.235 $X2=5.125 $Y2=0.36
r65 5 35 182 $w=1.7e-07 $l=3.68409e-07 $layer=licon1_NDIFF $count=1 $X=4.025
+ $Y=0.235 $X2=4.165 $Y2=0.54
r66 4 31 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.235 $X2=3.165 $Y2=0.7
r67 3 29 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=2.015
+ $Y=0.235 $X2=2.205 $Y2=0.7
r68 2 27 182 $w=1.7e-07 $l=5.30401e-07 $layer=licon1_NDIFF $count=1 $X=1.105
+ $Y=0.235 $X2=1.245 $Y2=0.7
r69 1 24 182 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_NDIFF $count=1 $X=0.16
+ $Y=0.235 $X2=0.285 $Y2=0.7
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_4%VGND 1 2 3 4 13 15 17 19 24 34 35 39 46 53
+ 60
r76 60 63 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=3.62 $Y=0 $X2=3.62
+ $Y2=0.36
r77 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r78 54 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r79 53 56 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.66 $Y=0 $X2=2.66
+ $Y2=0.36
r80 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r81 47 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r82 46 49 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=1.7 $Y=0 $X2=1.7
+ $Y2=0.36
r83 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r84 39 42 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.74 $Y=0 $X2=0.74
+ $Y2=0.36
r85 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r86 34 35 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r87 32 35 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=3.91 $Y=0 $X2=6.21
+ $Y2=0
r88 32 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=3.45
+ $Y2=0
r89 31 34 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=6.21
+ $Y2=0
r90 31 32 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r91 29 60 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.62
+ $Y2=0
r92 29 31 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.81 $Y=0 $X2=3.91
+ $Y2=0
r93 28 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r94 28 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r95 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r96 25 39 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=0.74
+ $Y2=0
r97 25 27 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=0.93 $Y=0 $X2=1.15
+ $Y2=0
r98 24 46 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.7
+ $Y2=0
r99 24 27 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r100 19 39 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.74
+ $Y2=0
r101 19 21 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.55 $Y=0 $X2=0.23
+ $Y2=0
r102 17 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r103 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r104 16 53 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.85 $Y=0 $X2=2.66
+ $Y2=0
r105 15 60 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=3.62
+ $Y2=0
r106 15 16 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.43 $Y=0 $X2=2.85
+ $Y2=0
r107 14 46 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.7
+ $Y2=0
r108 13 53 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=2.66
+ $Y2=0
r109 13 14 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.47 $Y=0 $X2=1.89
+ $Y2=0
r110 4 63 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.645 $Y2=0.36
r111 3 56 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=2.495
+ $Y=0.235 $X2=2.685 $Y2=0.36
r112 2 49 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.725 $Y2=0.36
r113 1 42 182 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=1 $X=0.625
+ $Y=0.235 $X2=0.765 $Y2=0.36
.ends

