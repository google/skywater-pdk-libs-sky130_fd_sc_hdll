* File: sky130_fd_sc_hdll__or4b_2.spice
* Created: Wed Sep  2 08:49:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4b_2.pex.spice"
.subckt sky130_fd_sc_hdll__or4b_2  VNB VPB D_N A B C VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* C	C
* B	B
* A	A
* D_N	D_N
* VPB	VPB
* VNB	VNB
MM1010 N_VGND_M1010_d N_D_N_M1010_g N_A_27_47#_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0787009 AS=0.1302 PD=0.773271 PS=1.46 NRD=8.568 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75003.2 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_186_21#_M1001_g N_VGND_M1010_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.121799 PD=0.97 PS=1.19673 NRD=8.304 NRS=4.608 M=1 R=4.33333
+ SA=75000.5 SB=75002 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1001_d N_A_186_21#_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.141542 PD=0.97 PS=1.25748 NRD=0 NRS=11.076 M=1 R=4.33333
+ SA=75001 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1009 N_A_186_21#_M1009_d N_A_M1009_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0914579 PD=0.8 PS=0.812523 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75001.7 A=0.063 P=1.14 MULT=1
MM1007 N_VGND_M1007_d N_B_M1007_g N_A_186_21#_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0798 PD=0.69 PS=0.8 NRD=0 NRS=15.708 M=1 R=2.8 SA=75002.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1011 N_A_186_21#_M1011_d N_C_M1011_g N_VGND_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75002.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_27_47#_M1002_g N_A_186_21#_M1011_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0777 PD=1.46 PS=0.79 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75003.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1004 N_VPWR_M1004_d N_D_N_M1004_g N_A_27_47#_M1004_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.109969 AS=0.1134 PD=0.928732 PS=1.38 NRD=97.0028 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90003.2 A=0.0756 P=1.2 MULT=1
MM1005 N_VPWR_M1004_d N_A_186_21#_M1005_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.261831 AS=0.145 PD=2.21127 PS=1.29 NRD=14.7553 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1012_d N_A_186_21#_M1012_g N_X_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.247113 AS=0.145 PD=2.1338 PS=1.29 NRD=14.7553 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90001 A=0.18 P=2.36 MULT=1
MM1000 A_425_297# N_A_M1000_g N_VPWR_M1012_d VPB PHIGHVT L=0.18 W=0.42 AD=0.0735
+ AS=0.103787 PD=0.77 PS=0.896197 NRD=56.2829 NRS=90.1078 M=1 R=2.33333
+ SA=90001.7 SB=90001.6 A=0.0756 P=1.2 MULT=1
MM1008 A_531_297# N_B_M1008_g A_425_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0504
+ AS=0.0735 PD=0.66 PS=0.77 NRD=30.4759 NRS=56.2829 M=1 R=2.33333 SA=90002.2
+ SB=90001.1 A=0.0756 P=1.2 MULT=1
MM1006 A_615_297# N_C_M1006_g A_531_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0714
+ AS=0.0504 PD=0.76 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333 SA=90002.7
+ SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1003 N_A_186_21#_M1003_d N_A_27_47#_M1003_g A_615_297# VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.0714 PD=1.38 PS=0.76 NRD=2.3443 NRS=53.9386 M=1
+ R=2.33333 SA=90003.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX15_noxref noxref_15 X X PROBETYPE=1
pX16_noxref noxref_16 A A PROBETYPE=1
pX17_noxref noxref_17 B B PROBETYPE=1
*
.include "sky130_fd_sc_hdll__or4b_2.pxi.spice"
*
.ends
*
*
