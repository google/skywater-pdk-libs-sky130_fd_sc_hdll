* File: sky130_fd_sc_hdll__inputiso1n_1.pxi.spice
* Created: Wed Sep  2 08:32:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%SLEEP_B N_SLEEP_B_c_59_n N_SLEEP_B_M1002_g
+ N_SLEEP_B_M1000_g SLEEP_B N_SLEEP_B_c_58_n SLEEP_B
+ PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%SLEEP_B
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_27_53# N_A_27_53#_M1000_s
+ N_A_27_53#_M1002_d N_A_27_53#_c_91_n N_A_27_53#_M1003_g N_A_27_53#_M1006_g
+ N_A_27_53#_c_85_n N_A_27_53#_c_86_n N_A_27_53#_c_87_n N_A_27_53#_c_92_n
+ N_A_27_53#_c_88_n N_A_27_53#_c_89_n N_A_27_53#_c_90_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_27_53#
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A N_A_c_136_n N_A_c_133_n N_A_c_134_n
+ N_A_c_137_n N_A_M1001_g N_A_M1005_g N_A_c_139_n A N_A_c_141_n A
+ PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_229_297# N_A_229_297#_M1006_d
+ N_A_229_297#_M1003_s N_A_229_297#_c_179_n N_A_229_297#_M1007_g
+ N_A_229_297#_c_180_n N_A_229_297#_M1004_g N_A_229_297#_c_188_n
+ N_A_229_297#_c_226_p N_A_229_297#_c_181_n N_A_229_297#_c_182_n
+ N_A_229_297#_c_183_n N_A_229_297#_c_186_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%A_229_297#
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VPWR N_VPWR_M1002_s N_VPWR_M1001_d
+ N_VPWR_c_238_n N_VPWR_c_239_n N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n
+ VPWR N_VPWR_c_243_n N_VPWR_c_237_n PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VPWR
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%X N_X_M1004_d N_X_M1007_d N_X_c_270_n
+ N_X_c_272_n N_X_c_271_n X PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%X
x_PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VGND N_VGND_M1000_d N_VGND_M1005_d
+ N_VGND_c_288_n VGND N_VGND_c_289_n N_VGND_c_290_n N_VGND_c_291_n
+ N_VGND_c_292_n N_VGND_c_293_n PM_SKY130_FD_SC_HDLL__INPUTISO1N_1%VGND
cc_1 VNB N_SLEEP_B_M1000_g 0.0401282f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.475
cc_2 VNB SLEEP_B 0.0092769f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_SLEEP_B_c_58_n 0.0431049f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_A_27_53#_M1006_g 0.0345946f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_5 VNB N_A_27_53#_c_85_n 0.0205152f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_6 VNB N_A_27_53#_c_86_n 0.00342105f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.2
cc_7 VNB N_A_27_53#_c_87_n 0.00940306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_53#_c_88_n 0.00460073f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_53#_c_89_n 0.0134238f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_53#_c_90_n 0.0392689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_c_133_n 0.00696033f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.695
cc_12 VNB N_A_c_134_n 0.0106821f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_13 VNB N_A_M1005_g 0.0288162f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_14 VNB N_A_229_297#_c_179_n 0.0290589f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_229_297#_c_180_n 0.020598f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_16 VNB N_A_229_297#_c_181_n 0.00233799f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_229_297#_c_182_n 0.00451202f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_229_297#_c_183_n 0.00113231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VPWR_c_237_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_270_n 0.0182958f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_21 VNB N_X_c_271_n 0.0273182f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_22 VNB N_VGND_c_288_n 0.0166718f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_289_n 0.024346f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.2
cc_24 VNB N_VGND_c_290_n 0.195305f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.19
cc_25 VNB N_VGND_c_291_n 0.018858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_292_n 0.0228528f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_293_n 0.0102968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VPB N_SLEEP_B_c_59_n 0.0238148f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_29 VPB SLEEP_B 8.85293e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_30 VPB N_SLEEP_B_c_58_n 0.0190244f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_31 VPB N_A_27_53#_c_91_n 0.0193758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A_27_53#_c_92_n 0.00464761f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_A_27_53#_c_88_n 0.00639441f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_27_53#_c_89_n 0.00350361f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_53#_c_90_n 0.0148363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_c_136_n 0.0406198f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB N_A_c_137_n 0.00661582f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.475
cc_38 VPB N_A_M1001_g 0.0122761f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_39 VPB N_A_c_139_n 0.0291674f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_40 VPB A 0.0292646f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_41 VPB N_A_c_141_n 0.0374051f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_229_297#_c_179_n 0.032959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_229_297#_c_183_n 0.00165371f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_229_297#_c_186_n 0.008297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_238_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_239_n 0.0554415f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_240_n 0.0121527f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_48 VPB N_VPWR_c_241_n 0.0450247f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_49 VPB N_VPWR_c_242_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_243_n 0.0242869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_237_n 0.0679987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_X_c_272_n 0.00970498f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_53 VPB N_X_c_271_n 0.00932001f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.2
cc_54 VPB X 0.0358702f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.19
cc_55 N_SLEEP_B_M1000_g N_A_27_53#_c_85_n 0.00300084f $X=0.52 $Y=0.475 $X2=0
+ $Y2=0
cc_56 N_SLEEP_B_M1000_g N_A_27_53#_c_86_n 0.0187886f $X=0.52 $Y=0.475 $X2=0
+ $Y2=0
cc_57 SLEEP_B N_A_27_53#_c_86_n 3.30304e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_58 N_SLEEP_B_c_58_n N_A_27_53#_c_86_n 0.00104773f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_59 SLEEP_B N_A_27_53#_c_87_n 0.0255233f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_60 N_SLEEP_B_c_58_n N_A_27_53#_c_87_n 0.00800665f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_61 N_SLEEP_B_c_59_n N_A_27_53#_c_92_n 0.00630275f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_62 N_SLEEP_B_c_58_n N_A_27_53#_c_92_n 0.00650453f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_63 N_SLEEP_B_M1000_g N_A_27_53#_c_89_n 0.00807875f $X=0.52 $Y=0.475 $X2=0
+ $Y2=0
cc_64 SLEEP_B N_A_27_53#_c_89_n 0.0159063f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_65 N_SLEEP_B_c_58_n N_A_27_53#_c_90_n 0.00528959f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_66 N_SLEEP_B_c_59_n A 0.00227571f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_67 N_SLEEP_B_c_58_n A 2.63734e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_68 N_SLEEP_B_c_59_n N_A_229_297#_c_186_n 0.00166948f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_69 N_SLEEP_B_c_59_n N_VPWR_c_239_n 0.00874982f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 SLEEP_B N_VPWR_c_239_n 0.0206483f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_71 N_SLEEP_B_c_58_n N_VPWR_c_239_n 0.00545118f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_72 N_SLEEP_B_c_59_n N_VPWR_c_241_n 0.00298464f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_SLEEP_B_c_59_n N_VPWR_c_237_n 0.0037574f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_SLEEP_B_M1000_g N_VGND_c_290_n 0.00754515f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_75 N_SLEEP_B_M1000_g N_VGND_c_291_n 0.00413798f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_76 N_SLEEP_B_M1000_g N_VGND_c_292_n 0.00505351f $X=0.52 $Y=0.475 $X2=0 $Y2=0
cc_77 N_A_27_53#_c_91_n N_A_c_136_n 0.010421f $X=1.505 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_27_53#_c_88_n N_A_c_133_n 0.00130319f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_27_53#_c_90_n N_A_c_133_n 0.0214081f $X=1.505 $Y=1.202 $X2=0 $Y2=0
cc_80 N_A_27_53#_c_91_n N_A_M1001_g 0.0281104f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_27_53#_M1006_g N_A_M1005_g 0.019627f $X=1.53 $Y=0.475 $X2=0 $Y2=0
cc_82 N_A_27_53#_c_91_n A 0.00205903f $X=1.505 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_27_53#_c_92_n A 0.0124285f $X=0.73 $Y=1.62 $X2=0 $Y2=0
cc_84 N_A_27_53#_c_91_n N_A_229_297#_c_188_n 0.0131318f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_85 N_A_27_53#_M1006_g N_A_229_297#_c_182_n 0.00459933f $X=1.53 $Y=0.475 $X2=0
+ $Y2=0
cc_86 N_A_27_53#_c_91_n N_A_229_297#_c_186_n 0.00939681f $X=1.505 $Y=1.41 $X2=0
+ $Y2=0
cc_87 N_A_27_53#_c_92_n N_A_229_297#_c_186_n 0.0253576f $X=0.73 $Y=1.62 $X2=0
+ $Y2=0
cc_88 N_A_27_53#_c_88_n N_A_229_297#_c_186_n 0.0267679f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_27_53#_c_90_n N_A_229_297#_c_186_n 0.006068f $X=1.505 $Y=1.202 $X2=0
+ $Y2=0
cc_90 N_A_27_53#_c_92_n N_VPWR_c_239_n 0.0192276f $X=0.73 $Y=1.62 $X2=0 $Y2=0
cc_91 N_A_27_53#_M1006_g N_VGND_c_288_n 0.00555245f $X=1.53 $Y=0.475 $X2=0 $Y2=0
cc_92 N_A_27_53#_M1006_g N_VGND_c_290_n 0.011632f $X=1.53 $Y=0.475 $X2=0 $Y2=0
cc_93 N_A_27_53#_c_85_n N_VGND_c_290_n 0.0117861f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_94 N_A_27_53#_c_86_n N_VGND_c_290_n 0.0050353f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_95 N_A_27_53#_c_89_n N_VGND_c_290_n 0.00105248f $X=0.77 $Y=0.82 $X2=0 $Y2=0
cc_96 N_A_27_53#_c_85_n N_VGND_c_291_n 0.0192939f $X=0.26 $Y=0.445 $X2=0 $Y2=0
cc_97 N_A_27_53#_c_86_n N_VGND_c_291_n 0.00299761f $X=0.645 $Y=0.82 $X2=0 $Y2=0
cc_98 N_A_27_53#_M1006_g N_VGND_c_292_n 0.0107462f $X=1.53 $Y=0.475 $X2=0 $Y2=0
cc_99 N_A_27_53#_c_88_n N_VGND_c_292_n 0.0202613f $X=1.27 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_27_53#_c_89_n N_VGND_c_292_n 0.0214575f $X=0.77 $Y=0.82 $X2=0 $Y2=0
cc_101 N_A_27_53#_c_90_n N_VGND_c_292_n 0.00471044f $X=1.505 $Y=1.202 $X2=0
+ $Y2=0
cc_102 N_A_27_53#_M1006_g N_VGND_c_293_n 6.0833e-19 $X=1.53 $Y=0.475 $X2=0 $Y2=0
cc_103 N_A_c_137_n N_A_229_297#_c_179_n 0.00275812f $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_M1001_g N_A_229_297#_c_179_n 0.0161769f $X=1.975 $Y=1.695 $X2=0 $Y2=0
cc_105 N_A_M1005_g N_A_229_297#_c_179_n 0.0216416f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_106 N_A_M1005_g N_A_229_297#_c_180_n 0.0189258f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_107 N_A_c_136_n N_A_229_297#_c_188_n 0.00104251f $X=1.875 $Y=2.34 $X2=0 $Y2=0
cc_108 N_A_M1001_g N_A_229_297#_c_188_n 0.0200197f $X=1.975 $Y=1.695 $X2=0 $Y2=0
cc_109 A N_A_229_297#_c_188_n 0.0152425f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_110 N_A_c_133_n N_A_229_297#_c_181_n 0.00149549f $X=1.975 $Y=1.115 $X2=0
+ $Y2=0
cc_111 N_A_M1005_g N_A_229_297#_c_181_n 0.0135334f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_112 N_A_c_137_n N_A_229_297#_c_183_n 0.00164174f $X=1.975 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_M1001_g N_A_229_297#_c_183_n 0.00161078f $X=1.975 $Y=1.695 $X2=0
+ $Y2=0
cc_114 N_A_M1005_g N_A_229_297#_c_183_n 0.00530858f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_115 N_A_c_136_n N_A_229_297#_c_186_n 9.83498e-19 $X=1.875 $Y=2.34 $X2=0 $Y2=0
cc_116 N_A_M1001_g N_A_229_297#_c_186_n 0.00115363f $X=1.975 $Y=1.695 $X2=0
+ $Y2=0
cc_117 A N_A_229_297#_c_186_n 0.0344364f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_118 N_A_c_141_n N_A_229_297#_c_186_n 0.00119166f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_119 A N_VPWR_c_239_n 0.0258572f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_120 N_A_c_141_n N_VPWR_c_239_n 9.23051e-19 $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_121 N_A_M1001_g N_VPWR_c_240_n 0.00448545f $X=1.975 $Y=1.695 $X2=0 $Y2=0
cc_122 N_A_c_139_n N_VPWR_c_240_n 0.00487993f $X=1.975 $Y=2.34 $X2=0 $Y2=0
cc_123 A N_VPWR_c_240_n 0.0216404f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_124 A N_VPWR_c_241_n 0.0666505f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_125 N_A_c_141_n N_VPWR_c_241_n 0.0251009f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_126 A N_VPWR_c_237_n 0.0490703f $X=1.12 $Y=2.125 $X2=0 $Y2=0
cc_127 N_A_c_141_n N_VPWR_c_237_n 0.0347738f $X=1.225 $Y=2.28 $X2=0 $Y2=0
cc_128 N_A_M1005_g N_VGND_c_288_n 0.00188229f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_129 N_A_M1005_g N_VGND_c_290_n 0.00261357f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_130 N_A_M1005_g N_VGND_c_293_n 0.0102417f $X=2 $Y=0.475 $X2=0 $Y2=0
cc_131 N_A_229_297#_c_188_n N_VPWR_M1001_d 0.00651861f $X=2.335 $Y=1.58 $X2=0
+ $Y2=0
cc_132 N_A_229_297#_c_179_n N_VPWR_c_240_n 0.00512739f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A_229_297#_c_188_n N_VPWR_c_240_n 0.0198977f $X=2.335 $Y=1.58 $X2=0
+ $Y2=0
cc_134 N_A_229_297#_c_186_n N_VPWR_c_240_n 0.00211805f $X=1.25 $Y=1.58 $X2=0
+ $Y2=0
cc_135 N_A_229_297#_c_179_n N_VPWR_c_243_n 0.00702461f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_229_297#_c_179_n N_VPWR_c_237_n 0.0148665f $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_229_297#_c_188_n A_319_297# 0.00596563f $X=2.335 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_138 N_A_229_297#_c_181_n N_X_c_270_n 0.00874309f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_139 N_A_229_297#_c_179_n N_X_c_272_n 0.0123985f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_229_297#_c_188_n N_X_c_272_n 0.0142209f $X=2.335 $Y=1.58 $X2=0 $Y2=0
cc_141 N_A_229_297#_c_179_n N_X_c_271_n 0.00159158f $X=2.515 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_229_297#_c_180_n N_X_c_271_n 0.0127184f $X=2.54 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_229_297#_c_181_n N_X_c_271_n 0.00269941f $X=2.335 $Y=0.74 $X2=0 $Y2=0
cc_144 N_A_229_297#_c_183_n N_X_c_271_n 0.0250104f $X=2.42 $Y=1.16 $X2=0 $Y2=0
cc_145 N_A_229_297#_c_181_n N_VGND_M1005_d 0.00650959f $X=2.335 $Y=0.74 $X2=0
+ $Y2=0
cc_146 N_A_229_297#_c_183_n N_VGND_M1005_d 7.32946e-19 $X=2.42 $Y=1.16 $X2=0
+ $Y2=0
cc_147 N_A_229_297#_c_226_p N_VGND_c_288_n 0.00861358f $X=1.74 $Y=0.47 $X2=0
+ $Y2=0
cc_148 N_A_229_297#_c_181_n N_VGND_c_288_n 0.00232988f $X=2.335 $Y=0.74 $X2=0
+ $Y2=0
cc_149 N_A_229_297#_c_180_n N_VGND_c_289_n 0.00543382f $X=2.54 $Y=0.995 $X2=0
+ $Y2=0
cc_150 N_A_229_297#_c_181_n N_VGND_c_289_n 0.00105918f $X=2.335 $Y=0.74 $X2=0
+ $Y2=0
cc_151 N_A_229_297#_c_180_n N_VGND_c_290_n 0.0110495f $X=2.54 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_229_297#_c_226_p N_VGND_c_290_n 0.00625722f $X=1.74 $Y=0.47 $X2=0
+ $Y2=0
cc_153 N_A_229_297#_c_181_n N_VGND_c_290_n 0.00843284f $X=2.335 $Y=0.74 $X2=0
+ $Y2=0
cc_154 N_A_229_297#_c_179_n N_VGND_c_293_n 4.00709e-19 $X=2.515 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_229_297#_c_180_n N_VGND_c_293_n 0.00498808f $X=2.54 $Y=0.995 $X2=0
+ $Y2=0
cc_156 N_A_229_297#_c_226_p N_VGND_c_293_n 0.0135697f $X=1.74 $Y=0.47 $X2=0
+ $Y2=0
cc_157 N_A_229_297#_c_181_n N_VGND_c_293_n 0.0273767f $X=2.335 $Y=0.74 $X2=0
+ $Y2=0
cc_158 N_VPWR_c_237_n N_X_M1007_d 0.00481197f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_159 N_VPWR_c_243_n X 0.0285921f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_160 N_VPWR_c_237_n X 0.0155202f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_161 N_X_c_270_n N_VGND_c_289_n 0.0134041f $X=2.995 $Y=0.587 $X2=0 $Y2=0
cc_162 N_X_M1004_d N_VGND_c_290_n 0.00454412f $X=2.615 $Y=0.235 $X2=0 $Y2=0
cc_163 N_X_c_270_n N_VGND_c_290_n 0.0138697f $X=2.995 $Y=0.587 $X2=0 $Y2=0
