* File: sky130_fd_sc_hdll__nand4bb_2.pxi.spice
* Created: Thu Aug 27 19:15:08 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%B_N N_B_N_c_107_n N_B_N_c_108_n N_B_N_M1002_g
+ N_B_N_c_102_n N_B_N_M1012_g N_B_N_c_103_n N_B_N_c_109_n B_N B_N N_B_N_c_105_n
+ N_B_N_c_106_n PM_SKY130_FD_SC_HDLL__NAND4BB_2%B_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_N N_A_N_c_148_n N_A_N_c_149_n N_A_N_M1013_g
+ N_A_N_M1000_g A_N A_N N_A_N_c_147_n PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_211_413# N_A_211_413#_M1000_d
+ N_A_211_413#_M1013_d N_A_211_413#_c_192_n N_A_211_413#_M1010_g
+ N_A_211_413#_c_186_n N_A_211_413#_M1003_g N_A_211_413#_c_193_n
+ N_A_211_413#_M1014_g N_A_211_413#_M1004_g N_A_211_413#_c_188_n
+ N_A_211_413#_c_189_n N_A_211_413#_c_190_n N_A_211_413#_c_196_n
+ N_A_211_413#_c_191_n PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_211_413#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_27_47# N_A_27_47#_M1012_s N_A_27_47#_M1002_s
+ N_A_27_47#_c_272_n N_A_27_47#_M1007_g N_A_27_47#_M1015_g N_A_27_47#_c_273_n
+ N_A_27_47#_M1016_g N_A_27_47#_M1018_g N_A_27_47#_c_265_n N_A_27_47#_c_274_n
+ N_A_27_47#_c_266_n N_A_27_47#_c_267_n N_A_27_47#_c_275_n N_A_27_47#_c_276_n
+ N_A_27_47#_c_268_n N_A_27_47#_c_269_n N_A_27_47#_c_270_n N_A_27_47#_c_271_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%C N_C_c_376_n N_C_M1001_g N_C_M1011_g
+ N_C_c_377_n N_C_M1017_g N_C_M1019_g C C N_C_c_375_n C C
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%C
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%D N_D_c_421_n N_D_M1005_g N_D_M1006_g
+ N_D_c_422_n N_D_M1009_g N_D_M1008_g D D N_D_c_420_n D D
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%D
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%VPWR N_VPWR_M1002_d N_VPWR_M1010_d
+ N_VPWR_M1014_d N_VPWR_M1016_s N_VPWR_M1017_s N_VPWR_M1009_d N_VPWR_c_462_n
+ N_VPWR_c_463_n N_VPWR_c_464_n N_VPWR_c_465_n N_VPWR_c_466_n N_VPWR_c_467_n
+ N_VPWR_c_468_n N_VPWR_c_469_n N_VPWR_c_470_n N_VPWR_c_471_n N_VPWR_c_472_n
+ N_VPWR_c_473_n N_VPWR_c_474_n VPWR N_VPWR_c_475_n N_VPWR_c_476_n
+ N_VPWR_c_477_n N_VPWR_c_478_n N_VPWR_c_479_n N_VPWR_c_461_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%Y N_Y_M1003_s N_Y_M1010_s N_Y_M1007_d
+ N_Y_M1001_d N_Y_M1005_s N_Y_c_568_n N_Y_c_574_n N_Y_c_562_n N_Y_c_578_n
+ N_Y_c_563_n N_Y_c_561_n N_Y_c_603_n N_Y_c_565_n N_Y_c_566_n N_Y_c_608_n
+ N_Y_c_579_n N_Y_c_567_n Y Y PM_SKY130_FD_SC_HDLL__NAND4BB_2%Y
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%VGND N_VGND_M1012_d N_VGND_M1006_s
+ N_VGND_c_660_n N_VGND_c_661_n N_VGND_c_662_n N_VGND_c_663_n VGND
+ N_VGND_c_664_n N_VGND_c_665_n N_VGND_c_666_n N_VGND_c_667_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_361_47# N_A_361_47#_M1003_d
+ N_A_361_47#_M1004_d N_A_361_47#_M1018_d N_A_361_47#_c_731_n
+ N_A_361_47#_c_736_n PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_361_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_641_47# N_A_641_47#_M1015_s
+ N_A_641_47#_M1011_s N_A_641_47#_c_756_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_641_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_841_47# N_A_841_47#_M1011_d
+ N_A_841_47#_M1019_d N_A_841_47#_M1008_d N_A_841_47#_c_780_n
+ N_A_841_47#_c_802_n N_A_841_47#_c_781_n N_A_841_47#_c_782_n
+ N_A_841_47#_c_783_n PM_SKY130_FD_SC_HDLL__NAND4BB_2%A_841_47#
cc_1 VNB N_B_N_c_102_n 0.0173166f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_2 VNB N_B_N_c_103_n 0.0250037f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_3 VNB B_N 0.00978855f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_B_N_c_105_n 0.0216679f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_5 VNB N_B_N_c_106_n 0.014785f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_6 VNB N_A_N_M1000_g 0.0422749f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.73
cc_7 VNB A_N 0.00478742f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_8 VNB N_A_N_c_147_n 0.0251862f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_211_413#_c_186_n 0.0197985f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_10 VNB N_A_211_413#_M1004_g 0.0182531f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_11 VNB N_A_211_413#_c_188_n 0.0476346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_211_413#_c_189_n 0.037689f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_13 VNB N_A_211_413#_c_190_n 0.00474714f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.4
cc_14 VNB N_A_211_413#_c_191_n 0.00881569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_M1015_g 0.0187423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_M1018_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_265_n 0.018767f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_18 VNB N_A_27_47#_c_266_n 0.0181957f $X=-0.19 $Y=-0.24 $X2=0.207 $Y2=1.53
cc_19 VNB N_A_27_47#_c_267_n 0.00786701f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_268_n 0.00653181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_269_n 0.00611781f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_270_n 0.00113736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_27_47#_c_271_n 0.0512939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C_M1011_g 0.023617f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_25 VNB N_C_M1019_g 0.0188422f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_26 VNB C 0.00526324f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.887
cc_27 VNB N_C_c_375_n 0.0461062f $X=-0.19 $Y=-0.24 $X2=0.242 $Y2=1.07
cc_28 VNB N_D_M1006_g 0.0186248f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.275
cc_29 VNB N_D_M1008_g 0.0235985f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_30 VNB D 0.010695f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.887
cc_31 VNB N_D_c_420_n 0.0605637f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.235
cc_32 VNB N_VPWR_c_461_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_561_n 0.00691848f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_660_n 0.00232623f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_35 VNB N_VGND_c_661_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.805
cc_36 VNB N_VGND_c_662_n 0.111658f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.887
cc_37 VNB N_VGND_c_663_n 0.00323991f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_38 VNB N_VGND_c_664_n 0.0144236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_665_n 0.018342f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_666_n 0.324638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_667_n 0.00420022f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_361_47#_c_731_n 0.00272806f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_641_47#_c_756_n 0.0195965f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=0.805
cc_44 VNB N_A_841_47#_c_780_n 0.00271098f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_45 VNB N_A_841_47#_c_781_n 0.00317287f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.887
cc_46 VNB N_A_841_47#_c_782_n 0.0122279f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.887
cc_47 VNB N_A_841_47#_c_783_n 0.0191373f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VPB N_B_N_c_107_n 0.0282622f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.785
cc_49 VPB N_B_N_c_108_n 0.0189637f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_50 VPB N_B_N_c_109_n 0.0313252f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.887
cc_51 VPB B_N 0.0124835f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_52 VPB N_B_N_c_105_n 0.0108199f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_53 VPB N_A_N_c_148_n 0.0326007f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.07
cc_54 VPB N_A_N_c_149_n 0.0267018f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=1.4
cc_55 VPB A_N 0.00485075f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_56 VPB N_A_N_c_147_n 0.0157889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_211_413#_c_192_n 0.0191727f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_58 VPB N_A_211_413#_c_193_n 0.0153522f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.805
cc_59 VPB N_A_211_413#_c_188_n 0.0247079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_211_413#_c_189_n 0.0127696f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_61 VPB N_A_211_413#_c_196_n 0.00482638f $X=-0.19 $Y=1.305 $X2=0.207 $Y2=1.53
cc_62 VPB N_A_211_413#_c_191_n 0.0157599f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_272_n 0.0159735f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_64 VPB N_A_27_47#_c_273_n 0.0194278f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_274_n 0.0185631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_275_n 0.0118838f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_276_n 0.00897929f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_268_n 0.0102175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_269_n 0.00827671f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_271_n 0.0140252f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_C_c_376_n 0.0193344f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.88
cc_72 VPB N_C_c_377_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_73 VPB N_C_c_375_n 0.0138223f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_74 VPB N_D_c_421_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.305 $Y2=0.88
cc_75 VPB N_D_c_422_n 0.0198539f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.73
cc_76 VPB N_D_c_420_n 0.0223491f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.235
cc_77 VPB N_VPWR_c_462_n 0.00237984f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.235
cc_78 VPB N_VPWR_c_463_n 0.00414143f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.4
cc_79 VPB N_VPWR_c_464_n 0.00231485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_465_n 0.00743936f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_466_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_467_n 0.0100141f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_468_n 0.0466691f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_469_n 0.0254917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_470_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_471_n 0.016313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_472_n 0.00426174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_473_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_474_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_475_n 0.0151232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_476_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_477_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_478_n 0.00392577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_479_n 0.0126657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_461_n 0.0506097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_562_n 0.00268483f $X=-0.19 $Y=1.305 $X2=0.242 $Y2=1.07
cc_97 VPB N_Y_c_563_n 0.00510867f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_561_n 0.00511202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_Y_c_565_n 0.00470447f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_Y_c_566_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_Y_c_567_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 N_B_N_c_107_n N_A_N_c_148_n 0.00603885f $X=0.305 $Y=1.785 $X2=0 $Y2=0
cc_103 N_B_N_c_109_n N_A_N_c_148_n 0.00973765f $X=0.305 $Y=1.887 $X2=0 $Y2=0
cc_104 N_B_N_c_108_n N_A_N_c_149_n 0.0139076f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_105 N_B_N_c_102_n N_A_N_M1000_g 0.0173062f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_106 N_B_N_c_106_n N_A_N_M1000_g 0.00310679f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_107 N_B_N_c_103_n A_N 2.4588e-19 $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_108 N_B_N_c_109_n A_N 8.59498e-19 $X=0.305 $Y=1.887 $X2=0 $Y2=0
cc_109 B_N A_N 0.0340681f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_110 N_B_N_c_105_n A_N 0.00416475f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_111 B_N N_A_N_c_147_n 3.41991e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B_N_c_105_n N_A_N_c_147_n 0.0154571f $X=0.245 $Y=1.235 $X2=0 $Y2=0
cc_113 N_B_N_c_102_n N_A_27_47#_c_265_n 0.00596875f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_114 N_B_N_c_108_n N_A_27_47#_c_274_n 0.00349167f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_115 N_B_N_c_109_n N_A_27_47#_c_274_n 4.17387e-19 $X=0.305 $Y=1.887 $X2=0
+ $Y2=0
cc_116 N_B_N_c_103_n N_A_27_47#_c_266_n 0.0129738f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_117 N_B_N_c_106_n N_A_27_47#_c_266_n 0.00156143f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_118 N_B_N_c_103_n N_A_27_47#_c_267_n 0.00675396f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_119 B_N N_A_27_47#_c_267_n 0.020875f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_120 N_B_N_c_105_n N_A_27_47#_c_267_n 9.79955e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_121 N_B_N_c_106_n N_A_27_47#_c_267_n 0.00273512f $X=0.242 $Y=1.07 $X2=0 $Y2=0
cc_122 N_B_N_c_109_n N_A_27_47#_c_275_n 0.0190734f $X=0.305 $Y=1.887 $X2=0 $Y2=0
cc_123 N_B_N_c_109_n N_A_27_47#_c_276_n 0.0111984f $X=0.305 $Y=1.887 $X2=0 $Y2=0
cc_124 B_N N_A_27_47#_c_276_n 0.0214513f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_125 N_B_N_c_105_n N_A_27_47#_c_276_n 6.00486e-19 $X=0.245 $Y=1.235 $X2=0
+ $Y2=0
cc_126 N_B_N_c_108_n N_VPWR_c_462_n 0.010811f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_127 N_B_N_c_108_n N_VPWR_c_475_n 0.00395083f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_128 N_B_N_c_108_n N_VPWR_c_461_n 0.00565038f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_129 N_B_N_c_109_n N_VPWR_c_461_n 2.51067e-19 $X=0.305 $Y=1.887 $X2=0 $Y2=0
cc_130 N_B_N_c_102_n N_VGND_c_660_n 0.0122159f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_131 N_B_N_c_102_n N_VGND_c_664_n 0.00203849f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_132 N_B_N_c_103_n N_VGND_c_664_n 0.00162345f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_133 N_B_N_c_102_n N_VGND_c_666_n 0.00378134f $X=0.52 $Y=0.73 $X2=0 $Y2=0
cc_134 N_B_N_c_103_n N_VGND_c_666_n 0.00236448f $X=0.52 $Y=0.805 $X2=0 $Y2=0
cc_135 N_A_N_M1000_g N_A_211_413#_c_188_n 0.00969224f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_136 N_A_N_M1000_g N_A_211_413#_c_190_n 0.00634903f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_137 N_A_N_c_149_n N_A_211_413#_c_196_n 0.00633362f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_138 N_A_N_c_148_n N_A_211_413#_c_191_n 0.00138999f $X=0.965 $Y=1.89 $X2=0
+ $Y2=0
cc_139 N_A_N_c_149_n N_A_211_413#_c_191_n 0.00425858f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_140 N_A_N_M1000_g N_A_211_413#_c_191_n 0.00400849f $X=0.99 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_N_M1000_g N_A_27_47#_c_266_n 0.0168269f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_142 A_N N_A_27_47#_c_266_n 0.0311488f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A_N_c_147_n N_A_27_47#_c_266_n 0.00182559f $X=0.99 $Y=1.255 $X2=0 $Y2=0
cc_144 N_A_N_c_148_n N_A_27_47#_c_275_n 0.0118029f $X=0.965 $Y=1.89 $X2=0 $Y2=0
cc_145 N_A_N_c_149_n N_A_27_47#_c_275_n 0.00842914f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_146 A_N N_A_27_47#_c_275_n 0.0309101f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_N_c_147_n N_A_27_47#_c_275_n 0.00101174f $X=0.99 $Y=1.255 $X2=0 $Y2=0
cc_148 N_A_N_M1000_g N_A_27_47#_c_268_n 0.0210704f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_149 A_N N_A_27_47#_c_268_n 0.0311332f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_150 N_A_N_M1000_g N_A_27_47#_c_269_n 0.00539107f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_151 A_N N_A_27_47#_c_269_n 0.00791211f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_152 N_A_N_c_149_n N_VPWR_c_462_n 0.00403433f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_153 N_A_N_c_149_n N_VPWR_c_469_n 0.00506137f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_154 N_A_N_c_149_n N_VPWR_c_461_n 0.00812584f $X=0.965 $Y=1.99 $X2=0 $Y2=0
cc_155 N_A_N_M1000_g N_VGND_c_660_n 0.00387396f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A_N_M1000_g N_VGND_c_662_n 0.00395516f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_157 N_A_N_M1000_g N_VGND_c_666_n 0.00713717f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_158 N_A_211_413#_c_193_n N_A_27_47#_c_272_n 0.0227106f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_159 N_A_211_413#_M1004_g N_A_27_47#_M1015_g 0.0215289f $X=2.66 $Y=0.56 $X2=0
+ $Y2=0
cc_160 N_A_211_413#_c_190_n N_A_27_47#_c_265_n 3.93796e-19 $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_161 N_A_211_413#_c_190_n N_A_27_47#_c_266_n 0.0238028f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_162 N_A_211_413#_c_191_n N_A_27_47#_c_266_n 0.0143865f $X=1.585 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_211_413#_c_196_n N_A_27_47#_c_275_n 0.0245034f $X=1.5 $Y=2.307 $X2=0
+ $Y2=0
cc_164 N_A_211_413#_c_191_n N_A_27_47#_c_275_n 0.0165021f $X=1.585 $Y=1.16 $X2=0
+ $Y2=0
cc_165 N_A_211_413#_c_188_n N_A_27_47#_c_268_n 0.00251018f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_166 N_A_211_413#_c_191_n N_A_27_47#_c_268_n 0.0645524f $X=1.585 $Y=1.16 $X2=0
+ $Y2=0
cc_167 N_A_211_413#_c_188_n N_A_27_47#_c_269_n 0.0251843f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_211_413#_c_189_n N_A_27_47#_c_269_n 0.0108919f $X=2.635 $Y=1.202
+ $X2=0 $Y2=0
cc_169 N_A_211_413#_c_190_n N_A_27_47#_c_269_n 0.00678325f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_170 N_A_211_413#_c_191_n N_A_27_47#_c_269_n 0.0305537f $X=1.585 $Y=1.16 $X2=0
+ $Y2=0
cc_171 N_A_211_413#_c_189_n N_A_27_47#_c_270_n 8.30797e-19 $X=2.635 $Y=1.202
+ $X2=0 $Y2=0
cc_172 N_A_211_413#_c_189_n N_A_27_47#_c_271_n 0.0248348f $X=2.635 $Y=1.202
+ $X2=0 $Y2=0
cc_173 N_A_211_413#_c_196_n N_VPWR_c_462_n 0.0219006f $X=1.5 $Y=2.307 $X2=0
+ $Y2=0
cc_174 N_A_211_413#_c_192_n N_VPWR_c_463_n 0.00592862f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_211_413#_c_188_n N_VPWR_c_463_n 0.00746613f $X=2.065 $Y=1.16 $X2=0
+ $Y2=0
cc_176 N_A_211_413#_c_196_n N_VPWR_c_463_n 0.026217f $X=1.5 $Y=2.307 $X2=0 $Y2=0
cc_177 N_A_211_413#_c_191_n N_VPWR_c_463_n 0.0485183f $X=1.585 $Y=1.16 $X2=0
+ $Y2=0
cc_178 N_A_211_413#_c_192_n N_VPWR_c_464_n 7.42159e-19 $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_211_413#_c_193_n N_VPWR_c_464_n 0.0151063f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_211_413#_c_196_n N_VPWR_c_469_n 0.0445542f $X=1.5 $Y=2.307 $X2=0
+ $Y2=0
cc_181 N_A_211_413#_c_192_n N_VPWR_c_471_n 0.00597712f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_211_413#_c_193_n N_VPWR_c_471_n 0.00427505f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_211_413#_M1013_d N_VPWR_c_461_n 0.00389718f $X=1.055 $Y=2.065 $X2=0
+ $Y2=0
cc_184 N_A_211_413#_c_192_n N_VPWR_c_461_n 0.0112769f $X=2.165 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_211_413#_c_193_n N_VPWR_c_461_n 0.00732977f $X=2.635 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_211_413#_c_196_n N_VPWR_c_461_n 0.0257855f $X=1.5 $Y=2.307 $X2=0
+ $Y2=0
cc_187 N_A_211_413#_c_192_n N_Y_c_568_n 0.00116523f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_211_413#_c_186_n N_Y_c_568_n 0.010297f $X=2.19 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_211_413#_c_193_n N_Y_c_568_n 0.0012025f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_211_413#_M1004_g N_Y_c_568_n 0.00954012f $X=2.66 $Y=0.56 $X2=0 $Y2=0
cc_191 N_A_211_413#_c_189_n N_Y_c_568_n 0.038801f $X=2.635 $Y=1.202 $X2=0 $Y2=0
cc_192 N_A_211_413#_c_191_n N_Y_c_568_n 0.0218681f $X=1.585 $Y=1.16 $X2=0 $Y2=0
cc_193 N_A_211_413#_c_192_n N_Y_c_574_n 0.0133529f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_211_413#_c_193_n N_Y_c_574_n 0.00416059f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_211_413#_c_193_n N_Y_c_562_n 0.00812043f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_211_413#_c_189_n N_Y_c_562_n 4.93319e-19 $X=2.635 $Y=1.202 $X2=0
+ $Y2=0
cc_197 N_A_211_413#_c_193_n N_Y_c_578_n 4.84481e-19 $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_211_413#_c_192_n N_Y_c_579_n 0.00541795f $X=2.165 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_211_413#_c_193_n N_Y_c_579_n 0.00784714f $X=2.635 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_211_413#_c_191_n N_Y_c_579_n 0.00173962f $X=1.585 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A_211_413#_c_190_n N_VGND_c_660_n 0.0236772f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_202 N_A_211_413#_c_186_n N_VGND_c_662_n 0.00357877f $X=2.19 $Y=0.995 $X2=0
+ $Y2=0
cc_203 N_A_211_413#_M1004_g N_VGND_c_662_n 0.00357877f $X=2.66 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_211_413#_c_190_n N_VGND_c_662_n 0.0445308f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_205 N_A_211_413#_M1000_d N_VGND_c_666_n 0.00382322f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_A_211_413#_c_186_n N_VGND_c_666_n 0.00668309f $X=2.19 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A_211_413#_M1004_g N_VGND_c_666_n 0.00550244f $X=2.66 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_211_413#_c_190_n N_VGND_c_666_n 0.0258015f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_209 N_A_211_413#_c_186_n N_A_361_47#_c_731_n 0.0103488f $X=2.19 $Y=0.995
+ $X2=0 $Y2=0
cc_210 N_A_211_413#_M1004_g N_A_361_47#_c_731_n 0.0107346f $X=2.66 $Y=0.56 $X2=0
+ $Y2=0
cc_211 N_A_211_413#_c_188_n N_A_361_47#_c_731_n 0.00206727f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_212 N_A_211_413#_c_189_n N_A_361_47#_c_731_n 4.65706e-19 $X=2.635 $Y=1.202
+ $X2=0 $Y2=0
cc_213 N_A_211_413#_c_188_n N_A_361_47#_c_736_n 0.00533162f $X=2.065 $Y=1.16
+ $X2=0 $Y2=0
cc_214 N_A_211_413#_c_190_n N_A_361_47#_c_736_n 0.027349f $X=1.5 $Y=0.407 $X2=0
+ $Y2=0
cc_215 N_A_211_413#_c_191_n N_A_361_47#_c_736_n 0.00175037f $X=1.585 $Y=1.16
+ $X2=0 $Y2=0
cc_216 N_A_211_413#_M1004_g N_A_641_47#_c_756_n 8.09376e-19 $X=2.66 $Y=0.56
+ $X2=0 $Y2=0
cc_217 N_A_27_47#_c_271_n C 7.28558e-19 $X=3.575 $Y=1.217 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_275_n N_VPWR_c_462_n 0.0155163f $X=1.16 $Y=1.882 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_269_n N_VPWR_c_463_n 0.00840714f $X=3.24 $Y=1.19 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_272_n N_VPWR_c_464_n 0.00519708f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_27_47#_c_273_n N_VPWR_c_465_n 0.0210968f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_275_n N_VPWR_c_469_n 0.00231103f $X=1.16 $Y=1.882 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_274_n N_VPWR_c_475_n 0.0165425f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_224 N_A_27_47#_c_275_n N_VPWR_c_475_n 0.00225651f $X=1.16 $Y=1.882 $X2=0
+ $Y2=0
cc_225 N_A_27_47#_c_272_n N_VPWR_c_476_n 0.00597712f $X=3.105 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_c_273_n N_VPWR_c_476_n 0.00673617f $X=3.575 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_M1002_s N_VPWR_c_461_n 0.002367f $X=0.135 $Y=2.065 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_272_n N_VPWR_c_461_n 0.0100198f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_273_n N_VPWR_c_461_n 0.0132531f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_274_n N_VPWR_c_461_n 0.0107554f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_275_n N_VPWR_c_461_n 0.00909208f $X=1.16 $Y=1.882 $X2=0
+ $Y2=0
cc_232 N_A_27_47#_M1015_g N_Y_c_568_n 0.0013554f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_269_n N_Y_c_568_n 0.0529413f $X=3.24 $Y=1.19 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_270_n N_Y_c_568_n 0.00634521f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_271_n N_Y_c_568_n 0.00151796f $X=3.575 $Y=1.217 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_272_n N_Y_c_562_n 0.0112758f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_269_n N_Y_c_562_n 0.0197089f $X=3.24 $Y=1.19 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_270_n N_Y_c_562_n 0.0111151f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_271_n N_Y_c_562_n 0.00131794f $X=3.575 $Y=1.217 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_272_n N_Y_c_578_n 0.0132741f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_273_n N_Y_c_578_n 0.0153658f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_272_n N_Y_c_561_n 0.00309425f $X=3.105 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_273_n N_Y_c_561_n 0.0197405f $X=3.575 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_269_n N_Y_c_561_n 0.0158211f $X=3.24 $Y=1.19 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_270_n N_Y_c_561_n 0.0267631f $X=3.11 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_271_n N_Y_c_561_n 0.0281276f $X=3.575 $Y=1.217 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_265_n N_VGND_c_660_n 0.0219468f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_266_n N_VGND_c_660_n 0.0191727f $X=1.16 $Y=0.815 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1015_g N_VGND_c_662_n 0.00357877f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A_27_47#_M1018_g N_VGND_c_662_n 0.00357877f $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_266_n N_VGND_c_662_n 0.00242914f $X=1.16 $Y=0.815 $X2=0
+ $Y2=0
cc_252 N_A_27_47#_c_265_n N_VGND_c_664_n 0.0181392f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_266_n N_VGND_c_664_n 0.00223864f $X=1.16 $Y=0.815 $X2=0
+ $Y2=0
cc_254 N_A_27_47#_M1012_s N_VGND_c_666_n 0.00303307f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_255 N_A_27_47#_M1015_g N_VGND_c_666_n 0.00550244f $X=3.13 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A_27_47#_M1018_g N_VGND_c_666_n 0.00668309f $X=3.6 $Y=0.56 $X2=0 $Y2=0
cc_257 N_A_27_47#_c_265_n N_VGND_c_666_n 0.00992225f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_266_n N_VGND_c_666_n 0.00956571f $X=1.16 $Y=0.815 $X2=0
+ $Y2=0
cc_259 N_A_27_47#_M1015_g N_A_361_47#_c_731_n 0.0104867f $X=3.13 $Y=0.56 $X2=0
+ $Y2=0
cc_260 N_A_27_47#_M1018_g N_A_361_47#_c_731_n 0.00958923f $X=3.6 $Y=0.56 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_269_n N_A_361_47#_c_731_n 0.0193573f $X=3.24 $Y=1.19 $X2=0
+ $Y2=0
cc_262 N_A_27_47#_c_270_n N_A_361_47#_c_731_n 0.00196923f $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_c_271_n N_A_361_47#_c_731_n 0.00178081f $X=3.575 $Y=1.217
+ $X2=0 $Y2=0
cc_264 N_A_27_47#_c_269_n N_A_361_47#_c_736_n 0.00575495f $X=3.24 $Y=1.19 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1015_g N_A_641_47#_c_756_n 0.00754593f $X=3.13 $Y=0.56 $X2=0
+ $Y2=0
cc_266 N_A_27_47#_M1018_g N_A_641_47#_c_756_n 0.0138307f $X=3.6 $Y=0.56 $X2=0
+ $Y2=0
cc_267 N_A_27_47#_c_269_n N_A_641_47#_c_756_n 0.00650261f $X=3.24 $Y=1.19 $X2=0
+ $Y2=0
cc_268 N_A_27_47#_c_270_n N_A_641_47#_c_756_n 0.0127136f $X=3.11 $Y=1.16 $X2=0
+ $Y2=0
cc_269 N_A_27_47#_c_271_n N_A_641_47#_c_756_n 0.00372917f $X=3.575 $Y=1.217
+ $X2=0 $Y2=0
cc_270 N_C_c_377_n N_D_c_421_n 0.0231619f $X=5.005 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_271 N_C_M1019_g N_D_M1006_g 0.011669f $X=5.03 $Y=0.56 $X2=0 $Y2=0
cc_272 C D 0.00905729f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_273 N_C_c_375_n D 8.65592e-19 $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_274 N_C_c_375_n N_D_c_420_n 0.0254816f $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_275 N_C_c_376_n N_VPWR_c_465_n 0.00758137f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_276 N_C_c_377_n N_VPWR_c_466_n 0.0052072f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_277 N_C_c_376_n N_VPWR_c_473_n 0.00597712f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_278 N_C_c_377_n N_VPWR_c_473_n 0.00673617f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_279 N_C_c_376_n N_VPWR_c_461_n 0.0112769f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_280 N_C_c_377_n N_VPWR_c_461_n 0.011869f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_281 N_C_c_376_n N_Y_c_563_n 0.0139912f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_282 C N_Y_c_563_n 0.0235651f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_283 N_C_c_375_n N_Y_c_563_n 2.74992e-19 $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_284 N_C_c_376_n N_Y_c_561_n 0.00109412f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_285 C N_Y_c_561_n 0.0166175f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_286 N_C_c_375_n N_Y_c_561_n 0.00546018f $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_287 N_C_c_376_n N_Y_c_603_n 0.0178402f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_288 N_C_c_377_n N_Y_c_603_n 0.0106251f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_289 N_C_c_377_n N_Y_c_565_n 0.0199378f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_290 C N_Y_c_565_n 0.00101487f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_291 N_C_c_375_n N_Y_c_565_n 4.93319e-19 $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_292 N_C_c_377_n N_Y_c_608_n 6.48386e-19 $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_293 N_C_c_376_n N_Y_c_567_n 0.00292783f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_294 N_C_c_377_n N_Y_c_567_n 0.00116723f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_295 C N_Y_c_567_n 0.0305808f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_296 N_C_c_375_n N_Y_c_567_n 0.0074788f $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_297 N_C_M1011_g N_VGND_c_662_n 0.00357877f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_298 N_C_M1019_g N_VGND_c_662_n 0.00357877f $X=5.03 $Y=0.56 $X2=0 $Y2=0
cc_299 N_C_M1011_g N_VGND_c_666_n 0.00668309f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_300 N_C_M1019_g N_VGND_c_666_n 0.00550244f $X=5.03 $Y=0.56 $X2=0 $Y2=0
cc_301 N_C_M1011_g N_A_641_47#_c_756_n 0.0138006f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_302 C N_A_641_47#_c_756_n 0.0520461f $X=4.74 $Y=1.105 $X2=0 $Y2=0
cc_303 N_C_c_375_n N_A_641_47#_c_756_n 0.00461919f $X=5.005 $Y=1.212 $X2=0 $Y2=0
cc_304 N_C_M1011_g N_A_841_47#_c_780_n 0.00958923f $X=4.56 $Y=0.56 $X2=0 $Y2=0
cc_305 N_C_M1019_g N_A_841_47#_c_780_n 0.0143475f $X=5.03 $Y=0.56 $X2=0 $Y2=0
cc_306 N_C_M1019_g N_A_841_47#_c_781_n 2.11779e-19 $X=5.03 $Y=0.56 $X2=0 $Y2=0
cc_307 N_D_c_421_n N_VPWR_c_466_n 0.004751f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_308 N_D_c_422_n N_VPWR_c_468_n 0.00950067f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_309 D N_VPWR_c_468_n 0.0164394f $X=6.05 $Y=1.105 $X2=0 $Y2=0
cc_310 N_D_c_420_n N_VPWR_c_468_n 0.00339068f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_311 N_D_c_421_n N_VPWR_c_477_n 0.00597712f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_312 N_D_c_422_n N_VPWR_c_477_n 0.00673617f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_313 N_D_c_421_n N_VPWR_c_461_n 0.0100198f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_314 N_D_c_422_n N_VPWR_c_461_n 0.0127552f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_315 N_D_c_421_n N_Y_c_603_n 6.24674e-19 $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_316 N_D_c_421_n N_Y_c_565_n 0.0113403f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_317 D N_Y_c_565_n 0.0128375f $X=6.05 $Y=1.105 $X2=0 $Y2=0
cc_318 N_D_c_420_n N_Y_c_565_n 0.00160364f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_319 N_D_c_421_n N_Y_c_566_n 0.00292783f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_320 N_D_c_422_n N_Y_c_566_n 0.00349846f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_321 D N_Y_c_566_n 0.0305808f $X=6.05 $Y=1.105 $X2=0 $Y2=0
cc_322 N_D_c_420_n N_Y_c_566_n 0.0074788f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_323 N_D_c_421_n N_Y_c_608_n 0.0130707f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_324 N_D_c_422_n N_Y_c_608_n 0.0100147f $X=5.945 $Y=1.41 $X2=0 $Y2=0
cc_325 N_D_M1006_g N_VGND_c_661_n 0.00276126f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_326 N_D_M1008_g N_VGND_c_661_n 0.00361688f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_327 N_D_M1006_g N_VGND_c_662_n 0.00439206f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_328 N_D_M1008_g N_VGND_c_665_n 0.00397237f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_329 N_D_M1006_g N_VGND_c_666_n 0.00618369f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_330 N_D_M1008_g N_VGND_c_666_n 0.00665354f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_331 D N_A_841_47#_c_781_n 0.00731021f $X=6.05 $Y=1.105 $X2=0 $Y2=0
cc_332 N_D_c_420_n N_A_841_47#_c_781_n 0.00225392f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_333 N_D_M1006_g N_A_841_47#_c_782_n 0.0106613f $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_334 N_D_M1008_g N_A_841_47#_c_782_n 0.00883457f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_335 D N_A_841_47#_c_782_n 0.0662999f $X=6.05 $Y=1.105 $X2=0 $Y2=0
cc_336 N_D_c_420_n N_A_841_47#_c_782_n 0.00849941f $X=5.97 $Y=1.212 $X2=0 $Y2=0
cc_337 N_D_M1006_g N_A_841_47#_c_783_n 5.85252e-19 $X=5.5 $Y=0.56 $X2=0 $Y2=0
cc_338 N_D_M1008_g N_A_841_47#_c_783_n 0.00864756f $X=5.97 $Y=0.56 $X2=0 $Y2=0
cc_339 N_VPWR_c_461_n N_Y_M1010_s 0.00439555f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_340 N_VPWR_c_461_n N_Y_M1007_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_341 N_VPWR_c_461_n N_Y_M1001_d 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_342 N_VPWR_c_461_n N_Y_M1005_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_343 N_VPWR_c_463_n N_Y_c_574_n 0.058597f $X=1.93 $Y=1.66 $X2=0 $Y2=0
cc_344 N_VPWR_c_464_n N_Y_c_574_n 0.048204f $X=2.87 $Y=2 $X2=0 $Y2=0
cc_345 N_VPWR_c_471_n N_Y_c_574_n 0.0187893f $X=2.655 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_461_n N_Y_c_574_n 0.0110885f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_347 N_VPWR_M1014_d N_Y_c_562_n 0.00184299f $X=2.725 $Y=1.485 $X2=0 $Y2=0
cc_348 N_VPWR_c_464_n N_Y_c_562_n 0.0188867f $X=2.87 $Y=2 $X2=0 $Y2=0
cc_349 N_VPWR_c_464_n N_Y_c_578_n 0.0490625f $X=2.87 $Y=2 $X2=0 $Y2=0
cc_350 N_VPWR_c_465_n N_Y_c_578_n 0.0428045f $X=4.25 $Y=2 $X2=0 $Y2=0
cc_351 N_VPWR_c_476_n N_Y_c_578_n 0.0223557f $X=3.725 $Y=2.72 $X2=0 $Y2=0
cc_352 N_VPWR_c_461_n N_Y_c_578_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_353 N_VPWR_M1016_s N_Y_c_563_n 0.00579147f $X=3.665 $Y=1.485 $X2=0 $Y2=0
cc_354 N_VPWR_c_465_n N_Y_c_563_n 0.0280298f $X=4.25 $Y=2 $X2=0 $Y2=0
cc_355 N_VPWR_M1016_s N_Y_c_561_n 0.00544937f $X=3.665 $Y=1.485 $X2=0 $Y2=0
cc_356 N_VPWR_c_465_n N_Y_c_561_n 0.028462f $X=4.25 $Y=2 $X2=0 $Y2=0
cc_357 N_VPWR_c_465_n N_Y_c_603_n 0.0521674f $X=4.25 $Y=2 $X2=0 $Y2=0
cc_358 N_VPWR_c_466_n N_Y_c_603_n 0.0385613f $X=5.24 $Y=2 $X2=0 $Y2=0
cc_359 N_VPWR_c_473_n N_Y_c_603_n 0.0223557f $X=5.155 $Y=2.72 $X2=0 $Y2=0
cc_360 N_VPWR_c_461_n N_Y_c_603_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_361 N_VPWR_M1017_s N_Y_c_565_n 0.00180012f $X=5.095 $Y=1.485 $X2=0 $Y2=0
cc_362 N_VPWR_c_466_n N_Y_c_565_n 0.0139097f $X=5.24 $Y=2 $X2=0 $Y2=0
cc_363 N_VPWR_c_468_n N_Y_c_566_n 0.0146106f $X=6.18 $Y=1.66 $X2=0 $Y2=0
cc_364 N_VPWR_c_466_n N_Y_c_608_n 0.0470327f $X=5.24 $Y=2 $X2=0 $Y2=0
cc_365 N_VPWR_c_468_n N_Y_c_608_n 0.0503631f $X=6.18 $Y=1.66 $X2=0 $Y2=0
cc_366 N_VPWR_c_477_n N_Y_c_608_n 0.0223557f $X=6.095 $Y=2.72 $X2=0 $Y2=0
cc_367 N_VPWR_c_461_n N_Y_c_608_n 0.0140101f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_368 N_VPWR_c_463_n N_Y_c_579_n 0.0133617f $X=1.93 $Y=1.66 $X2=0 $Y2=0
cc_369 N_VPWR_c_468_n N_A_841_47#_c_782_n 0.00204238f $X=6.18 $Y=1.66 $X2=0
+ $Y2=0
cc_370 N_Y_M1003_s N_VGND_c_666_n 0.00256987f $X=2.265 $Y=0.235 $X2=0 $Y2=0
cc_371 N_Y_M1003_s N_A_361_47#_c_731_n 0.00398387f $X=2.265 $Y=0.235 $X2=0 $Y2=0
cc_372 N_Y_c_568_n N_A_361_47#_c_731_n 0.0246284f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_373 N_Y_c_568_n N_A_641_47#_c_756_n 0.0084425f $X=2.4 $Y=0.74 $X2=0 $Y2=0
cc_374 N_Y_c_563_n N_A_641_47#_c_756_n 0.00690462f $X=4.555 $Y=1.555 $X2=0 $Y2=0
cc_375 N_Y_c_561_n N_A_641_47#_c_756_n 0.0509087f $X=4.045 $Y=1.555 $X2=0 $Y2=0
cc_376 N_Y_c_565_n N_A_841_47#_c_781_n 0.00613486f $X=5.495 $Y=1.555 $X2=0 $Y2=0
cc_377 N_VGND_c_666_n N_A_361_47#_M1003_d 0.00389198f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_378 N_VGND_c_666_n N_A_361_47#_M1004_d 0.00255381f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_666_n N_A_361_47#_M1018_d 0.00209344f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_662_n N_A_361_47#_c_736_n 0.123406f $X=5.625 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_666_n N_A_361_47#_c_736_n 0.0768867f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_382 N_VGND_c_666_n N_A_641_47#_M1015_s 0.00256987f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_383 N_VGND_c_666_n N_A_641_47#_M1011_s 0.00256987f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_662_n N_A_641_47#_c_756_n 0.00342407f $X=5.625 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_666_n N_A_641_47#_c_756_n 0.00851921f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_386 N_VGND_c_666_n N_A_841_47#_M1011_d 0.00225742f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_387 N_VGND_c_666_n N_A_841_47#_M1019_d 0.00265084f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_666_n N_A_841_47#_M1008_d 0.00209319f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_c_662_n N_A_841_47#_c_780_n 0.056955f $X=5.625 $Y=0 $X2=0 $Y2=0
cc_390 N_VGND_c_666_n N_A_841_47#_c_780_n 0.0356031f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_662_n N_A_841_47#_c_802_n 0.0159994f $X=5.625 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_666_n N_A_841_47#_c_802_n 0.00961652f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_M1006_s N_A_841_47#_c_782_n 0.00251598f $X=5.575 $Y=0.235 $X2=0
+ $Y2=0
cc_394 N_VGND_c_661_n N_A_841_47#_c_782_n 0.0127122f $X=5.71 $Y=0.4 $X2=0 $Y2=0
cc_395 N_VGND_c_662_n N_A_841_47#_c_782_n 0.00248202f $X=5.625 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_665_n N_A_841_47#_c_782_n 0.00194552f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_666_n N_A_841_47#_c_782_n 0.00966112f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_c_661_n N_A_841_47#_c_783_n 0.0231432f $X=5.71 $Y=0.4 $X2=0 $Y2=0
cc_399 N_VGND_c_665_n N_A_841_47#_c_783_n 0.024373f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_666_n N_A_841_47#_c_783_n 0.0141066f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_401 N_A_361_47#_c_731_n N_A_641_47#_M1015_s 0.00400026f $X=3.81 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_402 N_A_361_47#_M1018_d N_A_641_47#_c_756_n 0.00312742f $X=3.675 $Y=0.235
+ $X2=0 $Y2=0
cc_403 N_A_361_47#_c_731_n N_A_641_47#_c_756_n 0.0479647f $X=3.81 $Y=0.4 $X2=0
+ $Y2=0
cc_404 N_A_361_47#_c_731_n N_A_841_47#_c_780_n 0.0197364f $X=3.81 $Y=0.4 $X2=0
+ $Y2=0
cc_405 N_A_641_47#_c_756_n N_A_841_47#_M1011_d 0.00358914f $X=4.77 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_406 N_A_641_47#_M1011_s N_A_841_47#_c_780_n 0.00401739f $X=4.635 $Y=0.235
+ $X2=0 $Y2=0
cc_407 N_A_641_47#_c_756_n N_A_841_47#_c_780_n 0.0443916f $X=4.77 $Y=0.74 $X2=0
+ $Y2=0
cc_408 N_A_641_47#_c_756_n N_A_841_47#_c_781_n 0.00140356f $X=4.77 $Y=0.74 $X2=0
+ $Y2=0
