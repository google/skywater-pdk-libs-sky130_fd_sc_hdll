* File: sky130_fd_sc_hdll__nor3_1.pxi.spice
* Created: Thu Aug 27 19:16:11 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3_1%C N_C_c_38_n N_C_M1003_g N_C_c_35_n N_C_M1004_g C
+ N_C_c_37_n PM_SKY130_FD_SC_HDLL__NOR3_1%C
x_PM_SKY130_FD_SC_HDLL__NOR3_1%B N_B_c_65_n N_B_M1000_g N_B_c_66_n N_B_M1001_g
+ N_B_c_67_n B B PM_SKY130_FD_SC_HDLL__NOR3_1%B
x_PM_SKY130_FD_SC_HDLL__NOR3_1%A N_A_c_102_n N_A_M1002_g N_A_c_105_n N_A_M1005_g
+ A A A N_A_c_104_n PM_SKY130_FD_SC_HDLL__NOR3_1%A
x_PM_SKY130_FD_SC_HDLL__NOR3_1%Y N_Y_M1004_s N_Y_M1001_d N_Y_M1003_s N_Y_c_138_n
+ N_Y_c_141_n N_Y_c_154_n N_Y_c_133_n N_Y_c_134_n Y N_Y_c_136_n N_Y_c_137_n Y
+ PM_SKY130_FD_SC_HDLL__NOR3_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR3_1%VPWR N_VPWR_M1005_d N_VPWR_c_196_n N_VPWR_c_197_n
+ VPWR N_VPWR_c_198_n N_VPWR_c_195_n PM_SKY130_FD_SC_HDLL__NOR3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3_1%VGND N_VGND_M1004_d N_VGND_M1002_d N_VGND_c_219_n
+ VGND N_VGND_c_220_n N_VGND_c_221_n N_VGND_c_222_n N_VGND_c_223_n
+ N_VGND_c_224_n PM_SKY130_FD_SC_HDLL__NOR3_1%VGND
cc_1 VNB N_C_c_35_n 0.0221314f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB C 0.0146493f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_C_c_37_n 0.0365272f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_c_65_n 0.0229924f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_c_66_n 0.0169241f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B_c_67_n 0.00218519f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.16
cc_7 VNB N_A_c_102_n 0.018137f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB A 0.0283514f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_9 VNB N_A_c_104_n 0.0471122f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_Y_c_133_n 0.00287947f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_Y_c_134_n 0.017363f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_195_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_VGND_c_219_n 0.00214285f $X=-0.19 $Y=-0.24 $X2=0.26 $Y2=1.202
cc_14 VNB N_VGND_c_220_n 0.0149052f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_15 VNB N_VGND_c_221_n 0.0139729f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_222_n 0.00573782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_223_n 0.0344539f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_224_n 0.142854f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_C_c_38_n 0.0212409f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_20 VPB C 0.00356082f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_21 VPB N_C_c_37_n 0.0177787f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_22 VPB N_B_c_65_n 0.0274686f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_23 VPB N_B_c_67_n 6.11484e-19 $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_24 VPB B 0.00224805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_25 VPB N_A_c_105_n 0.0189903f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_26 VPB A 0.0176689f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_27 VPB N_A_c_104_n 0.0215864f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_Y_c_133_n 0.00137192f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_Y_c_136_n 0.00753565f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_Y_c_137_n 0.030912f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_196_n 0.0175109f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_32 VPB N_VPWR_c_197_n 0.0342222f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_33 VPB N_VPWR_c_198_n 0.0404685f $X=-0.19 $Y=1.305 $X2=0.26 $Y2=1.16
cc_34 VPB N_VPWR_c_195_n 0.0445202f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 N_C_c_38_n N_B_c_65_n 0.0499809f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_36 C N_B_c_65_n 2.18763e-19 $X=0.15 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_37 N_C_c_37_n N_B_c_65_n 0.0251016f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_38 N_C_c_35_n N_B_c_66_n 0.0212683f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_39 C N_B_c_67_n 0.0254977f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_40 N_C_c_37_n N_B_c_67_n 0.00285958f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_41 N_C_c_38_n B 0.00467476f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_42 N_C_c_37_n B 0.00241518f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_43 N_C_c_35_n N_Y_c_138_n 0.0151348f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_44 C N_Y_c_138_n 0.00454953f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_45 N_C_c_37_n N_Y_c_138_n 4.76291e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_46 N_C_c_38_n N_Y_c_141_n 0.0130498f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_47 N_C_c_35_n N_Y_c_134_n 5.27683e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_48 C N_Y_c_134_n 0.0204953f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_49 N_C_c_37_n N_Y_c_134_n 0.0016628f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_50 N_C_c_38_n N_Y_c_136_n 4.79874e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_C_c_38_n N_Y_c_137_n 0.0107395f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 C N_Y_c_137_n 0.0251904f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_53 N_C_c_37_n N_Y_c_137_n 0.00199455f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_54 N_C_c_38_n N_VPWR_c_198_n 0.00433173f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_C_c_38_n N_VPWR_c_195_n 0.00700698f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_56 N_C_c_35_n N_VGND_c_219_n 0.01594f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_57 N_C_c_35_n N_VGND_c_220_n 0.00199015f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 N_C_c_35_n N_VGND_c_224_n 0.00369362f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_59 N_B_c_66_n N_A_c_102_n 0.0229484f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_60 N_B_c_65_n N_A_c_105_n 0.049532f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_61 B N_A_c_105_n 5.2765e-19 $X=0.66 $Y=1.445 $X2=0 $Y2=0
cc_62 N_B_c_65_n N_A_c_104_n 0.0242211f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B_c_67_n N_A_c_104_n 3.12362e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B_c_65_n N_Y_c_138_n 0.00250966f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_65 N_B_c_66_n N_Y_c_138_n 0.0109919f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_66 N_B_c_67_n N_Y_c_138_n 0.0314391f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_65_n N_Y_c_141_n 0.0163163f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 B N_Y_c_141_n 0.00909094f $X=0.66 $Y=1.445 $X2=0 $Y2=0
cc_69 N_B_c_65_n N_Y_c_154_n 2.67351e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B_c_65_n N_Y_c_133_n 0.012736f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_71 N_B_c_66_n N_Y_c_133_n 0.00343469f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B_c_67_n N_Y_c_133_n 0.0254975f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_73 B N_Y_c_133_n 0.0277874f $X=0.66 $Y=1.445 $X2=0 $Y2=0
cc_74 N_B_c_65_n N_Y_c_137_n 0.00161399f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_75 B A_117_297# 0.00377224f $X=0.66 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_76 N_B_c_65_n N_VPWR_c_198_n 0.00433201f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B_c_65_n N_VPWR_c_195_n 0.00612629f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B_c_66_n N_VGND_c_219_n 0.0016282f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B_c_66_n N_VGND_c_221_n 0.00428022f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B_c_66_n N_VGND_c_223_n 8.80204e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_66_n N_VGND_c_224_n 0.00585784f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_105_n N_Y_c_141_n 0.00517469f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_c_102_n N_Y_c_154_n 0.00589126f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_84 A N_Y_c_154_n 0.00871801f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_c_102_n N_Y_c_133_n 0.00403226f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_c_105_n N_Y_c_133_n 0.0242279f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_87 A N_Y_c_133_n 0.0384861f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_c_104_n N_Y_c_133_n 0.0126098f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_89 A N_VPWR_M1005_d 0.00991436f $X=1.96 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_90 N_A_c_105_n N_VPWR_c_197_n 0.00780701f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_91 A N_VPWR_c_197_n 0.0391779f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_92 N_A_c_104_n N_VPWR_c_197_n 0.00568923f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_c_105_n N_VPWR_c_198_n 0.00597653f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_105_n N_VPWR_c_195_n 0.0113087f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_95 A N_VGND_M1002_d 0.0103562f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_96 N_A_c_102_n N_VGND_c_221_n 0.00382526f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_c_102_n N_VGND_c_223_n 0.0106627f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_98 A N_VGND_c_223_n 0.0375024f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_99 N_A_c_104_n N_VGND_c_223_n 0.00779123f $X=1.435 $Y=1.202 $X2=0 $Y2=0
cc_100 N_A_c_102_n N_VGND_c_224_n 0.00534016f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_101 A N_VGND_c_224_n 0.00297073f $X=1.96 $Y=0.765 $X2=0 $Y2=0
cc_102 N_Y_c_141_n A_117_297# 0.00403673f $X=1.245 $Y=2.365 $X2=-0.19 $Y2=-0.24
cc_103 N_Y_c_141_n A_211_297# 0.00674245f $X=1.245 $Y=2.365 $X2=-0.19 $Y2=-0.24
cc_104 N_Y_c_133_n A_211_297# 0.00923569f $X=1.33 $Y=2.28 $X2=-0.19 $Y2=-0.24
cc_105 N_Y_c_141_n N_VPWR_c_197_n 0.0146277f $X=1.245 $Y=2.365 $X2=0 $Y2=0
cc_106 N_Y_c_133_n N_VPWR_c_197_n 0.0345065f $X=1.33 $Y=2.28 $X2=0 $Y2=0
cc_107 N_Y_c_141_n N_VPWR_c_198_n 0.0513508f $X=1.245 $Y=2.365 $X2=0 $Y2=0
cc_108 N_Y_c_136_n N_VPWR_c_198_n 0.0196458f $X=0.257 $Y=2.28 $X2=0 $Y2=0
cc_109 N_Y_M1003_s N_VPWR_c_195_n 0.00218082f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_110 N_Y_c_141_n N_VPWR_c_195_n 0.0348664f $X=1.245 $Y=2.365 $X2=0 $Y2=0
cc_111 N_Y_c_136_n N_VPWR_c_195_n 0.0126395f $X=0.257 $Y=2.28 $X2=0 $Y2=0
cc_112 N_Y_c_138_n N_VGND_M1004_d 0.00418829f $X=1.115 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_113 N_Y_c_138_n N_VGND_c_219_n 0.0214497f $X=1.115 $Y=0.74 $X2=0 $Y2=0
cc_114 N_Y_c_134_n N_VGND_c_219_n 0.0076929f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_115 N_Y_c_138_n N_VGND_c_220_n 0.00232807f $X=1.115 $Y=0.74 $X2=0 $Y2=0
cc_116 N_Y_c_134_n N_VGND_c_220_n 0.00938511f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_117 N_Y_c_138_n N_VGND_c_221_n 0.0029785f $X=1.115 $Y=0.74 $X2=0 $Y2=0
cc_118 N_Y_c_154_n N_VGND_c_221_n 0.00790924f $X=1.33 $Y=0.825 $X2=0 $Y2=0
cc_119 N_Y_M1004_s N_VGND_c_224_n 0.00305109f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_120 N_Y_M1001_d N_VGND_c_224_n 0.00266592f $X=1.065 $Y=0.235 $X2=0 $Y2=0
cc_121 N_Y_c_138_n N_VGND_c_224_n 0.011334f $X=1.115 $Y=0.74 $X2=0 $Y2=0
cc_122 N_Y_c_154_n N_VGND_c_224_n 0.00944761f $X=1.33 $Y=0.825 $X2=0 $Y2=0
cc_123 N_Y_c_134_n N_VGND_c_224_n 0.00892296f $X=0.26 $Y=0.55 $X2=0 $Y2=0
cc_124 A_117_297# N_VPWR_c_195_n 0.00233531f $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_125 A_211_297# N_VPWR_c_195_n 0.00233512f $X=1.055 $Y=1.485 $X2=0.26 $Y2=0.55
