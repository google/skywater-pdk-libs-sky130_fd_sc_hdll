* File: sky130_fd_sc_hdll__nand2_12.pex.spice
* Created: Thu Aug 27 19:12:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%B 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61
+ 63 64 66 67 69 70 72 73 102 103
r252 103 104 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.665 $Y=1.202
+ $X2=5.69 $Y2=1.202
r253 101 103 8.53679 $w=3.67e-07 $l=6.5e-08 $layer=POLY_cond $X=5.6 $Y=1.202
+ $X2=5.665 $Y2=1.202
r254 101 102 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=5.6
+ $Y=1.16 $X2=5.6 $Y2=1.16
r255 99 101 53.1907 $w=3.67e-07 $l=4.05e-07 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.6 $Y2=1.202
r256 98 99 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.202
+ $X2=5.195 $Y2=1.202
r257 97 98 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=4.75 $Y=1.202
+ $X2=5.17 $Y2=1.202
r258 96 97 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.725 $Y=1.202
+ $X2=4.75 $Y2=1.202
r259 95 96 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.725 $Y2=1.202
r260 94 95 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.202
+ $X2=4.255 $Y2=1.202
r261 93 94 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=3.81 $Y=1.202
+ $X2=4.23 $Y2=1.202
r262 92 93 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=3.81 $Y2=1.202
r263 91 92 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.785 $Y2=1.202
r264 90 91 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.202
+ $X2=3.315 $Y2=1.202
r265 89 90 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=2.87 $Y=1.202
+ $X2=3.29 $Y2=1.202
r266 88 89 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=2.87 $Y2=1.202
r267 87 88 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.845 $Y2=1.202
r268 86 87 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r269 85 86 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=1.93 $Y=1.202
+ $X2=2.35 $Y2=1.202
r270 84 85 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.202
+ $X2=1.93 $Y2=1.202
r271 83 84 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.905 $Y2=1.202
r272 82 83 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.202
+ $X2=1.435 $Y2=1.202
r273 81 82 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.41 $Y2=1.202
r274 80 81 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r275 78 80 61.0708 $w=3.67e-07 $l=4.65e-07 $layer=POLY_cond $X=0.5 $Y=1.202
+ $X2=0.965 $Y2=1.202
r276 78 79 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=0.5
+ $Y=1.16 $X2=0.5 $Y2=1.16
r277 76 78 0.656676 $w=3.67e-07 $l=5e-09 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.5 $Y2=1.202
r278 75 76 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r279 73 102 111.403 $w=2.68e-07 $l=2.61e-06 $layer=LI1_cond $X=2.99 $Y=1.19
+ $X2=5.6 $Y2=1.19
r280 73 79 106.281 $w=2.68e-07 $l=2.49e-06 $layer=LI1_cond $X=2.99 $Y=1.19
+ $X2=0.5 $Y2=1.19
r281 70 104 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r282 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r283 67 103 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r284 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r285 64 99 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r286 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r287 61 98 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=1.202
r288 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.17 $Y=0.995
+ $X2=5.17 $Y2=0.56
r289 58 97 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=1.202
r290 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.75 $Y=0.995
+ $X2=4.75 $Y2=0.56
r291 55 96 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r292 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r293 52 95 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r294 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r295 49 94 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=1.202
r296 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.23 $Y=0.995
+ $X2=4.23 $Y2=0.56
r297 46 93 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=1.202
r298 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.81 $Y=0.995
+ $X2=3.81 $Y2=0.56
r299 43 92 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r300 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r301 40 91 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r302 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r303 37 90 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=1.202
r304 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.29 $Y=0.995
+ $X2=3.29 $Y2=0.56
r305 34 89 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=1.202
r306 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.87 $Y=0.995
+ $X2=2.87 $Y2=0.56
r307 31 88 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r308 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r309 28 87 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r310 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r311 25 86 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r312 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r313 22 85 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=1.202
r314 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r315 19 84 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.202
r316 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r317 16 83 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r318 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r319 13 82 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=1.202
r320 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.41 $Y=0.995
+ $X2=1.41 $Y2=0.56
r321 10 81 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r322 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r323 7 80 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r324 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r325 4 76 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r326 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r327 1 75 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r328 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61
+ 63 64 66 67 69 70 72 73 100 103
r195 103 104 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=11.305 $Y=1.202
+ $X2=11.33 $Y2=1.202
r196 102 103 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=10.835 $Y=1.202
+ $X2=11.305 $Y2=1.202
r197 101 102 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.81 $Y=1.202
+ $X2=10.835 $Y2=1.202
r198 99 101 36.7738 $w=3.67e-07 $l=2.8e-07 $layer=POLY_cond $X=10.53 $Y=1.202
+ $X2=10.81 $Y2=1.202
r199 99 100 24.2133 $w=1.7e-07 $l=1.02e-06 $layer=licon1_POLY $count=6 $X=10.53
+ $Y=1.16 $X2=10.53 $Y2=1.16
r200 97 99 18.3869 $w=3.67e-07 $l=1.4e-07 $layer=POLY_cond $X=10.39 $Y=1.202
+ $X2=10.53 $Y2=1.202
r201 96 97 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=10.365 $Y=1.202
+ $X2=10.39 $Y2=1.202
r202 95 96 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=9.895 $Y=1.202
+ $X2=10.365 $Y2=1.202
r203 94 95 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.87 $Y=1.202
+ $X2=9.895 $Y2=1.202
r204 93 94 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=9.425 $Y=1.202
+ $X2=9.87 $Y2=1.202
r205 92 93 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=9.4 $Y=1.202
+ $X2=9.425 $Y2=1.202
r206 91 92 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=8.955 $Y=1.202
+ $X2=9.4 $Y2=1.202
r207 90 91 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.93 $Y=1.202
+ $X2=8.955 $Y2=1.202
r208 89 90 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=8.51 $Y=1.202
+ $X2=8.93 $Y2=1.202
r209 88 89 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=8.485 $Y=1.202
+ $X2=8.51 $Y2=1.202
r210 87 88 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=8.015 $Y=1.202
+ $X2=8.485 $Y2=1.202
r211 86 87 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.99 $Y=1.202
+ $X2=8.015 $Y2=1.202
r212 85 86 55.1608 $w=3.67e-07 $l=4.2e-07 $layer=POLY_cond $X=7.57 $Y=1.202
+ $X2=7.99 $Y2=1.202
r213 84 85 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.545 $Y=1.202
+ $X2=7.57 $Y2=1.202
r214 83 84 61.7275 $w=3.67e-07 $l=4.7e-07 $layer=POLY_cond $X=7.075 $Y=1.202
+ $X2=7.545 $Y2=1.202
r215 82 83 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.202
+ $X2=7.075 $Y2=1.202
r216 80 82 34.1471 $w=3.67e-07 $l=2.6e-07 $layer=POLY_cond $X=6.79 $Y=1.202
+ $X2=7.05 $Y2=1.202
r217 80 81 24.2133 $w=1.7e-07 $l=1.02e-06 $layer=licon1_POLY $count=6 $X=6.79
+ $Y=1.16 $X2=6.79 $Y2=1.16
r218 78 80 24.297 $w=3.67e-07 $l=1.85e-07 $layer=POLY_cond $X=6.605 $Y=1.202
+ $X2=6.79 $Y2=1.202
r219 77 78 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.202
+ $X2=6.605 $Y2=1.202
r220 76 77 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=6.135 $Y=1.202
+ $X2=6.58 $Y2=1.202
r221 75 76 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.202
+ $X2=6.135 $Y2=1.202
r222 73 100 66.5856 $w=2.68e-07 $l=1.56e-06 $layer=LI1_cond $X=8.97 $Y=1.19
+ $X2=10.53 $Y2=1.19
r223 73 81 93.0491 $w=2.68e-07 $l=2.18e-06 $layer=LI1_cond $X=8.97 $Y=1.19
+ $X2=6.79 $Y2=1.19
r224 70 104 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=11.33 $Y=0.995
+ $X2=11.33 $Y2=1.202
r225 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=11.33 $Y=0.995
+ $X2=11.33 $Y2=0.56
r226 67 103 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.202
r227 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.305 $Y=1.41
+ $X2=11.305 $Y2=1.985
r228 64 102 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.202
r229 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.835 $Y=1.41
+ $X2=10.835 $Y2=1.985
r230 61 101 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.81 $Y=0.995
+ $X2=10.81 $Y2=1.202
r231 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.81 $Y=0.995
+ $X2=10.81 $Y2=0.56
r232 58 97 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.39 $Y=0.995
+ $X2=10.39 $Y2=1.202
r233 58 60 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.39 $Y=0.995
+ $X2=10.39 $Y2=0.56
r234 55 96 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.202
r235 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.985
r236 52 95 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.202
r237 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.985
r238 49 94 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.87 $Y=0.995
+ $X2=9.87 $Y2=1.202
r239 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.87 $Y=0.995
+ $X2=9.87 $Y2=0.56
r240 46 93 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.202
r241 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.985
r242 43 92 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.4 $Y=0.995 $X2=9.4
+ $Y2=1.202
r243 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.4 $Y=0.995
+ $X2=9.4 $Y2=0.56
r244 40 91 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.202
r245 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.985
r246 37 90 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.93 $Y=0.995
+ $X2=8.93 $Y2=1.202
r247 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.93 $Y=0.995
+ $X2=8.93 $Y2=0.56
r248 34 89 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.51 $Y=0.995
+ $X2=8.51 $Y2=1.202
r249 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.51 $Y=0.995
+ $X2=8.51 $Y2=0.56
r250 31 88 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.202
r251 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.985
r252 28 87 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.202
r253 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.985
r254 25 86 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.99 $Y=0.995
+ $X2=7.99 $Y2=1.202
r255 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.99 $Y=0.995
+ $X2=7.99 $Y2=0.56
r256 22 85 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=1.202
r257 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.57 $Y=0.995
+ $X2=7.57 $Y2=0.56
r258 19 84 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.202
r259 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r260 16 83 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.202
r261 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r262 13 82 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=1.202
r263 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.05 $Y=0.995
+ $X2=7.05 $Y2=0.56
r264 10 78 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.202
r265 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r266 7 77 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=1.202
r267 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.58 $Y=0.995
+ $X2=6.58 $Y2=0.56
r268 4 76 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.202
r269 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r270 1 75 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=1.202
r271 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.11 $Y=0.995
+ $X2=6.11 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 40 42
+ 48 50 54 56 60 62 66 68 72 76 80 84 88 92 96 100 105 106 108 109 111 112 114
+ 115 117 118 120 121 122 123 124 125 127 156 161 164 167 170 173
r175 173 174 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r176 171 174 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r177 170 171 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 168 171 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r179 167 168 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r180 165 168 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r181 164 165 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r182 162 165 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r183 161 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r184 155 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r185 153 156 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.27 $Y=2.72
+ $X2=11.73 $Y2=2.72
r186 152 153 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r187 150 153 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r188 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r189 147 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r190 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r191 144 147 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r192 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r193 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r194 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r195 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r196 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r197 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r198 135 174 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=4.83 $Y2=2.72
r199 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r200 132 173 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=4.96 $Y2=2.72
r201 132 134 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=5.095 $Y=2.72
+ $X2=5.75 $Y2=2.72
r202 131 162 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r203 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r204 128 158 4.1687 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r205 128 130 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r206 127 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=1.2 $Y2=2.72
r207 127 130 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.065 $Y=2.72
+ $X2=0.69 $Y2=2.72
r208 125 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r209 125 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r210 123 152 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=11.405 $Y=2.72
+ $X2=11.27 $Y2=2.72
r211 123 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.405 $Y=2.72
+ $X2=11.54 $Y2=2.72
r212 122 155 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=11.675 $Y=2.72
+ $X2=11.73 $Y2=2.72
r213 122 124 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=11.675 $Y=2.72
+ $X2=11.54 $Y2=2.72
r214 120 149 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.35 $Y2=2.72
r215 120 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.465 $Y=2.72
+ $X2=10.6 $Y2=2.72
r216 119 152 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=10.735 $Y=2.72
+ $X2=11.27 $Y2=2.72
r217 119 121 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=10.735 $Y=2.72
+ $X2=10.6 $Y2=2.72
r218 117 146 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.43 $Y2=2.72
r219 117 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.525 $Y=2.72
+ $X2=9.66 $Y2=2.72
r220 116 149 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=10.35 $Y2=2.72
r221 116 118 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=9.795 $Y=2.72
+ $X2=9.66 $Y2=2.72
r222 114 143 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=8.585 $Y=2.72
+ $X2=8.51 $Y2=2.72
r223 114 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.585 $Y=2.72
+ $X2=8.72 $Y2=2.72
r224 113 146 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=9.43 $Y2=2.72
r225 113 115 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.855 $Y=2.72
+ $X2=8.72 $Y2=2.72
r226 111 140 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.59 $Y2=2.72
r227 111 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.645 $Y=2.72
+ $X2=7.78 $Y2=2.72
r228 110 143 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=7.915 $Y=2.72
+ $X2=8.51 $Y2=2.72
r229 110 112 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.915 $Y=2.72
+ $X2=7.78 $Y2=2.72
r230 108 137 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.705 $Y=2.72
+ $X2=6.67 $Y2=2.72
r231 108 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.705 $Y=2.72
+ $X2=6.84 $Y2=2.72
r232 107 140 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=7.59 $Y2=2.72
r233 107 109 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.975 $Y=2.72
+ $X2=6.84 $Y2=2.72
r234 105 134 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.75 $Y2=2.72
r235 105 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.765 $Y=2.72
+ $X2=5.9 $Y2=2.72
r236 104 137 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r237 104 106 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.035 $Y=2.72
+ $X2=5.9 $Y2=2.72
r238 100 103 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=11.54 $Y=1.66
+ $X2=11.54 $Y2=2.34
r239 98 124 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=11.54 $Y=2.635
+ $X2=11.54 $Y2=2.72
r240 98 103 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.54 $Y=2.635
+ $X2=11.54 $Y2=2.34
r241 94 121 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2.72
r242 94 96 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2
r243 90 118 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r244 90 92 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2
r245 86 115 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2.72
r246 86 88 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2
r247 82 112 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.72
r248 82 84 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2
r249 78 109 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r250 78 80 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2
r251 74 106 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r252 74 76 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2
r253 70 173 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r254 70 72 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2
r255 69 170 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.02 $Y2=2.72
r256 68 173 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.96 $Y2=2.72
r257 68 69 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.825 $Y=2.72
+ $X2=4.155 $Y2=2.72
r258 64 170 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r259 64 66 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r260 63 167 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.08 $Y2=2.72
r261 62 170 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.02 $Y2=2.72
r262 62 63 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=3.215 $Y2=2.72
r263 58 167 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r264 58 60 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r265 57 164 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.14 $Y2=2.72
r266 56 167 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=3.08 $Y2=2.72
r267 56 57 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.945 $Y=2.72
+ $X2=2.275 $Y2=2.72
r268 52 164 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r269 52 54 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r270 51 161 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.2 $Y2=2.72
r271 50 164 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=2.14 $Y2=2.72
r272 50 51 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=2.72
+ $X2=1.335 $Y2=2.72
r273 46 161 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r274 46 48 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r275 42 45 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r276 40 158 3.116 $w=2.7e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.197 $Y2=2.72
r277 40 45 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r278 13 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=1.485 $X2=11.54 $Y2=2.34
r279 13 100 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=11.395
+ $Y=1.485 $X2=11.54 $Y2=1.66
r280 12 96 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.455
+ $Y=1.485 $X2=10.6 $Y2=2
r281 11 92 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.515
+ $Y=1.485 $X2=9.66 $Y2=2
r282 10 88 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=2
r283 9 84 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2
r284 8 80 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2
r285 7 76 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2
r286 6 72 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r287 5 66 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r288 4 60 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r289 3 54 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r290 2 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r291 1 45 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r292 1 42 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%Y 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 17 18 55 57 59 63 65 69 71 75 77 81 83 87 89 91 95 97 107 111 113 117 119 123
+ 125 129 131 135 137 140 144 146 148 150 152 155 159 161 163 165 167 170 171
+ 172 178 180
r252 175 180 1.96759 $w=4.08e-07 $l=7e-08 $layer=LI1_cond $X=6.25 $Y=1.26
+ $X2=6.25 $Y2=1.19
r253 172 180 0.224867 $w=4.08e-07 $l=8e-09 $layer=LI1_cond $X=6.25 $Y=1.182
+ $X2=6.25 $Y2=1.19
r254 172 178 4.42096 $w=4.08e-07 $l=1.27e-07 $layer=LI1_cond $X=6.25 $Y=1.182
+ $X2=6.25 $Y2=1.055
r255 172 175 0.196759 $w=4.08e-07 $l=7e-09 $layer=LI1_cond $X=6.25 $Y=1.267
+ $X2=6.25 $Y2=1.26
r256 170 171 6.87109 $w=4.68e-07 $l=2.7e-07 $layer=LI1_cond $X=11.2 $Y=1.055
+ $X2=11.2 $Y2=1.325
r257 153 172 6.40871 $w=4.08e-07 $l=2.28e-07 $layer=LI1_cond $X=6.25 $Y=1.495
+ $X2=6.25 $Y2=1.267
r258 153 155 1.06026 $w=4.1e-07 $l=1.03078e-07 $layer=LI1_cond $X=6.25 $Y=1.495
+ $X2=6.29 $Y2=1.58
r259 140 167 3.14896 $w=3e-07 $l=9.88686e-08 $layer=LI1_cond $X=11.1 $Y=1.495
+ $X2=11.07 $Y2=1.58
r260 140 171 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.1 $Y=1.495
+ $X2=11.1 $Y2=1.325
r261 137 169 3.28347 $w=2.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.1 $Y=0.885
+ $X2=11.1 $Y2=0.76
r262 137 170 7.25612 $w=2.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.1 $Y=0.885
+ $X2=11.1 $Y2=1.055
r263 133 167 3.14896 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.07 $Y=1.665
+ $X2=11.07 $Y2=1.58
r264 133 135 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=11.07 $Y=1.665
+ $X2=11.07 $Y2=2.34
r265 132 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.295 $Y=1.58
+ $X2=10.13 $Y2=1.58
r266 131 167 3.44808 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=10.905 $Y=1.58
+ $X2=11.07 $Y2=1.58
r267 131 132 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=10.905 $Y=1.58
+ $X2=10.295 $Y2=1.58
r268 127 165 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.13 $Y=1.665
+ $X2=10.13 $Y2=1.58
r269 127 129 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.13 $Y=1.665
+ $X2=10.13 $Y2=2.34
r270 126 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.355 $Y=1.58
+ $X2=9.19 $Y2=1.58
r271 125 165 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.965 $Y=1.58
+ $X2=10.13 $Y2=1.58
r272 125 126 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.965 $Y=1.58
+ $X2=9.355 $Y2=1.58
r273 121 163 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.19 $Y=1.665
+ $X2=9.19 $Y2=1.58
r274 121 123 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.19 $Y=1.665
+ $X2=9.19 $Y2=2.34
r275 120 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.415 $Y=1.58
+ $X2=8.25 $Y2=1.58
r276 119 163 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.025 $Y=1.58
+ $X2=9.19 $Y2=1.58
r277 119 120 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=9.025 $Y=1.58
+ $X2=8.415 $Y2=1.58
r278 115 161 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=8.25 $Y=1.665
+ $X2=8.25 $Y2=1.58
r279 115 117 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=8.25 $Y=1.665
+ $X2=8.25 $Y2=2.34
r280 114 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.475 $Y=1.58
+ $X2=7.31 $Y2=1.58
r281 113 161 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.085 $Y=1.58
+ $X2=8.25 $Y2=1.58
r282 113 114 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=8.085 $Y=1.58
+ $X2=7.475 $Y2=1.58
r283 109 159 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.31 $Y2=1.58
r284 109 111 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.31 $Y=1.665
+ $X2=7.31 $Y2=2.34
r285 108 155 5.68638 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=6.535 $Y=1.58
+ $X2=6.29 $Y2=1.58
r286 107 159 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=7.31 $Y2=1.58
r287 107 108 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.145 $Y=1.58
+ $X2=6.535 $Y2=1.58
r288 104 106 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=9.19 $Y=0.76
+ $X2=10.13 $Y2=0.76
r289 102 104 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=8.25 $Y=0.76
+ $X2=9.19 $Y2=0.76
r290 100 102 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=7.31 $Y=0.76
+ $X2=8.25 $Y2=0.76
r291 98 157 3.75819 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=6.455 $Y=0.76
+ $X2=6.305 $Y2=0.76
r292 98 100 39.4136 $w=2.48e-07 $l=8.55e-07 $layer=LI1_cond $X=6.455 $Y=0.76
+ $X2=7.31 $Y2=0.76
r293 97 169 3.54615 $w=2.5e-07 $l=1.35e-07 $layer=LI1_cond $X=10.965 $Y=0.76
+ $X2=11.1 $Y2=0.76
r294 97 106 38.4916 $w=2.48e-07 $l=8.35e-07 $layer=LI1_cond $X=10.965 $Y=0.76
+ $X2=10.13 $Y2=0.76
r295 93 155 1.06026 $w=3.3e-07 $l=1.18427e-07 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.29 $Y2=1.58
r296 93 95 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.37 $Y=1.665
+ $X2=6.37 $Y2=2.34
r297 91 157 3.13183 $w=3e-07 $l=1.25e-07 $layer=LI1_cond $X=6.305 $Y=0.885
+ $X2=6.305 $Y2=0.76
r298 91 178 6.53051 $w=2.98e-07 $l=1.7e-07 $layer=LI1_cond $X=6.305 $Y=0.885
+ $X2=6.305 $Y2=1.055
r299 90 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.595 $Y=1.58
+ $X2=5.43 $Y2=1.58
r300 89 155 5.68638 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=6.29 $Y2=1.58
r301 89 90 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=5.595 $Y2=1.58
r302 85 152 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=1.58
r303 85 87 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.43 $Y=1.665
+ $X2=5.43 $Y2=2.34
r304 84 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.655 $Y=1.58
+ $X2=4.49 $Y2=1.58
r305 83 152 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=5.43 $Y2=1.58
r306 83 84 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.265 $Y=1.58
+ $X2=4.655 $Y2=1.58
r307 79 150 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=1.58
r308 79 81 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.49 $Y=1.665
+ $X2=4.49 $Y2=2.34
r309 78 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.715 $Y=1.58
+ $X2=3.55 $Y2=1.58
r310 77 150 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=4.49 $Y2=1.58
r311 77 78 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.325 $Y=1.58
+ $X2=3.715 $Y2=1.58
r312 73 148 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=1.58
r313 73 75 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.55 $Y=1.665
+ $X2=3.55 $Y2=2.34
r314 72 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.775 $Y=1.58
+ $X2=2.61 $Y2=1.58
r315 71 148 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=3.55 $Y2=1.58
r316 71 72 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.385 $Y=1.58
+ $X2=2.775 $Y2=1.58
r317 67 146 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=1.58
r318 67 69 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.61 $Y=1.665
+ $X2=2.61 $Y2=2.34
r319 66 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.58
+ $X2=1.67 $Y2=1.58
r320 65 146 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=2.61 $Y2=1.58
r321 65 66 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.445 $Y=1.58
+ $X2=1.835 $Y2=1.58
r322 61 144 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=1.58
r323 61 63 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.67 $Y=1.665
+ $X2=1.67 $Y2=2.34
r324 60 142 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.73 $Y2=1.58
r325 59 144 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=1.67 $Y2=1.58
r326 59 60 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.505 $Y=1.58
+ $X2=0.895 $Y2=1.58
r327 55 142 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=1.58
r328 55 57 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=0.73 $Y=1.665
+ $X2=0.73 $Y2=2.34
r329 18 167 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.925
+ $Y=1.485 $X2=11.07 $Y2=1.66
r330 18 135 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.925
+ $Y=1.485 $X2=11.07 $Y2=2.34
r331 17 165 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=1.66
r332 17 129 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=2.34
r333 16 163 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=1.66
r334 16 123 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=2.34
r335 15 161 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=1.66
r336 15 117 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=2.34
r337 14 159 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.66
r338 14 111 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.34
r339 13 155 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.66
r340 13 95 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.34
r341 12 152 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.66
r342 12 87 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.34
r343 11 150 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.66
r344 11 81 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.34
r345 10 148 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.66
r346 10 75 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.34
r347 9 146 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.66
r348 9 69 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r349 8 144 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r350 8 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r351 7 142 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r352 7 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r353 6 169 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=10.885
+ $Y=0.235 $X2=11.07 $Y2=0.72
r354 5 106 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.13 $Y2=0.72
r355 4 104 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=9.005
+ $Y=0.235 $X2=9.19 $Y2=0.72
r356 3 102 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=8.065
+ $Y=0.235 $X2=8.25 $Y2=0.72
r357 2 100 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.72
r358 1 157 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 12 13 42
+ 44 45 48 50 54 56 60 62 66 68 72 74 76 77 78 90 92 94 95 96 97 98
r176 90 104 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=11.58 $Y=0.465
+ $X2=11.58 $Y2=0.36
r177 90 92 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.58 $Y=0.465
+ $X2=11.58 $Y2=0.72
r178 87 89 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=9.66 $Y=0.36
+ $X2=10.6 $Y2=0.36
r179 85 87 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=8.72 $Y=0.36
+ $X2=9.66 $Y2=0.36
r180 83 85 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=7.78 $Y=0.36
+ $X2=8.72 $Y2=0.36
r181 81 83 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=6.84 $Y=0.36
+ $X2=7.78 $Y2=0.36
r182 79 100 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.985 $Y=0.36
+ $X2=5.86 $Y2=0.36
r183 79 81 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=5.985 $Y=0.36
+ $X2=6.84 $Y2=0.36
r184 78 104 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=11.455 $Y=0.36
+ $X2=11.58 $Y2=0.36
r185 78 89 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=11.455 $Y=0.36
+ $X2=10.6 $Y2=0.36
r186 77 102 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.86 $Y=0.715
+ $X2=5.86 $Y2=0.8
r187 76 100 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.86 $Y=0.465
+ $X2=5.86 $Y2=0.36
r188 76 77 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=5.86 $Y=0.465
+ $X2=5.86 $Y2=0.715
r189 75 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0.8
+ $X2=4.96 $Y2=0.8
r190 74 102 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.735 $Y=0.8
+ $X2=5.86 $Y2=0.8
r191 74 75 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=0.8
+ $X2=5.125 $Y2=0.8
r192 70 98 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.715
+ $X2=4.96 $Y2=0.8
r193 70 72 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.96 $Y=0.715
+ $X2=4.96 $Y2=0.38
r194 69 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0.8
+ $X2=4.02 $Y2=0.8
r195 68 98 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0.8
+ $X2=4.96 $Y2=0.8
r196 68 69 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=0.8
+ $X2=4.185 $Y2=0.8
r197 64 97 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.715
+ $X2=4.02 $Y2=0.8
r198 64 66 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.02 $Y=0.715
+ $X2=4.02 $Y2=0.38
r199 63 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0.8
+ $X2=3.08 $Y2=0.8
r200 62 97 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0.8
+ $X2=4.02 $Y2=0.8
r201 62 63 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0.8
+ $X2=3.245 $Y2=0.8
r202 58 96 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.8
r203 58 60 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.08 $Y=0.715
+ $X2=3.08 $Y2=0.38
r204 57 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=0.8
+ $X2=2.14 $Y2=0.8
r205 56 96 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=3.08 $Y2=0.8
r206 56 57 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=0.8
+ $X2=2.305 $Y2=0.8
r207 52 95 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.8
r208 52 54 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=0.715
+ $X2=2.14 $Y2=0.38
r209 51 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=0.8
+ $X2=1.2 $Y2=0.8
r210 50 95 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=2.14 $Y2=0.8
r211 50 51 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.975 $Y=0.8
+ $X2=1.365 $Y2=0.8
r212 46 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.715 $X2=1.2
+ $Y2=0.8
r213 46 48 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=0.715
+ $X2=1.2 $Y2=0.38
r214 44 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=1.2 $Y2=0.8
r215 44 45 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=0.425 $Y2=0.8
r216 40 45 7.80856 $w=1.7e-07 $l=2.06165e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.425 $Y2=0.8
r217 40 42 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.257 $Y=0.715
+ $X2=0.257 $Y2=0.38
r218 13 104 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=11.405
+ $Y=0.235 $X2=11.54 $Y2=0.38
r219 13 92 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=11.405
+ $Y=0.235 $X2=11.54 $Y2=0.72
r220 12 89 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=10.465
+ $Y=0.235 $X2=10.6 $Y2=0.38
r221 11 87 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=9.475
+ $Y=0.235 $X2=9.66 $Y2=0.38
r222 10 85 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=8.585
+ $Y=0.235 $X2=8.72 $Y2=0.38
r223 9 83 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.645
+ $Y=0.235 $X2=7.78 $Y2=0.38
r224 8 81 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.38
r225 7 102 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.235 $X2=5.9 $Y2=0.72
r226 7 100 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.765
+ $Y=0.235 $X2=5.9 $Y2=0.38
r227 6 72 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.825
+ $Y=0.235 $X2=4.96 $Y2=0.38
r228 5 66 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.885
+ $Y=0.235 $X2=4.02 $Y2=0.38
r229 4 60 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.38
r230 3 54 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r231 2 48 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r232 1 42 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND2_12%VGND 1 2 3 4 5 6 21 23 27 29 33 35 39 41
+ 45 49 52 53 54 56 69 70 73 76 79 82 85
r147 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r148 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.37
+ $Y2=0
r149 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r150 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r151 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r152 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r153 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r154 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r155 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r156 69 70 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r157 67 70 1.70156 $w=4.8e-07 $l=5.98e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=11.73 $Y2=0
r158 66 69 390.139 $w=1.68e-07 $l=5.98e-06 $layer=LI1_cond $X=5.75 $Y=0
+ $X2=11.73 $Y2=0
r159 66 67 1.32857 $w=1.7e-07 $l=1.19e-06 $layer=mcon $count=7 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r160 64 67 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r161 64 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=4.37
+ $Y2=0
r162 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r163 61 85 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=4.49
+ $Y2=0
r164 61 63 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=4.625 $Y=0 $X2=5.29
+ $Y2=0
r165 56 73 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.73
+ $Y2=0
r166 56 58 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=0
+ $X2=0.23 $Y2=0
r167 54 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r168 54 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r169 52 63 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.29
+ $Y2=0
r170 52 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.295 $Y=0 $X2=5.43
+ $Y2=0
r171 51 66 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=5.75 $Y2=0
r172 51 53 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.43
+ $Y2=0
r173 47 53 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0
r174 47 49 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.43 $Y=0.085
+ $X2=5.43 $Y2=0.38
r175 43 85 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0
r176 43 45 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.49 $Y=0.085
+ $X2=4.49 $Y2=0.38
r177 42 82 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.55
+ $Y2=0
r178 41 85 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.49
+ $Y2=0
r179 41 42 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0
+ $X2=3.685 $Y2=0
r180 37 82 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0
r181 37 39 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.55 $Y=0.085
+ $X2=3.55 $Y2=0.38
r182 36 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.745 $Y=0 $X2=2.61
+ $Y2=0
r183 35 82 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0 $X2=3.55
+ $Y2=0
r184 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0
+ $X2=2.745 $Y2=0
r185 31 79 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r186 31 33 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.38
r187 30 76 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=0 $X2=1.67
+ $Y2=0
r188 29 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.61
+ $Y2=0
r189 29 30 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.475 $Y=0
+ $X2=1.805 $Y2=0
r190 25 76 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r191 25 27 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.38
r192 24 73 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.865 $Y=0 $X2=0.73
+ $Y2=0
r193 23 76 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=0 $X2=1.67
+ $Y2=0
r194 23 24 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=0
+ $X2=0.865 $Y2=0
r195 19 73 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r196 19 21 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r197 6 49 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.38
r198 5 45 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.38
r199 4 39 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.38
r200 3 33 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.38
r201 2 27 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.38
r202 1 21 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

