* File: sky130_fd_sc_hdll__a22o_1.pxi.spice
* Created: Wed Sep  2 08:18:30 2020
* 
x_PM_SKY130_FD_SC_HDLL__A22O_1%B2 N_B2_c_50_n N_B2_M1003_g N_B2_c_51_n
+ N_B2_M1009_g B2 N_B2_c_52_n PM_SKY130_FD_SC_HDLL__A22O_1%B2
x_PM_SKY130_FD_SC_HDLL__A22O_1%B1 N_B1_c_73_n N_B1_M1002_g N_B1_c_74_n
+ N_B1_M1000_g B1 B1 B1 PM_SKY130_FD_SC_HDLL__A22O_1%B1
x_PM_SKY130_FD_SC_HDLL__A22O_1%A1 N_A1_c_106_n N_A1_M1008_g N_A1_c_107_n
+ N_A1_M1004_g A1 A1 N_A1_c_109_n N_A1_c_110_n PM_SKY130_FD_SC_HDLL__A22O_1%A1
x_PM_SKY130_FD_SC_HDLL__A22O_1%A2 N_A2_c_141_n N_A2_M1005_g N_A2_c_142_n
+ N_A2_M1001_g A2 PM_SKY130_FD_SC_HDLL__A22O_1%A2
x_PM_SKY130_FD_SC_HDLL__A22O_1%A_27_297# N_A_27_297#_M1002_d N_A_27_297#_M1004_s
+ N_A_27_297#_M1003_s N_A_27_297#_M1000_d N_A_27_297#_c_176_n
+ N_A_27_297#_M1007_g N_A_27_297#_c_177_n N_A_27_297#_M1006_g
+ N_A_27_297#_c_181_n N_A_27_297#_c_182_n N_A_27_297#_c_178_n
+ N_A_27_297#_c_214_n N_A_27_297#_c_215_n N_A_27_297#_c_218_n
+ N_A_27_297#_c_179_n N_A_27_297#_c_184_n N_A_27_297#_c_185_n
+ PM_SKY130_FD_SC_HDLL__A22O_1%A_27_297#
x_PM_SKY130_FD_SC_HDLL__A22O_1%A_117_297# N_A_117_297#_M1003_d
+ N_A_117_297#_M1008_d N_A_117_297#_c_263_n N_A_117_297#_c_267_n
+ N_A_117_297#_c_268_n PM_SKY130_FD_SC_HDLL__A22O_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A22O_1%VPWR N_VPWR_M1008_s N_VPWR_M1005_d N_VPWR_c_285_n
+ N_VPWR_c_286_n N_VPWR_c_287_n N_VPWR_c_288_n VPWR N_VPWR_c_289_n
+ N_VPWR_c_290_n N_VPWR_c_284_n N_VPWR_c_292_n PM_SKY130_FD_SC_HDLL__A22O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A22O_1%X N_X_M1006_d N_X_M1007_d N_X_c_328_n X X X
+ PM_SKY130_FD_SC_HDLL__A22O_1%X
x_PM_SKY130_FD_SC_HDLL__A22O_1%VGND N_VGND_M1009_s N_VGND_M1001_d N_VGND_c_344_n
+ N_VGND_c_345_n N_VGND_c_346_n N_VGND_c_347_n N_VGND_c_348_n VGND
+ N_VGND_c_349_n N_VGND_c_350_n PM_SKY130_FD_SC_HDLL__A22O_1%VGND
cc_1 VNB N_B2_c_50_n 0.0277636f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B2_c_51_n 0.0206423f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_B2_c_52_n 0.0160638f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_4 VNB N_B1_c_73_n 0.0194095f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B1_c_74_n 0.0244535f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B1 0.00302118f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_7 VNB B1 0.00726178f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A1_c_106_n 0.0247457f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_9 VNB N_A1_c_107_n 0.020234f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_10 VNB A1 0.00598053f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_A1_c_109_n 0.00320017f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A1_c_110_n 0.00452669f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.175
cc_13 VNB N_A2_c_141_n 0.0217306f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_A2_c_142_n 0.0160288f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_15 VNB A2 0.00585232f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_16 VNB N_A_27_297#_c_176_n 0.0254815f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_177_n 0.0198493f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_178_n 0.0125385f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_297#_c_179_n 0.00111447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VPWR_c_284_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_328_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_22 VNB X 0.0313676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_344_n 0.0128325f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_24 VNB N_VGND_c_345_n 0.0286001f $X=-0.19 $Y=-0.24 $X2=0.46 $Y2=1.16
cc_25 VNB N_VGND_c_346_n 0.00561478f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_347_n 0.0472927f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_348_n 0.00631318f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_349_n 0.0234912f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_350_n 0.204275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VPB N_B2_c_50_n 0.0329415f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_31 VPB N_B1_c_74_n 0.0320744f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_32 VPB N_A1_c_106_n 0.0319244f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB N_A2_c_141_n 0.0260877f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_34 VPB N_A_27_297#_c_176_n 0.0283389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_297#_c_181_n 0.0097796f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_27_297#_c_182_n 0.0124552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_297#_c_179_n 0.0016874f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_297#_c_184_n 0.00889261f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_297#_c_185_n 0.0199249f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_117_297#_c_263_n 0.00769094f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_41 VPB N_VPWR_c_285_n 0.00710338f $X=-0.19 $Y=1.305 $X2=0.46 $Y2=1.16
cc_42 VPB N_VPWR_c_286_n 0.00285927f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_VPWR_c_287_n 0.0168749f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_VPWR_c_288_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_289_n 0.0435631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_290_n 0.0230131f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_284_n 0.0489369f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_292_n 0.005552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB X 0.0457201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 N_B2_c_51_n N_B1_c_73_n 0.0305731f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_51 N_B2_c_50_n N_B1_c_74_n 0.0681641f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_B2_c_52_n N_B1_c_74_n 6.85412e-19 $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_53 N_B2_c_50_n B1 3.65043e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_54 N_B2_c_50_n B1 9.41434e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_55 N_B2_c_52_n B1 0.016379f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_56 N_B2_c_50_n N_A_27_297#_c_181_n 4.82237e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_B2_c_52_n N_A_27_297#_c_181_n 0.0176967f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_58 N_B2_c_50_n N_A_27_297#_c_182_n 0.0162887f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_59 N_B2_c_52_n N_A_27_297#_c_182_n 0.0131715f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_60 N_B2_c_51_n N_A_27_297#_c_178_n 6.82958e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_61 N_B2_c_50_n N_A_27_297#_c_184_n 0.00470744f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_B2_c_50_n N_A_117_297#_c_263_n 0.00314906f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B2_c_50_n N_VPWR_c_289_n 0.00652245f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 N_B2_c_50_n N_VPWR_c_284_n 0.012299f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_B2_c_50_n N_VGND_c_345_n 0.00293084f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_66 N_B2_c_51_n N_VGND_c_345_n 0.0270304f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_67 N_B2_c_52_n N_VGND_c_345_n 0.0308276f $X=0.46 $Y=1.16 $X2=0 $Y2=0
cc_68 N_B2_c_51_n N_VGND_c_350_n 8.26999e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_69 N_B1_c_74_n N_A1_c_106_n 0.00499895f $X=0.965 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_70 B1 N_A1_c_106_n 5.82999e-19 $X=1.115 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_71 N_B1_c_74_n A1 2.13396e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_72 B1 A1 0.0236616f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_73 N_B1_c_74_n N_A1_c_110_n 7.79245e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_74 B1 N_A1_c_110_n 6.65477e-19 $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_75 B1 N_A1_c_110_n 0.0146486f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_76 B1 N_A_27_297#_M1002_d 0.00648477f $X=1.115 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_77 N_B1_c_74_n N_A_27_297#_c_182_n 0.0130286f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_78 B1 N_A_27_297#_c_182_n 0.0257002f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_79 N_B1_c_73_n N_A_27_297#_c_178_n 0.00947416f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B1_c_74_n N_A_27_297#_c_178_n 2.40258e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 B1 N_A_27_297#_c_178_n 0.0132859f $X=1.115 $Y=0.765 $X2=0 $Y2=0
cc_82 B1 N_A_27_297#_c_178_n 0.00416148f $X=1.115 $Y=1.105 $X2=0 $Y2=0
cc_83 N_B1_c_74_n N_A_27_297#_c_184_n 0.00102139f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B1_c_74_n N_A_117_297#_c_263_n 0.0146945f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B1_c_74_n N_VPWR_c_285_n 0.00839193f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B1_c_74_n N_VPWR_c_289_n 0.00510113f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B1_c_74_n N_VPWR_c_284_n 0.00819924f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B1_c_73_n N_VGND_c_345_n 0.00415884f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_89 N_B1_c_73_n N_VGND_c_347_n 0.00365461f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_90 N_B1_c_73_n N_VGND_c_350_n 0.0067644f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A1_c_106_n N_A2_c_141_n 0.0246624f $X=1.955 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_92 N_A1_c_107_n N_A2_c_141_n 0.0192306f $X=1.98 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_93 N_A1_c_109_n N_A2_c_141_n 7.83772e-19 $X=1.92 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_94 N_A1_c_107_n N_A2_c_142_n 0.0255838f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A1_c_106_n A2 7.20005e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A1_c_107_n A2 8.14688e-19 $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_97 A1 A2 0.0030604f $X=1.575 $Y=0.765 $X2=0 $Y2=0
cc_98 N_A1_c_109_n A2 0.017696f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_99 A1 N_A_27_297#_M1004_s 0.00661906f $X=1.575 $Y=0.765 $X2=0 $Y2=0
cc_100 N_A1_c_106_n N_A_27_297#_c_182_n 0.0187885f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A1_c_109_n N_A_27_297#_c_182_n 0.0177633f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_102 N_A1_c_110_n N_A_27_297#_c_182_n 0.0159326f $X=1.635 $Y=1.065 $X2=0 $Y2=0
cc_103 N_A1_c_106_n N_A_27_297#_c_178_n 0.00203364f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A1_c_107_n N_A_27_297#_c_178_n 0.0156626f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_105 A1 N_A_27_297#_c_178_n 0.0142092f $X=1.575 $Y=0.765 $X2=0 $Y2=0
cc_106 N_A1_c_109_n N_A_27_297#_c_178_n 0.00783329f $X=1.92 $Y=1.16 $X2=0 $Y2=0
cc_107 N_A1_c_106_n N_A_117_297#_c_263_n 0.0144021f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A1_c_106_n N_VPWR_c_285_n 0.00927816f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A1_c_106_n N_VPWR_c_287_n 0.00424386f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A1_c_106_n N_VPWR_c_284_n 0.0049917f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A1_c_107_n N_VGND_c_347_n 0.00357877f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A1_c_107_n N_VGND_c_350_n 0.00690424f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_113 N_A2_c_141_n N_A_27_297#_c_176_n 0.0414907f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_114 A2 N_A_27_297#_c_176_n 0.00191096f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A2_c_142_n N_A_27_297#_c_177_n 0.0187481f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_116 N_A2_c_141_n N_A_27_297#_c_182_n 0.0217691f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_117 A2 N_A_27_297#_c_182_n 0.018459f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_118 N_A2_c_142_n N_A_27_297#_c_178_n 0.00247262f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_119 N_A2_c_142_n N_A_27_297#_c_214_n 0.0033083f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_120 N_A2_c_141_n N_A_27_297#_c_215_n 0.00277363f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A2_c_142_n N_A_27_297#_c_215_n 0.0124213f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_122 A2 N_A_27_297#_c_215_n 0.0191785f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_123 A2 N_A_27_297#_c_218_n 3.82704e-19 $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_124 N_A2_c_141_n N_A_27_297#_c_179_n 0.00355601f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A2_c_142_n N_A_27_297#_c_179_n 0.00363279f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_126 A2 N_A_27_297#_c_179_n 0.0179114f $X=2.395 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A2_c_141_n N_A_117_297#_c_267_n 0.00268226f $X=2.475 $Y=1.41 $X2=0
+ $Y2=0
cc_128 N_A2_c_141_n N_A_117_297#_c_268_n 0.00399182f $X=2.475 $Y=1.41 $X2=0
+ $Y2=0
cc_129 N_A2_c_141_n N_VPWR_c_285_n 9.52784e-19 $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A2_c_141_n N_VPWR_c_286_n 0.00315802f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A2_c_141_n N_VPWR_c_287_n 0.00688798f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A2_c_141_n N_VPWR_c_284_n 0.0123702f $X=2.475 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A2_c_142_n N_VGND_c_346_n 0.00325341f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_134 N_A2_c_142_n N_VGND_c_347_n 0.00422112f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_135 N_A2_c_142_n N_VGND_c_350_n 0.00605887f $X=2.5 $Y=0.96 $X2=0 $Y2=0
cc_136 N_A_27_297#_c_182_n N_A_117_297#_M1003_d 0.00870057f $X=2.865 $Y=1.605
+ $X2=-0.19 $Y2=-0.24
cc_137 N_A_27_297#_c_182_n N_A_117_297#_M1008_d 0.00979537f $X=2.865 $Y=1.605
+ $X2=0 $Y2=0
cc_138 N_A_27_297#_M1000_d N_A_117_297#_c_263_n 0.00698008f $X=1.055 $Y=1.485
+ $X2=0 $Y2=0
cc_139 N_A_27_297#_c_182_n N_A_117_297#_c_263_n 0.0925814f $X=2.865 $Y=1.605
+ $X2=0 $Y2=0
cc_140 N_A_27_297#_c_185_n N_A_117_297#_c_263_n 0.0131144f $X=0.257 $Y=2.245
+ $X2=0 $Y2=0
cc_141 N_A_27_297#_c_182_n N_A_117_297#_c_267_n 0.0192007f $X=2.865 $Y=1.605
+ $X2=0 $Y2=0
cc_142 N_A_27_297#_c_182_n N_VPWR_M1008_s 0.00581464f $X=2.865 $Y=1.605
+ $X2=-0.19 $Y2=-0.24
cc_143 N_A_27_297#_c_182_n N_VPWR_M1005_d 0.0103454f $X=2.865 $Y=1.605 $X2=0
+ $Y2=0
cc_144 N_A_27_297#_c_176_n N_VPWR_c_286_n 0.0142059f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_27_297#_c_182_n N_VPWR_c_286_n 0.0160369f $X=2.865 $Y=1.605 $X2=0
+ $Y2=0
cc_146 N_A_27_297#_c_184_n N_VPWR_c_289_n 0.0213091f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_147 N_A_27_297#_c_176_n N_VPWR_c_290_n 0.00622633f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_27_297#_M1003_s N_VPWR_c_284_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_149 N_A_27_297#_M1000_d N_VPWR_c_284_n 0.00316822f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_A_27_297#_c_176_n N_VPWR_c_284_n 0.0115709f $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_27_297#_c_184_n N_VPWR_c_284_n 0.0125861f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_152 N_A_27_297#_c_177_n N_X_c_328_n 0.00890133f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_27_297#_c_176_n X 0.0245409f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_154 N_A_27_297#_c_177_n X 0.0162093f $X=3.01 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_27_297#_c_182_n X 0.0103522f $X=2.865 $Y=1.605 $X2=0 $Y2=0
cc_156 N_A_27_297#_c_215_n X 0.00799934f $X=2.865 $Y=0.7 $X2=0 $Y2=0
cc_157 N_A_27_297#_c_179_n X 0.0307752f $X=2.95 $Y=1.16 $X2=0 $Y2=0
cc_158 N_A_27_297#_c_215_n N_VGND_M1001_d 0.0100685f $X=2.865 $Y=0.7 $X2=0 $Y2=0
cc_159 N_A_27_297#_c_179_n N_VGND_M1001_d 0.00126198f $X=2.95 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_27_297#_c_178_n N_VGND_c_345_n 0.011643f $X=2.11 $Y=0.36 $X2=0 $Y2=0
cc_161 N_A_27_297#_c_176_n N_VGND_c_346_n 2.02589e-19 $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_27_297#_c_177_n N_VGND_c_346_n 0.00319032f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_163 N_A_27_297#_c_215_n N_VGND_c_346_n 0.0187192f $X=2.865 $Y=0.7 $X2=0 $Y2=0
cc_164 N_A_27_297#_c_178_n N_VGND_c_347_n 0.0861951f $X=2.11 $Y=0.36 $X2=0 $Y2=0
cc_165 N_A_27_297#_c_215_n N_VGND_c_347_n 0.00485617f $X=2.865 $Y=0.7 $X2=0
+ $Y2=0
cc_166 N_A_27_297#_c_177_n N_VGND_c_349_n 0.00476436f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_27_297#_c_215_n N_VGND_c_349_n 0.00207807f $X=2.865 $Y=0.7 $X2=0
+ $Y2=0
cc_168 N_A_27_297#_M1002_d N_VGND_c_350_n 0.00225742f $X=1.015 $Y=0.235 $X2=0
+ $Y2=0
cc_169 N_A_27_297#_M1004_s N_VGND_c_350_n 0.00275739f $X=1.565 $Y=0.235 $X2=0
+ $Y2=0
cc_170 N_A_27_297#_c_177_n N_VGND_c_350_n 0.00862093f $X=3.01 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_27_297#_c_178_n N_VGND_c_350_n 0.0514717f $X=2.11 $Y=0.36 $X2=0 $Y2=0
cc_172 N_A_27_297#_c_215_n N_VGND_c_350_n 0.0126247f $X=2.865 $Y=0.7 $X2=0 $Y2=0
cc_173 N_A_27_297#_c_178_n A_411_47# 0.00445489f $X=2.11 $Y=0.36 $X2=-0.19
+ $Y2=-0.24
cc_174 N_A_27_297#_c_214_n A_411_47# 0.00177177f $X=2.195 $Y=0.615 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_27_297#_c_215_n A_411_47# 0.00230977f $X=2.865 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_27_297#_c_218_n A_411_47# 0.00824921f $X=2.28 $Y=0.7 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_117_297#_c_263_n N_VPWR_M1008_s 0.00543138f $X=2.065 $Y=1.985
+ $X2=-0.19 $Y2=1.305
cc_178 N_A_117_297#_c_263_n N_VPWR_c_285_n 0.0227984f $X=2.065 $Y=1.985 $X2=0
+ $Y2=0
cc_179 N_A_117_297#_c_263_n N_VPWR_c_287_n 0.00265869f $X=2.065 $Y=1.985 $X2=0
+ $Y2=0
cc_180 N_A_117_297#_c_268_n N_VPWR_c_287_n 0.0195833f $X=2.23 $Y=2.36 $X2=0
+ $Y2=0
cc_181 N_A_117_297#_c_263_n N_VPWR_c_289_n 0.0158139f $X=2.065 $Y=1.985 $X2=0
+ $Y2=0
cc_182 N_A_117_297#_M1003_d N_VPWR_c_284_n 0.00338665f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_183 N_A_117_297#_M1008_d N_VPWR_c_284_n 0.00277539f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_184 N_A_117_297#_c_263_n N_VPWR_c_284_n 0.0324675f $X=2.065 $Y=1.985 $X2=0
+ $Y2=0
cc_185 N_A_117_297#_c_268_n N_VPWR_c_284_n 0.0124664f $X=2.23 $Y=2.36 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_284_n N_X_M1007_d 0.0103088f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_c_286_n X 0.0226961f $X=2.75 $Y=2.02 $X2=0 $Y2=0
cc_188 N_VPWR_c_290_n X 0.0182101f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_189 N_VPWR_c_284_n X 0.00993603f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_190 N_X_c_328_n N_VGND_c_349_n 0.0173041f $X=3.45 $Y=0.42 $X2=0 $Y2=0
cc_191 N_X_M1006_d N_VGND_c_350_n 0.00984512f $X=3.085 $Y=0.235 $X2=0 $Y2=0
cc_192 N_X_c_328_n N_VGND_c_350_n 0.00982816f $X=3.45 $Y=0.42 $X2=0 $Y2=0
cc_193 N_VGND_c_350_n A_119_47# 0.0114986f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_194 N_VGND_c_350_n A_411_47# 0.00345858f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
