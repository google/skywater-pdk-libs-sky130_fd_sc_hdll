* File: sky130_fd_sc_hdll__o2bb2a_4.pex.spice
* Created: Thu Aug 27 19:21:56 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%B1 1 3 4 6 7 9 10 12 13 16 21 25
c76 10 0 8.50955e-20 $X=1.93 $Y=0.995
r77 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r78 21 31 7.53086 $w=5.38e-07 $l=3.4e-07 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.53
r79 21 25 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=0.355 $Y=1.19
+ $X2=0.355 $Y2=1.16
r80 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.905 $Y=1.16
+ $X2=1.905 $Y2=1.53
r81 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r82 14 31 7.6426 $w=1.7e-07 $l=2.7e-07 $layer=LI1_cond $X=0.625 $Y=1.53
+ $X2=0.355 $Y2=1.53
r83 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=1.905 $Y2=1.53
r84 13 14 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.715 $Y=1.53
+ $X2=0.625 $Y2=1.53
r85 10 17 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.905 $Y2=1.16
r86 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.93 $Y=0.995
+ $X2=1.93 $Y2=0.56
r87 7 17 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.16
r88 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r89 4 24 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r90 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r91 1 24 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r92 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%B2 1 3 4 6 7 9 10 12 13 20
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r48 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=1.2 $Y=1.202
+ $X2=1.435 $Y2=1.202
r49 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=1.2 $Y2=1.202
r50 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.202
+ $X2=0.965 $Y2=1.202
r51 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2
+ $Y=1.16 $X2=1.2 $Y2=1.16
r52 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r53 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r54 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r55 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r56 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r57 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r58 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=0.94 $Y2=1.202
r59 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_455_21# 1 2 3 10 12 13 15 16 18 19 21
+ 22 28 30 32 33 34 35 39 40 46 47 50 54
c121 54 0 1.82401e-19 $X=2.845 $Y=1.202
c122 50 0 1.45256e-19 $X=5.01 $Y=1.96
c123 40 0 1.35552e-19 $X=4.07 $Y=1.875
c124 10 0 1.56657e-19 $X=2.35 $Y=0.995
c125 2 0 1.6626e-19 $X=3.925 $Y=1.485
r126 53 54 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r127 52 53 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.82 $Y2=1.202
r128 51 52 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.202
+ $X2=2.375 $Y2=1.202
r129 46 47 10.6316 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=4.54 $Y=0.775
+ $X2=4.325 $Y2=0.775
r130 40 43 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=1.875
+ $X2=4.07 $Y2=1.96
r131 36 40 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.195 $Y=1.875
+ $X2=4.07 $Y2=1.875
r132 35 50 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=4.885 $Y=1.875
+ $X2=5.01 $Y2=1.875
r133 35 36 42.5152 $w=1.78e-07 $l=6.9e-07 $layer=LI1_cond $X=4.885 $Y=1.875
+ $X2=4.195 $Y2=1.875
r134 33 40 2.6621 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=3.945 $Y=1.875
+ $X2=4.07 $Y2=1.875
r135 33 34 30.8081 $w=1.78e-07 $l=5e-07 $layer=LI1_cond $X=3.945 $Y=1.875
+ $X2=3.445 $Y2=1.875
r136 32 47 54.2222 $w=1.78e-07 $l=8.8e-07 $layer=LI1_cond $X=3.445 $Y=0.815
+ $X2=4.325 $Y2=0.815
r137 30 34 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.35 $Y=1.785
+ $X2=3.445 $Y2=1.875
r138 29 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=1.245
+ $X2=3.35 $Y2=1.16
r139 29 30 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=3.35 $Y=1.245
+ $X2=3.35 $Y2=1.785
r140 28 39 4.70473 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.35 $Y=1.075
+ $X2=3.35 $Y2=1.16
r141 27 32 6.82297 $w=1.8e-07 $l=1.32571e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.445 $Y2=0.815
r142 27 28 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=3.35 $Y=0.905
+ $X2=3.35 $Y2=1.075
r143 25 54 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=3.08 $Y=1.202
+ $X2=2.845 $Y2=1.202
r144 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.08
+ $Y=1.16 $X2=3.08 $Y2=1.16
r145 22 39 1.74598 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.255 $Y=1.16
+ $X2=3.35 $Y2=1.16
r146 22 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=3.255 $Y=1.16
+ $X2=3.08 $Y2=1.16
r147 19 54 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r148 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r149 16 53 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r150 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r151 13 52 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r152 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r153 10 51 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.202
r154 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=0.56
r155 3 50 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=1.96
r156 2 43 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=1.96
r157 1 46 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A1_N 1 3 4 6 7 9 10 12 13 16 21
c84 16 0 3.48661e-19 $X=3.78 $Y=1.16
c85 10 0 1.86002e-19 $X=5.27 $Y=0.995
c86 7 0 4.72997e-19 $X=5.245 $Y=1.41
c87 1 0 1.60193e-19 $X=3.835 $Y=1.41
r88 21 30 10.4001 $w=4.08e-07 $l=3.7e-07 $layer=LI1_cond $X=5.26 $Y=1.16
+ $X2=5.26 $Y2=1.53
r89 21 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.22
+ $Y=1.16 $X2=5.22 $Y2=1.16
r90 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=3.805 $Y=1.16
+ $X2=3.805 $Y2=1.53
r91 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.78
+ $Y=1.16 $X2=3.78 $Y2=1.16
r92 14 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.995 $Y=1.53
+ $X2=3.805 $Y2=1.53
r93 13 30 5.92876 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=5.055 $Y=1.53
+ $X2=5.26 $Y2=1.53
r94 13 14 69.1551 $w=1.68e-07 $l=1.06e-06 $layer=LI1_cond $X=5.055 $Y=1.53
+ $X2=3.995 $Y2=1.53
r95 10 25 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.245 $Y2=1.16
r96 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.27 $Y=0.995
+ $X2=5.27 $Y2=0.56
r97 7 25 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.16
r98 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.245 $Y=1.41
+ $X2=5.245 $Y2=1.985
r99 4 17 38.7084 $w=3.43e-07 $l=1.90526e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.805 $Y2=1.16
r100 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r101 1 17 45.964 $w=3.43e-07 $l=2.64575e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.805 $Y2=1.16
r102 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A2_N 1 3 4 6 7 9 10 12 13 19 20 25
c46 10 0 8.25269e-20 $X=4.8 $Y=0.995
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.202
+ $X2=4.8 $Y2=1.202
r48 19 25 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=4.545 $Y=1.175
+ $X2=4.44 $Y2=1.175
r49 18 20 29.1737 $w=3.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.545 $Y=1.202
+ $X2=4.775 $Y2=1.202
r50 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.545
+ $Y=1.16 $X2=4.545 $Y2=1.16
r51 16 18 30.4421 $w=3.8e-07 $l=2.4e-07 $layer=POLY_cond $X=4.305 $Y=1.202
+ $X2=4.545 $Y2=1.202
r52 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.305 $Y2=1.202
r53 13 25 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=4.33 $Y=1.175 $X2=4.44
+ $Y2=1.175
r54 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.8 $Y=0.995
+ $X2=4.8 $Y2=1.202
r55 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.8 $Y=0.995 $X2=4.8
+ $Y2=0.56
r56 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.202
r57 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r58 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.202
r59 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r60 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r61 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995 $X2=4.28
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_211_297# 1 2 3 10 12 13 15 16 18 19 21
+ 22 24 25 27 28 30 31 33 34 37 40 45 48 54 64 66 67 68 78 86
c154 68 0 2.4641e-20 $X=5.665 $Y=1.52
c155 66 0 1.53217e-19 $X=5.81 $Y=1.53
c156 54 0 8.50955e-20 $X=2.61 $Y=0.73
c157 40 0 1.74525e-19 $X=6.005 $Y=1.16
c158 28 0 1.46608e-19 $X=7.125 $Y=1.41
r159 84 86 2.06391 $w=5.32e-07 $l=9e-08 $layer=LI1_cond $X=2.565 $Y=1.87
+ $X2=2.565 $Y2=1.96
r160 78 79 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=7.125 $Y=1.202
+ $X2=7.15 $Y2=1.202
r161 75 76 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.63 $Y=1.202
+ $X2=6.655 $Y2=1.202
r162 74 75 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=6.185 $Y=1.202
+ $X2=6.63 $Y2=1.202
r163 73 74 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=6.16 $Y=1.202
+ $X2=6.185 $Y2=1.202
r164 70 71 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=5.69 $Y=1.202
+ $X2=5.715 $Y2=1.202
r165 66 68 0.113931 $w=2.5e-07 $l=1.45e-07 $layer=MET1_cond $X=5.81 $Y=1.52
+ $X2=5.665 $Y2=1.52
r166 66 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.81 $Y=1.53
+ $X2=5.81 $Y2=1.53
r167 64 68 3.3292 $w=1.4e-07 $l=2.69e-06 $layer=MET1_cond $X=2.975 $Y=1.53
+ $X2=5.665 $Y2=1.53
r168 62 84 8.02632 $w=5.32e-07 $l=3.5e-07 $layer=LI1_cond $X=2.565 $Y=1.52
+ $X2=2.565 $Y2=1.87
r169 61 64 0.143445 $w=2.5e-07 $l=1.95e-07 $layer=MET1_cond $X=2.78 $Y=1.51
+ $X2=2.975 $Y2=1.51
r170 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.78 $Y=1.52
+ $X2=2.78 $Y2=1.52
r171 57 67 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=5.835 $Y=1.245
+ $X2=5.835 $Y2=1.53
r172 54 56 3.12082 $w=3.78e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.73
+ $X2=2.585 $Y2=0.815
r173 48 51 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=1.2 $Y=1.87 $X2=1.2
+ $Y2=1.96
r174 46 78 34.336 $w=3.72e-07 $l=2.65e-07 $layer=POLY_cond $X=6.86 $Y=1.202
+ $X2=7.125 $Y2=1.202
r175 46 76 26.5618 $w=3.72e-07 $l=2.05e-07 $layer=POLY_cond $X=6.86 $Y=1.202
+ $X2=6.655 $Y2=1.202
r176 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.86
+ $Y=1.16 $X2=6.86 $Y2=1.16
r177 43 73 10.3656 $w=3.72e-07 $l=8e-08 $layer=POLY_cond $X=6.08 $Y=1.202
+ $X2=6.16 $Y2=1.202
r178 43 71 47.293 $w=3.72e-07 $l=3.65e-07 $layer=POLY_cond $X=6.08 $Y=1.202
+ $X2=5.715 $Y2=1.202
r179 42 45 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=6.08 $Y=1.16
+ $X2=6.86 $Y2=1.16
r180 42 43 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.08
+ $Y=1.16 $X2=6.08 $Y2=1.16
r181 40 57 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=6.005 $Y=1.16
+ $X2=5.835 $Y2=1.245
r182 40 42 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.005 $Y=1.16
+ $X2=6.08 $Y2=1.16
r183 37 62 12.5061 $w=5.32e-07 $l=4.5489e-07 $layer=LI1_cond $X=2.545 $Y=1.075
+ $X2=2.565 $Y2=1.52
r184 37 56 9.98784 $w=2.98e-07 $l=2.6e-07 $layer=LI1_cond $X=2.545 $Y=1.075
+ $X2=2.545 $Y2=0.815
r185 35 48 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.325 $Y=1.87
+ $X2=1.2 $Y2=1.87
r186 34 84 7.54793 $w=1.7e-07 $l=3e-07 $layer=LI1_cond $X=2.265 $Y=1.87
+ $X2=2.565 $Y2=1.87
r187 34 35 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=2.265 $Y=1.87
+ $X2=1.325 $Y2=1.87
r188 31 79 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=1.202
r189 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.15 $Y=0.995
+ $X2=7.15 $Y2=0.56
r190 28 78 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.202
r191 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.125 $Y=1.41
+ $X2=7.125 $Y2=1.985
r192 25 76 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.202
r193 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.655 $Y2=1.985
r194 22 75 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=1.202
r195 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.63 $Y=0.995
+ $X2=6.63 $Y2=0.56
r196 19 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.202
r197 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.185 $Y=1.41
+ $X2=6.185 $Y2=1.985
r198 16 73 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=1.202
r199 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.16 $Y=0.995
+ $X2=6.16 $Y2=0.56
r200 13 71 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.202
r201 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.715 $Y=1.41
+ $X2=5.715 $Y2=1.985
r202 10 70 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=1.202
r203 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.69 $Y=0.995
+ $X2=5.69 $Y2=0.56
r204 3 86 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.96
r205 3 62 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r206 2 51 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r207 1 54 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44
+ 47 48 50 51 53 54 56 57 58 60 84 85 91 96 99
r122 98 99 9.89763 $w=6.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.6 $Y=2.47
+ $X2=3.725 $Y2=2.47
r123 94 98 2.67779 $w=6.68e-07 $l=1.5e-07 $layer=LI1_cond $X=3.45 $Y=2.47
+ $X2=3.6 $Y2=2.47
r124 94 96 15.7888 $w=6.68e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=2.47
+ $X2=2.995 $Y2=2.47
r125 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r126 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 84 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r128 82 85 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r129 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r130 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r131 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r132 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r133 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r134 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r135 73 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.45 $Y2=2.72
r136 72 99 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=3.725 $Y2=2.72
r137 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r138 69 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r139 69 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r140 68 96 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.995 $Y2=2.72
r141 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r142 66 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.265 $Y=2.72
+ $X2=2.14 $Y2=2.72
r143 66 68 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=2.265 $Y=2.72
+ $X2=2.99 $Y2=2.72
r144 64 92 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 61 88 3.63617 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r147 61 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r148 60 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.14 $Y2=2.72
r149 60 63 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=0.69 $Y2=2.72
r150 58 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r151 58 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r152 56 81 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.13 $Y2=2.72
r153 56 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.235 $Y=2.72
+ $X2=7.36 $Y2=2.72
r154 55 84 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.59 $Y2=2.72
r155 55 57 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.485 $Y=2.72
+ $X2=7.36 $Y2=2.72
r156 53 78 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.21 $Y2=2.72
r157 53 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.295 $Y=2.72
+ $X2=6.42 $Y2=2.72
r158 52 81 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=7.13 $Y2=2.72
r159 52 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.545 $Y=2.72
+ $X2=6.42 $Y2=2.72
r160 50 75 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.29 $Y2=2.72
r161 50 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.355 $Y=2.72
+ $X2=5.48 $Y2=2.72
r162 49 78 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=6.21 $Y2=2.72
r163 49 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.605 $Y=2.72
+ $X2=5.48 $Y2=2.72
r164 47 72 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.37 $Y2=2.72
r165 47 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.415 $Y=2.72
+ $X2=4.54 $Y2=2.72
r166 46 75 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=4.665 $Y=2.72
+ $X2=5.29 $Y2=2.72
r167 46 48 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.665 $Y=2.72
+ $X2=4.54 $Y2=2.72
r168 42 57 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=2.72
r169 42 44 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=7.36 $Y=2.635
+ $X2=7.36 $Y2=1.99
r170 38 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.72
r171 38 40 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=2.635
+ $X2=6.42 $Y2=2.33
r172 34 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=2.72
r173 34 36 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=5.48 $Y=2.635
+ $X2=5.48 $Y2=1.96
r174 30 48 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.72
r175 30 32 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=4.54 $Y=2.635
+ $X2=4.54 $Y2=2.3
r176 26 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r177 26 28 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.3
r178 22 88 3.25784 $w=2.05e-07 $l=1.14782e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.172 $Y2=2.72
r179 22 24 36.5188 $w=2.03e-07 $l=6.75e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=1.96
r180 7 44 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=7.215
+ $Y=1.485 $X2=7.36 $Y2=1.99
r181 6 40 600 $w=1.7e-07 $l=9.14631e-07 $layer=licon1_PDIFF $count=1 $X=6.275
+ $Y=1.485 $X2=6.42 $Y2=2.33
r182 5 36 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.335
+ $Y=1.485 $X2=5.48 $Y2=1.96
r183 4 32 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.3
r184 3 98 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.6 $Y2=2.3
r185 2 28 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.3
r186 1 24 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_117_297# 1 2 9 11 12 14
r19 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=1.67 $Y=2.3 $X2=1.67
+ $Y2=2.38
r20 11 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.545 $Y=2.38
+ $X2=1.67 $Y2=2.38
r21 11 12 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.545 $Y=2.38
+ $X2=0.855 $Y2=2.38
r22 7 12 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=0.73 $Y=2.295
+ $X2=0.855 $Y2=2.38
r23 7 9 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=0.73 $Y=2.295
+ $X2=0.73 $Y2=1.96
r24 2 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.3
r25 1 9 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%X 1 2 3 4 15 19 21 22 23 24 27 31 33 35
+ 36 43 44 48
c79 43 0 1.46608e-19 $X=7.405 $Y=1.105
c80 24 0 9.79736e-20 $X=6.115 $Y=0.815
r81 44 48 3.06325 $w=3.05e-07 $l=1.2e-07 $layer=LI1_cond $X=7.557 $Y=1.535
+ $X2=7.557 $Y2=1.415
r82 43 48 8.50163 $w=3.03e-07 $l=2.25e-07 $layer=LI1_cond $X=7.557 $Y=1.19
+ $X2=7.557 $Y2=1.415
r83 42 43 10.7687 $w=3.03e-07 $l=2.85e-07 $layer=LI1_cond $X=7.557 $Y=0.905
+ $X2=7.557 $Y2=1.19
r84 40 41 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=6.89 $Y=1.62
+ $X2=6.89 $Y2=1.87
r85 37 44 11.9744 $w=4.08e-07 $l=3.9e-07 $layer=LI1_cond $X=7.015 $Y=1.535
+ $X2=7.405 $Y2=1.535
r86 36 40 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.535
+ $X2=6.89 $Y2=1.62
r87 36 37 0.964185 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=6.89 $Y=1.535
+ $X2=7.015 $Y2=1.535
r88 34 35 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.055 $Y=0.815
+ $X2=6.865 $Y2=0.815
r89 33 42 7.42255 $w=1.8e-07 $l=1.91792e-07 $layer=LI1_cond $X=7.405 $Y=0.815
+ $X2=7.557 $Y2=0.905
r90 33 34 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=7.405 $Y=0.815
+ $X2=7.055 $Y2=0.815
r91 29 41 3.91831 $w=2.48e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.955
+ $X2=6.89 $Y2=1.87
r92 29 31 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.89 $Y=1.955
+ $X2=6.89 $Y2=1.96
r93 25 35 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.815
r94 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.865 $Y=0.725
+ $X2=6.865 $Y2=0.39
r95 23 35 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.865 $Y2=0.815
r96 23 24 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.675 $Y=0.815
+ $X2=6.115 $Y2=0.815
r97 21 41 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.765 $Y=1.87
+ $X2=6.89 $Y2=1.87
r98 21 22 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.765 $Y=1.87
+ $X2=6.075 $Y2=1.87
r99 17 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.95 $Y=1.955
+ $X2=6.075 $Y2=1.87
r100 17 19 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=5.95 $Y=1.955
+ $X2=5.95 $Y2=1.96
r101 13 24 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=6.115 $Y2=0.815
r102 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.925 $Y=0.725
+ $X2=5.925 $Y2=0.39
r103 4 40 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.62
r104 4 31 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.745
+ $Y=1.485 $X2=6.89 $Y2=1.96
r105 3 19 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.805
+ $Y=1.485 $X2=5.95 $Y2=1.96
r106 2 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.705
+ $Y=0.235 $X2=6.89 $Y2=0.39
r107 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.765
+ $Y=0.235 $X2=5.95 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_27_47# 1 2 3 4 15 17 18 21 23 25 28 31
+ 33
c61 23 0 1.56657e-19 $X=1.925 $Y=0.82
r62 29 35 4.05488 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=2.075 $Y2=0.365
r63 29 31 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=2.225 $Y=0.365
+ $X2=3.08 $Y2=0.365
r64 26 28 0.192074 $w=2.98e-07 $l=5e-09 $layer=LI1_cond $X=2.075 $Y=0.735
+ $X2=2.075 $Y2=0.73
r65 25 35 2.97358 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=2.075 $Y=0.475
+ $X2=2.075 $Y2=0.365
r66 25 28 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=2.075 $Y=0.475
+ $X2=2.075 $Y2=0.73
r67 24 33 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=1.365 $Y=0.82
+ $X2=1.175 $Y2=0.815
r68 23 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=1.925 $Y=0.82
+ $X2=2.075 $Y2=0.735
r69 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.925 $Y=0.82
+ $X2=1.365 $Y2=0.82
r70 19 33 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.815
r71 19 21 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.175 $Y=0.725
+ $X2=1.175 $Y2=0.39
r72 17 33 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=1.175 $Y2=0.815
r73 17 18 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=0.985 $Y=0.815
+ $X2=0.425 $Y2=0.815
r74 13 18 7.61292 $w=1.8e-07 $l=2.05122e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.425 $Y2=0.815
r75 13 15 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.725
+ $X2=0.26 $Y2=0.39
r76 4 31 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.39
r77 3 35 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.39
r78 3 28 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.73
r79 2 21 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.39
r80 1 15 91 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%VGND 1 2 3 4 5 6 23 25 29 33 37 41 45 48
+ 49 51 52 54 55 57 58 59 81 82 85 88
r121 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r122 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r123 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r124 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r125 79 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r126 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r127 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r128 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r129 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r130 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r131 70 73 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=5.29 $Y2=0
r132 69 72 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=5.29
+ $Y2=0
r133 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r134 67 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r135 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r136 64 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.45 $Y2=0
r137 64 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r138 63 66 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r139 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r140 61 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=0 $X2=1.67
+ $Y2=0
r141 61 63 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=0
+ $X2=2.07 $Y2=0
r142 59 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r143 57 78 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.275 $Y=0
+ $X2=7.13 $Y2=0
r144 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.275 $Y=0 $X2=7.36
+ $Y2=0
r145 56 81 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=7.445 $Y=0
+ $X2=7.59 $Y2=0
r146 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0 $X2=7.36
+ $Y2=0
r147 54 75 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r148 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.335 $Y=0 $X2=6.42
+ $Y2=0
r149 53 78 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=6.505 $Y=0
+ $X2=7.13 $Y2=0
r150 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.505 $Y=0 $X2=6.42
+ $Y2=0
r151 51 72 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=0
+ $X2=5.29 $Y2=0
r152 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.395 $Y=0 $X2=5.48
+ $Y2=0
r153 50 75 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=5.565 $Y=0
+ $X2=6.21 $Y2=0
r154 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.565 $Y=0 $X2=5.48
+ $Y2=0
r155 48 66 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.45
+ $Y2=0
r156 48 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.515 $Y=0 $X2=3.6
+ $Y2=0
r157 47 69 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=3.685 $Y=0
+ $X2=3.91 $Y2=0
r158 47 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.685 $Y=0 $X2=3.6
+ $Y2=0
r159 43 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0
r160 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.36 $Y=0.085
+ $X2=7.36 $Y2=0.39
r161 39 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0
r162 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.42 $Y=0.085
+ $X2=6.42 $Y2=0.39
r163 35 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r164 35 37 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.39
r165 31 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.6 $Y=0.085 $X2=3.6
+ $Y2=0
r166 31 33 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.6 $Y=0.085
+ $X2=3.6 $Y2=0.39
r167 27 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0
r168 27 29 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.67 $Y=0.085
+ $X2=1.67 $Y2=0.39
r169 26 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r170 25 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.67
+ $Y2=0
r171 25 26 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.585 $Y=0
+ $X2=0.815 $Y2=0
r172 21 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r173 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.39
r174 6 45 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=7.225
+ $Y=0.235 $X2=7.36 $Y2=0.39
r175 5 41 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.235
+ $Y=0.235 $X2=6.42 $Y2=0.39
r176 4 37 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=5.345
+ $Y=0.235 $X2=5.48 $Y2=0.39
r177 3 33 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=3.475
+ $Y=0.235 $X2=3.6 $Y2=0.39
r178 2 29 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.39
r179 1 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2A_4%A_787_47# 1 2 7 11 13
c22 13 0 1.70555e-19 $X=5.01 $Y=0.73
r23 11 16 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.05 $Y=0.475
+ $X2=5.05 $Y2=0.39
r24 11 13 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=5.05 $Y=0.475
+ $X2=5.05 $Y2=0.73
r25 7 16 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.925 $Y=0.39
+ $X2=5.05 $Y2=0.39
r26 7 9 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=4.925 $Y=0.39
+ $X2=4.07 $Y2=0.39
r27 2 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.39
r28 2 13 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.73
r29 1 9 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.39
.ends

