* File: sky130_fd_sc_hdll__nor2_2.pxi.spice
* Created: Wed Sep  2 08:39:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2_2%A N_A_c_45_n N_A_M1003_g N_A_c_49_n N_A_M1000_g
+ N_A_c_50_n N_A_M1005_g N_A_c_46_n N_A_M1007_g A A N_A_c_48_n
+ PM_SKY130_FD_SC_HDLL__NOR2_2%A
x_PM_SKY130_FD_SC_HDLL__NOR2_2%B N_B_c_81_n N_B_M1004_g N_B_c_85_n N_B_M1001_g
+ N_B_c_86_n N_B_M1002_g N_B_c_82_n N_B_M1006_g B B N_B_c_84_n
+ PM_SKY130_FD_SC_HDLL__NOR2_2%B
x_PM_SKY130_FD_SC_HDLL__NOR2_2%A_27_297# N_A_27_297#_M1000_s N_A_27_297#_M1005_s
+ N_A_27_297#_M1002_d N_A_27_297#_c_129_n N_A_27_297#_c_130_n
+ N_A_27_297#_c_131_n N_A_27_297#_c_132_n N_A_27_297#_c_148_p
+ N_A_27_297#_c_133_n N_A_27_297#_c_134_n PM_SKY130_FD_SC_HDLL__NOR2_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR2_2%VPWR N_VPWR_M1000_d N_VPWR_c_169_n VPWR
+ N_VPWR_c_170_n N_VPWR_c_171_n N_VPWR_c_168_n N_VPWR_c_173_n
+ PM_SKY130_FD_SC_HDLL__NOR2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2_2%Y N_Y_M1003_d N_Y_M1004_s N_Y_M1001_s N_Y_c_207_n
+ N_Y_c_199_n N_Y_c_200_n N_Y_c_212_n N_Y_c_201_n N_Y_c_204_n N_Y_c_202_n
+ N_Y_c_203_n N_Y_c_206_n Y PM_SKY130_FD_SC_HDLL__NOR2_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR2_2%VGND N_VGND_M1003_s N_VGND_M1007_s N_VGND_M1006_d
+ N_VGND_c_260_n N_VGND_c_261_n N_VGND_c_262_n N_VGND_c_263_n N_VGND_c_264_n
+ N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n VGND N_VGND_c_268_n
+ N_VGND_c_269_n PM_SKY130_FD_SC_HDLL__NOR2_2%VGND
cc_1 VNB N_A_c_45_n 0.0222857f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_46_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB A 0.0164709f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.11
cc_4 VNB N_A_c_48_n 0.0430106f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_B_c_81_n 0.0169297f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_82_n 0.0200775f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB B 0.00630293f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.11
cc_8 VNB N_B_c_84_n 0.038927f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_9 VNB N_VPWR_c_168_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_10 VNB N_Y_c_199_n 0.00277197f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.11
cc_11 VNB N_Y_c_200_n 0.00296223f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_Y_c_201_n 0.00198035f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_13 VNB N_Y_c_202_n 0.0194803f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_203_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_260_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_16 VNB N_VGND_c_261_n 0.0334598f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.56
cc_17 VNB N_VGND_c_262_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.11
cc_18 VNB N_VGND_c_263_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_19 VNB N_VGND_c_264_n 0.0216754f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_20 VNB N_VGND_c_265_n 0.0110534f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=1.175
cc_21 VNB N_VGND_c_266_n 0.0211387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_267_n 0.00651182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_268_n 0.168353f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_269_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VPB N_A_c_49_n 0.0198936f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_26 VPB N_A_c_50_n 0.015934f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_27 VPB N_A_c_48_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_28 VPB N_B_c_85_n 0.0162445f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_29 VPB N_B_c_86_n 0.0191677f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_30 VPB N_B_c_84_n 0.0201102f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_31 VPB N_A_27_297#_c_129_n 0.0116385f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_32 VPB N_A_27_297#_c_130_n 0.0307403f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_33 VPB N_A_27_297#_c_131_n 0.00289118f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.11
cc_34 VPB N_A_27_297#_c_132_n 0.00184959f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_27_297#_c_133_n 0.00813676f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_36 VPB N_A_27_297#_c_134_n 0.0212257f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_37 VPB N_VPWR_c_169_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_38 VPB N_VPWR_c_170_n 0.015553f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_39 VPB N_VPWR_c_171_n 0.0478585f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_40 VPB N_VPWR_c_168_n 0.056403f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_41 VPB N_VPWR_c_173_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.175
cc_42 VPB N_Y_c_204_n 0.0105119f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_43 VPB N_Y_c_202_n 0.00680727f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_Y_c_206_n 0.00174301f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.175
cc_45 N_A_c_46_n N_B_c_81_n 0.024382f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_46 N_A_c_50_n N_B_c_85_n 0.00965769f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_47 A B 0.0167609f $X=0.6 $Y=1.11 $X2=0 $Y2=0
cc_48 N_A_c_48_n B 0.00766653f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_49 N_A_c_48_n N_B_c_84_n 0.024382f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_50 A N_A_27_297#_c_129_n 0.0225537f $X=0.6 $Y=1.11 $X2=0 $Y2=0
cc_51 N_A_c_49_n N_A_27_297#_c_131_n 0.0150902f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_c_50_n N_A_27_297#_c_131_n 0.0180389f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_53 A N_A_27_297#_c_131_n 0.0343628f $X=0.6 $Y=1.11 $X2=0 $Y2=0
cc_54 N_A_c_48_n N_A_27_297#_c_131_n 0.00813304f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_55 N_A_c_49_n N_VPWR_c_169_n 0.0171285f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A_c_50_n N_VPWR_c_169_n 0.0127351f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A_c_49_n N_VPWR_c_170_n 0.00427505f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_c_50_n N_VPWR_c_171_n 0.00622633f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_c_49_n N_VPWR_c_168_n 0.00825932f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_50_n N_VPWR_c_168_n 0.0104264f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_45_n N_Y_c_207_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_62 N_A_c_46_n N_Y_c_199_n 0.0117945f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_63 N_A_c_45_n N_Y_c_200_n 0.00269085f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_64 A N_Y_c_200_n 0.0262661f $X=0.6 $Y=1.11 $X2=0 $Y2=0
cc_65 N_A_c_48_n N_Y_c_200_n 0.00486271f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_66 N_A_c_46_n N_Y_c_212_n 5.32212e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_c_45_n N_VGND_c_261_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_68 A N_VGND_c_261_n 0.0233158f $X=0.6 $Y=1.11 $X2=0 $Y2=0
cc_69 N_A_c_45_n N_VGND_c_262_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_70 N_A_c_46_n N_VGND_c_262_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_c_46_n N_VGND_c_263_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_72 N_A_c_45_n N_VGND_c_268_n 0.0107167f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_73 N_A_c_46_n N_VGND_c_268_n 0.00615622f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_74 B N_A_27_297#_c_131_n 0.0073868f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_75 N_B_c_85_n N_A_27_297#_c_132_n 9.32325e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_76 B N_A_27_297#_c_132_n 0.0139423f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_77 N_B_c_85_n N_A_27_297#_c_133_n 0.0122476f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_78 N_B_c_86_n N_A_27_297#_c_133_n 0.0111074f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B_c_85_n N_VPWR_c_169_n 0.00100567f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_80 N_B_c_85_n N_VPWR_c_171_n 0.00429453f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B_c_86_n N_VPWR_c_171_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B_c_85_n N_VPWR_c_168_n 0.00609021f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_86_n N_VPWR_c_168_n 0.00734734f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B_c_81_n N_Y_c_199_n 0.00865686f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_85 B N_Y_c_199_n 0.0327042f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_86 N_B_c_81_n N_Y_c_212_n 0.00644736f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_87 N_B_c_82_n N_Y_c_201_n 0.0132459f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_88 B N_Y_c_201_n 0.00312628f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_89 N_B_c_86_n N_Y_c_204_n 0.0156341f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_90 B N_Y_c_204_n 0.00311514f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_91 N_B_c_84_n N_Y_c_204_n 3.62813e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_92 N_B_c_86_n N_Y_c_202_n 0.00134694f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_82_n N_Y_c_202_n 0.0190155f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_94 B N_Y_c_202_n 0.0145026f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_95 N_B_c_81_n N_Y_c_203_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_96 B N_Y_c_203_n 0.0307352f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_97 N_B_c_84_n N_Y_c_203_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_98 N_B_c_85_n N_Y_c_206_n 0.00464547f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_86_n N_Y_c_206_n 0.00115273f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_100 B N_Y_c_206_n 0.0305798f $X=1.52 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B_c_84_n N_Y_c_206_n 0.00764372f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_102 N_B_c_85_n Y 0.00738283f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B_c_86_n Y 0.0112727f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_81_n N_VGND_c_263_n 0.00268723f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B_c_82_n N_VGND_c_264_n 0.0115613f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_106 N_B_c_81_n N_VGND_c_266_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_107 N_B_c_82_n N_VGND_c_266_n 0.00439206f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B_c_81_n N_VGND_c_268_n 0.00598581f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B_c_82_n N_VGND_c_268_n 0.00769806f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_27_297#_c_131_n N_VPWR_M1000_d 0.00188315f $X=1.135 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_111 N_A_27_297#_c_130_n N_VPWR_c_169_n 0.0487409f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_112 N_A_27_297#_c_131_n N_VPWR_c_169_n 0.0212439f $X=1.135 $Y=1.56 $X2=0
+ $Y2=0
cc_113 N_A_27_297#_c_148_p N_VPWR_c_169_n 0.0397472f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_114 N_A_27_297#_c_130_n N_VPWR_c_170_n 0.019258f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_115 N_A_27_297#_c_148_p N_VPWR_c_171_n 0.0119545f $X=1.22 $Y=2.295 $X2=0
+ $Y2=0
cc_116 N_A_27_297#_c_133_n N_VPWR_c_171_n 0.0626043f $X=2.075 $Y=2.38 $X2=0
+ $Y2=0
cc_117 N_A_27_297#_M1000_s N_VPWR_c_168_n 0.00442207f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_118 N_A_27_297#_M1005_s N_VPWR_c_168_n 0.00436089f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_119 N_A_27_297#_M1002_d N_VPWR_c_168_n 0.00217523f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_120 N_A_27_297#_c_130_n N_VPWR_c_168_n 0.0105137f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_121 N_A_27_297#_c_148_p N_VPWR_c_168_n 0.006547f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_122 N_A_27_297#_c_133_n N_VPWR_c_168_n 0.0384086f $X=2.075 $Y=2.38 $X2=0
+ $Y2=0
cc_123 N_A_27_297#_c_133_n N_Y_M1001_s 0.00352392f $X=2.075 $Y=2.38 $X2=0 $Y2=0
cc_124 N_A_27_297#_c_131_n N_Y_c_199_n 0.00309388f $X=1.135 $Y=1.56 $X2=0 $Y2=0
cc_125 N_A_27_297#_c_131_n N_Y_c_200_n 0.00199016f $X=1.135 $Y=1.56 $X2=0 $Y2=0
cc_126 N_A_27_297#_M1002_d N_Y_c_204_n 0.00319213f $X=2.015 $Y=1.485 $X2=0 $Y2=0
cc_127 N_A_27_297#_c_133_n N_Y_c_204_n 0.00374545f $X=2.075 $Y=2.38 $X2=0 $Y2=0
cc_128 N_A_27_297#_c_134_n N_Y_c_204_n 0.0208421f $X=2.16 $Y=2 $X2=0 $Y2=0
cc_129 N_A_27_297#_c_132_n N_Y_c_206_n 0.0184068f $X=1.22 $Y=1.665 $X2=0 $Y2=0
cc_130 N_A_27_297#_c_148_p Y 0.0342667f $X=1.22 $Y=2.295 $X2=0 $Y2=0
cc_131 N_A_27_297#_c_133_n Y 0.0196128f $X=2.075 $Y=2.38 $X2=0 $Y2=0
cc_132 N_A_27_297#_c_134_n Y 0.0185225f $X=2.16 $Y=2 $X2=0 $Y2=0
cc_133 N_VPWR_c_168_n N_Y_M1001_s 0.00232895f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_134 N_Y_c_199_n N_VGND_M1007_s 0.00162089f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_135 N_Y_c_201_n N_VGND_M1006_d 0.0106573f $X=2.095 $Y=0.82 $X2=0 $Y2=0
cc_136 N_Y_c_200_n N_VGND_c_261_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_137 N_Y_c_207_n N_VGND_c_262_n 0.0231806f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_138 N_Y_c_199_n N_VGND_c_262_n 0.00254521f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_139 N_Y_c_199_n N_VGND_c_263_n 0.0122559f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_140 N_Y_c_201_n N_VGND_c_264_n 0.0139372f $X=2.095 $Y=0.82 $X2=0 $Y2=0
cc_141 N_Y_c_199_n N_VGND_c_266_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_142 N_Y_c_212_n N_VGND_c_266_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_143 N_Y_c_201_n N_VGND_c_266_n 0.00342158f $X=2.095 $Y=0.82 $X2=0 $Y2=0
cc_144 N_Y_M1003_d N_VGND_c_268_n 0.00304143f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_145 N_Y_M1004_s N_VGND_c_268_n 0.00304426f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_146 N_Y_c_207_n N_VGND_c_268_n 0.0143352f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_147 N_Y_c_199_n N_VGND_c_268_n 0.0094839f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_148 N_Y_c_212_n N_VGND_c_268_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_149 N_Y_c_201_n N_VGND_c_268_n 0.00752724f $X=2.095 $Y=0.82 $X2=0 $Y2=0
