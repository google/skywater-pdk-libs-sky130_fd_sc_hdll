* File: sky130_fd_sc_hdll__diode_6.pex.spice
* Created: Wed Sep  2 08:28:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DIODE_6%DIODE 1 4 10 54
r7 52 54 3.75385 $w=2.208e-06 $l=6.8e-07 $layer=LI1_cond $X=1.735 $Y=1.36
+ $X2=2.415 $Y2=1.36
r8 50 52 1.02127 $w=2.208e-06 $l=1.85e-07 $layer=LI1_cond $X=1.55 $Y=1.36
+ $X2=1.735 $Y2=1.36
r9 48 50 0.855656 $w=2.208e-06 $l=1.55e-07 $layer=LI1_cond $X=1.395 $Y=1.36
+ $X2=1.55 $Y2=1.36
r10 46 48 1.87692 $w=2.208e-06 $l=3.4e-07 $layer=LI1_cond $X=1.055 $Y=1.36
+ $X2=1.395 $Y2=1.36
r11 10 46 2.01493 $w=2.208e-06 $l=3.65e-07 $layer=LI1_cond $X=0.69 $Y=1.36
+ $X2=1.055 $Y2=1.36
r12 10 37 1.73891 $w=2.208e-06 $l=3.15e-07 $layer=LI1_cond $X=0.69 $Y=1.36
+ $X2=0.375 $Y2=1.36
r13 4 37 0.800452 $w=2.208e-06 $l=1.45e-07 $layer=LI1_cond $X=0.23 $Y=1.36
+ $X2=0.375 $Y2=1.36
r14 1 54 60.6667 $w=1.7e-07 $l=2.36588e-06 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=2.415 $Y2=0.37
r15 1 52 60.6667 $w=1.7e-07 $l=1.68523e-06 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=1.735 $Y2=0.37
r16 1 50 45.5 $w=1.7e-07 $l=1.79222e-06 $layer=licon1_NDIFF $count=4 $X=0.135
+ $Y=0.195 $X2=1.55 $Y2=1.05
r17 1 48 91 $w=1.7e-07 $l=1.34466e-06 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.195 $X2=1.395 $Y2=0.37
r18 1 46 60.6667 $w=1.7e-07 $l=1.00369e-06 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=1.055 $Y2=0.37
r19 1 37 60.6667 $w=1.7e-07 $l=3.15595e-07 $layer=licon1_NDIFF $count=3 $X=0.135
+ $Y=0.195 $X2=0.375 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__DIODE_6%VGND 1 8 9
r5 8 9 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r6 4 8 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r7 1 9 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=2.53
+ $Y2=0
r8 1 4 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
.ends

.subckt PM_SKY130_FD_SC_HDLL__DIODE_6%VPWR 1 8 9
r5 8 9 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72 $X2=2.53
+ $Y2=2.72
r6 4 8 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r7 1 9 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=0.23 $Y=2.72 $X2=2.53
+ $Y2=2.72
r8 1 4 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72 $X2=0.23
+ $Y2=2.72
.ends

