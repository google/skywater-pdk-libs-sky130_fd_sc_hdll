* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
X0 a_436_413# a_211_363# a_534_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 Q a_1323_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_1330_413# a_1323_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X3 VPWR a_1323_21# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_1237_47# a_1323_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X5 VPWR RESET_B a_649_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X6 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X7 a_436_413# a_27_47# a_534_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X8 Q a_1323_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_649_413# a_751_289# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 a_1128_47# a_211_363# a_1330_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 a_534_47# a_211_363# a_642_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X12 a_751_289# a_211_363# a_1128_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X13 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_751_289# a_27_47# a_1128_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X15 VGND D a_436_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 VPWR D a_436_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X17 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X18 a_805_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_1128_47# a_27_47# a_1237_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X20 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X21 VPWR a_534_47# a_751_289# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X22 VPWR RESET_B a_1323_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X23 VGND a_534_47# a_751_289# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 a_1323_21# a_1128_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X25 a_1542_47# a_1128_47# a_1323_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 a_534_47# a_27_47# a_649_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X27 VGND RESET_B a_1542_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_642_47# a_751_289# a_805_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VGND a_1323_21# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
