* File: sky130_fd_sc_hdll__clkinv_8.pex.spice
* Created: Wed Sep  2 08:26:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKINV_8%A 1 3 4 6 7 9 12 14 16 19 21 23 26 28 30
+ 33 35 37 40 42 44 47 49 51 54 56 58 61 63 65 66 68 69 70 71 72 73 74 75 76 77
+ 109 110 114 117 121 125 129 133 137 140 143
c170 109 0 1.51599e-19 $X=5.35 $Y=1.16
r171 109 111 38.7248 $w=5.85e-07 $l=4.7e-07 $layer=POLY_cond $X=5.35 $Y=1.11
+ $X2=5.82 $Y2=1.11
r172 109 110 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=5.35
+ $Y=1.16 $X2=5.35 $Y2=1.16
r173 107 109 26.7778 $w=5.85e-07 $l=3.25e-07 $layer=POLY_cond $X=5.025 $Y=1.11
+ $X2=5.35 $Y2=1.11
r174 106 107 16.0667 $w=5.85e-07 $l=1.95e-07 $layer=POLY_cond $X=4.83 $Y=1.11
+ $X2=5.025 $Y2=1.11
r175 105 106 27.6017 $w=5.85e-07 $l=3.35e-07 $layer=POLY_cond $X=4.495 $Y=1.11
+ $X2=4.83 $Y2=1.11
r176 104 105 15.2427 $w=5.85e-07 $l=1.85e-07 $layer=POLY_cond $X=4.31 $Y=1.11
+ $X2=4.495 $Y2=1.11
r177 103 104 28.4256 $w=5.85e-07 $l=3.45e-07 $layer=POLY_cond $X=3.965 $Y=1.11
+ $X2=4.31 $Y2=1.11
r178 102 103 14.4188 $w=5.85e-07 $l=1.75e-07 $layer=POLY_cond $X=3.79 $Y=1.11
+ $X2=3.965 $Y2=1.11
r179 101 102 29.2496 $w=5.85e-07 $l=3.55e-07 $layer=POLY_cond $X=3.435 $Y=1.11
+ $X2=3.79 $Y2=1.11
r180 100 101 9.47521 $w=5.85e-07 $l=1.15e-07 $layer=POLY_cond $X=3.32 $Y=1.11
+ $X2=3.435 $Y2=1.11
r181 99 100 30.0735 $w=5.85e-07 $l=3.65e-07 $layer=POLY_cond $X=2.955 $Y=1.11
+ $X2=3.32 $Y2=1.11
r182 98 99 8.65128 $w=5.85e-07 $l=1.05e-07 $layer=POLY_cond $X=2.85 $Y=1.11
+ $X2=2.955 $Y2=1.11
r183 97 98 30.8974 $w=5.85e-07 $l=3.75e-07 $layer=POLY_cond $X=2.475 $Y=1.11
+ $X2=2.85 $Y2=1.11
r184 96 97 7.82735 $w=5.85e-07 $l=9.5e-08 $layer=POLY_cond $X=2.38 $Y=1.11
+ $X2=2.475 $Y2=1.11
r185 95 96 31.7214 $w=5.85e-07 $l=3.85e-07 $layer=POLY_cond $X=1.995 $Y=1.11
+ $X2=2.38 $Y2=1.11
r186 94 95 7.00342 $w=5.85e-07 $l=8.5e-08 $layer=POLY_cond $X=1.91 $Y=1.11
+ $X2=1.995 $Y2=1.11
r187 93 94 32.5453 $w=5.85e-07 $l=3.95e-07 $layer=POLY_cond $X=1.515 $Y=1.11
+ $X2=1.91 $Y2=1.11
r188 92 93 6.17949 $w=5.85e-07 $l=7.5e-08 $layer=POLY_cond $X=1.44 $Y=1.11
+ $X2=1.515 $Y2=1.11
r189 91 92 39.1368 $w=5.85e-07 $l=4.75e-07 $layer=POLY_cond $X=0.965 $Y=1.11
+ $X2=1.44 $Y2=1.11
r190 89 91 28.4256 $w=5.85e-07 $l=3.45e-07 $layer=POLY_cond $X=0.62 $Y=1.11
+ $X2=0.965 $Y2=1.11
r191 89 114 22.3508 $w=1.7e-07 $l=1.105e-06 $layer=licon1_POLY $count=6 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r192 87 89 10.2991 $w=5.85e-07 $l=1.25e-07 $layer=POLY_cond $X=0.495 $Y=1.11
+ $X2=0.62 $Y2=1.11
r193 77 110 23.2748 $w=2.53e-07 $l=5.15e-07 $layer=LI1_cond $X=4.835 $Y=1.162
+ $X2=5.35 $Y2=1.162
r194 77 143 20.7892 $w=2.53e-07 $l=4.6e-07 $layer=LI1_cond $X=4.835 $Y=1.162
+ $X2=4.375 $Y2=1.162
r195 76 143 0.451938 $w=2.53e-07 $l=1e-08 $layer=LI1_cond $X=4.365 $Y=1.162
+ $X2=4.375 $Y2=1.162
r196 76 140 20.3372 $w=2.53e-07 $l=4.5e-07 $layer=LI1_cond $X=4.365 $Y=1.162
+ $X2=3.915 $Y2=1.162
r197 75 140 0.903877 $w=2.53e-07 $l=2e-08 $layer=LI1_cond $X=3.895 $Y=1.162
+ $X2=3.915 $Y2=1.162
r198 75 137 19.8853 $w=2.53e-07 $l=4.4e-07 $layer=LI1_cond $X=3.895 $Y=1.162
+ $X2=3.455 $Y2=1.162
r199 74 137 0.225969 $w=2.53e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.162
+ $X2=3.455 $Y2=1.162
r200 74 133 20.5632 $w=2.53e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.162
+ $X2=2.995 $Y2=1.162
r201 73 133 9.49071 $w=2.53e-07 $l=2.1e-07 $layer=LI1_cond $X=2.785 $Y=1.162
+ $X2=2.995 $Y2=1.162
r202 73 129 11.2985 $w=2.53e-07 $l=2.5e-07 $layer=LI1_cond $X=2.785 $Y=1.162
+ $X2=2.535 $Y2=1.162
r203 72 129 11.7504 $w=2.53e-07 $l=2.6e-07 $layer=LI1_cond $X=2.275 $Y=1.162
+ $X2=2.535 $Y2=1.162
r204 72 125 9.03877 $w=2.53e-07 $l=2e-07 $layer=LI1_cond $X=2.275 $Y=1.162
+ $X2=2.075 $Y2=1.162
r205 71 125 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=1.765 $Y=1.162
+ $X2=2.075 $Y2=1.162
r206 71 121 6.77908 $w=2.53e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.162
+ $X2=1.615 $Y2=1.162
r207 70 121 16.2698 $w=2.53e-07 $l=3.6e-07 $layer=LI1_cond $X=1.255 $Y=1.162
+ $X2=1.615 $Y2=1.162
r208 70 117 4.51938 $w=2.53e-07 $l=1e-07 $layer=LI1_cond $X=1.255 $Y=1.162
+ $X2=1.155 $Y2=1.162
r209 69 117 18.5295 $w=2.53e-07 $l=4.1e-07 $layer=LI1_cond $X=0.745 $Y=1.162
+ $X2=1.155 $Y2=1.162
r210 69 114 5.64923 $w=2.53e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.162
+ $X2=0.62 $Y2=1.162
r211 66 111 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.11
r212 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.82 $Y=1.41
+ $X2=5.82 $Y2=1.985
r213 63 109 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.11
r214 63 65 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.35 $Y=1.41
+ $X2=5.35 $Y2=1.985
r215 59 107 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=5.025 $Y=0.81
+ $X2=5.025 $Y2=1.11
r216 59 61 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=5.025 $Y=0.81
+ $X2=5.025 $Y2=0.445
r217 56 106 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=4.83 $Y=1.41
+ $X2=4.83 $Y2=1.11
r218 56 58 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.83 $Y=1.41
+ $X2=4.83 $Y2=1.985
r219 52 105 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=4.495 $Y=0.81
+ $X2=4.495 $Y2=1.11
r220 52 54 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=4.495 $Y=0.81
+ $X2=4.495 $Y2=0.445
r221 49 104 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=4.31 $Y=1.41
+ $X2=4.31 $Y2=1.11
r222 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.31 $Y=1.41
+ $X2=4.31 $Y2=1.985
r223 45 103 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.965 $Y=0.81
+ $X2=3.965 $Y2=1.11
r224 45 47 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.965 $Y=0.81
+ $X2=3.965 $Y2=0.445
r225 42 102 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.79 $Y=1.41
+ $X2=3.79 $Y2=1.11
r226 42 44 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.79 $Y=1.41
+ $X2=3.79 $Y2=1.985
r227 38 101 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=3.435 $Y=0.81
+ $X2=3.435 $Y2=1.11
r228 38 40 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=3.435 $Y=0.81
+ $X2=3.435 $Y2=0.445
r229 35 100 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=3.32 $Y=1.41
+ $X2=3.32 $Y2=1.11
r230 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.32 $Y=1.41
+ $X2=3.32 $Y2=1.985
r231 31 99 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.955 $Y=0.81
+ $X2=2.955 $Y2=1.11
r232 31 33 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.955 $Y=0.81
+ $X2=2.955 $Y2=0.445
r233 28 98 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=2.85 $Y=1.41 $X2=2.85
+ $Y2=1.11
r234 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.85 $Y=1.41
+ $X2=2.85 $Y2=1.985
r235 24 97 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=2.475 $Y=0.81
+ $X2=2.475 $Y2=1.11
r236 24 26 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=2.475 $Y=0.81
+ $X2=2.475 $Y2=0.445
r237 21 96 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=2.38 $Y=1.41 $X2=2.38
+ $Y2=1.11
r238 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.38 $Y=1.41
+ $X2=2.38 $Y2=1.985
r239 17 95 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.995 $Y=0.81
+ $X2=1.995 $Y2=1.11
r240 17 19 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.995 $Y=0.81
+ $X2=1.995 $Y2=0.445
r241 14 94 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.91 $Y=1.41 $X2=1.91
+ $Y2=1.11
r242 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.91 $Y=1.41
+ $X2=1.91 $Y2=1.985
r243 10 93 35.4195 $w=1.5e-07 $l=3e-07 $layer=POLY_cond $X=1.515 $Y=0.81
+ $X2=1.515 $Y2=1.11
r244 10 12 187.16 $w=1.5e-07 $l=3.65e-07 $layer=POLY_cond $X=1.515 $Y=0.81
+ $X2=1.515 $Y2=0.445
r245 7 92 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=1.44 $Y=1.41 $X2=1.44
+ $Y2=1.11
r246 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.44 $Y=1.41
+ $X2=1.44 $Y2=1.985
r247 4 91 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.11
r248 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r249 1 87 30.7696 $w=1.8e-07 $l=3e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.11
r250 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_8%VPWR 1 2 3 4 5 6 7 22 24 26 30 32 36 38
+ 42 44 48 52 54 56 59 60 61 67 75 78 81 84 88
r94 87 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r95 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r96 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r97 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r98 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r99 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r100 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r101 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r102 70 88 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r103 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r104 67 87 3.90794 $w=1.7e-07 $l=2.57e-07 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=6.182 $Y2=2.72
r105 67 69 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=5.925 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 66 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r107 66 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=3.91 $Y2=2.72
r108 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r109 63 84 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.2 $Y=2.72
+ $X2=4.047 $Y2=2.72
r110 63 65 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=4.2 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 61 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r112 61 72 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 59 65 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.945 $Y=2.72
+ $X2=4.83 $Y2=2.72
r114 59 60 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.945 $Y=2.72
+ $X2=5.095 $Y2=2.72
r115 58 69 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=5.245 $Y=2.72
+ $X2=5.75 $Y2=2.72
r116 58 60 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.245 $Y=2.72
+ $X2=5.095 $Y2=2.72
r117 54 87 3.26929 $w=2.55e-07 $l=1.67183e-07 $layer=LI1_cond $X=6.052 $Y=2.635
+ $X2=6.182 $Y2=2.72
r118 54 56 30.2799 $w=2.53e-07 $l=6.7e-07 $layer=LI1_cond $X=6.052 $Y=2.635
+ $X2=6.052 $Y2=1.965
r119 50 60 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.095 $Y=2.635
+ $X2=5.095 $Y2=2.72
r120 50 52 25.7379 $w=2.98e-07 $l=6.7e-07 $layer=LI1_cond $X=5.095 $Y=2.635
+ $X2=5.095 $Y2=1.965
r121 46 84 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.047 $Y=2.635
+ $X2=4.047 $Y2=2.72
r122 46 48 25.316 $w=3.03e-07 $l=6.7e-07 $layer=LI1_cond $X=4.047 $Y=2.635
+ $X2=4.047 $Y2=1.965
r123 45 81 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.21 $Y=2.72
+ $X2=3.087 $Y2=2.72
r124 44 84 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=4.047 $Y2=2.72
r125 44 45 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.895 $Y=2.72
+ $X2=3.21 $Y2=2.72
r126 40 81 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=2.72
r127 40 42 31.5158 $w=2.43e-07 $l=6.7e-07 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=1.965
r128 39 78 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.145 $Y2=2.72
r129 38 81 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=3.087 $Y2=2.72
r130 38 39 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.965 $Y=2.72
+ $X2=2.275 $Y2=2.72
r131 34 78 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=2.72
r132 34 36 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=2.145 $Y=2.635
+ $X2=2.145 $Y2=1.965
r133 33 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.205 $Y2=2.72
r134 32 78 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=2.145 $Y2=2.72
r135 32 33 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.015 $Y=2.72
+ $X2=1.335 $Y2=2.72
r136 28 75 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=2.635
+ $X2=1.205 $Y2=2.72
r137 28 30 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=1.205 $Y=2.635
+ $X2=1.205 $Y2=1.965
r138 27 72 4.06843 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r139 26 75 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=1.205 $Y2=2.72
r140 26 27 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=1.075 $Y=2.72
+ $X2=0.395 $Y2=2.72
r141 22 72 3.14379 $w=2.6e-07 $l=1.14039e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.197 $Y2=2.72
r142 22 24 29.6976 $w=2.58e-07 $l=6.7e-07 $layer=LI1_cond $X=0.265 $Y=2.635
+ $X2=0.265 $Y2=1.965
r143 7 56 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=5.91
+ $Y=1.485 $X2=6.055 $Y2=1.965
r144 6 52 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=4.92
+ $Y=1.485 $X2=5.065 $Y2=1.965
r145 5 48 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=3.88
+ $Y=1.485 $X2=4.025 $Y2=1.965
r146 4 42 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=2.94
+ $Y=1.485 $X2=3.085 $Y2=1.965
r147 3 36 300 $w=1.7e-07 $l=5.47723e-07 $layer=licon1_PDIFF $count=2 $X=2
+ $Y=1.485 $X2=2.145 $Y2=1.965
r148 2 30 300 $w=1.7e-07 $l=5.49909e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.205 $Y2=1.965
r149 1 24 300 $w=1.7e-07 $l=5.38888e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.965
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_8%Y 1 2 3 4 5 6 7 8 9 10 32 33 34 35 36 39
+ 41 45 49 51 53 57 61 63 65 69 73 75 77 81 85 87 89 93 95 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 115 116
r185 109 116 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=1.545
+ $X2=6.195 $Y2=1.46
r186 109 116 0.341465 $w=2.68e-07 $l=8e-09 $layer=LI1_cond $X=6.195 $Y=1.452
+ $X2=6.195 $Y2=1.46
r187 108 109 11.183 $w=2.68e-07 $l=2.62e-07 $layer=LI1_cond $X=6.195 $Y=1.19
+ $X2=6.195 $Y2=1.452
r188 107 115 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=0.78
+ $X2=6.195 $Y2=0.865
r189 107 108 12.3781 $w=2.68e-07 $l=2.9e-07 $layer=LI1_cond $X=6.195 $Y=0.9
+ $X2=6.195 $Y2=1.19
r190 107 115 1.49391 $w=2.68e-07 $l=3.5e-08 $layer=LI1_cond $X=6.195 $Y=0.9
+ $X2=6.195 $Y2=0.865
r191 96 106 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.705 $Y=1.545
+ $X2=5.585 $Y2=1.545
r192 95 109 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.06 $Y=1.545
+ $X2=6.195 $Y2=1.545
r193 95 96 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=6.06 $Y=1.545
+ $X2=5.705 $Y2=1.545
r194 91 106 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=5.585 $Y=1.63
+ $X2=5.585 $Y2=1.545
r195 91 93 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=5.585 $Y=1.63
+ $X2=5.585 $Y2=1.83
r196 90 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.855 $Y=0.78
+ $X2=4.76 $Y2=0.78
r197 89 107 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=6.06 $Y=0.78
+ $X2=6.195 $Y2=0.78
r198 89 90 78.615 $w=1.68e-07 $l=1.205e-06 $layer=LI1_cond $X=6.06 $Y=0.78
+ $X2=4.855 $Y2=0.78
r199 88 104 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=4.725 $Y=1.545
+ $X2=4.572 $Y2=1.545
r200 87 106 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=5.465 $Y=1.545
+ $X2=5.585 $Y2=1.545
r201 87 88 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=5.465 $Y=1.545
+ $X2=4.725 $Y2=1.545
r202 83 105 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.76 $Y=0.695
+ $X2=4.76 $Y2=0.78
r203 83 85 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=4.76 $Y=0.695
+ $X2=4.76 $Y2=0.445
r204 79 104 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=4.572 $Y=1.63
+ $X2=4.572 $Y2=1.545
r205 79 81 7.557 $w=3.03e-07 $l=2e-07 $layer=LI1_cond $X=4.572 $Y=1.63 $X2=4.572
+ $Y2=1.83
r206 78 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.795 $Y=0.78
+ $X2=3.7 $Y2=0.78
r207 77 105 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=4.665 $Y=0.78
+ $X2=4.76 $Y2=0.78
r208 77 78 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.665 $Y=0.78
+ $X2=3.795 $Y2=0.78
r209 76 102 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=3.675 $Y=1.545
+ $X2=3.552 $Y2=1.545
r210 75 104 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.42 $Y=1.545
+ $X2=4.572 $Y2=1.545
r211 75 76 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=4.42 $Y=1.545
+ $X2=3.675 $Y2=1.545
r212 71 103 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=3.7 $Y=0.695
+ $X2=3.7 $Y2=0.78
r213 71 73 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=3.7 $Y=0.695
+ $X2=3.7 $Y2=0.445
r214 67 102 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=3.552 $Y=1.63
+ $X2=3.552 $Y2=1.545
r215 67 69 9.4077 $w=2.43e-07 $l=2e-07 $layer=LI1_cond $X=3.552 $Y=1.63
+ $X2=3.552 $Y2=1.83
r216 66 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.835 $Y=0.78
+ $X2=2.74 $Y2=0.78
r217 65 103 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=3.605 $Y=0.78
+ $X2=3.7 $Y2=0.78
r218 65 66 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.605 $Y=0.78
+ $X2=2.835 $Y2=0.78
r219 64 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.745 $Y=1.545
+ $X2=2.62 $Y2=1.545
r220 63 102 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=3.43 $Y=1.545
+ $X2=3.552 $Y2=1.545
r221 63 64 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=3.43 $Y=1.545
+ $X2=2.745 $Y2=1.545
r222 59 101 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.74 $Y=0.695
+ $X2=2.74 $Y2=0.78
r223 59 61 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=2.74 $Y=0.695
+ $X2=2.74 $Y2=0.445
r224 55 100 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.62 $Y=1.63
+ $X2=2.62 $Y2=1.545
r225 55 57 9.21954 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=2.62 $Y=1.63 $X2=2.62
+ $Y2=1.83
r226 54 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.875 $Y=0.78
+ $X2=1.78 $Y2=0.78
r227 53 101 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.645 $Y=0.78
+ $X2=2.74 $Y2=0.78
r228 53 54 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.645 $Y=0.78
+ $X2=1.875 $Y2=0.78
r229 52 98 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.795 $Y=1.545
+ $X2=1.675 $Y2=1.545
r230 51 100 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.495 $Y=1.545
+ $X2=2.62 $Y2=1.545
r231 51 52 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.495 $Y=1.545
+ $X2=1.795 $Y2=1.545
r232 47 99 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.78 $Y=0.695
+ $X2=1.78 $Y2=0.78
r233 47 49 14.5933 $w=1.88e-07 $l=2.5e-07 $layer=LI1_cond $X=1.78 $Y=0.695
+ $X2=1.78 $Y2=0.445
r234 43 98 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=1.63
+ $X2=1.675 $Y2=1.545
r235 43 45 9.60369 $w=2.38e-07 $l=2e-07 $layer=LI1_cond $X=1.675 $Y=1.63
+ $X2=1.675 $Y2=1.83
r236 42 97 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.855 $Y=1.545
+ $X2=0.735 $Y2=1.545
r237 41 98 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.555 $Y=1.545
+ $X2=1.675 $Y2=1.545
r238 41 42 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.555 $Y=1.545
+ $X2=0.855 $Y2=1.545
r239 37 97 0.135687 $w=2.4e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=1.63
+ $X2=0.735 $Y2=1.545
r240 37 39 14.4055 $w=2.38e-07 $l=3e-07 $layer=LI1_cond $X=0.735 $Y=1.63
+ $X2=0.735 $Y2=1.93
r241 35 97 6.81202 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=0.615 $Y=1.545
+ $X2=0.735 $Y2=1.545
r242 35 36 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.615 $Y=1.545
+ $X2=0.285 $Y2=1.545
r243 33 99 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.685 $Y=0.78
+ $X2=1.78 $Y2=0.78
r244 33 34 91.3369 $w=1.68e-07 $l=1.4e-06 $layer=LI1_cond $X=1.685 $Y=0.78
+ $X2=0.285 $Y2=0.78
r245 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=1.46
+ $X2=0.285 $Y2=1.545
r246 31 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.285 $Y2=0.78
r247 31 32 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=0.2 $Y=0.865
+ $X2=0.2 $Y2=1.46
r248 10 93 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=5.44
+ $Y=1.485 $X2=5.585 $Y2=1.83
r249 9 81 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=4.4
+ $Y=1.485 $X2=4.545 $Y2=1.83
r250 8 69 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=3.41
+ $Y=1.485 $X2=3.555 $Y2=1.83
r251 7 57 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=2.47
+ $Y=1.485 $X2=2.615 $Y2=1.83
r252 6 45 300 $w=1.7e-07 $l=4.11157e-07 $layer=licon1_PDIFF $count=2 $X=1.53
+ $Y=1.485 $X2=1.675 $Y2=1.83
r253 5 39 300 $w=1.7e-07 $l=5.12396e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.93
r254 4 85 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.57
+ $Y=0.235 $X2=4.76 $Y2=0.445
r255 3 73 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.51
+ $Y=0.235 $X2=3.7 $Y2=0.445
r256 2 61 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.55
+ $Y=0.235 $X2=2.74 $Y2=0.445
r257 1 49 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=1.59
+ $Y=0.235 $X2=1.78 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKINV_8%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 45 47 62 68 69 72 75
c94 69 0 1.51599e-19 $X=6.21 $Y=0
r95 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r96 72 73 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r97 69 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.29
+ $Y2=0
r98 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r99 66 75 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.505 $Y=0 $X2=5.29
+ $Y2=0
r100 66 68 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.505 $Y=0
+ $X2=6.21 $Y2=0
r101 65 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.29
+ $Y2=0
r102 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r103 62 75 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=5.075 $Y=0 $X2=5.29
+ $Y2=0
r104 62 64 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=5.075 $Y=0 $X2=4.83
+ $Y2=0
r105 61 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r106 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r107 58 61 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r108 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r109 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r110 55 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r111 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r112 52 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.465 $Y=0 $X2=1.3
+ $Y2=0
r113 52 54 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=1.465 $Y=0
+ $X2=2.07 $Y2=0
r114 47 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.3
+ $Y2=0
r115 47 49 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.135 $Y=0
+ $X2=0.23 $Y2=0
r116 45 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r117 45 49 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r118 43 60 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=4.015 $Y=0
+ $X2=3.91 $Y2=0
r119 43 44 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.015 $Y=0 $X2=4.23
+ $Y2=0
r120 42 64 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=4.445 $Y=0
+ $X2=4.83 $Y2=0
r121 42 44 10.2816 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.445 $Y=0 $X2=4.23
+ $Y2=0
r122 40 57 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=0 $X2=2.99
+ $Y2=0
r123 40 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.055 $Y=0 $X2=3.245
+ $Y2=0
r124 39 60 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=3.435 $Y=0
+ $X2=3.91 $Y2=0
r125 39 41 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.435 $Y=0 $X2=3.245
+ $Y2=0
r126 37 54 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.07
+ $Y2=0
r127 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.095 $Y=0 $X2=2.26
+ $Y2=0
r128 36 57 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.99
+ $Y2=0
r129 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0 $X2=2.26
+ $Y2=0
r130 32 75 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0
r131 32 34 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=5.29 $Y=0.085
+ $X2=5.29 $Y2=0.39
r132 28 44 1.67165 $w=4.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0
r133 28 30 8.1743 $w=4.28e-07 $l=3.05e-07 $layer=LI1_cond $X=4.23 $Y=0.085
+ $X2=4.23 $Y2=0.39
r134 24 41 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0
r135 24 26 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0.39
r136 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0
r137 20 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.26 $Y=0.085
+ $X2=2.26 $Y2=0.39
r138 16 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.3 $Y=0.085 $X2=1.3
+ $Y2=0
r139 16 18 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.3 $Y=0.085
+ $X2=1.3 $Y2=0.39
r140 5 34 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=5.1
+ $Y=0.235 $X2=5.29 $Y2=0.39
r141 4 30 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=4.04
+ $Y=0.235 $X2=4.23 $Y2=0.39
r142 3 26 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=3.03
+ $Y=0.235 $X2=3.22 $Y2=0.39
r143 2 22 182 $w=1.7e-07 $l=2.56027e-07 $layer=licon1_NDIFF $count=1 $X=2.07
+ $Y=0.235 $X2=2.26 $Y2=0.39
r144 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.39
.ends

