* File: sky130_fd_sc_hdll__or2_1.spice
* Created: Thu Aug 27 19:23:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or2_1.pex.spice"
.subckt sky130_fd_sc_hdll__or2_1  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1002 N_A_38_297#_M1002_d N_B_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.1092 PD=0.73 PS=1.36 NRD=9.996 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_38_297#_M1002_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0869439 AS=0.0651 PD=0.812523 PS=0.73 NRD=30 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1003 N_X_M1003_d N_A_38_297#_M1003_g N_VGND_M1004_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.134556 PD=1.92 PS=1.25748 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.8 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 A_128_297# N_B_M1001_g N_A_38_297#_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.1134 PD=0.65 PS=1.38 NRD=28.1316 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_128_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.0483 PD=0.801549 PS=0.65 NRD=35.1645 NRS=28.1316 M=1
+ R=2.33333 SA=90000.6 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1005 N_X_M1005_d N_A_38_297#_M1005_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1
+ AD=0.35 AS=0.215282 PD=2.7 PS=1.90845 NRD=16.7253 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.3 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_10 X X PROBETYPE=1
c_148 A_128_297# 0 9.99956e-20 $X=0.64 $Y=1.485
*
.include "sky130_fd_sc_hdll__or2_1.pxi.spice"
*
.ends
*
*
