* File: sky130_fd_sc_hdll__dlygate4sd3_1.pxi.spice
* Created: Wed Sep  2 08:30:29 2020
* 
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A N_A_M1002_g N_A_M1004_g A A N_A_c_64_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_27_47# N_A_27_47#_M1004_s
+ N_A_27_47#_M1002_s N_A_27_47#_M1003_g N_A_27_47#_M1007_g N_A_27_47#_c_101_n
+ N_A_27_47#_c_95_n N_A_27_47#_c_96_n N_A_27_47#_c_97_n N_A_27_47#_c_102_n
+ N_A_27_47#_c_103_n N_A_27_47#_c_104_n N_A_27_47#_c_126_p N_A_27_47#_c_98_n
+ N_A_27_47#_c_99_n PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_273_47# N_A_273_47#_M1003_d
+ N_A_273_47#_M1007_d N_A_273_47#_c_164_n N_A_273_47#_M1006_g
+ N_A_273_47#_M1000_g N_A_273_47#_c_165_n N_A_273_47#_c_166_n
+ N_A_273_47#_c_167_n N_A_273_47#_c_168_n N_A_273_47#_c_172_n
+ N_A_273_47#_c_169_n PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_273_47#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_379_93# N_A_379_93#_M1006_s
+ N_A_379_93#_M1000_s N_A_379_93#_M1001_g N_A_379_93#_M1005_g
+ N_A_379_93#_c_233_n N_A_379_93#_c_227_n N_A_379_93#_c_228_n
+ N_A_379_93#_c_221_n N_A_379_93#_c_222_n N_A_379_93#_c_230_n
+ N_A_379_93#_c_223_n N_A_379_93#_c_224_n N_A_379_93#_c_225_n
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%A_379_93#
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VPWR N_VPWR_M1002_d N_VPWR_M1000_d
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_281_n N_VPWR_c_282_n VPWR
+ N_VPWR_c_283_n N_VPWR_c_284_n N_VPWR_c_278_n N_VPWR_c_286_n VPWR
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VPWR
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%X N_X_M1005_d N_X_M1001_d X X X X X X X
+ N_X_c_319_n X PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%X
x_PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VGND N_VGND_M1004_d N_VGND_M1006_d
+ N_VGND_c_337_n N_VGND_c_338_n N_VGND_c_339_n N_VGND_c_340_n VGND
+ N_VGND_c_341_n N_VGND_c_342_n N_VGND_c_343_n N_VGND_c_344_n VGND
+ PM_SKY130_FD_SC_HDLL__DLYGATE4SD3_1%VGND
cc_1 VNB N_A_M1004_g 0.035522f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.445
cc_2 VNB A 0.0126787f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_3 VNB N_A_c_64_n 0.0334471f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.16
cc_4 VNB N_A_27_47#_M1003_g 0.0617273f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_5 VNB N_A_27_47#_c_95_n 0.0185706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_96_n 0.00913047f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.53
cc_7 VNB N_A_27_47#_c_97_n 0.00974844f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_98_n 0.0340688f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_99_n 0.00456744f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_273_47#_c_164_n 0.115096f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.445
cc_11 VNB N_A_273_47#_c_165_n 0.0107825f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_12 VNB N_A_273_47#_c_166_n 5.20958e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_273_47#_c_167_n 0.00658895f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_273_47#_c_168_n 0.00599379f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_273_47#_c_169_n 0.00177789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_379_93#_c_221_n 0.00248029f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.16
cc_17 VNB N_A_379_93#_c_222_n 0.00580676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_379_93#_c_223_n 0.00155374f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_379_93#_c_224_n 0.0273706f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_379_93#_c_225_n 0.0205286f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VPWR_c_278_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.0242902f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_X_c_319_n 0.0250158f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_337_n 0.00496928f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_25 VNB N_VGND_c_338_n 0.00817934f $X=-0.19 $Y=-0.24 $X2=0.31 $Y2=1.16
cc_26 VNB N_VGND_c_339_n 0.0515939f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_340_n 0.00631673f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.16
cc_28 VNB N_VGND_c_341_n 0.0177317f $X=-0.19 $Y=-0.24 $X2=0.345 $Y2=1.16
cc_29 VNB N_VGND_c_342_n 0.019232f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_343_n 0.211217f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_344_n 0.00410791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_A_M1002_g 0.0641083f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.275
cc_33 VPB A 0.0179142f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_34 VPB N_A_c_64_n 0.00821038f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_35 VPB N_A_27_47#_M1007_g 0.0985814f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_36 VPB N_A_27_47#_c_101_n 0.0188184f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.16
cc_37 VPB N_A_27_47#_c_102_n 0.00923338f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A_27_47#_c_103_n 0.0123946f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_104_n 0.00339742f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_98_n 0.00603539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_273_47#_c_164_n 0.120666f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.445
cc_42 VPB N_A_273_47#_c_166_n 0.0200526f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_273_47#_c_172_n 0.00620265f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_379_93#_M1001_g 0.0263455f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_45 VPB N_A_379_93#_c_227_n 0.00131442f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_46 VPB N_A_379_93#_c_228_n 0.00296707f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_379_93#_c_222_n 5.80315e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_379_93#_c_230_n 0.00274824f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.53
cc_49 VPB N_A_379_93#_c_224_n 0.00609669f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_279_n 0.00516546f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_51 VPB N_VPWR_c_280_n 0.0096412f $X=-0.19 $Y=1.305 $X2=0.31 $Y2=1.16
cc_52 VPB N_VPWR_c_281_n 0.0528193f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_53 VPB N_VPWR_c_282_n 0.00631825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_283_n 0.0177778f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_284_n 0.019232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_278_n 0.057119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_286_n 0.00478085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB X 0.0333747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB X 0.00949268f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB X 0.00857108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 N_A_M1004_g N_A_27_47#_M1003_g 0.0259108f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_62 N_A_M1002_g N_A_27_47#_M1007_g 0.0440108f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_63 A N_A_27_47#_M1007_g 8.8619e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_64 N_A_M1002_g N_A_27_47#_c_101_n 0.00381471f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_65 N_A_M1004_g N_A_27_47#_c_95_n 0.00358272f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_66 N_A_M1004_g N_A_27_47#_c_96_n 0.0130662f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_67 A N_A_27_47#_c_96_n 0.0171114f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_c_64_n N_A_27_47#_c_96_n 0.00144656f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_97_n 0.0252593f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_70 N_A_c_64_n N_A_27_47#_c_97_n 0.00511105f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_M1002_g N_A_27_47#_c_102_n 0.0176995f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_102_n 0.017423f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_73 A N_A_27_47#_c_103_n 0.0271506f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_64_n N_A_27_47#_c_103_n 8.59854e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_75 N_A_M1002_g N_A_27_47#_c_104_n 0.00424788f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_76 A N_A_27_47#_c_98_n 9.17263e-19 $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_77 N_A_c_64_n N_A_27_47#_c_98_n 0.0214298f $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_M1004_g N_A_27_47#_c_99_n 0.00359569f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_79 A N_A_27_47#_c_99_n 0.0460051f $X=0.14 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A_c_64_n N_A_27_47#_c_99_n 8.10742e-19 $X=0.51 $Y=1.16 $X2=0 $Y2=0
cc_81 N_A_M1002_g N_VPWR_c_279_n 0.00299091f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_82 N_A_M1002_g N_VPWR_c_283_n 0.00523784f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_83 N_A_M1002_g N_VPWR_c_278_n 0.00778046f $X=0.495 $Y=2.275 $X2=0 $Y2=0
cc_84 N_A_M1004_g N_VGND_c_337_n 0.00296217f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_85 N_A_M1004_g N_VGND_c_341_n 0.00436487f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_86 N_A_M1004_g N_VGND_c_343_n 0.00689889f $X=0.51 $Y=0.445 $X2=0 $Y2=0
cc_87 N_A_27_47#_c_126_p N_A_273_47#_c_164_n 2.10632e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_88 N_A_27_47#_c_98_n N_A_273_47#_c_164_n 0.00792752f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_89 N_A_27_47#_M1003_g N_A_273_47#_c_165_n 0.0135846f $X=1.115 $Y=0.445 $X2=0
+ $Y2=0
cc_90 N_A_27_47#_c_126_p N_A_273_47#_c_165_n 0.00607815f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_91 N_A_27_47#_c_98_n N_A_273_47#_c_165_n 7.17975e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_92 N_A_27_47#_c_99_n N_A_273_47#_c_165_n 0.0074409f $X=0.86 $Y=0.8 $X2=0
+ $Y2=0
cc_93 N_A_27_47#_M1007_g N_A_273_47#_c_166_n 0.0246818f $X=1.115 $Y=2.275 $X2=0
+ $Y2=0
cc_94 N_A_27_47#_c_102_n N_A_273_47#_c_166_n 0.00644317f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_95 N_A_27_47#_c_126_p N_A_273_47#_c_166_n 0.00375564f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_96 N_A_27_47#_c_98_n N_A_273_47#_c_166_n 4.49636e-19 $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_97 N_A_27_47#_c_99_n N_A_273_47#_c_166_n 0.0122032f $X=0.86 $Y=0.8 $X2=0
+ $Y2=0
cc_98 N_A_27_47#_M1003_g N_A_273_47#_c_168_n 0.00979252f $X=1.115 $Y=0.445 $X2=0
+ $Y2=0
cc_99 N_A_27_47#_c_126_p N_A_273_47#_c_168_n 0.00260624f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_M1007_g N_A_273_47#_c_172_n 0.0109054f $X=1.115 $Y=2.275 $X2=0
+ $Y2=0
cc_101 N_A_27_47#_c_126_p N_A_273_47#_c_169_n 0.0173287f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_102 N_A_27_47#_c_98_n N_A_273_47#_c_169_n 0.00196291f $X=1.27 $Y=1.16 $X2=0
+ $Y2=0
cc_103 N_A_27_47#_M1007_g N_VPWR_c_279_n 0.00312244f $X=1.115 $Y=2.275 $X2=0
+ $Y2=0
cc_104 N_A_27_47#_c_102_n N_VPWR_c_279_n 0.0168533f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_105 N_A_27_47#_M1007_g N_VPWR_c_281_n 0.0178079f $X=1.115 $Y=2.275 $X2=0
+ $Y2=0
cc_106 N_A_27_47#_c_102_n N_VPWR_c_281_n 0.00136391f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_107 N_A_27_47#_c_101_n N_VPWR_c_283_n 0.0195913f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_108 N_A_27_47#_c_102_n N_VPWR_c_283_n 0.0032011f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_109 N_A_27_47#_M1002_s N_VPWR_c_278_n 0.00229573f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_110 N_A_27_47#_M1007_g N_VPWR_c_278_n 0.0287032f $X=1.115 $Y=2.275 $X2=0
+ $Y2=0
cc_111 N_A_27_47#_c_101_n N_VPWR_c_278_n 0.0112839f $X=0.26 $Y=2.21 $X2=0 $Y2=0
cc_112 N_A_27_47#_c_102_n N_VPWR_c_278_n 0.00821595f $X=0.775 $Y=1.895 $X2=0
+ $Y2=0
cc_113 N_A_27_47#_M1003_g N_VGND_c_337_n 0.00284427f $X=1.115 $Y=0.445 $X2=0
+ $Y2=0
cc_114 N_A_27_47#_c_96_n N_VGND_c_337_n 0.0119788f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_99_n N_VGND_c_337_n 0.00307236f $X=0.86 $Y=0.8 $X2=0 $Y2=0
cc_116 N_A_27_47#_M1003_g N_VGND_c_339_n 0.0178179f $X=1.115 $Y=0.445 $X2=0
+ $Y2=0
cc_117 N_A_27_47#_c_99_n N_VGND_c_339_n 0.00204972f $X=0.86 $Y=0.8 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_95_n N_VGND_c_341_n 0.019808f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_96_n N_VGND_c_341_n 0.00312415f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_120 N_A_27_47#_M1004_s N_VGND_c_343_n 0.00268635f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_121 N_A_27_47#_M1003_g N_VGND_c_343_n 0.0288352f $X=1.115 $Y=0.445 $X2=0
+ $Y2=0
cc_122 N_A_27_47#_c_95_n N_VGND_c_343_n 0.0108719f $X=0.26 $Y=0.51 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_96_n N_VGND_c_343_n 0.00573599f $X=0.775 $Y=0.8 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_99_n N_VGND_c_343_n 0.0033826f $X=0.86 $Y=0.8 $X2=0 $Y2=0
cc_125 N_A_273_47#_c_164_n N_A_379_93#_M1001_g 0.0277062f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_126 N_A_273_47#_c_166_n N_A_379_93#_c_233_n 0.02522f $X=1.655 $Y=2.175 $X2=0
+ $Y2=0
cc_127 N_A_273_47#_c_164_n N_A_379_93#_c_227_n 0.046608f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_128 N_A_273_47#_c_167_n N_A_379_93#_c_227_n 0.0151066f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_273_47#_c_164_n N_A_379_93#_c_228_n 0.00497758f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_130 N_A_273_47#_c_166_n N_A_379_93#_c_228_n 0.0142871f $X=1.655 $Y=2.175
+ $X2=0 $Y2=0
cc_131 N_A_273_47#_c_167_n N_A_379_93#_c_228_n 0.0114696f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_132 N_A_273_47#_c_164_n N_A_379_93#_c_221_n 0.0333611f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_133 N_A_273_47#_c_167_n N_A_379_93#_c_221_n 0.0230499f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_134 N_A_273_47#_c_164_n N_A_379_93#_c_222_n 0.00719164f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_135 N_A_273_47#_c_167_n N_A_379_93#_c_222_n 0.0100466f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_136 N_A_273_47#_c_164_n N_A_379_93#_c_230_n 0.00604455f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_137 N_A_273_47#_c_164_n N_A_379_93#_c_223_n 0.0062773f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_138 N_A_273_47#_c_165_n N_A_379_93#_c_223_n 0.0272617f $X=1.655 $Y=1.075
+ $X2=0 $Y2=0
cc_139 N_A_273_47#_c_167_n N_A_379_93#_c_223_n 0.0177566f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_140 N_A_273_47#_c_168_n N_A_379_93#_c_223_n 0.00278075f $X=1.655 $Y=0.4 $X2=0
+ $Y2=0
cc_141 N_A_273_47#_c_164_n N_A_379_93#_c_224_n 0.0218228f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_142 N_A_273_47#_c_164_n N_A_379_93#_c_225_n 0.0235188f $X=2.405 $Y=0.995
+ $X2=0 $Y2=0
cc_143 N_A_273_47#_c_164_n N_VPWR_c_280_n 0.0157874f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_144 N_A_273_47#_c_164_n N_VPWR_c_281_n 0.0195128f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_A_273_47#_c_172_n N_VPWR_c_281_n 0.0268116f $X=1.655 $Y=2.32 $X2=0
+ $Y2=0
cc_146 N_A_273_47#_M1007_d N_VPWR_c_278_n 0.00209344f $X=1.365 $Y=2.065 $X2=0
+ $Y2=0
cc_147 N_A_273_47#_c_164_n N_VPWR_c_278_n 0.0338754f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_273_47#_c_172_n N_VPWR_c_278_n 0.0160449f $X=1.655 $Y=2.32 $X2=0
+ $Y2=0
cc_149 N_A_273_47#_c_164_n X 9.81975e-19 $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A_273_47#_c_164_n N_X_c_319_n 0.00102685f $X=2.405 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_273_47#_c_164_n N_VGND_c_338_n 0.0111736f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_152 N_A_273_47#_c_164_n N_VGND_c_339_n 0.0146402f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_153 N_A_273_47#_c_168_n N_VGND_c_339_n 0.0268432f $X=1.655 $Y=0.4 $X2=0 $Y2=0
cc_154 N_A_273_47#_M1003_d N_VGND_c_343_n 0.00209344f $X=1.365 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_273_47#_c_164_n N_VGND_c_343_n 0.0183107f $X=2.405 $Y=0.995 $X2=0
+ $Y2=0
cc_156 N_A_273_47#_c_168_n N_VGND_c_343_n 0.0160493f $X=1.655 $Y=0.4 $X2=0 $Y2=0
cc_157 N_A_379_93#_c_227_n N_VPWR_M1000_d 0.00570539f $X=2.81 $Y=1.66 $X2=0
+ $Y2=0
cc_158 N_A_379_93#_c_230_n N_VPWR_M1000_d 0.00157589f $X=2.915 $Y=1.575 $X2=0
+ $Y2=0
cc_159 N_A_379_93#_M1001_g N_VPWR_c_280_n 0.00329194f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_160 N_A_379_93#_c_227_n N_VPWR_c_280_n 0.0225879f $X=2.81 $Y=1.66 $X2=0 $Y2=0
cc_161 N_A_379_93#_c_224_n N_VPWR_c_280_n 4.55026e-19 $X=3.03 $Y=1.16 $X2=0
+ $Y2=0
cc_162 N_A_379_93#_c_233_n N_VPWR_c_281_n 0.00379879f $X=2.02 $Y=1.915 $X2=0
+ $Y2=0
cc_163 N_A_379_93#_M1001_g N_VPWR_c_284_n 0.00673617f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_164 N_A_379_93#_M1001_g N_VPWR_c_278_n 0.0128984f $X=3.12 $Y=1.985 $X2=0
+ $Y2=0
cc_165 N_A_379_93#_c_233_n N_VPWR_c_278_n 0.00644579f $X=2.02 $Y=1.915 $X2=0
+ $Y2=0
cc_166 N_A_379_93#_M1001_g X 0.00996615f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_167 N_A_379_93#_c_222_n X 0.0320535f $X=2.915 $Y=1.325 $X2=0 $Y2=0
cc_168 N_A_379_93#_c_230_n X 0.0063006f $X=2.915 $Y=1.575 $X2=0 $Y2=0
cc_169 N_A_379_93#_c_225_n X 0.0133381f $X=3.037 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_379_93#_c_225_n N_X_c_319_n 0.00806966f $X=3.037 $Y=0.995 $X2=0 $Y2=0
cc_171 N_A_379_93#_M1001_g X 0.00265072f $X=3.12 $Y=1.985 $X2=0 $Y2=0
cc_172 N_A_379_93#_c_221_n N_VGND_M1006_d 0.00100734f $X=2.81 $Y=0.82 $X2=0
+ $Y2=0
cc_173 N_A_379_93#_c_222_n N_VGND_M1006_d 0.00283033f $X=2.915 $Y=1.325 $X2=0
+ $Y2=0
cc_174 N_A_379_93#_c_221_n N_VGND_c_338_n 0.00765622f $X=2.81 $Y=0.82 $X2=0
+ $Y2=0
cc_175 N_A_379_93#_c_222_n N_VGND_c_338_n 0.016733f $X=2.915 $Y=1.325 $X2=0
+ $Y2=0
cc_176 N_A_379_93#_c_224_n N_VGND_c_338_n 6.50133e-19 $X=3.03 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_379_93#_c_225_n N_VGND_c_338_n 0.00509206f $X=3.037 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_379_93#_c_221_n N_VGND_c_339_n 0.0069179f $X=2.81 $Y=0.82 $X2=0 $Y2=0
cc_179 N_A_379_93#_c_223_n N_VGND_c_339_n 0.00524776f $X=2.02 $Y=0.675 $X2=0
+ $Y2=0
cc_180 N_A_379_93#_c_225_n N_VGND_c_342_n 0.0055654f $X=3.037 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_379_93#_c_221_n N_VGND_c_343_n 0.012399f $X=2.81 $Y=0.82 $X2=0 $Y2=0
cc_182 N_A_379_93#_c_222_n N_VGND_c_343_n 8.88378e-19 $X=2.915 $Y=1.325 $X2=0
+ $Y2=0
cc_183 N_A_379_93#_c_223_n N_VGND_c_343_n 0.00734212f $X=2.02 $Y=0.675 $X2=0
+ $Y2=0
cc_184 N_A_379_93#_c_225_n N_VGND_c_343_n 0.0112765f $X=3.037 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_278_n N_X_M1001_d 0.00217517f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_186 N_VPWR_c_284_n X 0.0264367f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_187 N_VPWR_c_278_n X 0.0153609f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_188 N_X_c_319_n N_VGND_c_342_n 0.0263689f $X=3.355 $Y=0.38 $X2=0 $Y2=0
cc_189 N_X_M1005_d N_VGND_c_343_n 0.00217517f $X=3.21 $Y=0.235 $X2=0 $Y2=0
cc_190 N_X_c_319_n N_VGND_c_343_n 0.0153377f $X=3.355 $Y=0.38 $X2=0 $Y2=0
