* File: sky130_fd_sc_hdll__o31ai_2.pex.spice
* Created: Thu Aug 27 19:22:32 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A1 1 3 6 8 10 13 15 16 17 29 36 40
c48 29 0 1.90595e-19 $X=0.985 $Y=1.217
r49 29 30 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.217
+ $X2=1.01 $Y2=1.217
r50 28 40 12.1647 $w=2.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.87 $Y=1.19
+ $X2=1.155 $Y2=1.19
r51 27 29 16.848 $w=3.29e-07 $l=1.15e-07 $layer=POLY_cond $X=0.87 $Y=1.217
+ $X2=0.985 $Y2=1.217
r52 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.87
+ $Y=1.16 $X2=0.87 $Y2=1.16
r53 25 27 48.3465 $w=3.29e-07 $l=3.3e-07 $layer=POLY_cond $X=0.54 $Y=1.217
+ $X2=0.87 $Y2=1.217
r54 24 25 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.217
+ $X2=0.54 $Y2=1.217
r55 23 36 9.17686 $w=2.68e-07 $l=2.15e-07 $layer=LI1_cond $X=0.48 $Y=1.19
+ $X2=0.695 $Y2=1.19
r56 22 24 5.12766 $w=3.29e-07 $l=3.5e-08 $layer=POLY_cond $X=0.48 $Y=1.217
+ $X2=0.515 $Y2=1.217
r57 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.48
+ $Y=1.16 $X2=0.48 $Y2=1.16
r58 17 40 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=1.16 $Y=1.19
+ $X2=1.155 $Y2=1.19
r59 16 28 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.19
+ $X2=0.87 $Y2=1.19
r60 16 36 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=0.745 $Y=1.19
+ $X2=0.695 $Y2=1.19
r61 15 23 10.4574 $w=2.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.235 $Y=1.19
+ $X2=0.48 $Y2=1.19
r62 11 30 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.01 $Y=1.025
+ $X2=1.01 $Y2=1.217
r63 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.01 $Y=1.025
+ $X2=1.01 $Y2=0.56
r64 8 29 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.217
r65 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r66 4 25 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.54 $Y=1.025
+ $X2=0.54 $Y2=1.217
r67 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.54 $Y=1.025
+ $X2=0.54 $Y2=0.56
r68 1 24 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.217
r69 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A2 3 5 7 8 10 13 15 16 26 30 36
c48 36 0 1.90595e-19 $X=2.075 $Y=1.19
r49 26 28 34.6486 $w=3.13e-07 $l=2.25e-07 $layer=POLY_cond $X=2.115 $Y=1.217
+ $X2=2.34 $Y2=1.217
r50 26 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.115
+ $Y=1.16 $X2=2.115 $Y2=1.16
r51 24 26 29.2588 $w=3.13e-07 $l=1.9e-07 $layer=POLY_cond $X=1.925 $Y=1.217
+ $X2=2.115 $Y2=1.217
r52 22 24 30.7987 $w=3.13e-07 $l=2e-07 $layer=POLY_cond $X=1.725 $Y=1.217
+ $X2=1.925 $Y2=1.217
r53 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r54 20 22 41.5783 $w=3.13e-07 $l=2.7e-07 $layer=POLY_cond $X=1.455 $Y=1.217
+ $X2=1.725 $Y2=1.217
r55 19 20 3.84984 $w=3.13e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.217
+ $X2=1.455 $Y2=1.217
r56 16 36 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=1.19
+ $X2=2.075 $Y2=1.19
r57 16 23 14.7257 $w=2.68e-07 $l=3.45e-07 $layer=LI1_cond $X=2.07 $Y=1.19
+ $X2=1.725 $Y2=1.19
r58 15 23 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=1.635 $Y=1.19
+ $X2=1.725 $Y2=1.19
r59 15 30 0.853661 $w=2.68e-07 $l=2e-08 $layer=LI1_cond $X=1.635 $Y=1.19
+ $X2=1.615 $Y2=1.19
r60 11 28 19.9686 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.34 $Y=1.025
+ $X2=2.34 $Y2=1.217
r61 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.34 $Y=1.025
+ $X2=2.34 $Y2=0.56
r62 8 24 15.7022 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.217
r63 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r64 5 20 15.7022 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.217
r65 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r66 1 19 19.9686 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.43 $Y=1.025
+ $X2=1.43 $Y2=1.217
r67 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.43 $Y=1.025
+ $X2=1.43 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A3 3 5 7 8 10 13 15 16 27
c55 3 0 1.21354e-19 $X=2.86 $Y=0.56
r56 27 28 3.66261 $w=3.29e-07 $l=2.5e-08 $layer=POLY_cond $X=3.455 $Y=1.217
+ $X2=3.48 $Y2=1.217
r57 25 27 16.848 $w=3.29e-07 $l=1.15e-07 $layer=POLY_cond $X=3.34 $Y=1.217
+ $X2=3.455 $Y2=1.217
r58 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.34
+ $Y=1.16 $X2=3.34 $Y2=1.16
r59 23 25 52.0091 $w=3.29e-07 $l=3.55e-07 $layer=POLY_cond $X=2.985 $Y=1.217
+ $X2=3.34 $Y2=1.217
r60 21 23 5.12766 $w=3.29e-07 $l=3.5e-08 $layer=POLY_cond $X=2.95 $Y=1.217
+ $X2=2.985 $Y2=1.217
r61 19 21 13.1854 $w=3.29e-07 $l=9e-08 $layer=POLY_cond $X=2.86 $Y=1.217
+ $X2=2.95 $Y2=1.217
r62 16 26 4.26831 $w=2.68e-07 $l=1e-07 $layer=LI1_cond $X=3.44 $Y=1.19 $X2=3.34
+ $Y2=1.19
r63 15 26 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=2.95 $Y=1.19
+ $X2=3.34 $Y2=1.19
r64 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r65 11 28 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.48 $Y=1.025
+ $X2=3.48 $Y2=1.217
r66 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.48 $Y=1.025
+ $X2=3.48 $Y2=0.56
r67 8 27 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.455 $Y2=1.217
r68 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.455 $Y=1.41
+ $X2=3.455 $Y2=1.985
r69 5 23 16.8611 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.217
r70 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.985
r71 1 19 21.1507 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.86 $Y=1.025
+ $X2=2.86 $Y2=1.217
r72 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.86 $Y=1.025
+ $X2=2.86 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%B1 1 3 4 6 7 9 11 12 14 15 16 17 21
c53 17 0 7.9412e-20 $X=4.83 $Y=0.85
r54 21 23 39.279 $w=3.62e-07 $l=2.95e-07 $layer=POLY_cond $X=4.515 $Y=1.202
+ $X2=4.81 $Y2=1.202
r55 20 21 3.32873 $w=3.62e-07 $l=2.5e-08 $layer=POLY_cond $X=4.49 $Y=1.202
+ $X2=4.515 $Y2=1.202
r56 16 17 10.5076 $w=3.38e-07 $l=3.1e-07 $layer=LI1_cond $X=4.8 $Y=1.16 $X2=4.8
+ $Y2=0.85
r57 16 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.81
+ $Y=1.16 $X2=4.81 $Y2=1.16
r58 12 21 19.0988 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.515 $Y=1.41
+ $X2=4.515 $Y2=1.202
r59 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.515 $Y=1.41
+ $X2=4.515 $Y2=1.985
r60 9 20 23.4391 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.49 $Y=0.995
+ $X2=4.49 $Y2=1.202
r61 9 11 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.49 $Y=0.995
+ $X2=4.49 $Y2=0.56
r62 8 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=4.025 $Y=1.16
+ $X2=3.925 $Y2=1.202
r63 7 20 10.4561 $w=3.62e-07 $l=9.3675e-08 $layer=POLY_cond $X=4.415 $Y=1.16
+ $X2=4.49 $Y2=1.202
r64 7 8 68.1959 $w=3.3e-07 $l=3.9e-07 $layer=POLY_cond $X=4.415 $Y=1.16
+ $X2=4.025 $Y2=1.16
r65 4 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.202
r66 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.925 $Y=1.41
+ $X2=3.925 $Y2=1.985
r67 1 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.9 $Y=0.995
+ $X2=3.925 $Y2=1.202
r68 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.9 $Y=0.995 $X2=3.9
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_297# 1 2 3 12 16 17 20 24 28 30
r49 26 28 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.135 $Y=1.665
+ $X2=2.135 $Y2=1.68
r50 25 30 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=1.58
+ $X2=1.195 $Y2=1.58
r51 24 26 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=1.945 $Y=1.58
+ $X2=2.135 $Y2=1.665
r52 24 25 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.945 $Y=1.58
+ $X2=1.385 $Y2=1.58
r53 20 22 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.195 $Y=1.68
+ $X2=1.195 $Y2=2.36
r54 18 30 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=1.58
r55 18 20 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.195 $Y=1.665
+ $X2=1.195 $Y2=1.68
r56 16 30 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=1.58
+ $X2=1.195 $Y2=1.58
r57 16 17 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=1.58
+ $X2=0.445 $Y2=1.58
r58 12 14 22.075 $w=3.53e-07 $l=6.8e-07 $layer=LI1_cond $X=0.267 $Y=1.68
+ $X2=0.267 $Y2=2.36
r59 10 17 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=1.665
+ $X2=0.445 $Y2=1.58
r60 10 12 0.486948 $w=3.53e-07 $l=1.5e-08 $layer=LI1_cond $X=0.267 $Y=1.665
+ $X2=0.267 $Y2=1.68
r61 3 28 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.68
r62 2 22 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.36
r63 2 20 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.68
r64 1 14 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.36
r65 1 12 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%VPWR 1 2 11 15 18 19 20 30 31 34 37
r56 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r57 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r58 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r59 27 28 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 25 28 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r61 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r62 24 27 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r63 24 25 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r64 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.75 $Y2=2.72
r65 22 24 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 20 35 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 20 37 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r68 18 27 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 18 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.075 $Y=2.72
+ $X2=4.24 $Y2=2.72
r70 17 30 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.83 $Y2=2.72
r71 17 19 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.405 $Y=2.72
+ $X2=4.24 $Y2=2.72
r72 13 19 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.24 $Y=2.635
+ $X2=4.24 $Y2=2.72
r73 13 15 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=4.24 $Y=2.635
+ $X2=4.24 $Y2=2.02
r74 9 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635 $X2=0.75
+ $Y2=2.72
r75 9 11 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2
r76 2 15 300 $w=1.7e-07 $l=6.37652e-07 $layer=licon1_PDIFF $count=2 $X=4.015
+ $Y=1.485 $X2=4.24 $Y2=2.02
r77 1 11 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A_309_297# 1 2 9 11 12 15
r31 13 15 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.22 $Y=2.295
+ $X2=3.22 $Y2=2.135
r32 11 13 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.135 $Y=2.38
+ $X2=3.22 $Y2=2.295
r33 11 12 88.7273 $w=1.68e-07 $l=1.36e-06 $layer=LI1_cond $X=3.135 $Y=2.38
+ $X2=1.775 $Y2=2.38
r34 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.69 $Y=2.295
+ $X2=1.775 $Y2=2.38
r35 7 9 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=1.69 $Y=2.295 $X2=1.69
+ $Y2=2.135
r36 2 15 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=3.075
+ $Y=1.485 $X2=3.22 $Y2=2.135
r37 1 9 600 $w=1.7e-07 $l=7.18853e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=2.135
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%Y 1 2 3 4 13 14 17 21 24 25 26 27 28 29 30
+ 39 45 52 54
r66 52 54 3.38954 $w=3.38e-07 $l=1e-07 $layer=LI1_cond $X=4.795 $Y=1.665
+ $X2=4.795 $Y2=1.765
r67 29 30 11.5244 $w=3.38e-07 $l=3.4e-07 $layer=LI1_cond $X=4.795 $Y=1.87
+ $X2=4.795 $Y2=2.21
r68 29 54 3.55902 $w=3.38e-07 $l=1.05e-07 $layer=LI1_cond $X=4.795 $Y=1.87
+ $X2=4.795 $Y2=1.765
r69 28 52 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.315 $Y=1.58
+ $X2=4.795 $Y2=1.58
r70 28 43 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.315 $Y=1.58
+ $X2=4.265 $Y2=1.58
r71 28 43 0.758186 $w=3.78e-07 $l=2.5e-08 $layer=LI1_cond $X=4.265 $Y=1.47
+ $X2=4.265 $Y2=1.495
r72 27 28 8.49168 $w=3.78e-07 $l=2.8e-07 $layer=LI1_cond $X=4.265 $Y=1.19
+ $X2=4.265 $Y2=1.47
r73 26 27 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=4.265 $Y=0.85
+ $X2=4.265 $Y2=1.19
r74 26 45 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=4.265 $Y=0.85
+ $X2=4.265 $Y2=0.755
r75 25 39 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=2.75 $Y=1.87
+ $X2=2.75 $Y2=1.68
r76 23 39 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.75 $Y=1.665
+ $X2=2.75 $Y2=1.68
r77 22 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=1.58
+ $X2=3.665 $Y2=1.58
r78 21 43 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.075 $Y=1.58
+ $X2=4.265 $Y2=1.58
r79 21 22 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.075 $Y=1.58
+ $X2=3.855 $Y2=1.58
r80 17 19 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.665 $Y=1.68
+ $X2=3.665 $Y2=2.36
r81 15 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=1.665
+ $X2=3.665 $Y2=1.58
r82 15 17 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.665 $Y=1.665
+ $X2=3.665 $Y2=1.68
r83 14 23 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.915 $Y=1.58
+ $X2=2.75 $Y2=1.665
r84 13 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.475 $Y=1.58
+ $X2=3.665 $Y2=1.58
r85 13 14 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.475 $Y=1.58
+ $X2=2.915 $Y2=1.58
r86 4 54 300 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=2 $X=4.605
+ $Y=1.485 $X2=4.75 $Y2=1.765
r87 3 19 400 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=1.485 $X2=3.69 $Y2=2.36
r88 3 17 400 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=1 $X=3.545
+ $Y=1.485 $X2=3.69 $Y2=1.68
r89 2 39 300 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_PDIFF $count=2 $X=2.605
+ $Y=1.485 $X2=2.75 $Y2=1.68
r90 1 45 182 $w=1.7e-07 $l=6.38905e-07 $layer=licon1_NDIFF $count=1 $X=3.975
+ $Y=0.235 $X2=4.24 $Y2=0.755
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%A_27_47# 1 2 3 4 5 18 20 21 24 26 30 32 34
+ 35 36 38 39
c82 34 0 1.21354e-19 $X=3.665 $Y=0.425
r83 37 41 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.855 $Y=0.34
+ $X2=3.665 $Y2=0.34
r84 36 45 2.7521 $w=3.33e-07 $l=8e-08 $layer=LI1_cond $X=4.797 $Y=0.34 $X2=4.797
+ $Y2=0.42
r85 36 37 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=4.63 $Y=0.34
+ $X2=3.855 $Y2=0.34
r86 34 41 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.665 $Y2=0.34
r87 34 35 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=3.665 $Y=0.425
+ $X2=3.665 $Y2=0.715
r88 33 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.755 $Y=0.8
+ $X2=2.59 $Y2=0.8
r89 32 35 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.475 $Y=0.8
+ $X2=3.665 $Y2=0.715
r90 32 33 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=3.475 $Y=0.8
+ $X2=2.755 $Y2=0.8
r91 28 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.59 $Y=0.715
+ $X2=2.59 $Y2=0.8
r92 28 30 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.59 $Y=0.715
+ $X2=2.59 $Y2=0.36
r93 27 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.385 $Y=0.8
+ $X2=1.195 $Y2=0.8
r94 26 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=2.59 $Y2=0.8
r95 26 27 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=2.425 $Y=0.8
+ $X2=1.385 $Y2=0.8
r96 22 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.715
+ $X2=1.195 $Y2=0.8
r97 22 24 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=1.195 $Y=0.715
+ $X2=1.195 $Y2=0.36
r98 20 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.005 $Y=0.8
+ $X2=1.195 $Y2=0.8
r99 20 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.005 $Y=0.8
+ $X2=0.445 $Y2=0.8
r100 16 21 7.97992 $w=1.7e-07 $l=2.16365e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.445 $Y2=0.8
r101 16 18 11.5244 $w=3.53e-07 $l=3.55e-07 $layer=LI1_cond $X=0.267 $Y=0.715
+ $X2=0.267 $Y2=0.36
r102 5 45 182 $w=1.7e-07 $l=2.66927e-07 $layer=licon1_NDIFF $count=1 $X=4.565
+ $Y=0.235 $X2=4.755 $Y2=0.42
r103 4 41 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=3.555
+ $Y=0.235 $X2=3.69 $Y2=0.36
r104 3 30 91 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=2 $X=2.415
+ $Y=0.235 $X2=2.59 $Y2=0.36
r105 2 24 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.36
r106 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__O31AI_2%VGND 1 2 3 14 18 22 24 31 32 35 40 46 48
+ 51
c68 31 0 7.9412e-20 $X=4.83 $Y=0
r69 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r70 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r71 44 46 9.02273 $w=6.28e-07 $l=9.5e-08 $layer=LI1_cond $X=2.07 $Y=0.23
+ $X2=2.165 $Y2=0.23
r72 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 42 44 0.759415 $w=6.28e-07 $l=4e-08 $layer=LI1_cond $X=2.03 $Y=0.23 $X2=2.07
+ $Y2=0.23
r74 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r75 38 42 7.97386 $w=6.28e-07 $l=4.2e-07 $layer=LI1_cond $X=1.61 $Y=0.23
+ $X2=2.03 $Y2=0.23
r76 38 40 7.31405 $w=6.28e-07 $l=5e-09 $layer=LI1_cond $X=1.61 $Y=0.23 $X2=1.605
+ $Y2=0.23
r77 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r78 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r79 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r80 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r81 29 32 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r82 29 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r83 28 31 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.45 $Y=0 $X2=4.83
+ $Y2=0
r84 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r85 26 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.115
+ $Y2=0
r86 26 28 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.305 $Y=0 $X2=3.45
+ $Y2=0
r87 24 36 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r88 24 51 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0 $X2=0.23
+ $Y2=0
r89 20 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0
r90 20 22 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=3.115 $Y=0.085
+ $X2=3.115 $Y2=0.36
r91 18 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=3.115
+ $Y2=0
r92 18 46 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=2.925 $Y=0 $X2=2.165
+ $Y2=0
r93 17 35 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.75
+ $Y2=0
r94 17 40 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=1.605
+ $Y2=0
r95 12 35 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0
r96 12 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r97 3 22 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.935
+ $Y=0.235 $X2=3.14 $Y2=0.36
r98 2 42 91 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=2.03 $Y2=0.38
r99 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.38
.ends

