* File: sky130_fd_sc_hdll__a221oi_1.pxi.spice
* Created: Wed Sep  2 08:18:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__A221OI_1%C1 N_C1_c_58_n N_C1_M1006_g N_C1_c_55_n
+ N_C1_M1008_g C1 N_C1_c_57_n PM_SKY130_FD_SC_HDLL__A221OI_1%C1
x_PM_SKY130_FD_SC_HDLL__A221OI_1%B2 N_B2_c_84_n N_B2_M1000_g N_B2_c_85_n
+ N_B2_M1002_g B2 N_B2_c_86_n B2 PM_SKY130_FD_SC_HDLL__A221OI_1%B2
x_PM_SKY130_FD_SC_HDLL__A221OI_1%B1 N_B1_c_110_n N_B1_M1003_g N_B1_c_111_n
+ N_B1_M1009_g B1 B1 N_B1_c_113_n B1 PM_SKY130_FD_SC_HDLL__A221OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A221OI_1%A1 N_A1_c_147_n N_A1_M1007_g N_A1_c_148_n
+ N_A1_M1005_g A1 A1 N_A1_c_150_n PM_SKY130_FD_SC_HDLL__A221OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A221OI_1%A2 N_A2_c_182_n N_A2_M1001_g N_A2_c_183_n
+ N_A2_M1004_g A2 A2 PM_SKY130_FD_SC_HDLL__A221OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A221OI_1%Y N_Y_M1008_s N_Y_M1003_d N_Y_M1005_s
+ N_Y_M1006_s N_Y_c_223_n N_Y_c_224_n N_Y_c_213_n N_Y_c_214_n N_Y_c_218_n
+ N_Y_c_215_n N_Y_c_248_n N_Y_c_256_n N_Y_c_263_n N_Y_c_264_n N_Y_c_267_n
+ N_Y_c_219_n N_Y_c_220_n Y Y Y N_Y_c_216_n N_Y_c_221_n Y
+ PM_SKY130_FD_SC_HDLL__A221OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A221OI_1%A_117_297# N_A_117_297#_M1006_d
+ N_A_117_297#_M1009_d N_A_117_297#_c_324_n N_A_117_297#_c_325_n
+ N_A_117_297#_c_327_n N_A_117_297#_c_323_n N_A_117_297#_c_326_n
+ PM_SKY130_FD_SC_HDLL__A221OI_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_1%A_211_297# N_A_211_297#_M1000_d
+ N_A_211_297#_M1007_d N_A_211_297#_c_348_n N_A_211_297#_c_351_n
+ N_A_211_297#_c_357_n N_A_211_297#_c_368_p N_A_211_297#_c_358_n
+ N_A_211_297#_c_349_n PM_SKY130_FD_SC_HDLL__A221OI_1%A_211_297#
x_PM_SKY130_FD_SC_HDLL__A221OI_1%VPWR N_VPWR_M1007_s N_VPWR_M1001_d
+ N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n VPWR
+ N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_377_n N_VPWR_c_385_n
+ PM_SKY130_FD_SC_HDLL__A221OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A221OI_1%VGND N_VGND_M1008_d N_VGND_M1004_d
+ N_VGND_c_427_n N_VGND_c_428_n N_VGND_c_429_n N_VGND_c_430_n VGND
+ N_VGND_c_431_n N_VGND_c_432_n N_VGND_c_433_n N_VGND_c_434_n
+ PM_SKY130_FD_SC_HDLL__A221OI_1%VGND
cc_1 VNB N_C1_c_55_n 0.0221052f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB C1 0.00922438f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_3 VNB N_C1_c_57_n 0.0424358f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B2_c_84_n 0.022309f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B2_c_85_n 0.0165758f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B2_c_86_n 0.00681607f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_7 VNB N_B1_c_110_n 0.0186714f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B1_c_111_n 0.026851f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB B1 0.00452296f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_10 VNB N_B1_c_113_n 0.00446396f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_147_n 0.0314769f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_A1_c_148_n 0.0203575f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_13 VNB A1 0.00500472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_150_n 0.00266387f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_15 VNB N_A2_c_182_n 0.0267005f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB N_A2_c_183_n 0.0196504f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_17 VNB A2 0.00594509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_213_n 0.006204f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_214_n 0.0018549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_Y_c_215_n 0.0114766f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_216_n 0.010692f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB Y 0.0253239f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_377_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_427_n 0.0028208f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_25 VNB N_VGND_c_428_n 0.0123943f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_26 VNB N_VGND_c_429_n 0.0493159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_430_n 0.00510247f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_431_n 0.0152294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_432_n 0.0115819f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_433_n 0.207858f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_434_n 0.00574292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VPB N_C1_c_58_n 0.020476f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB N_C1_c_57_n 0.0192397f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_34 VPB N_B2_c_84_n 0.0260529f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_35 VPB N_B1_c_111_n 0.0335055f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_36 VPB N_A1_c_147_n 0.0349005f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB N_A2_c_182_n 0.0302282f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_38 VPB A2 0.00116981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_218_n 0.00228382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_219_n 0.0204715f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_Y_c_220_n 2.05929e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_Y_c_221_n 0.0150917f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB Y 0.0106235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_117_297#_c_323_n 0.0025657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_211_297#_c_348_n 0.00782532f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_46 VPB N_A_211_297#_c_349_n 4.02524e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_378_n 0.00604461f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.202
cc_48 VPB N_VPWR_c_379_n 0.0295145f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_49 VPB N_VPWR_c_380_n 0.0176023f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_VPWR_c_381_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_382_n 0.0514066f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_383_n 0.011849f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_377_n 0.0562988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_385_n 0.00513322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 N_C1_c_58_n N_B2_c_84_n 0.0223835f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_56 N_C1_c_57_n N_B2_c_84_n 0.0271764f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_57 N_C1_c_55_n N_B2_c_85_n 0.0206527f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 C1 N_B2_c_86_n 0.0173048f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_59 N_C1_c_57_n N_B2_c_86_n 0.00180909f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_60 N_C1_c_55_n N_Y_c_223_n 0.00597802f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_61 N_C1_c_58_n N_Y_c_224_n 0.0103066f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_62 N_C1_c_55_n N_Y_c_213_n 0.0144197f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_63 C1 N_Y_c_213_n 0.00646022f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_64 N_C1_c_57_n N_Y_c_213_n 0.00269443f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_65 C1 N_Y_c_214_n 0.0143329f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_66 N_C1_c_57_n N_Y_c_214_n 0.00447564f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_67 C1 N_Y_c_218_n 0.0139774f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_68 N_C1_c_57_n N_Y_c_218_n 0.00415326f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_69 N_C1_c_58_n N_Y_c_219_n 0.0154002f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 C1 N_Y_c_219_n 0.00635212f $X=0.145 $Y=1.105 $X2=0 $Y2=0
cc_71 N_C1_c_57_n N_Y_c_219_n 0.00179908f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_72 N_C1_c_58_n N_A_117_297#_c_324_n 0.00822051f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_73 N_C1_c_58_n N_A_117_297#_c_325_n 0.00305463f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_74 N_C1_c_58_n N_VPWR_c_382_n 0.00596194f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C1_c_58_n N_VPWR_c_377_n 0.0109919f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_76 N_C1_c_55_n N_VGND_c_427_n 0.0129524f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_77 N_C1_c_55_n N_VGND_c_431_n 0.0020416f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_78 N_C1_c_55_n N_VGND_c_433_n 0.00378724f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_79 N_B2_c_85_n N_B1_c_110_n 0.037701f $X=1.05 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_80 N_B2_c_84_n N_B1_c_111_n 0.0799632f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_81 N_B2_c_86_n N_B1_c_111_n 7.29268e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_82 N_B2_c_84_n B1 3.79007e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B2_c_84_n N_B1_c_113_n 6.80936e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B2_c_86_n N_B1_c_113_n 0.0187077f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_85 N_B2_c_84_n N_Y_c_213_n 0.00463168f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B2_c_85_n N_Y_c_213_n 0.0122525f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_87 N_B2_c_86_n N_Y_c_213_n 0.040285f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_88 N_B2_c_84_n N_Y_c_219_n 0.0182032f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B2_c_86_n N_Y_c_219_n 0.0401733f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_90 N_B2_c_84_n N_A_117_297#_c_326_n 0.0115669f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B2_c_84_n N_VPWR_c_382_n 0.00429453f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B2_c_84_n N_VPWR_c_377_n 0.00611639f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B2_c_85_n N_VGND_c_427_n 0.00650448f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_94 N_B2_c_85_n N_VGND_c_429_n 0.00439206f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_95 N_B2_c_85_n N_VGND_c_433_n 0.00622536f $X=1.05 $Y=0.995 $X2=0 $Y2=0
cc_96 N_B1_c_111_n N_A1_c_147_n 0.00839899f $X=1.435 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_97 B1 N_A1_c_147_n 2.25452e-19 $X=1.535 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_98 N_B1_c_113_n N_A1_c_147_n 6.25636e-19 $X=1.67 $Y=1.075 $X2=-0.19 $Y2=-0.24
cc_99 N_B1_c_111_n A1 2.30532e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_100 B1 A1 0.0331978f $X=1.535 $Y=0.765 $X2=0 $Y2=0
cc_101 N_B1_c_111_n N_A1_c_150_n 6.20584e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B1_c_113_n N_A1_c_150_n 0.0183174f $X=1.67 $Y=1.075 $X2=0 $Y2=0
cc_103 B1 N_Y_M1003_d 0.00457458f $X=1.535 $Y=0.765 $X2=0 $Y2=0
cc_104 N_B1_c_110_n N_Y_c_213_n 0.00144078f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_105 B1 N_Y_c_213_n 0.00726661f $X=1.535 $Y=0.765 $X2=0 $Y2=0
cc_106 N_B1_c_113_n N_Y_c_213_n 8.53788e-19 $X=1.67 $Y=1.075 $X2=0 $Y2=0
cc_107 N_B1_c_110_n N_Y_c_215_n 0.0087337f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B1_c_111_n N_Y_c_215_n 5.39066e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_109 B1 N_Y_c_215_n 0.020856f $X=1.535 $Y=0.765 $X2=0 $Y2=0
cc_110 N_B1_c_113_n N_Y_c_215_n 0.00446876f $X=1.67 $Y=1.075 $X2=0 $Y2=0
cc_111 N_B1_c_110_n N_Y_c_248_n 0.00151997f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_112 N_B1_c_111_n N_Y_c_219_n 0.0178525f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_113_n N_Y_c_219_n 0.0354842f $X=1.67 $Y=1.075 $X2=0 $Y2=0
cc_114 N_B1_c_111_n N_A_117_297#_c_327_n 0.00365738f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_115 N_B1_c_111_n N_A_117_297#_c_326_n 0.00652054f $X=1.435 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_B1_c_111_n N_A_211_297#_c_348_n 0.0155679f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_117 N_B1_c_111_n N_VPWR_c_378_n 0.00234693f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B1_c_111_n N_VPWR_c_382_n 0.00429453f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B1_c_111_n N_VPWR_c_377_n 0.00737353f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_110_n N_VGND_c_429_n 0.00357877f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_110_n N_VGND_c_433_n 0.00641668f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A1_c_147_n N_A2_c_182_n 0.0528384f $X=2.425 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_123 N_A1_c_150_n N_A2_c_182_n 2.02422e-19 $X=2.26 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_124 N_A1_c_148_n N_A2_c_183_n 0.0253675f $X=2.45 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A1_c_147_n A2 0.00317888f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_126 A1 A2 0.00398621f $X=2.035 $Y=0.765 $X2=0 $Y2=0
cc_127 N_A1_c_150_n A2 0.0131758f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_128 A1 N_Y_M1005_s 0.00460924f $X=2.035 $Y=0.765 $X2=0 $Y2=0
cc_129 N_A1_c_147_n N_Y_c_215_n 7.73318e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A1_c_148_n N_Y_c_215_n 0.0136475f $X=2.45 $Y=0.995 $X2=0 $Y2=0
cc_131 A1 N_Y_c_215_n 0.0264394f $X=2.035 $Y=0.765 $X2=0 $Y2=0
cc_132 N_A1_c_150_n N_Y_c_215_n 0.00159807f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A1_c_147_n N_Y_c_256_n 0.00706514f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A1_c_147_n N_Y_c_219_n 0.00469821f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_150_n N_Y_c_219_n 0.0346364f $X=2.26 $Y=1.16 $X2=0 $Y2=0
cc_136 N_A1_c_147_n N_Y_c_220_n 0.0118577f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A1_c_147_n N_A_211_297#_c_351_n 0.015093f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_147_n N_A_211_297#_c_349_n 0.00164897f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A1_c_147_n N_VPWR_c_378_n 0.00938435f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A1_c_147_n N_VPWR_c_380_n 0.00458874f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A1_c_147_n N_VPWR_c_377_n 0.00540268f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A1_c_148_n N_VGND_c_428_n 0.00116008f $X=2.45 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A1_c_148_n N_VGND_c_429_n 0.00357877f $X=2.45 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A1_c_148_n N_VGND_c_433_n 0.00683557f $X=2.45 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A2_c_183_n N_Y_c_215_n 0.00279221f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A2_c_182_n N_Y_c_256_n 0.0219746f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_147 A2 N_Y_c_256_n 0.0266579f $X=2.955 $Y=1.19 $X2=0 $Y2=0
cc_148 N_A2_c_183_n N_Y_c_263_n 0.00351199f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_182_n N_Y_c_264_n 0.00284378f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A2_c_183_n N_Y_c_264_n 0.0136059f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_151 A2 N_Y_c_264_n 0.018668f $X=2.955 $Y=1.19 $X2=0 $Y2=0
cc_152 N_A2_c_182_n N_Y_c_267_n 0.00104119f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_153 A2 N_Y_c_267_n 0.0092235f $X=2.955 $Y=1.19 $X2=0 $Y2=0
cc_154 N_A2_c_182_n N_Y_c_220_n 2.0783e-19 $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A2_c_182_n Y 0.00835417f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A2_c_183_n Y 0.00598562f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_157 A2 Y 0.0264328f $X=2.955 $Y=1.19 $X2=0 $Y2=0
cc_158 N_A2_c_182_n N_VPWR_c_378_n 0.00102791f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A2_c_182_n N_VPWR_c_379_n 0.00501204f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A2_c_182_n N_VPWR_c_380_n 0.00700684f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_161 N_A2_c_182_n N_VPWR_c_377_n 0.0136557f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A2_c_183_n N_VGND_c_428_n 0.00935634f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A2_c_183_n N_VGND_c_429_n 0.00355956f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A2_c_183_n N_VGND_c_433_n 0.0044548f $X=2.98 $Y=0.995 $X2=0 $Y2=0
cc_165 N_Y_c_219_n N_A_117_297#_M1006_d 0.00182839f $X=2.3 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_166 N_Y_c_219_n N_A_117_297#_M1009_d 0.00296218f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_167 N_Y_c_224_n N_A_117_297#_c_324_n 0.0366092f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_168 N_Y_c_219_n N_A_117_297#_c_324_n 0.0191842f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_169 N_Y_c_224_n N_A_117_297#_c_325_n 0.0133617f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_170 N_Y_c_219_n N_A_117_297#_c_326_n 0.00398242f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_171 N_Y_c_219_n N_A_211_297#_M1000_d 0.00184351f $X=2.3 $Y=1.56 $X2=-0.19
+ $Y2=-0.24
cc_172 N_Y_c_256_n N_A_211_297#_M1007_d 0.00588744f $X=3.255 $Y=1.58 $X2=0 $Y2=0
cc_173 N_Y_c_219_n N_A_211_297#_c_351_n 0.00646916f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_174 N_Y_c_220_n N_A_211_297#_c_351_n 0.0125708f $X=2.45 $Y=1.56 $X2=0 $Y2=0
cc_175 N_Y_c_256_n N_A_211_297#_c_357_n 0.0188393f $X=3.255 $Y=1.58 $X2=0 $Y2=0
cc_176 N_Y_c_219_n N_A_211_297#_c_358_n 0.0708204f $X=2.3 $Y=1.56 $X2=0 $Y2=0
cc_177 N_Y_c_219_n N_VPWR_M1007_s 0.00306703f $X=2.3 $Y=1.56 $X2=-0.19 $Y2=-0.24
cc_178 N_Y_c_256_n N_VPWR_M1001_d 0.00508168f $X=3.255 $Y=1.58 $X2=0 $Y2=0
cc_179 N_Y_c_221_n N_VPWR_M1001_d 0.00171163f $X=3.395 $Y=1.495 $X2=0 $Y2=0
cc_180 N_Y_c_256_n N_VPWR_c_379_n 0.0106054f $X=3.255 $Y=1.58 $X2=0 $Y2=0
cc_181 N_Y_c_221_n N_VPWR_c_379_n 0.00926531f $X=3.395 $Y=1.495 $X2=0 $Y2=0
cc_182 N_Y_c_224_n N_VPWR_c_382_n 0.0118139f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_183 N_Y_M1006_s N_VPWR_c_377_n 0.00568146f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_184 N_Y_c_224_n N_VPWR_c_377_n 0.00646998f $X=0.26 $Y=1.65 $X2=0 $Y2=0
cc_185 N_Y_c_213_n N_VGND_M1008_d 0.003124f $X=1.165 $Y=0.82 $X2=-0.19 $Y2=-0.24
cc_186 N_Y_c_264_n N_VGND_M1004_d 0.00447954f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_187 N_Y_c_216_n N_VGND_M1004_d 0.00170795f $X=3.395 $Y=0.825 $X2=0 $Y2=0
cc_188 Y N_VGND_M1004_d 0.00101661f $X=3.355 $Y=0.85 $X2=0 $Y2=0
cc_189 N_Y_c_223_n N_VGND_c_427_n 0.0231923f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_190 N_Y_c_213_n N_VGND_c_427_n 0.0247522f $X=1.165 $Y=0.82 $X2=0 $Y2=0
cc_191 N_Y_c_215_n N_VGND_c_428_n 0.0141175f $X=2.58 $Y=0.38 $X2=0 $Y2=0
cc_192 N_Y_c_264_n N_VGND_c_428_n 0.0126282f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_193 N_Y_c_216_n N_VGND_c_428_n 0.00888209f $X=3.395 $Y=0.825 $X2=0 $Y2=0
cc_194 N_Y_c_213_n N_VGND_c_429_n 0.00301812f $X=1.165 $Y=0.82 $X2=0 $Y2=0
cc_195 N_Y_c_215_n N_VGND_c_429_n 0.0894211f $X=2.58 $Y=0.38 $X2=0 $Y2=0
cc_196 N_Y_c_248_n N_VGND_c_429_n 0.00935408f $X=1.335 $Y=0.38 $X2=0 $Y2=0
cc_197 N_Y_c_264_n N_VGND_c_429_n 0.00360532f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_198 N_Y_c_223_n N_VGND_c_431_n 0.0121253f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_199 N_Y_c_213_n N_VGND_c_431_n 0.00193889f $X=1.165 $Y=0.82 $X2=0 $Y2=0
cc_200 N_Y_c_216_n N_VGND_c_432_n 0.00340165f $X=3.395 $Y=0.825 $X2=0 $Y2=0
cc_201 N_Y_M1008_s N_VGND_c_433_n 0.00429029f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_202 N_Y_M1003_d N_VGND_c_433_n 0.00250339f $X=1.485 $Y=0.235 $X2=0 $Y2=0
cc_203 N_Y_M1005_s N_VGND_c_433_n 0.00250339f $X=2.065 $Y=0.235 $X2=0 $Y2=0
cc_204 N_Y_c_223_n N_VGND_c_433_n 0.00665463f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_205 N_Y_c_213_n N_VGND_c_433_n 0.0118775f $X=1.165 $Y=0.82 $X2=0 $Y2=0
cc_206 N_Y_c_215_n N_VGND_c_433_n 0.0529023f $X=2.58 $Y=0.38 $X2=0 $Y2=0
cc_207 N_Y_c_248_n N_VGND_c_433_n 0.00653924f $X=1.335 $Y=0.38 $X2=0 $Y2=0
cc_208 N_Y_c_264_n N_VGND_c_433_n 0.0073263f $X=3.255 $Y=0.74 $X2=0 $Y2=0
cc_209 N_Y_c_216_n N_VGND_c_433_n 0.0057408f $X=3.395 $Y=0.825 $X2=0 $Y2=0
cc_210 N_Y_c_248_n A_225_47# 9.37539e-19 $X=1.335 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_211 N_Y_c_215_n A_505_47# 0.00544883f $X=2.58 $Y=0.38 $X2=-0.19 $Y2=-0.24
cc_212 N_Y_c_263_n A_505_47# 0.00186816f $X=2.68 $Y=0.655 $X2=-0.19 $Y2=-0.24
cc_213 N_Y_c_264_n A_505_47# 0.00175614f $X=3.255 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_214 N_Y_c_267_n A_505_47# 0.00394575f $X=2.78 $Y=0.74 $X2=-0.19 $Y2=-0.24
cc_215 N_A_117_297#_c_326_n N_A_211_297#_M1000_d 0.00349652f $X=1.455 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_216 N_A_117_297#_M1009_d N_A_211_297#_c_348_n 0.00583435f $X=1.525 $Y=1.485
+ $X2=0 $Y2=0
cc_217 N_A_117_297#_c_327_n N_A_211_297#_c_348_n 0.0192438f $X=1.56 $Y=2.36
+ $X2=0 $Y2=0
cc_218 N_A_117_297#_c_326_n N_A_211_297#_c_348_n 0.00504187f $X=1.455 $Y=2.36
+ $X2=0 $Y2=0
cc_219 N_A_117_297#_c_324_n N_A_211_297#_c_358_n 0.0178745f $X=0.73 $Y=1.96
+ $X2=0 $Y2=0
cc_220 N_A_117_297#_c_326_n N_A_211_297#_c_358_n 0.0124153f $X=1.455 $Y=2.36
+ $X2=0 $Y2=0
cc_221 N_A_117_297#_c_323_n N_VPWR_c_378_n 0.0168662f $X=1.67 $Y=2.34 $X2=0
+ $Y2=0
cc_222 N_A_117_297#_c_325_n N_VPWR_c_382_n 0.0188769f $X=0.815 $Y=2.38 $X2=0
+ $Y2=0
cc_223 N_A_117_297#_c_326_n N_VPWR_c_382_n 0.0577415f $X=1.455 $Y=2.36 $X2=0
+ $Y2=0
cc_224 N_A_117_297#_M1006_d N_VPWR_c_377_n 0.00231266f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_225 N_A_117_297#_M1009_d N_VPWR_c_377_n 0.00217543f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_226 N_A_117_297#_c_325_n N_VPWR_c_377_n 0.0111519f $X=0.815 $Y=2.38 $X2=0
+ $Y2=0
cc_227 N_A_117_297#_c_326_n N_VPWR_c_377_n 0.0362574f $X=1.455 $Y=2.36 $X2=0
+ $Y2=0
cc_228 N_A_211_297#_c_351_n N_VPWR_M1007_s 0.00211943f $X=2.575 $Y=1.94
+ $X2=-0.19 $Y2=1.305
cc_229 N_A_211_297#_c_349_n N_VPWR_M1007_s 0.00403427f $X=2.175 $Y=1.92
+ $X2=-0.19 $Y2=1.305
cc_230 N_A_211_297#_c_348_n N_VPWR_c_378_n 0.0212636f $X=2.05 $Y=1.92 $X2=0
+ $Y2=0
cc_231 N_A_211_297#_c_368_p N_VPWR_c_378_n 0.0155816f $X=2.66 $Y=2.3 $X2=0 $Y2=0
cc_232 N_A_211_297#_c_351_n N_VPWR_c_380_n 0.00293617f $X=2.575 $Y=1.94 $X2=0
+ $Y2=0
cc_233 N_A_211_297#_c_368_p N_VPWR_c_380_n 0.0167911f $X=2.66 $Y=2.3 $X2=0 $Y2=0
cc_234 N_A_211_297#_c_348_n N_VPWR_c_382_n 0.00327883f $X=2.05 $Y=1.92 $X2=0
+ $Y2=0
cc_235 N_A_211_297#_M1000_d N_VPWR_c_377_n 0.00232895f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_A_211_297#_M1007_d N_VPWR_c_377_n 0.00446736f $X=2.515 $Y=1.485 $X2=0
+ $Y2=0
cc_237 N_A_211_297#_c_348_n N_VPWR_c_377_n 0.00785752f $X=2.05 $Y=1.92 $X2=0
+ $Y2=0
cc_238 N_A_211_297#_c_351_n N_VPWR_c_377_n 0.00525741f $X=2.575 $Y=1.94 $X2=0
+ $Y2=0
cc_239 N_A_211_297#_c_368_p N_VPWR_c_377_n 0.0095318f $X=2.66 $Y=2.3 $X2=0 $Y2=0
cc_240 N_VGND_c_433_n A_225_47# 0.0018911f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
cc_241 N_VGND_c_433_n A_505_47# 0.00354367f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
