* File: sky130_fd_sc_hdll__muxb4to1_1.pex.spice
* Created: Thu Aug 27 19:11:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[0] 1 3 4 6 8 13 15
c28 4 0 5.33021e-20 $X=0.495 $Y=1.41
r29 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=0.69 $Y=0.51
+ $X2=0.645 $Y2=0.51
r30 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=0.5 $Y=1.19
+ $X2=0.645 $Y2=1.19
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.5
+ $Y=1.16 $X2=0.5 $Y2=1.16
r32 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.645 $Y=1.055
+ $X2=0.645 $Y2=1.19
r33 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=0.51
r34 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=0.645 $Y=0.625
+ $X2=0.645 $Y2=1.055
r35 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.5 $Y2=1.16
r36 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r37 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.5 $Y2=1.16
r38 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995 $X2=0.47
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_184_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=1.545 $Y=1.405
+ $X2=1.775 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=1.325 $Y=1.34
+ $X2=1.02 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=1.325 $Y=1.405
+ $X2=1.545 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.325
+ $Y=1.34 $X2=1.325 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=1.775 $Y=2.31
+ $X2=1.775 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=1.545 $Y=1.175
+ $X2=1.545 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.775 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=1.545 $Y=0.755
+ $X2=1.545 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.02 $Y=1.475
+ $X2=1.02 $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.02 $Y=1.475 $X2=1.02
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.65
+ $Y=1.485 $X2=1.775 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=1.65
+ $Y=0.235 $X2=1.775 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[0] 1 3 4 5 6 8 9 11 12 17
r46 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.975
+ $Y=1.03 $X2=1.975 $Y2=1.03
r47 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=1.975 $Y=0.905
+ $X2=1.975 $Y2=1.03
r48 12 17 5.26831 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=1.98 $Y=1.19
+ $X2=1.98 $Y2=1.03
r49 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=1.975 $Y2=0.905
r50 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.01 $Y=0.83
+ $X2=2.01 $Y2=0.495
r51 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.01 $Y=1.41
+ $X2=1.975 $Y2=1.03
r52 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.01 $Y=1.41 $X2=2.01
+ $Y2=1.985
r53 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.84 $Y=0.905
+ $X2=1.975 $Y2=0.905
r54 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=1.84 $Y=0.905 $X2=1.02
+ $Y2=0.905
r55 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=1.02 $Y2=0.905
r56 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=0.945 $Y=0.83
+ $X2=0.945 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[1] 1 3 4 6 7 9 11 12 17
r44 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.625
+ $Y=1.03 $X2=2.625 $Y2=1.03
r45 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=2.625 $Y=0.905
+ $X2=2.625 $Y2=1.03
r46 12 17 5.26831 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=2.62 $Y=1.19
+ $X2=2.62 $Y2=1.03
r47 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.655 $Y=0.83
+ $X2=3.655 $Y2=0.495
r48 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.76 $Y=0.905
+ $X2=2.625 $Y2=0.905
r49 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.58 $Y=0.905
+ $X2=3.655 $Y2=0.83
r50 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=3.58 $Y=0.905 $X2=2.76
+ $Y2=0.905
r51 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=2.59 $Y=0.83
+ $X2=2.625 $Y2=0.905
r52 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.59 $Y=0.83 $X2=2.59
+ $Y2=0.495
r53 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=2.59 $Y=1.41
+ $X2=2.625 $Y2=1.03
r54 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.59 $Y=1.41 $X2=2.59
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_533_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=3.275 $Y=1.34
+ $X2=3.58 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.275
+ $Y=1.34 $X2=3.275 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=3.055 $Y=1.405
+ $X2=3.275 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=2.825 $Y=1.63
+ $X2=3.055 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.055 $Y=1.175
+ $X2=3.055 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=2.825 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=3.055 $Y=0.755
+ $X2=3.055 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.825 $Y=2.31
+ $X2=2.825 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=3.58 $Y=1.475
+ $X2=3.58 $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=3.58 $Y=1.475 $X2=3.58
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.68
+ $Y=1.485 $X2=2.825 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=2.665
+ $Y=0.235 $X2=2.825 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[1] 1 3 4 6 8 12 15 21
c37 8 0 1.78369e-19 $X=3.955 $Y=1.055
c38 1 0 2.31671e-19 $X=4.105 $Y=1.41
r39 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=3.91 $Y=0.51
+ $X2=3.955 $Y2=0.51
r40 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.1
+ $Y=1.16 $X2=4.1 $Y2=1.16
r41 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.955 $Y=1.19
+ $X2=4.1 $Y2=1.19
r42 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.955 $Y=1.055
+ $X2=3.955 $Y2=1.19
r43 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.955 $Y=0.625
+ $X2=3.955 $Y2=1.055
r45 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.13 $Y=0.995
+ $X2=4.1 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.13 $Y=0.995 $X2=4.13
+ $Y2=0.56
r47 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.1 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.105 $Y=1.41
+ $X2=4.105 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[2] 1 3 4 6 8 13 15
c37 8 0 1.78369e-19 $X=4.785 $Y=1.055
c38 4 0 2.31671e-19 $X=4.635 $Y=1.41
r39 15 18 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=4.83 $Y=0.51
+ $X2=4.785 $Y2=0.51
r40 10 13 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.64 $Y=1.19
+ $X2=4.785 $Y2=1.19
r41 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.64
+ $Y=1.16 $X2=4.64 $Y2=1.16
r42 8 13 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.785 $Y=1.055
+ $X2=4.785 $Y2=1.19
r43 7 18 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=0.51
r44 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=4.785 $Y=0.625
+ $X2=4.785 $Y2=1.055
r45 4 11 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.64 $Y2=1.16
r46 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.635 $Y=1.41
+ $X2=4.635 $Y2=1.985
r47 1 11 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=4.61 $Y=0.995
+ $X2=4.64 $Y2=1.16
r48 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.61 $Y=0.995 $X2=4.61
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1012_265# 1 2 9 11 12 15 22 26
r56 20 22 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=5.685 $Y=1.405
+ $X2=5.915 $Y2=1.63
r57 19 26 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=5.465 $Y=1.34
+ $X2=5.16 $Y2=1.34
r58 18 20 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=5.465 $Y=1.405
+ $X2=5.685 $Y2=1.405
r59 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.465
+ $Y=1.34 $X2=5.465 $Y2=1.34
r60 15 22 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.915 $Y=2.31
+ $X2=5.915 $Y2=1.635
r61 12 20 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=5.685 $Y=1.175
+ $X2=5.685 $Y2=1.405
r62 11 25 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.915 $Y2=0.542
r63 11 12 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=5.685 $Y=0.755
+ $X2=5.685 $Y2=1.175
r64 7 26 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.16 $Y=1.475
+ $X2=5.16 $Y2=1.34
r65 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=5.16 $Y=1.475 $X2=5.16
+ $Y2=2.075
r66 2 22 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=1.63
r67 2 15 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=5.79
+ $Y=1.485 $X2=5.915 $Y2=2.31
r68 1 25 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=5.79
+ $Y=0.235 $X2=5.915 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[2] 1 3 4 5 6 8 9 11 12 17
r47 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.115
+ $Y=1.03 $X2=6.115 $Y2=1.03
r48 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.115 $Y=0.905
+ $X2=6.115 $Y2=1.03
r49 12 17 5.26831 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=6.12 $Y=1.19
+ $X2=6.12 $Y2=1.03
r50 9 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.115 $Y2=0.905
r51 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.15 $Y=0.83
+ $X2=6.15 $Y2=0.495
r52 6 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.15 $Y=1.41
+ $X2=6.115 $Y2=1.03
r53 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.15 $Y=1.41 $X2=6.15
+ $Y2=1.985
r54 4 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.98 $Y=0.905
+ $X2=6.115 $Y2=0.905
r55 4 5 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=5.98 $Y=0.905 $X2=5.16
+ $Y2=0.905
r56 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.16 $Y2=0.905
r57 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=5.085 $Y=0.83
+ $X2=5.085 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%S[3] 1 3 4 6 7 9 11 12 17
r43 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.765
+ $Y=1.03 $X2=6.765 $Y2=1.03
r44 14 16 24.8967 $w=2.42e-07 $l=1.25e-07 $layer=POLY_cond $X=6.765 $Y=0.905
+ $X2=6.765 $Y2=1.03
r45 12 17 5.26831 $w=3.48e-07 $l=1.6e-07 $layer=LI1_cond $X=6.76 $Y=1.19
+ $X2=6.76 $Y2=1.03
r46 9 11 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=7.795 $Y=0.83
+ $X2=7.795 $Y2=0.495
r47 8 14 13.9682 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.9 $Y=0.905
+ $X2=6.765 $Y2=0.905
r48 7 9 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.72 $Y=0.905
+ $X2=7.795 $Y2=0.83
r49 7 8 420.468 $w=1.5e-07 $l=8.2e-07 $layer=POLY_cond $X=7.72 $Y=0.905 $X2=6.9
+ $Y2=0.905
r50 4 14 21.8618 $w=2.42e-07 $l=9.08295e-08 $layer=POLY_cond $X=6.73 $Y=0.83
+ $X2=6.765 $Y2=0.905
r51 4 6 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=6.73 $Y=0.83 $X2=6.73
+ $Y2=0.495
r52 1 16 78.9522 $w=2.42e-07 $l=3.97115e-07 $layer=POLY_cond $X=6.73 $Y=1.41
+ $X2=6.765 $Y2=1.03
r53 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.73 $Y=1.41 $X2=6.73
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%A_1361_47# 1 2 9 13 16 19 22 24
r55 22 27 67.1279 $w=2.19e-07 $l=3.05e-07 $layer=POLY_cond $X=7.415 $Y=1.34
+ $X2=7.72 $Y2=1.34
r56 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.415
+ $Y=1.34 $X2=7.415 $Y2=1.34
r57 19 21 9.25517 $w=2.9e-07 $l=2.2e-07 $layer=LI1_cond $X=7.195 $Y=1.405
+ $X2=7.415 $Y2=1.405
r58 18 19 9.67586 $w=2.9e-07 $l=3.23497e-07 $layer=LI1_cond $X=6.965 $Y=1.63
+ $X2=7.195 $Y2=1.405
r59 16 19 3.86198 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=7.195 $Y=1.175
+ $X2=7.195 $Y2=1.405
r60 15 24 8.93631 $w=3.14e-07 $l=3.19202e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=6.965 $Y2=0.542
r61 15 16 27.4011 $w=1.68e-07 $l=4.2e-07 $layer=LI1_cond $X=7.195 $Y=0.755
+ $X2=7.195 $Y2=1.175
r62 13 18 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.965 $Y=2.31
+ $X2=6.965 $Y2=1.635
r63 7 27 7.45852 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.72 $Y=1.475
+ $X2=7.72 $Y2=1.34
r64 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.72 $Y=1.475 $X2=7.72
+ $Y2=2.075
r65 2 18 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=1.63
r66 2 13 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.82
+ $Y=1.485 $X2=6.965 $Y2=2.31
r67 1 24 182 $w=1.7e-07 $l=3.30454e-07 $layer=licon1_NDIFF $count=1 $X=6.805
+ $Y=0.235 $X2=6.965 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%D[3] 1 3 4 6 8 12 15 21
c28 1 0 5.33021e-20 $X=8.245 $Y=1.41
r29 15 21 2.25478 $w=2.28e-07 $l=4.5e-08 $layer=LI1_cond $X=8.05 $Y=0.51
+ $X2=8.095 $Y2=0.51
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.24
+ $Y=1.16 $X2=8.24 $Y2=1.16
r31 9 12 6.18905 $w=2.68e-07 $l=1.45e-07 $layer=LI1_cond $X=8.095 $Y=1.19
+ $X2=8.24 $Y2=1.19
r32 8 9 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.095 $Y=1.055
+ $X2=8.095 $Y2=1.19
r33 7 21 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=0.51
r34 7 8 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=8.095 $Y=0.625
+ $X2=8.095 $Y2=1.055
r35 4 13 39.2931 $w=2.55e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.27 $Y=0.995
+ $X2=8.24 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.27 $Y=0.995 $X2=8.27
+ $Y2=0.56
r37 1 13 51.486 $w=2.55e-07 $l=2.52488e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.24 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.245 $Y=1.41
+ $X2=8.245 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VPWR 1 2 3 4 5 16 18 24 30 36 40 42 47
+ 48 50 51 52 61 75 86 90
r131 89 90 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r132 86 87 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r133 81 90 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.51 $Y2=2.72
r134 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r135 78 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r136 77 80 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.05 $Y2=2.72
r137 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r138 75 89 4.78613 $w=1.7e-07 $l=2.12e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.527 $Y2=2.72
r139 75 80 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=8.315 $Y=2.72
+ $X2=8.05 $Y2=2.72
r140 74 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r141 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r142 71 74 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r143 71 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r144 70 73 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r145 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r146 68 86 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.37 $Y2=2.72
r147 68 70 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.565 $Y=2.72
+ $X2=4.83 $Y2=2.72
r148 67 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r149 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r150 64 67 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r151 63 66 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r152 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r153 61 86 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=4.37 $Y2=2.72
r154 61 66 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.175 $Y=2.72
+ $X2=3.91 $Y2=2.72
r155 60 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r156 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r157 57 60 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r158 56 59 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r160 54 83 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r161 54 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.69 $Y2=2.72
r162 52 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r163 52 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r164 50 73 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.21 $Y2=2.72
r165 50 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.275 $Y=2.72
+ $X2=6.425 $Y2=2.72
r166 49 77 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.67 $Y2=2.72
r167 49 51 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.575 $Y=2.72
+ $X2=6.425 $Y2=2.72
r168 47 59 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.07 $Y2=2.72
r169 47 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.165 $Y=2.72
+ $X2=2.315 $Y2=2.72
r170 46 63 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.53 $Y2=2.72
r171 46 48 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.315 $Y2=2.72
r172 42 45 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=8.48 $Y=1.66
+ $X2=8.48 $Y2=2.34
r173 40 89 2.98004 $w=3.3e-07 $l=1.05924e-07 $layer=LI1_cond $X=8.48 $Y=2.635
+ $X2=8.527 $Y2=2.72
r174 40 45 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=8.48 $Y=2.635
+ $X2=8.48 $Y2=2.34
r175 36 39 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=6.425 $Y=1.63
+ $X2=6.425 $Y2=2.31
r176 34 51 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.425 $Y=2.635
+ $X2=6.425 $Y2=2.72
r177 34 39 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=6.425 $Y=2.635
+ $X2=6.425 $Y2=2.31
r178 30 33 20.0939 $w=3.88e-07 $l=6.8e-07 $layer=LI1_cond $X=4.37 $Y=1.66
+ $X2=4.37 $Y2=2.34
r179 28 86 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.72
r180 28 33 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=2.635
+ $X2=4.37 $Y2=2.34
r181 24 27 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=2.315 $Y=1.63
+ $X2=2.315 $Y2=2.31
r182 22 48 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=2.72
r183 22 27 12.4848 $w=2.98e-07 $l=3.25e-07 $layer=LI1_cond $X=2.315 $Y=2.635
+ $X2=2.315 $Y2=2.31
r184 18 21 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r185 16 83 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.212 $Y2=2.72
r186 16 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r187 5 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.48 $Y2=2.34
r188 5 42 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=8.335
+ $Y=1.485 $X2=8.48 $Y2=1.66
r189 4 39 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=2.31
r190 4 36 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=6.24
+ $Y=1.485 $X2=6.44 $Y2=1.63
r191 3 33 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=2.34
r192 3 30 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=4.195
+ $Y=1.485 $X2=4.37 $Y2=1.66
r193 2 27 400 $w=1.7e-07 $l=9.19579e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=2.31
r194 2 24 400 $w=1.7e-07 $l=2.62678e-07 $layer=licon1_PDIFF $count=1 $X=2.1
+ $Y=1.485 $X2=2.3 $Y2=1.63
r195 1 21 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r196 1 18 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%Z 1 2 3 4 5 6 7 8 26 27 29 33 37 41 44
+ 46 47 49 53 57 61 64 71 79 81 82 83 84 85 86 89 92 94 95 97 101
c230 79 0 5.33021e-20 $X=7.755 $Y=0.92
c231 71 0 5.33021e-20 $X=3.615 $Y=0.92
c232 47 0 5.33021e-20 $X=5.307 $Y=0.835
c233 27 0 5.33021e-20 $X=1.167 $Y=0.835
r234 99 101 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=0.985 $Y=1.87
+ $X2=1.15 $Y2=1.87
r235 97 101 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=1.87
+ $X2=1.15 $Y2=1.87
r236 95 112 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=7.59 $Y=1.87
+ $X2=7.755 $Y2=1.87
r237 94 95 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=1.87
+ $X2=7.59 $Y2=1.87
r238 92 107 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=5.29 $Y=1.87
+ $X2=5.125 $Y2=1.87
r239 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=1.87
+ $X2=5.29 $Y2=1.87
r240 89 106 9.2765 $w=2.17e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=1.87
+ $X2=3.615 $Y2=1.87
r241 88 89 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=1.87
+ $X2=3.45 $Y2=1.87
r242 86 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.435 $Y=1.87
+ $X2=5.29 $Y2=1.87
r243 85 94 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=7.59 $Y2=1.87
r244 85 86 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=7.445 $Y=1.87
+ $X2=5.435 $Y2=1.87
r245 84 88 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.595 $Y=1.87
+ $X2=3.45 $Y2=1.87
r246 83 91 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=5.29 $Y2=1.87
r247 83 84 1.91831 $w=1.4e-07 $l=1.55e-06 $layer=MET1_cond $X=5.145 $Y=1.87
+ $X2=3.595 $Y2=1.87
r248 82 97 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.295 $Y=1.87
+ $X2=1.15 $Y2=1.87
r249 81 88 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=3.45 $Y2=1.87
r250 81 82 2.48762 $w=1.4e-07 $l=2.01e-06 $layer=MET1_cond $X=3.305 $Y=1.87
+ $X2=1.295 $Y2=1.87
r251 64 112 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=7.755 $Y=1.755
+ $X2=7.755 $Y2=1.87
r252 63 79 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=0.92
r253 63 64 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=7.755 $Y=1.005
+ $X2=7.755 $Y2=1.755
r254 59 79 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=7.572 $Y=0.92
+ $X2=7.755 $Y2=0.92
r255 59 61 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=7.572 $Y=0.835
+ $X2=7.572 $Y2=0.495
r256 55 95 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=7.485 $Y=1.87
+ $X2=7.59 $Y2=1.87
r257 55 57 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=7.485 $Y=1.985
+ $X2=7.485 $Y2=2
r258 51 92 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=5.395 $Y=1.87
+ $X2=5.29 $Y2=1.87
r259 51 53 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=5.395 $Y=1.985
+ $X2=5.395 $Y2=2
r260 47 73 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=5.307 $Y=0.92
+ $X2=5.125 $Y2=0.92
r261 47 49 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=5.307 $Y=0.835
+ $X2=5.307 $Y2=0.495
r262 46 107 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=5.125 $Y=1.755
+ $X2=5.125 $Y2=1.87
r263 45 73 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=0.92
r264 45 46 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.125 $Y=1.005
+ $X2=5.125 $Y2=1.755
r265 44 106 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.615 $Y=1.755
+ $X2=3.615 $Y2=1.87
r266 43 71 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=0.92
r267 43 44 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=3.615 $Y=1.005
+ $X2=3.615 $Y2=1.755
r268 39 71 11.939 $w=1.68e-07 $l=1.83e-07 $layer=LI1_cond $X=3.432 $Y=0.92
+ $X2=3.615 $Y2=0.92
r269 39 41 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=3.432 $Y=0.835
+ $X2=3.432 $Y2=0.495
r270 35 89 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=1.87
+ $X2=3.45 $Y2=1.87
r271 35 37 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=3.345 $Y=1.985
+ $X2=3.345 $Y2=2
r272 31 101 5.90323 $w=2.17e-07 $l=1.05e-07 $layer=LI1_cond $X=1.255 $Y=1.87
+ $X2=1.15 $Y2=1.87
r273 31 33 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.255 $Y=1.985
+ $X2=1.255 $Y2=2
r274 27 65 11.8738 $w=1.68e-07 $l=1.82e-07 $layer=LI1_cond $X=1.167 $Y=0.92
+ $X2=0.985 $Y2=0.92
r275 27 29 15.9931 $w=2.43e-07 $l=3.4e-07 $layer=LI1_cond $X=1.167 $Y=0.835
+ $X2=1.167 $Y2=0.495
r276 26 99 2.16928 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.985 $Y=1.755
+ $X2=0.985 $Y2=1.87
r277 25 65 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=0.92
r278 25 26 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=0.985 $Y=1.005
+ $X2=0.985 $Y2=1.755
r279 8 57 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=7.36
+ $Y=1.665 $X2=7.485 $Y2=2
r280 7 53 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=5.25
+ $Y=1.665 $X2=5.395 $Y2=2
r281 6 37 300 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_PDIFF $count=2 $X=3.22
+ $Y=1.665 $X2=3.345 $Y2=2
r282 5 33 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.665 $X2=1.255 $Y2=2
r283 4 61 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.585 $Y2=0.495
r284 3 49 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=5.16
+ $Y=0.235 $X2=5.295 $Y2=0.495
r285 2 41 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=3.32
+ $Y=0.235 $X2=3.445 $Y2=0.495
r286 1 29 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.155 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB4TO1_1%VGND 1 2 3 4 5 16 18 22 26 30 32 34 37
+ 38 40 41 42 51 65 76 80
r106 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r107 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r108 71 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.51
+ $Y2=0
r109 70 71 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r110 68 71 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.05 $Y2=0
r111 67 70 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=6.67 $Y=0 $X2=8.05
+ $Y2=0
r112 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r113 65 79 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.545
+ $Y2=0
r114 65 70 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=8.35 $Y=0 $X2=8.05
+ $Y2=0
r115 64 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r116 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r117 61 64 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r118 61 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r119 60 63 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r120 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r121 58 76 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.37
+ $Y2=0
r122 58 60 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.53 $Y=0 $X2=4.83
+ $Y2=0
r123 57 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r124 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r125 54 57 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r126 53 56 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r127 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r128 51 76 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=4.37
+ $Y2=0
r129 51 56 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=4.21 $Y=0 $X2=3.91
+ $Y2=0
r130 50 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r131 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r132 47 50 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r133 46 49 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r134 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r135 44 73 4.07647 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.195
+ $Y2=0
r136 44 46 19.5722 $w=1.68e-07 $l=3e-07 $layer=LI1_cond $X=0.39 $Y=0 $X2=0.69
+ $Y2=0
r137 42 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r138 42 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r139 40 63 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.21
+ $Y2=0
r140 40 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.275 $Y=0 $X2=6.44
+ $Y2=0
r141 39 67 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.67
+ $Y2=0
r142 39 41 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.605 $Y=0 $X2=6.44
+ $Y2=0
r143 37 49 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.07
+ $Y2=0
r144 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.135 $Y=0 $X2=2.3
+ $Y2=0
r145 36 53 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.53
+ $Y2=0
r146 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0 $X2=2.3
+ $Y2=0
r147 32 79 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=8.48 $Y=0.085
+ $X2=8.545 $Y2=0
r148 32 34 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=8.48 $Y=0.085
+ $X2=8.48 $Y2=0.38
r149 28 41 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0
r150 28 30 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=6.44 $Y=0.085
+ $X2=6.44 $Y2=0.495
r151 24 76 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0
r152 24 26 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=4.37 $Y=0.085
+ $X2=4.37 $Y2=0.38
r153 20 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.085 $X2=2.3
+ $Y2=0
r154 20 22 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=2.3 $Y=0.085
+ $X2=2.3 $Y2=0.495
r155 16 73 3.13575 $w=2.6e-07 $l=1.12916e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.195 $Y2=0
r156 16 18 13.0758 $w=2.58e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r157 5 34 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=8.345
+ $Y=0.235 $X2=8.48 $Y2=0.38
r158 4 30 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=6.225
+ $Y=0.235 $X2=6.44 $Y2=0.495
r159 3 26 91 $w=1.7e-07 $l=2.26164e-07 $layer=licon1_NDIFF $count=2 $X=4.205
+ $Y=0.235 $X2=4.37 $Y2=0.38
r160 2 22 182 $w=1.7e-07 $l=3.51426e-07 $layer=licon1_NDIFF $count=1 $X=2.085
+ $Y=0.235 $X2=2.3 $Y2=0.495
r161 1 18 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

