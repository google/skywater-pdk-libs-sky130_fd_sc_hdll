* File: sky130_fd_sc_hdll__nor2_1.spice
* Created: Thu Aug 27 19:15:22 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor2_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor2_1  VNB VPB B A Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1003 N_Y_M1003_d N_B_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1001 N_VGND_M1001_d N_A_M1001_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65 AD=0.39
+ AS=0.08775 PD=2.5 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7 SB=75000.5
+ A=0.0975 P=1.6 MULT=1
MM1002 A_117_297# N_B_M1002_g N_Y_M1002_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.27 PD=1.29 PS=2.54 NRD=17.7103 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.61
+ AS=0.145 PD=3.22 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90000.6
+ SB=90000.5 A=0.18 P=2.36 MULT=1
DX4_noxref VNB VPB NWDIODE A=3.5631 P=7.65
pX5_noxref noxref_9 A A PROBETYPE=1
c_113 A_117_297# 0 1.00411e-19 $X=0.585 $Y=1.485
*
.include "sky130_fd_sc_hdll__nor2_1.pxi.spice"
*
.ends
*
*
