* File: sky130_fd_sc_hdll__nor4bb_2.pxi.spice
* Created: Wed Sep  2 08:42:03 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%D_N N_D_N_M1019_g N_D_N_c_103_n N_D_N_c_104_n
+ N_D_N_M1008_g D_N D_N N_D_N_c_100_n N_D_N_c_101_n N_D_N_c_102_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%C_N N_C_N_c_133_n N_C_N_M1002_g N_C_N_c_134_n
+ N_C_N_M1013_g C_N C_N PM_SKY130_FD_SC_HDLL__NOR4BB_2%C_N
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_216_93# N_A_216_93#_M1002_d
+ N_A_216_93#_M1013_d N_A_216_93#_c_172_n N_A_216_93#_M1003_g
+ N_A_216_93#_c_164_n N_A_216_93#_M1000_g N_A_216_93#_c_173_n
+ N_A_216_93#_M1018_g N_A_216_93#_c_165_n N_A_216_93#_M1012_g
+ N_A_216_93#_c_174_n N_A_216_93#_c_166_n N_A_216_93#_c_167_n
+ N_A_216_93#_c_168_n N_A_216_93#_c_169_n N_A_216_93#_c_170_n
+ N_A_216_93#_c_171_n PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_216_93#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_27_93# N_A_27_93#_M1019_s N_A_27_93#_M1008_s
+ N_A_27_93#_c_241_n N_A_27_93#_M1006_g N_A_27_93#_c_249_n N_A_27_93#_M1011_g
+ N_A_27_93#_c_250_n N_A_27_93#_M1017_g N_A_27_93#_c_242_n N_A_27_93#_M1010_g
+ N_A_27_93#_c_243_n N_A_27_93#_c_252_n N_A_27_93#_c_253_n N_A_27_93#_c_269_n
+ N_A_27_93#_c_254_n N_A_27_93#_c_255_n N_A_27_93#_c_244_n N_A_27_93#_c_245_n
+ N_A_27_93#_c_246_n N_A_27_93#_c_247_n N_A_27_93#_c_257_n N_A_27_93#_c_248_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_27_93#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%B N_B_c_341_n N_B_M1004_g N_B_c_345_n
+ N_B_M1009_g N_B_c_346_n N_B_M1015_g N_B_c_342_n N_B_M1016_g B N_B_c_343_n
+ N_B_c_344_n B PM_SKY130_FD_SC_HDLL__NOR4BB_2%B
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A N_A_c_386_n N_A_M1005_g N_A_c_390_n
+ N_A_M1001_g N_A_c_391_n N_A_M1007_g N_A_c_387_n N_A_M1014_g A N_A_c_389_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%A
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%VPWR N_VPWR_M1008_d N_VPWR_M1001_s
+ N_VPWR_c_423_n N_VPWR_c_424_n N_VPWR_c_425_n N_VPWR_c_426_n VPWR
+ N_VPWR_c_427_n N_VPWR_c_428_n N_VPWR_c_422_n N_VPWR_c_430_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_343_297# N_A_343_297#_M1003_s
+ N_A_343_297#_M1018_s N_A_343_297#_M1017_d N_A_343_297#_c_484_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_343_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_433_297# N_A_433_297#_M1003_d
+ N_A_433_297#_M1009_s N_A_433_297#_c_508_n N_A_433_297#_c_519_n
+ N_A_433_297#_c_509_n PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_433_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%Y N_Y_M1000_d N_Y_M1006_s N_Y_M1004_s
+ N_Y_M1005_d N_Y_M1011_s N_Y_c_554_n N_Y_c_543_n N_Y_c_544_n N_Y_c_562_n
+ N_Y_c_545_n N_Y_c_546_n N_Y_c_585_n N_Y_c_547_n N_Y_c_588_n N_Y_c_548_n
+ N_Y_c_549_n N_Y_c_550_n Y Y N_Y_c_553_n Y PM_SKY130_FD_SC_HDLL__NOR4BB_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_823_297# N_A_823_297#_M1009_d
+ N_A_823_297#_M1015_d N_A_823_297#_M1007_d N_A_823_297#_c_647_n
+ N_A_823_297#_c_648_n N_A_823_297#_c_666_n N_A_823_297#_c_649_n
+ N_A_823_297#_c_650_n PM_SKY130_FD_SC_HDLL__NOR4BB_2%A_823_297#
x_PM_SKY130_FD_SC_HDLL__NOR4BB_2%VGND N_VGND_M1019_d N_VGND_M1000_s
+ N_VGND_M1012_s N_VGND_M1010_d N_VGND_M1004_d N_VGND_M1016_d N_VGND_M1014_s
+ N_VGND_c_684_n N_VGND_c_685_n N_VGND_c_686_n N_VGND_c_687_n N_VGND_c_688_n
+ N_VGND_c_689_n N_VGND_c_690_n N_VGND_c_691_n N_VGND_c_692_n N_VGND_c_693_n
+ N_VGND_c_694_n VGND N_VGND_c_695_n N_VGND_c_696_n N_VGND_c_697_n
+ N_VGND_c_698_n N_VGND_c_699_n N_VGND_c_700_n
+ PM_SKY130_FD_SC_HDLL__NOR4BB_2%VGND
cc_1 VNB N_D_N_c_100_n 0.0249711f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_2 VNB N_D_N_c_101_n 0.00893562f $X=-0.19 $Y=-0.24 $X2=0.53 $Y2=1.16
cc_3 VNB N_D_N_c_102_n 0.0215629f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_4 VNB N_C_N_c_133_n 0.0197086f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_5 VNB N_C_N_c_134_n 0.0331548f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.325
cc_6 VNB N_A_216_93#_c_164_n 0.0201184f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_7 VNB N_A_216_93#_c_165_n 0.0164985f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_8 VNB N_A_216_93#_c_166_n 0.0064227f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_216_93#_c_167_n 0.00125585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_216_93#_c_168_n 0.00556811f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_216_93#_c_169_n 0.0113595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_216_93#_c_170_n 0.0020035f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_216_93#_c_171_n 0.0542007f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_93#_c_241_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=2.26
cc_15 VNB N_A_27_93#_c_242_n 0.0202308f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=0.995
cc_16 VNB N_A_27_93#_c_243_n 0.0219616f $X=-0.19 $Y=-0.24 $X2=0.627 $Y2=1.19
cc_17 VNB N_A_27_93#_c_244_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_93#_c_245_n 0.00320416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_93#_c_246_n 0.00410515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_93#_c_247_n 0.0181399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_93#_c_248_n 0.0398472f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_B_c_341_n 0.0201516f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_23 VNB N_B_c_342_n 0.0169151f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_24 VNB N_B_c_343_n 0.00701525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_B_c_344_n 0.0392451f $X=-0.19 $Y=-0.24 $X2=0.627 $Y2=1.19
cc_26 VNB N_A_c_386_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_27 VNB N_A_c_387_n 0.0223809f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.445
cc_28 VNB A 0.0171554f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.16
cc_29 VNB N_A_c_389_n 0.04422f $X=-0.19 $Y=-0.24 $X2=0.627 $Y2=1.19
cc_30 VNB N_VPWR_c_422_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_543_n 0.00303118f $X=-0.19 $Y=-0.24 $X2=0.627 $Y2=1.19
cc_32 VNB N_Y_c_544_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_545_n 0.00294903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_546_n 0.00567378f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_547_n 0.00570013f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_548_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_549_n 0.00424437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_550_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB Y 0.0128392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_684_n 0.0151641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_685_n 0.0211891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_686_n 0.0119652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_687_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_688_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_689_n 0.0109994f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_690_n 0.0336326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_691_n 0.0199148f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_692_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_693_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_694_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_695_n 0.0201171f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_696_n 0.0247769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_697_n 0.00631201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_698_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_699_n 0.0270892f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_700_n 0.337542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VPB N_D_N_c_103_n 0.0337057f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.875
cc_58 VPB N_D_N_c_104_n 0.0283679f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.975
cc_59 VPB N_D_N_c_100_n 0.00418278f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_60 VPB N_D_N_c_101_n 0.00237191f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_61 VPB N_C_N_c_134_n 0.0302306f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_62 VPB N_A_216_93#_c_172_n 0.0192053f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_63 VPB N_A_216_93#_c_173_n 0.0156053f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_64 VPB N_A_216_93#_c_174_n 0.00654754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_216_93#_c_167_n 0.00539386f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_216_93#_c_171_n 0.0249797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_93#_c_249_n 0.0161563f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.445
cc_68 VPB N_A_27_93#_c_250_n 0.0191622f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_69 VPB N_A_27_93#_c_243_n 0.0272067f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.19
cc_70 VPB N_A_27_93#_c_252_n 0.0155282f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_93#_c_253_n 0.0195829f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_93#_c_254_n 0.00330088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_27_93#_c_255_n 0.00163568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_27_93#_c_244_n 0.00190486f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_27_93#_c_257_n 0.011274f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_27_93#_c_248_n 0.0200389f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_B_c_345_n 0.0192127f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_78 VPB N_B_c_346_n 0.016292f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_79 VPB N_B_c_344_n 0.0204488f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.19
cc_80 VPB N_A_c_390_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.325
cc_81 VPB N_A_c_391_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_82 VPB N_A_c_389_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.19
cc_83 VPB N_VPWR_c_423_n 0.0130131f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_84 VPB N_VPWR_c_424_n 0.00491015f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_85 VPB N_VPWR_c_425_n 0.110609f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=0.995
cc_86 VPB N_VPWR_c_426_n 0.00401008f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.325
cc_87 VPB N_VPWR_c_427_n 0.0144832f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.19
cc_88 VPB N_VPWR_c_428_n 0.0202461f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_422_n 0.0610631f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_430_n 0.00593536f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_A_343_297#_c_484_n 0.013599f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=0.995
cc_92 VPB N_A_433_297#_c_508_n 0.00750102f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=2.26
cc_93 VPB N_A_433_297#_c_509_n 0.0019668f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.16
cc_94 VPB Y 0.0108553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_553_n 0.0045976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_A_823_297#_c_647_n 0.00254845f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.445
cc_97 VPB N_A_823_297#_c_648_n 0.00244172f $X=-0.19 $Y=1.305 $X2=0.53 $Y2=1.16
cc_98 VPB N_A_823_297#_c_649_n 0.0120871f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=0.995
cc_99 VPB N_A_823_297#_c_650_n 0.0327326f $X=-0.19 $Y=1.305 $X2=0.627 $Y2=1.19
cc_100 N_D_N_c_102_n N_C_N_c_133_n 0.0122079f $X=0.545 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_101 N_D_N_c_103_n N_C_N_c_134_n 0.0219501f $X=0.495 $Y=1.875 $X2=0 $Y2=0
cc_102 N_D_N_c_104_n N_C_N_c_134_n 0.00196013f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_103 N_D_N_c_100_n N_C_N_c_134_n 0.0178271f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_104 N_D_N_c_101_n N_C_N_c_134_n 0.00657742f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_105 N_D_N_c_100_n C_N 2.9088e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_106 N_D_N_c_101_n C_N 0.026141f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_107 N_D_N_c_103_n N_A_216_93#_c_174_n 2.29988e-19 $X=0.495 $Y=1.875 $X2=0
+ $Y2=0
cc_108 N_D_N_c_101_n N_A_216_93#_c_174_n 0.0116234f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_109 N_D_N_c_101_n N_A_216_93#_c_167_n 0.00650379f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_110 N_D_N_c_101_n N_A_27_93#_c_243_n 0.0534049f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_111 N_D_N_c_102_n N_A_27_93#_c_243_n 0.0276355f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_112 N_D_N_c_104_n N_A_27_93#_c_252_n 0.00541304f $X=0.495 $Y=1.975 $X2=0
+ $Y2=0
cc_113 N_D_N_c_104_n N_A_27_93#_c_253_n 0.0166237f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_114 N_D_N_c_100_n N_A_27_93#_c_253_n 3.24788e-19 $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_115 N_D_N_c_101_n N_A_27_93#_c_253_n 0.0296016f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_116 N_D_N_c_101_n N_A_27_93#_c_247_n 0.00314948f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_117 N_D_N_c_102_n N_A_27_93#_c_247_n 0.00855468f $X=0.545 $Y=0.995 $X2=0
+ $Y2=0
cc_118 N_D_N_c_101_n N_VPWR_M1008_d 0.00455541f $X=0.53 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_119 N_D_N_c_104_n N_VPWR_c_423_n 0.0122933f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_120 N_D_N_c_104_n N_VPWR_c_427_n 0.00308256f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_121 N_D_N_c_104_n N_VPWR_c_422_n 0.00457045f $X=0.495 $Y=1.975 $X2=0 $Y2=0
cc_122 N_D_N_c_101_n N_VGND_c_684_n 0.0131343f $X=0.53 $Y=1.16 $X2=0 $Y2=0
cc_123 N_D_N_c_102_n N_VGND_c_684_n 0.0054831f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_124 N_D_N_c_102_n N_VGND_c_696_n 0.00446966f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_125 N_D_N_c_102_n N_VGND_c_700_n 0.00512902f $X=0.545 $Y=0.995 $X2=0 $Y2=0
cc_126 N_C_N_c_134_n N_A_216_93#_c_174_n 0.00928798f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_127 C_N N_A_216_93#_c_174_n 0.0126971f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_128 N_C_N_c_133_n N_A_216_93#_c_166_n 0.00431395f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_129 N_C_N_c_134_n N_A_216_93#_c_166_n 7.45304e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_130 C_N N_A_216_93#_c_166_n 0.00583896f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_131 N_C_N_c_134_n N_A_216_93#_c_167_n 0.00419246f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_132 C_N N_A_216_93#_c_167_n 0.00583896f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_133 N_C_N_c_133_n N_A_216_93#_c_169_n 0.00216441f $X=1.005 $Y=0.995 $X2=0
+ $Y2=0
cc_134 N_C_N_c_134_n N_A_216_93#_c_169_n 0.00386344f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_135 C_N N_A_216_93#_c_169_n 0.00906071f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_136 N_C_N_c_134_n N_A_216_93#_c_170_n 0.00173423f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_137 C_N N_A_216_93#_c_170_n 0.0142121f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_138 N_C_N_c_134_n N_A_216_93#_c_171_n 0.0062984f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_139 N_C_N_c_134_n N_A_27_93#_c_253_n 0.0156347f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_140 C_N N_A_27_93#_c_253_n 0.00120587f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_141 N_C_N_c_134_n N_A_27_93#_c_269_n 0.00240615f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_142 N_C_N_c_134_n N_VPWR_c_425_n 6.57516e-19 $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_143 N_C_N_c_133_n N_VGND_c_684_n 0.00455897f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_144 N_C_N_c_133_n N_VGND_c_685_n 0.00510437f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_145 N_C_N_c_133_n N_VGND_c_686_n 0.00302957f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_146 N_C_N_c_133_n N_VGND_c_700_n 0.00512902f $X=1.005 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_216_93#_c_165_n N_A_27_93#_c_241_n 0.0231417f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_148 N_A_216_93#_c_173_n N_A_27_93#_c_249_n 0.037944f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_216_93#_M1013_d N_A_27_93#_c_253_n 0.00223951f $X=1.12 $Y=1.485 $X2=0
+ $Y2=0
cc_150 N_A_216_93#_c_174_n N_A_27_93#_c_253_n 0.0387178f $X=1.44 $Y=1.62 $X2=0
+ $Y2=0
cc_151 N_A_216_93#_c_168_n N_A_27_93#_c_253_n 0.00495382f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_152 N_A_216_93#_c_174_n N_A_27_93#_c_269_n 0.0106046f $X=1.44 $Y=1.62 $X2=0
+ $Y2=0
cc_153 N_A_216_93#_c_172_n N_A_27_93#_c_254_n 0.0153203f $X=2.075 $Y=1.41 $X2=0
+ $Y2=0
cc_154 N_A_216_93#_c_173_n N_A_27_93#_c_254_n 0.0140186f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_155 N_A_216_93#_c_168_n N_A_27_93#_c_254_n 0.0367613f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_156 N_A_216_93#_c_171_n N_A_27_93#_c_254_n 0.009123f $X=2.545 $Y=1.202 $X2=0
+ $Y2=0
cc_157 N_A_216_93#_c_174_n N_A_27_93#_c_255_n 0.00543966f $X=1.44 $Y=1.62 $X2=0
+ $Y2=0
cc_158 N_A_216_93#_c_167_n N_A_27_93#_c_255_n 0.00918172f $X=1.525 $Y=1.525
+ $X2=0 $Y2=0
cc_159 N_A_216_93#_c_168_n N_A_27_93#_c_255_n 0.0136617f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_160 N_A_216_93#_c_171_n N_A_27_93#_c_255_n 0.00422084f $X=2.545 $Y=1.202
+ $X2=0 $Y2=0
cc_161 N_A_216_93#_c_171_n N_A_27_93#_c_244_n 0.00331682f $X=2.545 $Y=1.202
+ $X2=0 $Y2=0
cc_162 N_A_216_93#_c_168_n N_A_27_93#_c_245_n 0.0123234f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_163 N_A_216_93#_c_171_n N_A_27_93#_c_245_n 0.00288841f $X=2.545 $Y=1.202
+ $X2=0 $Y2=0
cc_164 N_A_216_93#_c_171_n N_A_27_93#_c_248_n 0.0231417f $X=2.545 $Y=1.202 $X2=0
+ $Y2=0
cc_165 N_A_216_93#_c_172_n N_VPWR_c_425_n 0.00429453f $X=2.075 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_A_216_93#_c_173_n N_VPWR_c_425_n 0.00429453f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_216_93#_c_172_n N_VPWR_c_422_n 0.00734734f $X=2.075 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_216_93#_c_173_n N_VPWR_c_422_n 0.00609021f $X=2.545 $Y=1.41 $X2=0
+ $Y2=0
cc_169 N_A_216_93#_c_172_n N_A_343_297#_c_484_n 0.0133276f $X=2.075 $Y=1.41
+ $X2=0 $Y2=0
cc_170 N_A_216_93#_c_173_n N_A_343_297#_c_484_n 0.0110437f $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_171 N_A_216_93#_c_172_n N_A_433_297#_c_508_n 0.00257937f $X=2.075 $Y=1.41
+ $X2=0 $Y2=0
cc_172 N_A_216_93#_c_173_n N_A_433_297#_c_508_n 0.0106257f $X=2.545 $Y=1.41
+ $X2=0 $Y2=0
cc_173 N_A_216_93#_c_164_n N_Y_c_554_n 0.0139042f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_216_93#_c_169_n N_Y_c_554_n 0.0026118f $X=1.24 $Y=0.66 $X2=0 $Y2=0
cc_175 N_A_216_93#_c_165_n N_Y_c_543_n 0.0122714f $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_216_93#_c_164_n N_Y_c_544_n 0.00540497f $X=2.1 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_216_93#_c_166_n N_Y_c_544_n 0.00287206f $X=1.525 $Y=1.075 $X2=0 $Y2=0
cc_178 N_A_216_93#_c_168_n N_Y_c_544_n 0.030184f $X=2.31 $Y=1.16 $X2=0 $Y2=0
cc_179 N_A_216_93#_c_169_n N_Y_c_544_n 0.00391381f $X=1.24 $Y=0.66 $X2=0 $Y2=0
cc_180 N_A_216_93#_c_171_n N_Y_c_544_n 0.00358305f $X=2.545 $Y=1.202 $X2=0 $Y2=0
cc_181 N_A_216_93#_c_165_n N_Y_c_562_n 5.32212e-19 $X=2.57 $Y=0.995 $X2=0 $Y2=0
cc_182 N_A_216_93#_c_173_n N_Y_c_553_n 7.0686e-19 $X=2.545 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_216_93#_c_169_n N_VGND_c_684_n 0.0187732f $X=1.24 $Y=0.66 $X2=0 $Y2=0
cc_184 N_A_216_93#_c_169_n N_VGND_c_685_n 0.0105281f $X=1.24 $Y=0.66 $X2=0 $Y2=0
cc_185 N_A_216_93#_c_164_n N_VGND_c_686_n 0.00968298f $X=2.1 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_216_93#_c_168_n N_VGND_c_686_n 0.00982788f $X=2.31 $Y=1.16 $X2=0
+ $Y2=0
cc_187 N_A_216_93#_c_169_n N_VGND_c_686_n 0.00304964f $X=1.24 $Y=0.66 $X2=0
+ $Y2=0
cc_188 N_A_216_93#_c_171_n N_VGND_c_686_n 0.00261712f $X=2.545 $Y=1.202 $X2=0
+ $Y2=0
cc_189 N_A_216_93#_c_165_n N_VGND_c_687_n 0.00268723f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_190 N_A_216_93#_c_164_n N_VGND_c_691_n 0.00465454f $X=2.1 $Y=0.995 $X2=0
+ $Y2=0
cc_191 N_A_216_93#_c_165_n N_VGND_c_691_n 0.00437852f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_216_93#_c_164_n N_VGND_c_700_n 0.00935497f $X=2.1 $Y=0.995 $X2=0
+ $Y2=0
cc_193 N_A_216_93#_c_165_n N_VGND_c_700_n 0.00604088f $X=2.57 $Y=0.995 $X2=0
+ $Y2=0
cc_194 N_A_216_93#_c_169_n N_VGND_c_700_n 0.0137666f $X=1.24 $Y=0.66 $X2=0 $Y2=0
cc_195 N_A_27_93#_c_253_n N_VPWR_M1008_d 0.00607135f $X=1.78 $Y=1.97 $X2=-0.19
+ $Y2=-0.24
cc_196 N_A_27_93#_c_252_n N_VPWR_c_423_n 0.0165638f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_197 N_A_27_93#_c_253_n N_VPWR_c_423_n 0.0226765f $X=1.78 $Y=1.97 $X2=0 $Y2=0
cc_198 N_A_27_93#_c_249_n N_VPWR_c_425_n 0.00429453f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_27_93#_c_250_n N_VPWR_c_425_n 0.00429453f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A_27_93#_c_253_n N_VPWR_c_425_n 0.0133812f $X=1.78 $Y=1.97 $X2=0 $Y2=0
cc_201 N_A_27_93#_c_252_n N_VPWR_c_427_n 0.0170401f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_202 N_A_27_93#_c_253_n N_VPWR_c_427_n 0.00221427f $X=1.78 $Y=1.97 $X2=0 $Y2=0
cc_203 N_A_27_93#_c_249_n N_VPWR_c_422_n 0.00609021f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_27_93#_c_250_n N_VPWR_c_422_n 0.00734734f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_27_93#_c_252_n N_VPWR_c_422_n 0.00987287f $X=0.26 $Y=2.29 $X2=0 $Y2=0
cc_206 N_A_27_93#_c_253_n N_VPWR_c_422_n 0.027617f $X=1.78 $Y=1.97 $X2=0 $Y2=0
cc_207 N_A_27_93#_c_253_n N_A_343_297#_M1003_s 0.0054897f $X=1.78 $Y=1.97
+ $X2=-0.19 $Y2=-0.24
cc_208 N_A_27_93#_c_269_n N_A_343_297#_M1003_s 0.00544591f $X=1.865 $Y=1.885
+ $X2=-0.19 $Y2=-0.24
cc_209 N_A_27_93#_c_255_n N_A_343_297#_M1003_s 0.00115536f $X=1.95 $Y=1.5
+ $X2=-0.19 $Y2=-0.24
cc_210 N_A_27_93#_c_254_n N_A_343_297#_M1018_s 0.00345892f $X=2.695 $Y=1.5 $X2=0
+ $Y2=0
cc_211 N_A_27_93#_c_249_n N_A_343_297#_c_484_n 0.0110437f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_27_93#_c_250_n N_A_343_297#_c_484_n 0.0110437f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_27_93#_c_253_n N_A_343_297#_c_484_n 0.0192171f $X=1.78 $Y=1.97 $X2=0
+ $Y2=0
cc_214 N_A_27_93#_c_254_n N_A_343_297#_c_484_n 0.00368504f $X=2.695 $Y=1.5 $X2=0
+ $Y2=0
cc_215 N_A_27_93#_c_254_n N_A_433_297#_M1003_d 0.00239437f $X=2.695 $Y=1.5
+ $X2=-0.19 $Y2=-0.24
cc_216 N_A_27_93#_c_249_n N_A_433_297#_c_508_n 0.0134136f $X=3.015 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_27_93#_c_250_n N_A_433_297#_c_508_n 0.01396f $X=3.485 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_27_93#_c_254_n N_A_433_297#_c_508_n 0.0266119f $X=2.695 $Y=1.5 $X2=0
+ $Y2=0
cc_219 N_A_27_93#_c_246_n N_A_433_297#_c_508_n 0.00361241f $X=3.44 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A_27_93#_c_241_n N_Y_c_543_n 0.00865686f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_221 N_A_27_93#_c_254_n N_Y_c_543_n 0.00656431f $X=2.695 $Y=1.5 $X2=0 $Y2=0
cc_222 N_A_27_93#_c_245_n N_Y_c_543_n 0.0140787f $X=2.865 $Y=1.175 $X2=0 $Y2=0
cc_223 N_A_27_93#_c_246_n N_Y_c_543_n 0.0120283f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A_27_93#_c_241_n N_Y_c_562_n 0.00644736f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_27_93#_c_242_n N_Y_c_545_n 0.01289f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_27_93#_c_246_n N_Y_c_545_n 0.0159687f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_93#_c_241_n N_Y_c_548_n 0.00119564f $X=2.99 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_27_93#_c_246_n N_Y_c_548_n 0.0307352f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_229 N_A_27_93#_c_248_n N_Y_c_548_n 0.00486271f $X=3.485 $Y=1.202 $X2=0 $Y2=0
cc_230 N_A_27_93#_c_250_n Y 0.00123534f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_27_93#_c_242_n Y 0.0066531f $X=3.51 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_27_93#_c_246_n Y 0.0178203f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_233 N_A_27_93#_c_248_n Y 0.00660105f $X=3.485 $Y=1.202 $X2=0 $Y2=0
cc_234 N_A_27_93#_c_249_n N_Y_c_553_n 0.0071848f $X=3.015 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_27_93#_c_250_n N_Y_c_553_n 0.0159102f $X=3.485 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_27_93#_c_254_n N_Y_c_553_n 0.0122169f $X=2.695 $Y=1.5 $X2=0 $Y2=0
cc_237 N_A_27_93#_c_246_n N_Y_c_553_n 0.0445277f $X=3.44 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_27_93#_c_248_n N_Y_c_553_n 0.00775718f $X=3.485 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A_27_93#_c_247_n N_VGND_c_684_n 0.0229402f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_240 N_A_27_93#_c_241_n N_VGND_c_687_n 0.00268723f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_241 N_A_27_93#_c_247_n N_VGND_c_696_n 0.01138f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_242 N_A_27_93#_c_241_n N_VGND_c_698_n 0.00423334f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_243 N_A_27_93#_c_242_n N_VGND_c_698_n 0.00437852f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_244 N_A_27_93#_c_242_n N_VGND_c_699_n 0.00482606f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_27_93#_c_241_n N_VGND_c_700_n 0.00598581f $X=2.99 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_27_93#_c_242_n N_VGND_c_700_n 0.00745263f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_247 N_A_27_93#_c_247_n N_VGND_c_700_n 0.0126704f $X=0.26 $Y=0.66 $X2=0 $Y2=0
cc_248 N_B_c_342_n N_A_c_386_n 0.024293f $X=4.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_249 N_B_c_346_n N_A_c_390_n 0.00971835f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_343_n A 0.0175712f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B_c_343_n N_A_c_389_n 0.00196293f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_252 N_B_c_344_n N_A_c_389_n 0.024293f $X=4.965 $Y=1.202 $X2=0 $Y2=0
cc_253 N_B_c_345_n N_VPWR_c_425_n 0.00429453f $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_346_n N_VPWR_c_425_n 0.00429453f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_345_n N_VPWR_c_422_n 0.00734734f $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_346_n N_VPWR_c_422_n 0.00609021f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_345_n N_A_433_297#_c_508_n 0.0142129f $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_343_n N_A_433_297#_c_508_n 0.00464791f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B_c_346_n N_A_433_297#_c_519_n 0.00225067f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B_c_345_n N_A_433_297#_c_509_n 3.42233e-19 $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B_c_346_n N_A_433_297#_c_509_n 0.00544851f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B_c_343_n N_A_433_297#_c_509_n 0.0221391f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_263 N_B_c_344_n N_A_433_297#_c_509_n 0.00693986f $X=4.965 $Y=1.202 $X2=0
+ $Y2=0
cc_264 N_B_c_341_n N_Y_c_546_n 0.0110736f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_265 N_B_c_343_n N_Y_c_546_n 0.00789367f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_266 N_B_c_341_n N_Y_c_585_n 0.0110728f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_267 N_B_c_342_n N_Y_c_547_n 0.0106151f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_268 N_B_c_343_n N_Y_c_547_n 0.0293687f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_269 N_B_c_342_n N_Y_c_588_n 5.32212e-19 $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_270 N_B_c_341_n N_Y_c_550_n 0.00119564f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_271 N_B_c_343_n N_Y_c_550_n 0.0307352f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_272 N_B_c_344_n N_Y_c_550_n 0.00486271f $X=4.965 $Y=1.202 $X2=0 $Y2=0
cc_273 N_B_c_341_n Y 0.0180465f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_274 N_B_c_345_n Y 0.00765311f $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B_c_343_n Y 0.0169224f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_276 N_B_c_345_n N_A_823_297#_c_647_n 0.0112654f $X=4.495 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B_c_346_n N_A_823_297#_c_647_n 0.0164047f $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B_c_346_n N_A_823_297#_c_648_n 9.55966e-19 $X=4.965 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_343_n N_A_823_297#_c_648_n 0.0147624f $X=4.745 $Y=1.16 $X2=0 $Y2=0
cc_280 N_B_c_342_n N_VGND_c_688_n 0.00268723f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_281 N_B_c_341_n N_VGND_c_693_n 0.00423334f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_282 N_B_c_342_n N_VGND_c_693_n 0.00437852f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_283 N_B_c_341_n N_VGND_c_699_n 0.00482606f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_284 N_B_c_341_n N_VGND_c_700_n 0.00728222f $X=4.47 $Y=0.995 $X2=0 $Y2=0
cc_285 N_B_c_342_n N_VGND_c_700_n 0.00615622f $X=4.99 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_c_390_n N_VPWR_c_424_n 0.00295479f $X=5.435 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A_c_391_n N_VPWR_c_424_n 0.00502706f $X=5.905 $Y=1.41 $X2=0 $Y2=0
cc_288 N_A_c_390_n N_VPWR_c_425_n 0.00702461f $X=5.435 $Y=1.41 $X2=0 $Y2=0
cc_289 N_A_c_391_n N_VPWR_c_428_n 0.00597712f $X=5.905 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A_c_390_n N_VPWR_c_422_n 0.0124344f $X=5.435 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A_c_391_n N_VPWR_c_422_n 0.0109412f $X=5.905 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_c_386_n N_Y_c_547_n 0.011403f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_c_387_n N_Y_c_547_n 2.15189e-19 $X=5.93 $Y=0.995 $X2=0 $Y2=0
cc_294 A N_Y_c_547_n 0.0300441f $X=5.59 $Y=1.105 $X2=0 $Y2=0
cc_295 N_A_c_389_n N_Y_c_547_n 0.00485909f $X=5.905 $Y=1.202 $X2=0 $Y2=0
cc_296 N_A_c_386_n N_Y_c_588_n 0.00644736f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A_c_390_n N_A_823_297#_c_649_n 0.0170656f $X=5.435 $Y=1.41 $X2=0 $Y2=0
cc_298 N_A_c_391_n N_A_823_297#_c_649_n 0.0128395f $X=5.905 $Y=1.41 $X2=0 $Y2=0
cc_299 A N_A_823_297#_c_649_n 0.0619907f $X=5.59 $Y=1.105 $X2=0 $Y2=0
cc_300 N_A_c_389_n N_A_823_297#_c_649_n 0.00799226f $X=5.905 $Y=1.202 $X2=0
+ $Y2=0
cc_301 N_A_c_390_n N_A_823_297#_c_650_n 6.6798e-19 $X=5.435 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_c_391_n N_A_823_297#_c_650_n 0.0137341f $X=5.905 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_c_386_n N_VGND_c_688_n 0.00268723f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_c_387_n N_VGND_c_690_n 0.00498331f $X=5.93 $Y=0.995 $X2=0 $Y2=0
cc_305 A N_VGND_c_690_n 0.0234299f $X=5.59 $Y=1.105 $X2=0 $Y2=0
cc_306 N_A_c_386_n N_VGND_c_695_n 0.00423334f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_c_387_n N_VGND_c_695_n 0.00585385f $X=5.93 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_386_n N_VGND_c_700_n 0.00598581f $X=5.41 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_c_387_n N_VGND_c_700_n 0.0117699f $X=5.93 $Y=0.995 $X2=0 $Y2=0
cc_310 N_VPWR_c_422_n N_A_343_297#_M1003_s 0.00217543f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_311 N_VPWR_c_422_n N_A_343_297#_M1018_s 0.00231289f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_422_n N_A_343_297#_M1017_d 0.00217543f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_313 N_VPWR_c_425_n N_A_343_297#_c_484_n 0.12847f $X=5.545 $Y=2.72 $X2=0 $Y2=0
cc_314 N_VPWR_c_422_n N_A_343_297#_c_484_n 0.079368f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_422_n N_A_433_297#_M1003_d 0.00232895f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_316 N_VPWR_c_422_n N_A_433_297#_M1009_s 0.00232895f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_317 N_VPWR_c_425_n N_A_433_297#_c_508_n 0.00353234f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_318 N_VPWR_c_422_n N_A_433_297#_c_508_n 0.00975247f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_319 N_VPWR_c_422_n N_Y_M1011_s 0.00232895f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_422_n N_A_823_297#_M1009_d 0.00233941f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_321 N_VPWR_c_422_n N_A_823_297#_M1015_d 0.00297226f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_322 N_VPWR_c_422_n N_A_823_297#_M1007_d 0.00229814f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_323 N_VPWR_c_425_n N_A_823_297#_c_647_n 0.0587492f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_324 N_VPWR_c_422_n N_A_823_297#_c_647_n 0.0365159f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_425_n N_A_823_297#_c_666_n 0.0134783f $X=5.545 $Y=2.72 $X2=0
+ $Y2=0
cc_326 N_VPWR_c_422_n N_A_823_297#_c_666_n 0.00808747f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_327 N_VPWR_M1001_s N_A_823_297#_c_649_n 0.00182839f $X=5.525 $Y=1.485 $X2=0
+ $Y2=0
cc_328 N_VPWR_c_424_n N_A_823_297#_c_649_n 0.0139937f $X=5.67 $Y=1.96 $X2=0
+ $Y2=0
cc_329 N_VPWR_c_424_n N_A_823_297#_c_650_n 0.0508019f $X=5.67 $Y=1.96 $X2=0
+ $Y2=0
cc_330 N_VPWR_c_428_n N_A_823_297#_c_650_n 0.0244479f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_331 N_VPWR_c_422_n N_A_823_297#_c_650_n 0.0141694f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_332 N_A_343_297#_c_484_n N_A_433_297#_M1003_d 0.00361214f $X=3.72 $Y=2.31
+ $X2=-0.19 $Y2=1.305
cc_333 N_A_343_297#_M1018_s N_A_433_297#_c_508_n 0.00413606f $X=2.635 $Y=1.485
+ $X2=0 $Y2=0
cc_334 N_A_343_297#_M1017_d N_A_433_297#_c_508_n 0.0053555f $X=3.575 $Y=1.485
+ $X2=0 $Y2=0
cc_335 N_A_343_297#_c_484_n N_A_433_297#_c_508_n 0.0883876f $X=3.72 $Y=2.31
+ $X2=0 $Y2=0
cc_336 N_A_343_297#_c_484_n N_Y_M1011_s 0.00361214f $X=3.72 $Y=2.31 $X2=0 $Y2=0
cc_337 N_A_343_297#_M1017_d Y 8.14469e-19 $X=3.575 $Y=1.485 $X2=0 $Y2=0
cc_338 N_A_343_297#_M1017_d N_Y_c_553_n 0.00256556f $X=3.575 $Y=1.485 $X2=0
+ $Y2=0
cc_339 N_A_343_297#_c_484_n N_A_823_297#_c_647_n 0.0191977f $X=3.72 $Y=2.31
+ $X2=0 $Y2=0
cc_340 N_A_433_297#_c_508_n N_Y_M1011_s 0.00355096f $X=4.605 $Y=1.96 $X2=0 $Y2=0
cc_341 N_A_433_297#_c_508_n Y 0.0350081f $X=4.605 $Y=1.96 $X2=0 $Y2=0
cc_342 N_A_433_297#_c_509_n Y 0.00698829f $X=4.73 $Y=1.62 $X2=0 $Y2=0
cc_343 N_A_433_297#_c_508_n N_Y_c_553_n 0.0439624f $X=4.605 $Y=1.96 $X2=0 $Y2=0
cc_344 N_A_433_297#_c_508_n N_A_823_297#_M1009_d 0.00915276f $X=4.605 $Y=1.96
+ $X2=-0.19 $Y2=1.305
cc_345 N_A_433_297#_M1009_s N_A_823_297#_c_647_n 0.00356605f $X=4.585 $Y=1.485
+ $X2=0 $Y2=0
cc_346 N_A_433_297#_c_508_n N_A_823_297#_c_647_n 0.03012f $X=4.605 $Y=1.96 $X2=0
+ $Y2=0
cc_347 N_A_433_297#_c_519_n N_A_823_297#_c_647_n 0.0152922f $X=4.75 $Y=1.875
+ $X2=0 $Y2=0
cc_348 N_A_433_297#_c_509_n N_A_823_297#_c_648_n 0.0114601f $X=4.73 $Y=1.62
+ $X2=0 $Y2=0
cc_349 N_A_433_297#_c_519_n N_A_823_297#_c_666_n 0.0111041f $X=4.75 $Y=1.875
+ $X2=0 $Y2=0
cc_350 N_A_433_297#_c_509_n N_A_823_297#_c_666_n 0.0151665f $X=4.73 $Y=1.62
+ $X2=0 $Y2=0
cc_351 Y N_A_823_297#_M1009_d 0.00534861f $X=4.06 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_352 N_Y_c_547_n N_A_823_297#_c_648_n 0.00112383f $X=5.455 $Y=0.815 $X2=0
+ $Y2=0
cc_353 N_Y_c_547_n N_A_823_297#_c_649_n 0.00377384f $X=5.455 $Y=0.815 $X2=0
+ $Y2=0
cc_354 N_Y_c_543_n N_VGND_M1012_s 0.00162089f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_355 N_Y_c_545_n N_VGND_M1010_d 0.00212652f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_356 N_Y_c_549_n N_VGND_M1010_d 6.88755e-19 $X=4.02 $Y=0.815 $X2=0 $Y2=0
cc_357 N_Y_c_546_n N_VGND_M1004_d 0.00111439f $X=4.515 $Y=0.815 $X2=0 $Y2=0
cc_358 N_Y_c_549_n N_VGND_M1004_d 0.00213021f $X=4.02 $Y=0.815 $X2=0 $Y2=0
cc_359 N_Y_c_547_n N_VGND_M1016_d 0.00162089f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_360 N_Y_c_554_n N_VGND_c_686_n 0.0176499f $X=2.31 $Y=0.39 $X2=0 $Y2=0
cc_361 N_Y_c_543_n N_VGND_c_687_n 0.0122559f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_362 N_Y_c_547_n N_VGND_c_688_n 0.0122559f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_363 N_Y_c_547_n N_VGND_c_690_n 0.00138214f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_364 N_Y_c_554_n N_VGND_c_691_n 0.023074f $X=2.31 $Y=0.39 $X2=0 $Y2=0
cc_365 N_Y_c_543_n N_VGND_c_691_n 0.00254521f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_366 N_Y_c_546_n N_VGND_c_693_n 0.00198695f $X=4.515 $Y=0.815 $X2=0 $Y2=0
cc_367 N_Y_c_585_n N_VGND_c_693_n 0.0231806f $X=4.73 $Y=0.39 $X2=0 $Y2=0
cc_368 N_Y_c_547_n N_VGND_c_693_n 0.00254521f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_369 N_Y_c_547_n N_VGND_c_695_n 0.00198695f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_370 N_Y_c_588_n N_VGND_c_695_n 0.0231806f $X=5.67 $Y=0.39 $X2=0 $Y2=0
cc_371 N_Y_c_543_n N_VGND_c_698_n 0.00198695f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_372 N_Y_c_562_n N_VGND_c_698_n 0.0231806f $X=3.25 $Y=0.39 $X2=0 $Y2=0
cc_373 N_Y_c_545_n N_VGND_c_698_n 0.00254521f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_374 N_Y_c_545_n N_VGND_c_699_n 0.0130966f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_375 N_Y_c_546_n N_VGND_c_699_n 0.00840711f $X=4.515 $Y=0.815 $X2=0 $Y2=0
cc_376 N_Y_c_549_n N_VGND_c_699_n 0.0370461f $X=4.02 $Y=0.815 $X2=0 $Y2=0
cc_377 N_Y_M1000_d N_VGND_c_700_n 0.00263993f $X=2.175 $Y=0.235 $X2=0 $Y2=0
cc_378 N_Y_M1006_s N_VGND_c_700_n 0.00304143f $X=3.065 $Y=0.235 $X2=0 $Y2=0
cc_379 N_Y_M1004_s N_VGND_c_700_n 0.00304143f $X=4.545 $Y=0.235 $X2=0 $Y2=0
cc_380 N_Y_M1005_d N_VGND_c_700_n 0.00364931f $X=5.485 $Y=0.235 $X2=0 $Y2=0
cc_381 N_Y_c_554_n N_VGND_c_700_n 0.0141066f $X=2.31 $Y=0.39 $X2=0 $Y2=0
cc_382 N_Y_c_543_n N_VGND_c_700_n 0.0094839f $X=3.035 $Y=0.815 $X2=0 $Y2=0
cc_383 N_Y_c_562_n N_VGND_c_700_n 0.0143352f $X=3.25 $Y=0.39 $X2=0 $Y2=0
cc_384 N_Y_c_545_n N_VGND_c_700_n 0.00563527f $X=3.81 $Y=0.815 $X2=0 $Y2=0
cc_385 N_Y_c_546_n N_VGND_c_700_n 0.00427976f $X=4.515 $Y=0.815 $X2=0 $Y2=0
cc_386 N_Y_c_585_n N_VGND_c_700_n 0.0143352f $X=4.73 $Y=0.39 $X2=0 $Y2=0
cc_387 N_Y_c_547_n N_VGND_c_700_n 0.0094839f $X=5.455 $Y=0.815 $X2=0 $Y2=0
cc_388 N_Y_c_588_n N_VGND_c_700_n 0.0143352f $X=5.67 $Y=0.39 $X2=0 $Y2=0
cc_389 N_Y_c_549_n N_VGND_c_700_n 0.00181962f $X=4.02 $Y=0.815 $X2=0 $Y2=0
