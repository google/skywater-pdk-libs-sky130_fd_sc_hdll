* File: sky130_fd_sc_hdll__nor4_8.pxi.spice
* Created: Thu Aug 27 19:17:21 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4_8%A N_A_c_218_n N_A_M1000_g N_A_c_209_n N_A_M1018_g
+ N_A_c_210_n N_A_M1019_g N_A_c_219_n N_A_M1003_g N_A_c_220_n N_A_M1008_g
+ N_A_c_211_n N_A_M1031_g N_A_c_212_n N_A_M1038_g N_A_c_221_n N_A_M1016_g
+ N_A_c_222_n N_A_M1026_g N_A_c_213_n N_A_M1045_g N_A_c_214_n N_A_M1051_g
+ N_A_c_223_n N_A_M1032_g N_A_c_224_n N_A_M1040_g N_A_c_215_n N_A_M1057_g
+ N_A_c_216_n N_A_M1062_g N_A_c_225_n N_A_M1056_g A N_A_c_229_p N_A_c_217_n
+ PM_SKY130_FD_SC_HDLL__NOR4_8%A
x_PM_SKY130_FD_SC_HDLL__NOR4_8%B N_B_c_363_n N_B_M1005_g N_B_c_354_n N_B_M1002_g
+ N_B_c_355_n N_B_M1012_g N_B_c_364_n N_B_M1009_g N_B_c_365_n N_B_M1014_g
+ N_B_c_356_n N_B_M1020_g N_B_c_357_n N_B_M1024_g N_B_c_366_n N_B_M1035_g
+ N_B_c_367_n N_B_M1043_g N_B_c_358_n N_B_M1039_g N_B_c_359_n N_B_M1041_g
+ N_B_c_368_n N_B_M1047_g N_B_c_369_n N_B_M1053_g N_B_c_360_n N_B_M1052_g
+ N_B_c_361_n N_B_M1061_g N_B_c_370_n N_B_M1058_g B N_B_c_374_n N_B_c_362_n
+ PM_SKY130_FD_SC_HDLL__NOR4_8%B
x_PM_SKY130_FD_SC_HDLL__NOR4_8%C N_C_c_509_n N_C_M1001_g N_C_c_500_n N_C_M1004_g
+ N_C_c_501_n N_C_M1007_g N_C_c_510_n N_C_M1013_g N_C_c_511_n N_C_M1017_g
+ N_C_c_502_n N_C_M1015_g N_C_c_503_n N_C_M1028_g N_C_c_512_n N_C_M1021_g
+ N_C_c_513_n N_C_M1025_g N_C_c_504_n N_C_M1046_g N_C_c_505_n N_C_M1054_g
+ N_C_c_514_n N_C_M1034_g N_C_c_515_n N_C_M1050_g N_C_c_506_n N_C_M1055_g
+ N_C_c_507_n N_C_M1063_g N_C_c_516_n N_C_M1059_g C N_C_c_520_p N_C_c_508_n
+ PM_SKY130_FD_SC_HDLL__NOR4_8%C
x_PM_SKY130_FD_SC_HDLL__NOR4_8%D N_D_c_658_n N_D_M1006_g N_D_c_649_n N_D_M1010_g
+ N_D_c_650_n N_D_M1022_g N_D_c_659_n N_D_M1011_g N_D_c_660_n N_D_M1023_g
+ N_D_c_651_n N_D_M1027_g N_D_c_652_n N_D_M1030_g N_D_c_661_n N_D_M1029_g
+ N_D_c_662_n N_D_M1036_g N_D_c_653_n N_D_M1033_g N_D_c_654_n N_D_M1042_g
+ N_D_c_663_n N_D_M1037_g N_D_c_664_n N_D_M1044_g N_D_c_655_n N_D_M1048_g
+ N_D_c_656_n N_D_M1049_g N_D_c_665_n N_D_M1060_g D N_D_c_704_p N_D_c_657_n
+ PM_SKY130_FD_SC_HDLL__NOR4_8%D
x_PM_SKY130_FD_SC_HDLL__NOR4_8%A_27_297# N_A_27_297#_M1000_d N_A_27_297#_M1003_d
+ N_A_27_297#_M1016_d N_A_27_297#_M1032_d N_A_27_297#_M1056_d
+ N_A_27_297#_M1009_d N_A_27_297#_M1035_d N_A_27_297#_M1047_d
+ N_A_27_297#_M1058_d N_A_27_297#_c_789_n N_A_27_297#_c_790_n
+ N_A_27_297#_c_791_n N_A_27_297#_c_842_p N_A_27_297#_c_792_n
+ N_A_27_297#_c_844_p N_A_27_297#_c_793_n N_A_27_297#_c_846_p
+ N_A_27_297#_c_794_n N_A_27_297#_c_795_n N_A_27_297#_c_849_p
+ N_A_27_297#_c_829_n N_A_27_297#_c_884_p N_A_27_297#_c_831_n
+ N_A_27_297#_c_888_p N_A_27_297#_c_833_n N_A_27_297#_c_892_p
+ N_A_27_297#_c_796_n N_A_27_297#_c_797_n N_A_27_297#_c_798_n
+ N_A_27_297#_c_799_n N_A_27_297#_c_800_n N_A_27_297#_c_854_p
+ N_A_27_297#_c_855_p N_A_27_297#_c_856_p PM_SKY130_FD_SC_HDLL__NOR4_8%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_8%VPWR N_VPWR_M1000_s N_VPWR_M1008_s N_VPWR_M1026_s
+ N_VPWR_M1040_s N_VPWR_c_908_n N_VPWR_c_909_n N_VPWR_c_910_n N_VPWR_c_911_n
+ N_VPWR_c_912_n N_VPWR_c_913_n N_VPWR_c_914_n VPWR N_VPWR_c_915_n
+ N_VPWR_c_916_n N_VPWR_c_907_n N_VPWR_c_918_n N_VPWR_c_919_n N_VPWR_c_920_n
+ N_VPWR_c_921_n VPWR PM_SKY130_FD_SC_HDLL__NOR4_8%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4_8%A_869_297# N_A_869_297#_M1005_s
+ N_A_869_297#_M1014_s N_A_869_297#_M1043_s N_A_869_297#_M1053_s
+ N_A_869_297#_M1001_d N_A_869_297#_M1017_d N_A_869_297#_M1025_d
+ N_A_869_297#_M1050_d N_A_869_297#_c_1090_n N_A_869_297#_c_1091_n
+ N_A_869_297#_c_1092_n N_A_869_297#_c_1093_n N_A_869_297#_c_1094_n
+ N_A_869_297#_c_1095_n N_A_869_297#_c_1096_n N_A_869_297#_c_1097_n
+ N_A_869_297#_c_1098_n N_A_869_297#_c_1099_n N_A_869_297#_c_1100_n
+ N_A_869_297#_c_1101_n N_A_869_297#_c_1102_n N_A_869_297#_c_1103_n
+ N_A_869_297#_c_1104_n PM_SKY130_FD_SC_HDLL__NOR4_8%A_869_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_8%A_1635_297# N_A_1635_297#_M1001_s
+ N_A_1635_297#_M1013_s N_A_1635_297#_M1021_s N_A_1635_297#_M1034_s
+ N_A_1635_297#_M1059_s N_A_1635_297#_M1011_d N_A_1635_297#_M1029_d
+ N_A_1635_297#_M1037_d N_A_1635_297#_M1060_d N_A_1635_297#_c_1210_n
+ N_A_1635_297#_c_1215_n N_A_1635_297#_c_1211_n N_A_1635_297#_c_1217_n
+ N_A_1635_297#_c_1219_n N_A_1635_297#_c_1296_n N_A_1635_297#_c_1221_n
+ N_A_1635_297#_c_1301_n N_A_1635_297#_c_1223_n N_A_1635_297#_c_1212_n
+ N_A_1635_297#_c_1228_n N_A_1635_297#_c_1313_p N_A_1635_297#_c_1230_n
+ N_A_1635_297#_c_1317_p N_A_1635_297#_c_1232_n N_A_1635_297#_c_1321_p
+ N_A_1635_297#_c_1234_n N_A_1635_297#_c_1213_n N_A_1635_297#_c_1214_n
+ N_A_1635_297#_c_1226_n N_A_1635_297#_c_1270_n N_A_1635_297#_c_1272_n
+ N_A_1635_297#_c_1274_n N_A_1635_297#_c_1276_n N_A_1635_297#_c_1278_n
+ N_A_1635_297#_c_1280_n PM_SKY130_FD_SC_HDLL__NOR4_8%A_1635_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_8%Y N_Y_M1018_s N_Y_M1031_s N_Y_M1045_s N_Y_M1057_s
+ N_Y_M1002_d N_Y_M1020_d N_Y_M1039_d N_Y_M1052_d N_Y_M1004_d N_Y_M1015_d
+ N_Y_M1046_d N_Y_M1055_d N_Y_M1010_d N_Y_M1027_d N_Y_M1033_d N_Y_M1048_d
+ N_Y_M1006_s N_Y_M1023_s N_Y_M1036_s N_Y_M1044_s N_Y_c_1368_n N_Y_c_1330_n
+ N_Y_c_1331_n N_Y_c_1379_n N_Y_c_1332_n N_Y_c_1387_n N_Y_c_1333_n N_Y_c_1395_n
+ N_Y_c_1334_n N_Y_c_1401_n N_Y_c_1335_n N_Y_c_1425_n N_Y_c_1336_n N_Y_c_1433_n
+ N_Y_c_1337_n N_Y_c_1441_n N_Y_c_1338_n N_Y_c_1466_n N_Y_c_1339_n N_Y_c_1473_n
+ N_Y_c_1340_n N_Y_c_1481_n N_Y_c_1341_n N_Y_c_1489_n N_Y_c_1342_n N_Y_c_1495_n
+ N_Y_c_1343_n N_Y_c_1361_n N_Y_c_1527_n N_Y_c_1362_n N_Y_c_1344_n N_Y_c_1539_n
+ N_Y_c_1363_n N_Y_c_1345_n N_Y_c_1552_n N_Y_c_1346_n N_Y_c_1347_n N_Y_c_1348_n
+ N_Y_c_1349_n N_Y_c_1350_n N_Y_c_1351_n N_Y_c_1352_n N_Y_c_1353_n N_Y_c_1354_n
+ N_Y_c_1355_n N_Y_c_1356_n N_Y_c_1357_n N_Y_c_1557_n N_Y_c_1358_n N_Y_c_1364_n
+ N_Y_c_1359_n N_Y_c_1365_n N_Y_c_1366_n Y PM_SKY130_FD_SC_HDLL__NOR4_8%Y
x_PM_SKY130_FD_SC_HDLL__NOR4_8%VGND N_VGND_M1018_d N_VGND_M1019_d N_VGND_M1038_d
+ N_VGND_M1051_d N_VGND_M1062_d N_VGND_M1012_s N_VGND_M1024_s N_VGND_M1041_s
+ N_VGND_M1061_s N_VGND_M1007_s N_VGND_M1028_s N_VGND_M1054_s N_VGND_M1063_s
+ N_VGND_M1022_s N_VGND_M1030_s N_VGND_M1042_s N_VGND_M1049_s N_VGND_c_1738_n
+ N_VGND_c_1739_n N_VGND_c_1740_n N_VGND_c_1741_n N_VGND_c_1742_n
+ N_VGND_c_1743_n N_VGND_c_1744_n N_VGND_c_1745_n N_VGND_c_1746_n
+ N_VGND_c_1747_n N_VGND_c_1748_n N_VGND_c_1749_n N_VGND_c_1750_n
+ N_VGND_c_1751_n N_VGND_c_1752_n N_VGND_c_1753_n N_VGND_c_1754_n
+ N_VGND_c_1755_n N_VGND_c_1756_n N_VGND_c_1757_n N_VGND_c_1758_n
+ N_VGND_c_1759_n N_VGND_c_1760_n N_VGND_c_1761_n N_VGND_c_1762_n
+ N_VGND_c_1763_n N_VGND_c_1764_n N_VGND_c_1765_n N_VGND_c_1766_n
+ N_VGND_c_1767_n N_VGND_c_1768_n N_VGND_c_1769_n N_VGND_c_1770_n
+ N_VGND_c_1771_n N_VGND_c_1772_n N_VGND_c_1773_n N_VGND_c_1774_n
+ N_VGND_c_1775_n N_VGND_c_1776_n N_VGND_c_1777_n VGND N_VGND_c_1778_n
+ N_VGND_c_1779_n N_VGND_c_1780_n N_VGND_c_1781_n N_VGND_c_1782_n
+ N_VGND_c_1783_n N_VGND_c_1784_n N_VGND_c_1785_n N_VGND_c_1786_n
+ N_VGND_c_1787_n PM_SKY130_FD_SC_HDLL__NOR4_8%VGND
cc_1 VNB N_A_c_209_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_c_210_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_3 VNB N_A_c_211_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_A_c_212_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_5 VNB N_A_c_213_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_6 VNB N_A_c_214_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_7 VNB N_A_c_215_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=3.34 $Y2=0.995
cc_8 VNB N_A_c_216_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.995
cc_9 VNB N_A_c_217_n 0.163659f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.202
cc_10 VNB N_B_c_354_n 0.0168874f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_11 VNB N_B_c_355_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_12 VNB N_B_c_356_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_13 VNB N_B_c_357_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_14 VNB N_B_c_358_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_15 VNB N_B_c_359_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_16 VNB N_B_c_360_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=3.34 $Y2=0.995
cc_17 VNB N_B_c_361_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.995
cc_18 VNB N_B_c_362_n 0.162173f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.202
cc_19 VNB N_C_c_500_n 0.0214896f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_20 VNB N_C_c_501_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_21 VNB N_C_c_502_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_22 VNB N_C_c_503_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_23 VNB N_C_c_504_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_24 VNB N_C_c_505_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_25 VNB N_C_c_506_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=3.34 $Y2=0.995
cc_26 VNB N_C_c_507_n 0.0168583f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.995
cc_27 VNB N_C_c_508_n 0.16218f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.202
cc_28 VNB N_D_c_649_n 0.0168604f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_29 VNB N_D_c_650_n 0.0163313f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.995
cc_30 VNB N_D_c_651_n 0.0166841f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_31 VNB N_D_c_652_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.995
cc_32 VNB N_D_c_653_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.4 $Y2=0.995
cc_33 VNB N_D_c_654_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=0.995
cc_34 VNB N_D_c_655_n 0.0167214f $X=-0.19 $Y=-0.24 $X2=3.34 $Y2=0.995
cc_35 VNB N_D_c_656_n 0.0213647f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.995
cc_36 VNB N_D_c_657_n 0.164137f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.202
cc_37 VNB N_VPWR_c_907_n 0.668254f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_38 VNB N_Y_c_1330_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.202
cc_39 VNB N_Y_c_1331_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.202
cc_40 VNB N_Y_c_1332_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=1.202
cc_41 VNB N_Y_c_1333_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=3.63 $Y2=1.18
cc_42 VNB N_Y_c_1334_n 0.005207f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_1335_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_Y_c_1336_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_Y_c_1337_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_Y_c_1338_n 0.0130165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_Y_c_1339_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_Y_c_1340_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_Y_c_1341_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_Y_c_1342_n 0.005457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_Y_c_1343_n 0.00328943f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_Y_c_1344_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_Y_c_1345_n 0.00569435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_Y_c_1346_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_Y_c_1347_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_Y_c_1348_n 0.00222524f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_Y_c_1349_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_Y_c_1350_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_Y_c_1351_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_Y_c_1352_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_Y_c_1353_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_Y_c_1354_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_Y_c_1355_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_Y_c_1356_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_Y_c_1357_n 4.05044e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_Y_c_1358_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_Y_c_1359_n 0.00222525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB Y 8.94272e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_1738_n 0.011505f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_70 VNB N_VGND_c_1739_n 0.00967f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.16
cc_71 VNB N_VGND_c_1740_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.202
cc_72 VNB N_VGND_c_1741_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.202
cc_73 VNB N_VGND_c_1742_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=2.82 $Y2=1.202
cc_74 VNB N_VGND_c_1743_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.202
cc_75 VNB N_VGND_c_1744_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=3.63 $Y2=1.16
cc_76 VNB N_VGND_c_1745_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.202
cc_77 VNB N_VGND_c_1746_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1747_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1748_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1749_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1750_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1751_n 0.00413904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1752_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1753_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1754_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1755_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1756_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1757_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1758_n 0.0118897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1759_n 0.0342987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1760_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1761_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1762_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1763_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1764_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1765_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1766_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1767_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1768_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1769_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1770_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1771_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1772_n 0.0166675f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1773_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1774_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1775_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1776_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1777_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1778_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1779_n 0.0173087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1780_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1781_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1782_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1783_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1784_n 0.00515916f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1785_n 0.0166684f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_VGND_c_1786_n 0.0222052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_VGND_c_1787_n 0.716369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VPB N_A_c_218_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_120 VPB N_A_c_219_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_121 VPB N_A_c_220_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_122 VPB N_A_c_221_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_123 VPB N_A_c_222_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_124 VPB N_A_c_223_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_125 VPB N_A_c_224_n 0.0159747f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_126 VPB N_A_c_225_n 0.0161064f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_127 VPB N_A_c_217_n 0.0999345f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.202
cc_128 VPB N_B_c_363_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_129 VPB N_B_c_364_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_130 VPB N_B_c_365_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_131 VPB N_B_c_366_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_132 VPB N_B_c_367_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_133 VPB N_B_c_368_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_134 VPB N_B_c_369_n 0.0159747f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_135 VPB N_B_c_370_n 0.0203443f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_136 VPB N_B_c_362_n 0.100818f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.202
cc_137 VPB N_C_c_509_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_138 VPB N_C_c_510_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_139 VPB N_C_c_511_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_140 VPB N_C_c_512_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_141 VPB N_C_c_513_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_142 VPB N_C_c_514_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_143 VPB N_C_c_515_n 0.0159747f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_144 VPB N_C_c_516_n 0.0164209f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_145 VPB N_C_c_508_n 0.100813f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.202
cc_146 VPB N_D_c_658_n 0.0164077f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_147 VPB N_D_c_659_n 0.015773f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_148 VPB N_D_c_660_n 0.0159513f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_149 VPB N_D_c_661_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_150 VPB N_D_c_662_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_151 VPB N_D_c_663_n 0.0159747f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_152 VPB N_D_c_664_n 0.0159747f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_153 VPB N_D_c_665_n 0.0205492f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_154 VPB N_D_c_657_n 0.102316f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=1.202
cc_155 VPB N_A_27_297#_c_789_n 0.0327625f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.56
cc_156 VPB N_A_27_297#_c_790_n 0.0018222f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_157 VPB N_A_27_297#_c_791_n 0.0130892f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_158 VPB N_A_27_297#_c_792_n 0.00193318f $X=-0.19 $Y=1.305 $X2=3.34 $Y2=0.995
cc_159 VPB N_A_27_297#_c_793_n 0.00193318f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_160 VPB N_A_27_297#_c_794_n 0.00204701f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_161 VPB N_A_27_297#_c_795_n 0.00416602f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.16
cc_162 VPB N_A_27_297#_c_796_n 0.00180756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_A_27_297#_c_797_n 0.00482315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_A_27_297#_c_798_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_A_27_297#_c_799_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_27_297#_c_800_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_908_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_168 VPB N_VPWR_c_909_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_169 VPB N_VPWR_c_910_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.56
cc_170 VPB N_VPWR_c_911_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_171 VPB N_VPWR_c_912_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.985
cc_172 VPB N_VPWR_c_913_n 0.0195604f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.56
cc_173 VPB N_VPWR_c_914_n 0.00516582f $X=-0.19 $Y=1.305 $X2=2.82 $Y2=0.56
cc_174 VPB N_VPWR_c_915_n 0.0181841f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_175 VPB N_VPWR_c_916_n 0.282246f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.985
cc_176 VPB N_VPWR_c_907_n 0.0553493f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.985
cc_177 VPB N_VPWR_c_918_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_178 VPB N_VPWR_c_919_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.16
cc_179 VPB N_VPWR_c_920_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_180 VPB N_VPWR_c_921_n 0.0047828f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.202
cc_181 VPB N_A_869_297#_c_1090_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.375
+ $Y2=1.985
cc_182 VPB N_A_869_297#_c_1091_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.82
+ $Y2=0.995
cc_183 VPB N_A_869_297#_c_1092_n 0.00193318f $X=-0.19 $Y=1.305 $X2=2.845
+ $Y2=1.985
cc_184 VPB N_A_869_297#_c_1093_n 0.0215869f $X=-0.19 $Y=1.305 $X2=3.315
+ $Y2=1.985
cc_185 VPB N_A_869_297#_c_1094_n 0.00193318f $X=-0.19 $Y=1.305 $X2=3.76
+ $Y2=0.995
cc_186 VPB N_A_869_297#_c_1095_n 0.00193318f $X=-0.19 $Y=1.305 $X2=3.785
+ $Y2=1.985
cc_187 VPB N_A_869_297#_c_1096_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0.495
+ $Y2=1.202
cc_188 VPB N_A_869_297#_c_1097_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0.94
+ $Y2=1.202
cc_189 VPB N_A_869_297#_c_1098_n 0.00149756f $X=-0.19 $Y=1.305 $X2=1.435
+ $Y2=1.202
cc_190 VPB N_A_869_297#_c_1099_n 0.00149756f $X=-0.19 $Y=1.305 $X2=1.88
+ $Y2=1.202
cc_191 VPB N_A_869_297#_c_1100_n 0.00149756f $X=-0.19 $Y=1.305 $X2=2.375
+ $Y2=1.202
cc_192 VPB N_A_869_297#_c_1101_n 0.00149756f $X=-0.19 $Y=1.305 $X2=2.82
+ $Y2=1.202
cc_193 VPB N_A_869_297#_c_1102_n 0.00149756f $X=-0.19 $Y=1.305 $X2=3.315
+ $Y2=1.202
cc_194 VPB N_A_869_297#_c_1103_n 0.00149756f $X=-0.19 $Y=1.305 $X2=3.63
+ $Y2=1.202
cc_195 VPB N_A_869_297#_c_1104_n 0.00175152f $X=-0.19 $Y=1.305 $X2=3.63 $Y2=1.16
cc_196 VPB N_A_1635_297#_c_1210_n 0.00482315f $X=-0.19 $Y=1.305 $X2=2.4 $Y2=0.56
cc_197 VPB N_A_1635_297#_c_1211_n 0.00180756f $X=-0.19 $Y=1.305 $X2=2.82
+ $Y2=0.56
cc_198 VPB N_A_1635_297#_c_1212_n 0.0044883f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=1.16
cc_199 VPB N_A_1635_297#_c_1213_n 0.00746643f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_1635_297#_c_1214_n 0.037497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_Y_c_1361_n 0.00208662f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_Y_c_1362_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_Y_c_1363_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_Y_c_1364_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_Y_c_1365_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_Y_c_1366_n 0.00201963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB Y 0.00129652f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 N_A_c_225_n N_B_c_363_n 0.00971598f $X=3.785 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_209 N_A_c_216_n N_B_c_354_n 0.0179509f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_210 N_A_c_229_p N_B_c_374_n 0.00795414f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_211 N_A_c_217_n N_B_c_374_n 8.31714e-19 $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_212 N_A_c_229_p N_B_c_362_n 8.31714e-19 $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A_c_217_n N_B_c_362_n 0.0237215f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_214 N_A_c_218_n N_A_27_297#_c_789_n 0.0106975f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_c_219_n N_A_27_297#_c_789_n 6.18277e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_216 N_A_c_218_n N_A_27_297#_c_790_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_219_n N_A_27_297#_c_790_n 0.0156273f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_229_p N_A_27_297#_c_790_n 0.0458726f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_c_217_n N_A_27_297#_c_790_n 0.00827579f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_220 N_A_c_218_n N_A_27_297#_c_791_n 0.001185f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_c_229_p N_A_27_297#_c_791_n 0.001546f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_222 N_A_c_217_n N_A_27_297#_c_791_n 5.21847e-19 $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_223 N_A_c_220_n N_A_27_297#_c_792_n 0.0156273f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_221_n N_A_27_297#_c_792_n 0.0156273f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_229_p N_A_27_297#_c_792_n 0.0486996f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_226 N_A_c_217_n N_A_27_297#_c_792_n 0.00885494f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_227 N_A_c_222_n N_A_27_297#_c_793_n 0.0156273f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_223_n N_A_27_297#_c_793_n 0.0156273f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_c_229_p N_A_27_297#_c_793_n 0.0486996f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_230 N_A_c_217_n N_A_27_297#_c_793_n 0.00885494f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_231 N_A_c_224_n N_A_27_297#_c_794_n 0.0156273f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_c_225_n N_A_27_297#_c_794_n 0.0164448f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_c_229_p N_A_27_297#_c_794_n 0.0417725f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_234 N_A_c_217_n N_A_27_297#_c_794_n 0.00859761f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_235 N_A_c_229_p N_A_27_297#_c_798_n 0.0204509f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_c_217_n N_A_27_297#_c_798_n 0.00635938f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_237 N_A_c_229_p N_A_27_297#_c_799_n 0.0204509f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_c_217_n N_A_27_297#_c_799_n 0.00635938f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_239 N_A_c_229_p N_A_27_297#_c_800_n 0.0204509f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_c_217_n N_A_27_297#_c_800_n 0.00635938f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_c_218_n N_VPWR_c_908_n 0.00300743f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_c_219_n N_VPWR_c_908_n 0.00300743f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_c_219_n N_VPWR_c_909_n 0.00702461f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_c_220_n N_VPWR_c_909_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_c_220_n N_VPWR_c_910_n 0.00300743f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_221_n N_VPWR_c_910_n 0.00300743f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_221_n N_VPWR_c_911_n 0.00702461f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_248 N_A_c_222_n N_VPWR_c_911_n 0.00702461f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A_c_222_n N_VPWR_c_912_n 0.00300743f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_c_223_n N_VPWR_c_912_n 0.00300743f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_c_223_n N_VPWR_c_913_n 0.00702461f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_224_n N_VPWR_c_913_n 0.00702461f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_224_n N_VPWR_c_914_n 0.00300743f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_254 N_A_c_225_n N_VPWR_c_914_n 0.00300743f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_c_218_n N_VPWR_c_915_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_c_225_n N_VPWR_c_916_n 0.00702461f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_c_218_n N_VPWR_c_907_n 0.0126549f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_219_n N_VPWR_c_907_n 0.0124092f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_c_220_n N_VPWR_c_907_n 0.0124092f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_221_n N_VPWR_c_907_n 0.0124092f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_222_n N_VPWR_c_907_n 0.0124092f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_223_n N_VPWR_c_907_n 0.0124092f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_224_n N_VPWR_c_907_n 0.0124092f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_225_n N_VPWR_c_907_n 0.0124344f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_209_n N_Y_c_1368_n 0.00539651f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_c_210_n N_Y_c_1368_n 0.00671723f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_211_n N_Y_c_1368_n 5.24636e-19 $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_c_210_n N_Y_c_1330_n 0.00929182f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_c_211_n N_Y_c_1330_n 0.00929182f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_c_229_p N_Y_c_1330_n 0.0435408f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_c_217_n N_Y_c_1330_n 0.00468948f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_272 N_A_c_209_n N_Y_c_1331_n 0.00262807f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_c_210_n N_Y_c_1331_n 0.00113286f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_c_229_p N_Y_c_1331_n 0.0266272f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_c_217_n N_Y_c_1331_n 0.00230339f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_276 N_A_c_210_n N_Y_c_1379_n 5.24636e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_277 N_A_c_211_n N_Y_c_1379_n 0.00671723f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_278 N_A_c_212_n N_Y_c_1379_n 0.00671723f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_279 N_A_c_213_n N_Y_c_1379_n 5.24636e-19 $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_280 N_A_c_212_n N_Y_c_1332_n 0.00929182f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_281 N_A_c_213_n N_Y_c_1332_n 0.00929182f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_282 N_A_c_229_p N_Y_c_1332_n 0.0435408f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_c_217_n N_Y_c_1332_n 0.00468948f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_284 N_A_c_212_n N_Y_c_1387_n 5.24636e-19 $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_285 N_A_c_213_n N_Y_c_1387_n 0.00671723f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_286 N_A_c_214_n N_Y_c_1387_n 0.00671723f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_287 N_A_c_215_n N_Y_c_1387_n 5.24636e-19 $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_288 N_A_c_214_n N_Y_c_1333_n 0.00929182f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_289 N_A_c_215_n N_Y_c_1333_n 0.00929182f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_290 N_A_c_229_p N_Y_c_1333_n 0.0435408f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_291 N_A_c_217_n N_Y_c_1333_n 0.00468948f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_292 N_A_c_214_n N_Y_c_1395_n 5.24636e-19 $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A_c_215_n N_Y_c_1395_n 0.00671723f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A_c_216_n N_Y_c_1395_n 0.00671723f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A_c_216_n N_Y_c_1334_n 0.00972073f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A_c_229_p N_Y_c_1334_n 0.00550176f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_297 N_A_c_217_n N_Y_c_1334_n 0.00164699f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_298 N_A_c_216_n N_Y_c_1401_n 5.24636e-19 $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A_c_211_n N_Y_c_1346_n 0.00113286f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A_c_212_n N_Y_c_1346_n 0.00113286f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_301 N_A_c_229_p N_Y_c_1346_n 0.0266272f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_302 N_A_c_217_n N_Y_c_1346_n 0.00230339f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_303 N_A_c_213_n N_Y_c_1347_n 0.00113286f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A_c_214_n N_Y_c_1347_n 0.00113286f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_c_229_p N_Y_c_1347_n 0.0266272f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_306 N_A_c_217_n N_Y_c_1347_n 0.00230339f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_307 N_A_c_215_n N_Y_c_1348_n 0.00113286f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_216_n N_Y_c_1348_n 0.00113286f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_c_229_p N_Y_c_1348_n 0.0266272f $X=3.63 $Y=1.16 $X2=0 $Y2=0
cc_310 N_A_c_217_n N_Y_c_1348_n 0.00230339f $X=3.76 $Y=1.202 $X2=0 $Y2=0
cc_311 N_A_c_209_n N_VGND_c_1739_n 0.00366155f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A_c_210_n N_VGND_c_1740_n 0.00166854f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A_c_211_n N_VGND_c_1740_n 0.00166854f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_c_211_n N_VGND_c_1741_n 0.00423334f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A_c_212_n N_VGND_c_1741_n 0.00423334f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_c_212_n N_VGND_c_1742_n 0.00166854f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_c_213_n N_VGND_c_1742_n 0.00166854f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A_c_213_n N_VGND_c_1743_n 0.00423334f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_214_n N_VGND_c_1743_n 0.00423334f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_214_n N_VGND_c_1744_n 0.00166854f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_c_215_n N_VGND_c_1744_n 0.00166854f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_c_215_n N_VGND_c_1745_n 0.00423334f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_c_216_n N_VGND_c_1745_n 0.00423334f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_c_216_n N_VGND_c_1746_n 0.00166854f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_c_209_n N_VGND_c_1778_n 0.00541359f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_c_210_n N_VGND_c_1778_n 0.00423334f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_c_209_n N_VGND_c_1787_n 0.0105004f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_c_210_n N_VGND_c_1787_n 0.00595861f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_c_211_n N_VGND_c_1787_n 0.00595861f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_c_212_n N_VGND_c_1787_n 0.00595861f $X=1.88 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_c_213_n N_VGND_c_1787_n 0.00595861f $X=2.4 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_c_214_n N_VGND_c_1787_n 0.00595861f $X=2.82 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_c_215_n N_VGND_c_1787_n 0.00595861f $X=3.34 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_c_216_n N_VGND_c_1787_n 0.00596967f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_363_n N_A_27_297#_c_795_n 2.98195e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_336 N_B_c_363_n N_A_27_297#_c_829_n 0.0143578f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_337 N_B_c_364_n N_A_27_297#_c_829_n 0.01161f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_338 N_B_c_365_n N_A_27_297#_c_831_n 0.01161f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_339 N_B_c_366_n N_A_27_297#_c_831_n 0.01161f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_340 N_B_c_367_n N_A_27_297#_c_833_n 0.01161f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_341 N_B_c_368_n N_A_27_297#_c_833_n 0.01161f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_342 N_B_c_369_n N_A_27_297#_c_796_n 0.01161f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_343 N_B_c_370_n N_A_27_297#_c_796_n 0.01161f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_344 N_B_c_363_n N_VPWR_c_916_n 0.00429453f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_345 N_B_c_364_n N_VPWR_c_916_n 0.00429453f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_346 N_B_c_365_n N_VPWR_c_916_n 0.00429453f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_347 N_B_c_366_n N_VPWR_c_916_n 0.00429453f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_348 N_B_c_367_n N_VPWR_c_916_n 0.00429453f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_349 N_B_c_368_n N_VPWR_c_916_n 0.00429453f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_350 N_B_c_369_n N_VPWR_c_916_n 0.00429453f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_351 N_B_c_370_n N_VPWR_c_916_n 0.00429453f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_352 N_B_c_363_n N_VPWR_c_907_n 0.00609021f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_353 N_B_c_364_n N_VPWR_c_907_n 0.00606499f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_354 N_B_c_365_n N_VPWR_c_907_n 0.00606499f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_355 N_B_c_366_n N_VPWR_c_907_n 0.00606499f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_356 N_B_c_367_n N_VPWR_c_907_n 0.00606499f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_357 N_B_c_368_n N_VPWR_c_907_n 0.00606499f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_358 N_B_c_369_n N_VPWR_c_907_n 0.00606499f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_359 N_B_c_370_n N_VPWR_c_907_n 0.00734734f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_360 N_B_c_364_n N_A_869_297#_c_1090_n 0.0128188f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_361 N_B_c_365_n N_A_869_297#_c_1090_n 0.0128795f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_362 N_B_c_374_n N_A_869_297#_c_1090_n 0.0486996f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_363 N_B_c_362_n N_A_869_297#_c_1090_n 0.00844349f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_364 N_B_c_366_n N_A_869_297#_c_1091_n 0.0128795f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_365 N_B_c_367_n N_A_869_297#_c_1091_n 0.0128795f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_366 N_B_c_374_n N_A_869_297#_c_1091_n 0.0486996f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_367 N_B_c_362_n N_A_869_297#_c_1091_n 0.00844349f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_368 N_B_c_368_n N_A_869_297#_c_1092_n 0.0128795f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_369 N_B_c_369_n N_A_869_297#_c_1092_n 0.0128795f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_370 N_B_c_374_n N_A_869_297#_c_1092_n 0.0486996f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_371 N_B_c_362_n N_A_869_297#_c_1092_n 0.00844349f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_372 N_B_c_370_n N_A_869_297#_c_1093_n 0.0148794f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_373 N_B_c_374_n N_A_869_297#_c_1093_n 0.0138171f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_374 N_B_c_362_n N_A_869_297#_c_1093_n 9.00973e-19 $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_375 N_B_c_363_n N_A_869_297#_c_1097_n 2.98195e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_376 N_B_c_374_n N_A_869_297#_c_1097_n 0.0204252f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_377 N_B_c_362_n N_A_869_297#_c_1097_n 0.00675794f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_378 N_B_c_374_n N_A_869_297#_c_1098_n 0.0204252f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_379 N_B_c_362_n N_A_869_297#_c_1098_n 0.00675794f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_380 N_B_c_374_n N_A_869_297#_c_1099_n 0.0204252f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_381 N_B_c_362_n N_A_869_297#_c_1099_n 0.00675794f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_382 N_B_c_374_n N_A_869_297#_c_1100_n 0.0204252f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_383 N_B_c_362_n N_A_869_297#_c_1100_n 0.00675794f $X=7.52 $Y=1.202 $X2=0
+ $Y2=0
cc_384 N_B_c_354_n N_Y_c_1395_n 5.24636e-19 $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_385 N_B_c_354_n N_Y_c_1334_n 0.0104562f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_386 N_B_c_374_n N_Y_c_1334_n 0.00550176f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B_c_362_n N_Y_c_1334_n 0.00224539f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_388 N_B_c_354_n N_Y_c_1401_n 0.00671723f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_389 N_B_c_355_n N_Y_c_1401_n 0.00671723f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_390 N_B_c_356_n N_Y_c_1401_n 5.24636e-19 $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_391 N_B_c_355_n N_Y_c_1335_n 0.00929182f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_392 N_B_c_356_n N_Y_c_1335_n 0.00929182f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_393 N_B_c_374_n N_Y_c_1335_n 0.0435408f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_394 N_B_c_362_n N_Y_c_1335_n 0.00468948f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_395 N_B_c_355_n N_Y_c_1425_n 5.24636e-19 $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_396 N_B_c_356_n N_Y_c_1425_n 0.00671723f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_397 N_B_c_357_n N_Y_c_1425_n 0.00671723f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_398 N_B_c_358_n N_Y_c_1425_n 5.24636e-19 $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B_c_357_n N_Y_c_1336_n 0.00929182f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_400 N_B_c_358_n N_Y_c_1336_n 0.00929182f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_401 N_B_c_374_n N_Y_c_1336_n 0.0435408f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_402 N_B_c_362_n N_Y_c_1336_n 0.00468948f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_403 N_B_c_357_n N_Y_c_1433_n 5.24636e-19 $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_404 N_B_c_358_n N_Y_c_1433_n 0.00671723f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_405 N_B_c_359_n N_Y_c_1433_n 0.00671723f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_406 N_B_c_360_n N_Y_c_1433_n 5.24636e-19 $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B_c_359_n N_Y_c_1337_n 0.00929182f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_408 N_B_c_360_n N_Y_c_1337_n 0.00929182f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_409 N_B_c_374_n N_Y_c_1337_n 0.0435408f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_410 N_B_c_362_n N_Y_c_1337_n 0.00468948f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_411 N_B_c_359_n N_Y_c_1441_n 5.24636e-19 $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_412 N_B_c_360_n N_Y_c_1441_n 0.00671723f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_413 N_B_c_361_n N_Y_c_1441_n 0.0109565f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_414 N_B_c_361_n N_Y_c_1338_n 0.0109318f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_415 N_B_c_374_n N_Y_c_1338_n 0.0111883f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_416 N_B_c_362_n N_Y_c_1338_n 0.00146367f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_417 N_B_c_354_n N_Y_c_1349_n 0.00113286f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_418 N_B_c_355_n N_Y_c_1349_n 0.00113286f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_419 N_B_c_374_n N_Y_c_1349_n 0.0266272f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_420 N_B_c_362_n N_Y_c_1349_n 0.00230339f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_421 N_B_c_356_n N_Y_c_1350_n 0.00113286f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_422 N_B_c_357_n N_Y_c_1350_n 0.00113286f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_423 N_B_c_374_n N_Y_c_1350_n 0.0266272f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_424 N_B_c_362_n N_Y_c_1350_n 0.00230339f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_425 N_B_c_358_n N_Y_c_1351_n 0.00113286f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_426 N_B_c_359_n N_Y_c_1351_n 0.00113286f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_427 N_B_c_374_n N_Y_c_1351_n 0.0266272f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_428 N_B_c_362_n N_Y_c_1351_n 0.00230339f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_429 N_B_c_360_n N_Y_c_1352_n 0.00113286f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_430 N_B_c_361_n N_Y_c_1352_n 0.00113286f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_431 N_B_c_374_n N_Y_c_1352_n 0.0266272f $X=7.47 $Y=1.16 $X2=0 $Y2=0
cc_432 N_B_c_362_n N_Y_c_1352_n 0.00230339f $X=7.52 $Y=1.202 $X2=0 $Y2=0
cc_433 N_B_c_354_n N_VGND_c_1746_n 0.00166854f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_434 N_B_c_354_n N_VGND_c_1747_n 0.00423334f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_355_n N_VGND_c_1747_n 0.00423334f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_436 N_B_c_355_n N_VGND_c_1748_n 0.00166854f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_356_n N_VGND_c_1748_n 0.00166854f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_438 N_B_c_357_n N_VGND_c_1749_n 0.00166854f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_358_n N_VGND_c_1749_n 0.00166854f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B_c_359_n N_VGND_c_1750_n 0.00166854f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_360_n N_VGND_c_1750_n 0.00166738f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_356_n N_VGND_c_1760_n 0.00423334f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_357_n N_VGND_c_1760_n 0.00423334f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_444 N_B_c_358_n N_VGND_c_1762_n 0.00423334f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_359_n N_VGND_c_1762_n 0.00423334f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_446 N_B_c_360_n N_VGND_c_1785_n 0.00423334f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_c_361_n N_VGND_c_1785_n 0.00423334f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_448 N_B_c_361_n N_VGND_c_1786_n 0.00336547f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_449 N_B_c_354_n N_VGND_c_1787_n 0.00596967f $X=4.28 $Y=0.995 $X2=0 $Y2=0
cc_450 N_B_c_355_n N_VGND_c_1787_n 0.00595861f $X=4.7 $Y=0.995 $X2=0 $Y2=0
cc_451 N_B_c_356_n N_VGND_c_1787_n 0.00595861f $X=5.22 $Y=0.995 $X2=0 $Y2=0
cc_452 N_B_c_357_n N_VGND_c_1787_n 0.00595861f $X=5.64 $Y=0.995 $X2=0 $Y2=0
cc_453 N_B_c_358_n N_VGND_c_1787_n 0.00595861f $X=6.16 $Y=0.995 $X2=0 $Y2=0
cc_454 N_B_c_359_n N_VGND_c_1787_n 0.00595861f $X=6.58 $Y=0.995 $X2=0 $Y2=0
cc_455 N_B_c_360_n N_VGND_c_1787_n 0.00595861f $X=7.1 $Y=0.995 $X2=0 $Y2=0
cc_456 N_B_c_361_n N_VGND_c_1787_n 0.0070399f $X=7.52 $Y=0.995 $X2=0 $Y2=0
cc_457 N_C_c_516_n N_D_c_658_n 0.00937092f $X=11.825 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_458 N_C_c_507_n N_D_c_649_n 0.0175129f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_459 N_C_c_520_p N_D_c_657_n 8.6651e-19 $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_460 N_C_c_508_n N_D_c_657_n 0.0229666f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_461 N_C_c_509_n N_VPWR_c_916_n 0.00429453f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_462 N_C_c_510_n N_VPWR_c_916_n 0.00429425f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_463 N_C_c_511_n N_VPWR_c_916_n 0.00429453f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_464 N_C_c_512_n N_VPWR_c_916_n 0.00429453f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_465 N_C_c_513_n N_VPWR_c_916_n 0.00429453f $X=10.415 $Y=1.41 $X2=0 $Y2=0
cc_466 N_C_c_514_n N_VPWR_c_916_n 0.00429453f $X=10.885 $Y=1.41 $X2=0 $Y2=0
cc_467 N_C_c_515_n N_VPWR_c_916_n 0.00429453f $X=11.355 $Y=1.41 $X2=0 $Y2=0
cc_468 N_C_c_516_n N_VPWR_c_916_n 0.00429453f $X=11.825 $Y=1.41 $X2=0 $Y2=0
cc_469 N_C_c_509_n N_VPWR_c_907_n 0.00734734f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_470 N_C_c_510_n N_VPWR_c_907_n 0.00606497f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_471 N_C_c_511_n N_VPWR_c_907_n 0.00606499f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_472 N_C_c_512_n N_VPWR_c_907_n 0.00606499f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_473 N_C_c_513_n N_VPWR_c_907_n 0.00606499f $X=10.415 $Y=1.41 $X2=0 $Y2=0
cc_474 N_C_c_514_n N_VPWR_c_907_n 0.00606499f $X=10.885 $Y=1.41 $X2=0 $Y2=0
cc_475 N_C_c_515_n N_VPWR_c_907_n 0.00606499f $X=11.355 $Y=1.41 $X2=0 $Y2=0
cc_476 N_C_c_516_n N_VPWR_c_907_n 0.00609021f $X=11.825 $Y=1.41 $X2=0 $Y2=0
cc_477 N_C_c_509_n N_A_869_297#_c_1093_n 0.0148794f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_478 N_C_c_520_p N_A_869_297#_c_1093_n 0.0138171f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_479 N_C_c_508_n N_A_869_297#_c_1093_n 9.00973e-19 $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_480 N_C_c_510_n N_A_869_297#_c_1094_n 0.0125613f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_481 N_C_c_511_n N_A_869_297#_c_1094_n 0.0128795f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_482 N_C_c_520_p N_A_869_297#_c_1094_n 0.0486996f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_483 N_C_c_508_n N_A_869_297#_c_1094_n 0.00844349f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_484 N_C_c_512_n N_A_869_297#_c_1095_n 0.0128795f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_485 N_C_c_513_n N_A_869_297#_c_1095_n 0.0128795f $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_486 N_C_c_520_p N_A_869_297#_c_1095_n 0.0486996f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_487 N_C_c_508_n N_A_869_297#_c_1095_n 0.00844349f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_488 N_C_c_514_n N_A_869_297#_c_1096_n 0.0128795f $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_489 N_C_c_515_n N_A_869_297#_c_1096_n 0.0128188f $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_490 N_C_c_520_p N_A_869_297#_c_1096_n 0.0486996f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_491 N_C_c_508_n N_A_869_297#_c_1096_n 0.00844349f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_492 N_C_c_520_p N_A_869_297#_c_1101_n 0.0204252f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_493 N_C_c_508_n N_A_869_297#_c_1101_n 0.00675794f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_494 N_C_c_520_p N_A_869_297#_c_1102_n 0.0204252f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_495 N_C_c_508_n N_A_869_297#_c_1102_n 0.00675794f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_496 N_C_c_520_p N_A_869_297#_c_1103_n 0.0204252f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_497 N_C_c_508_n N_A_869_297#_c_1103_n 0.00675794f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_498 N_C_c_516_n N_A_869_297#_c_1104_n 2.98817e-19 $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_499 N_C_c_520_p N_A_869_297#_c_1104_n 0.0204252f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_500 N_C_c_508_n N_A_869_297#_c_1104_n 0.00675794f $X=11.8 $Y=1.202 $X2=0
+ $Y2=0
cc_501 N_C_c_509_n N_A_1635_297#_c_1215_n 0.01161f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_502 N_C_c_510_n N_A_1635_297#_c_1215_n 0.0105438f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_503 N_C_c_509_n N_A_1635_297#_c_1217_n 5.289e-19 $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_504 N_C_c_510_n N_A_1635_297#_c_1217_n 0.00714881f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_505 N_C_c_511_n N_A_1635_297#_c_1219_n 0.01161f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_506 N_C_c_512_n N_A_1635_297#_c_1219_n 0.01161f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_507 N_C_c_513_n N_A_1635_297#_c_1221_n 0.01161f $X=10.415 $Y=1.41 $X2=0 $Y2=0
cc_508 N_C_c_514_n N_A_1635_297#_c_1221_n 0.01161f $X=10.885 $Y=1.41 $X2=0 $Y2=0
cc_509 N_C_c_515_n N_A_1635_297#_c_1223_n 0.01161f $X=11.355 $Y=1.41 $X2=0 $Y2=0
cc_510 N_C_c_516_n N_A_1635_297#_c_1223_n 0.0143578f $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_511 N_C_c_516_n N_A_1635_297#_c_1212_n 2.65342e-19 $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_512 N_C_c_510_n N_A_1635_297#_c_1226_n 4.58352e-19 $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_513 N_C_c_500_n N_Y_c_1338_n 0.0109318f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_514 N_C_c_520_p N_Y_c_1338_n 0.0111883f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_515 N_C_c_508_n N_Y_c_1338_n 0.00146367f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_516 N_C_c_500_n N_Y_c_1466_n 0.0109565f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_517 N_C_c_501_n N_Y_c_1466_n 0.00671723f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_518 N_C_c_502_n N_Y_c_1466_n 5.24636e-19 $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_519 N_C_c_501_n N_Y_c_1339_n 0.00929182f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_520 N_C_c_502_n N_Y_c_1339_n 0.00929182f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_521 N_C_c_520_p N_Y_c_1339_n 0.0435408f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_522 N_C_c_508_n N_Y_c_1339_n 0.00468948f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_523 N_C_c_501_n N_Y_c_1473_n 5.24636e-19 $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_524 N_C_c_502_n N_Y_c_1473_n 0.00671723f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_525 N_C_c_503_n N_Y_c_1473_n 0.00671723f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_526 N_C_c_504_n N_Y_c_1473_n 5.24636e-19 $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_527 N_C_c_503_n N_Y_c_1340_n 0.00929182f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_528 N_C_c_504_n N_Y_c_1340_n 0.00929182f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_529 N_C_c_520_p N_Y_c_1340_n 0.0435408f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_530 N_C_c_508_n N_Y_c_1340_n 0.00468948f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_531 N_C_c_503_n N_Y_c_1481_n 5.24636e-19 $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_532 N_C_c_504_n N_Y_c_1481_n 0.00671723f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_533 N_C_c_505_n N_Y_c_1481_n 0.00671723f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_534 N_C_c_506_n N_Y_c_1481_n 5.24636e-19 $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_535 N_C_c_505_n N_Y_c_1341_n 0.00929182f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_536 N_C_c_506_n N_Y_c_1341_n 0.00929182f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_537 N_C_c_520_p N_Y_c_1341_n 0.0435408f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_538 N_C_c_508_n N_Y_c_1341_n 0.00468948f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_539 N_C_c_505_n N_Y_c_1489_n 5.24636e-19 $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_540 N_C_c_506_n N_Y_c_1489_n 0.00671723f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_541 N_C_c_507_n N_Y_c_1489_n 0.00671723f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_542 N_C_c_507_n N_Y_c_1342_n 0.0104562f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_543 N_C_c_520_p N_Y_c_1342_n 0.00550176f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_544 N_C_c_508_n N_Y_c_1342_n 0.00224539f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_545 N_C_c_507_n N_Y_c_1495_n 5.24636e-19 $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_546 N_C_c_500_n N_Y_c_1353_n 0.00113286f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_547 N_C_c_501_n N_Y_c_1353_n 0.00113286f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_548 N_C_c_520_p N_Y_c_1353_n 0.0266272f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_549 N_C_c_508_n N_Y_c_1353_n 0.00230339f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_550 N_C_c_502_n N_Y_c_1354_n 0.00113286f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_551 N_C_c_503_n N_Y_c_1354_n 0.00113286f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_552 N_C_c_520_p N_Y_c_1354_n 0.0266272f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_553 N_C_c_508_n N_Y_c_1354_n 0.00230339f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_554 N_C_c_504_n N_Y_c_1355_n 0.00113286f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_555 N_C_c_505_n N_Y_c_1355_n 0.00113286f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_556 N_C_c_520_p N_Y_c_1355_n 0.0266272f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_557 N_C_c_508_n N_Y_c_1355_n 0.00230339f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_558 N_C_c_506_n N_Y_c_1356_n 0.00113286f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_559 N_C_c_507_n N_Y_c_1356_n 0.00113286f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_560 N_C_c_520_p N_Y_c_1356_n 0.0266272f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_561 N_C_c_508_n N_Y_c_1356_n 0.00230339f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_562 N_C_c_520_p Y 0.00620594f $X=11.67 $Y=1.16 $X2=0 $Y2=0
cc_563 N_C_c_508_n Y 0.00129488f $X=11.8 $Y=1.202 $X2=0 $Y2=0
cc_564 N_C_c_501_n N_VGND_c_1751_n 0.00166738f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_565 N_C_c_502_n N_VGND_c_1751_n 0.00166854f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_566 N_C_c_503_n N_VGND_c_1752_n 0.00166854f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_567 N_C_c_504_n N_VGND_c_1752_n 0.00166854f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_568 N_C_c_505_n N_VGND_c_1753_n 0.00166854f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_569 N_C_c_506_n N_VGND_c_1753_n 0.00166854f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_570 N_C_c_507_n N_VGND_c_1754_n 0.00166854f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_571 N_C_c_500_n N_VGND_c_1764_n 0.00423334f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_572 N_C_c_501_n N_VGND_c_1764_n 0.00423334f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_573 N_C_c_502_n N_VGND_c_1766_n 0.00423334f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_574 N_C_c_503_n N_VGND_c_1766_n 0.00423334f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_575 N_C_c_504_n N_VGND_c_1768_n 0.00423334f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_576 N_C_c_505_n N_VGND_c_1768_n 0.00423334f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_577 N_C_c_506_n N_VGND_c_1770_n 0.00423334f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_578 N_C_c_507_n N_VGND_c_1770_n 0.00423334f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_579 N_C_c_500_n N_VGND_c_1786_n 0.00336547f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_580 N_C_c_500_n N_VGND_c_1787_n 0.0070399f $X=8.56 $Y=0.995 $X2=0 $Y2=0
cc_581 N_C_c_501_n N_VGND_c_1787_n 0.00595861f $X=8.98 $Y=0.995 $X2=0 $Y2=0
cc_582 N_C_c_502_n N_VGND_c_1787_n 0.00595861f $X=9.5 $Y=0.995 $X2=0 $Y2=0
cc_583 N_C_c_503_n N_VGND_c_1787_n 0.00595861f $X=9.92 $Y=0.995 $X2=0 $Y2=0
cc_584 N_C_c_504_n N_VGND_c_1787_n 0.00595861f $X=10.44 $Y=0.995 $X2=0 $Y2=0
cc_585 N_C_c_505_n N_VGND_c_1787_n 0.00595861f $X=10.86 $Y=0.995 $X2=0 $Y2=0
cc_586 N_C_c_506_n N_VGND_c_1787_n 0.00595861f $X=11.38 $Y=0.995 $X2=0 $Y2=0
cc_587 N_C_c_507_n N_VGND_c_1787_n 0.00596967f $X=11.8 $Y=0.995 $X2=0 $Y2=0
cc_588 N_D_c_658_n N_VPWR_c_916_n 0.00429453f $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_589 N_D_c_659_n N_VPWR_c_916_n 0.00429453f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_590 N_D_c_660_n N_VPWR_c_916_n 0.00429453f $X=13.235 $Y=1.41 $X2=0 $Y2=0
cc_591 N_D_c_661_n N_VPWR_c_916_n 0.00429453f $X=13.705 $Y=1.41 $X2=0 $Y2=0
cc_592 N_D_c_662_n N_VPWR_c_916_n 0.00429453f $X=14.175 $Y=1.41 $X2=0 $Y2=0
cc_593 N_D_c_663_n N_VPWR_c_916_n 0.00429453f $X=14.645 $Y=1.41 $X2=0 $Y2=0
cc_594 N_D_c_664_n N_VPWR_c_916_n 0.00429453f $X=15.115 $Y=1.41 $X2=0 $Y2=0
cc_595 N_D_c_665_n N_VPWR_c_916_n 0.00429453f $X=15.585 $Y=1.41 $X2=0 $Y2=0
cc_596 N_D_c_658_n N_VPWR_c_907_n 0.00609021f $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_597 N_D_c_659_n N_VPWR_c_907_n 0.00606499f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_598 N_D_c_660_n N_VPWR_c_907_n 0.00606499f $X=13.235 $Y=1.41 $X2=0 $Y2=0
cc_599 N_D_c_661_n N_VPWR_c_907_n 0.00606499f $X=13.705 $Y=1.41 $X2=0 $Y2=0
cc_600 N_D_c_662_n N_VPWR_c_907_n 0.00606499f $X=14.175 $Y=1.41 $X2=0 $Y2=0
cc_601 N_D_c_663_n N_VPWR_c_907_n 0.00606499f $X=14.645 $Y=1.41 $X2=0 $Y2=0
cc_602 N_D_c_664_n N_VPWR_c_907_n 0.00606499f $X=15.115 $Y=1.41 $X2=0 $Y2=0
cc_603 N_D_c_665_n N_VPWR_c_907_n 0.00699455f $X=15.585 $Y=1.41 $X2=0 $Y2=0
cc_604 N_D_c_658_n N_A_1635_297#_c_1212_n 2.65342e-19 $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_605 N_D_c_658_n N_A_1635_297#_c_1228_n 0.0143578f $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_606 N_D_c_659_n N_A_1635_297#_c_1228_n 0.0115695f $X=12.765 $Y=1.41 $X2=0
+ $Y2=0
cc_607 N_D_c_660_n N_A_1635_297#_c_1230_n 0.01161f $X=13.235 $Y=1.41 $X2=0 $Y2=0
cc_608 N_D_c_661_n N_A_1635_297#_c_1230_n 0.01161f $X=13.705 $Y=1.41 $X2=0 $Y2=0
cc_609 N_D_c_662_n N_A_1635_297#_c_1232_n 0.01161f $X=14.175 $Y=1.41 $X2=0 $Y2=0
cc_610 N_D_c_663_n N_A_1635_297#_c_1232_n 0.01161f $X=14.645 $Y=1.41 $X2=0 $Y2=0
cc_611 N_D_c_664_n N_A_1635_297#_c_1234_n 0.01161f $X=15.115 $Y=1.41 $X2=0 $Y2=0
cc_612 N_D_c_665_n N_A_1635_297#_c_1234_n 0.0143578f $X=15.585 $Y=1.41 $X2=0
+ $Y2=0
cc_613 N_D_c_665_n N_A_1635_297#_c_1214_n 4.96615e-19 $X=15.585 $Y=1.41 $X2=0
+ $Y2=0
cc_614 N_D_c_649_n N_Y_c_1489_n 5.24636e-19 $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_615 N_D_c_649_n N_Y_c_1342_n 0.0128895f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_616 N_D_c_657_n N_Y_c_1342_n 0.00224539f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_617 N_D_c_649_n N_Y_c_1495_n 0.00671723f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_618 N_D_c_650_n N_Y_c_1495_n 0.00671723f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_619 N_D_c_651_n N_Y_c_1495_n 5.24636e-19 $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_620 N_D_c_651_n N_Y_c_1343_n 0.00929182f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_621 N_D_c_704_p N_Y_c_1343_n 0.0228649f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_622 N_D_c_657_n N_Y_c_1343_n 0.00505612f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_623 N_D_c_659_n N_Y_c_1361_n 0.00480023f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_624 N_D_c_660_n N_Y_c_1361_n 0.0128795f $X=13.235 $Y=1.41 $X2=0 $Y2=0
cc_625 N_D_c_704_p N_Y_c_1361_n 0.0254394f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_626 N_D_c_657_n N_Y_c_1361_n 0.00841805f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_627 N_D_c_650_n N_Y_c_1527_n 5.24636e-19 $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_628 N_D_c_651_n N_Y_c_1527_n 0.00671723f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_629 N_D_c_652_n N_Y_c_1527_n 0.00671723f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_630 N_D_c_653_n N_Y_c_1527_n 5.24636e-19 $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_631 N_D_c_661_n N_Y_c_1362_n 0.0128795f $X=13.705 $Y=1.41 $X2=0 $Y2=0
cc_632 N_D_c_662_n N_Y_c_1362_n 0.0128795f $X=14.175 $Y=1.41 $X2=0 $Y2=0
cc_633 N_D_c_704_p N_Y_c_1362_n 0.0486996f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_634 N_D_c_657_n N_Y_c_1362_n 0.00844349f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_635 N_D_c_652_n N_Y_c_1344_n 0.00929182f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_636 N_D_c_653_n N_Y_c_1344_n 0.00929182f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_637 N_D_c_704_p N_Y_c_1344_n 0.0435408f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_638 N_D_c_657_n N_Y_c_1344_n 0.00468948f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_639 N_D_c_652_n N_Y_c_1539_n 5.24636e-19 $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_640 N_D_c_653_n N_Y_c_1539_n 0.00671723f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_641 N_D_c_654_n N_Y_c_1539_n 0.00671723f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_642 N_D_c_655_n N_Y_c_1539_n 5.24636e-19 $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_643 N_D_c_663_n N_Y_c_1363_n 0.0128795f $X=14.645 $Y=1.41 $X2=0 $Y2=0
cc_644 N_D_c_664_n N_Y_c_1363_n 0.0128188f $X=15.115 $Y=1.41 $X2=0 $Y2=0
cc_645 N_D_c_704_p N_Y_c_1363_n 0.0486996f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_646 N_D_c_657_n N_Y_c_1363_n 0.00844349f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_647 N_D_c_654_n N_Y_c_1345_n 0.00929182f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_648 N_D_c_655_n N_Y_c_1345_n 0.0104247f $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_649 N_D_c_656_n N_Y_c_1345_n 0.00367582f $X=15.56 $Y=0.995 $X2=0 $Y2=0
cc_650 N_D_c_704_p N_Y_c_1345_n 0.0572618f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_651 N_D_c_657_n N_Y_c_1345_n 0.00723932f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_652 N_D_c_654_n N_Y_c_1552_n 5.24636e-19 $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_653 N_D_c_655_n N_Y_c_1552_n 0.00671723f $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_654 N_D_c_656_n N_Y_c_1552_n 0.00539651f $X=15.56 $Y=0.995 $X2=0 $Y2=0
cc_655 N_D_c_649_n N_Y_c_1357_n 0.00218061f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_656 N_D_c_650_n N_Y_c_1357_n 0.00846356f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_657 N_D_c_658_n N_Y_c_1557_n 2.98817e-19 $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_658 N_D_c_659_n N_Y_c_1557_n 0.00677148f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_659 N_D_c_651_n N_Y_c_1358_n 0.00113286f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_660 N_D_c_652_n N_Y_c_1358_n 0.00113286f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_661 N_D_c_704_p N_Y_c_1358_n 0.0266272f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_662 N_D_c_657_n N_Y_c_1358_n 0.00230339f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_663 N_D_c_704_p N_Y_c_1364_n 0.0204252f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_664 N_D_c_657_n N_Y_c_1364_n 0.00675794f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_665 N_D_c_653_n N_Y_c_1359_n 0.00113286f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_666 N_D_c_654_n N_Y_c_1359_n 0.00113286f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_667 N_D_c_704_p N_Y_c_1359_n 0.0266272f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_668 N_D_c_657_n N_Y_c_1359_n 0.00230339f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_669 N_D_c_704_p N_Y_c_1365_n 0.0204252f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_670 N_D_c_657_n N_Y_c_1365_n 0.00675794f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_671 N_D_c_665_n N_Y_c_1366_n 5.31299e-19 $X=15.585 $Y=1.41 $X2=0 $Y2=0
cc_672 N_D_c_704_p N_Y_c_1366_n 0.0106211f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_673 N_D_c_657_n N_Y_c_1366_n 0.00745007f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_674 N_D_c_658_n Y 0.0013148f $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_675 N_D_c_649_n Y 0.00264975f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_676 N_D_c_650_n Y 0.00341687f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_677 N_D_c_659_n Y 0.00164342f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_678 N_D_c_660_n Y 2.526e-19 $X=13.235 $Y=1.41 $X2=0 $Y2=0
cc_679 N_D_c_651_n Y 5.17693e-19 $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_680 N_D_c_704_p Y 0.0168684f $X=15.19 $Y=1.16 $X2=0 $Y2=0
cc_681 N_D_c_657_n Y 0.0426768f $X=15.56 $Y=1.202 $X2=0 $Y2=0
cc_682 N_D_c_649_n N_VGND_c_1754_n 0.00166854f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_683 N_D_c_650_n N_VGND_c_1755_n 0.00166854f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_684 N_D_c_651_n N_VGND_c_1755_n 0.00166854f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_685 N_D_c_652_n N_VGND_c_1756_n 0.00166854f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_686 N_D_c_653_n N_VGND_c_1756_n 0.00166854f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_687 N_D_c_654_n N_VGND_c_1757_n 0.00166854f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_688 N_D_c_655_n N_VGND_c_1757_n 0.00166854f $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_689 N_D_c_656_n N_VGND_c_1759_n 0.0036723f $X=15.56 $Y=0.995 $X2=0 $Y2=0
cc_690 N_D_c_649_n N_VGND_c_1772_n 0.00423334f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_691 N_D_c_650_n N_VGND_c_1772_n 0.00423225f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_692 N_D_c_651_n N_VGND_c_1774_n 0.00423334f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_693 N_D_c_652_n N_VGND_c_1774_n 0.00423334f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_694 N_D_c_653_n N_VGND_c_1776_n 0.00423334f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_695 N_D_c_654_n N_VGND_c_1776_n 0.00423334f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_696 N_D_c_655_n N_VGND_c_1779_n 0.00423334f $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_697 N_D_c_656_n N_VGND_c_1779_n 0.00541359f $X=15.56 $Y=0.995 $X2=0 $Y2=0
cc_698 N_D_c_649_n N_VGND_c_1787_n 0.00596967f $X=12.32 $Y=0.995 $X2=0 $Y2=0
cc_699 N_D_c_650_n N_VGND_c_1787_n 0.00595664f $X=12.74 $Y=0.995 $X2=0 $Y2=0
cc_700 N_D_c_651_n N_VGND_c_1787_n 0.00595861f $X=13.26 $Y=0.995 $X2=0 $Y2=0
cc_701 N_D_c_652_n N_VGND_c_1787_n 0.00595861f $X=13.68 $Y=0.995 $X2=0 $Y2=0
cc_702 N_D_c_653_n N_VGND_c_1787_n 0.00595861f $X=14.2 $Y=0.995 $X2=0 $Y2=0
cc_703 N_D_c_654_n N_VGND_c_1787_n 0.00595861f $X=14.62 $Y=0.995 $X2=0 $Y2=0
cc_704 N_D_c_655_n N_VGND_c_1787_n 0.00595861f $X=15.14 $Y=0.995 $X2=0 $Y2=0
cc_705 N_D_c_656_n N_VGND_c_1787_n 0.0105165f $X=15.56 $Y=0.995 $X2=0 $Y2=0
cc_706 N_A_27_297#_c_790_n N_VPWR_M1000_s 0.00187091f $X=1.075 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_707 N_A_27_297#_c_792_n N_VPWR_M1008_s 0.00187091f $X=2.015 $Y=1.54 $X2=0
+ $Y2=0
cc_708 N_A_27_297#_c_793_n N_VPWR_M1026_s 0.00187091f $X=2.955 $Y=1.54 $X2=0
+ $Y2=0
cc_709 N_A_27_297#_c_794_n N_VPWR_M1040_s 0.00187091f $X=3.895 $Y=1.54 $X2=0
+ $Y2=0
cc_710 N_A_27_297#_c_790_n N_VPWR_c_908_n 0.0143191f $X=1.075 $Y=1.54 $X2=0
+ $Y2=0
cc_711 N_A_27_297#_c_842_p N_VPWR_c_909_n 0.0149311f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_712 N_A_27_297#_c_792_n N_VPWR_c_910_n 0.0143191f $X=2.015 $Y=1.54 $X2=0
+ $Y2=0
cc_713 N_A_27_297#_c_844_p N_VPWR_c_911_n 0.0149311f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_714 N_A_27_297#_c_793_n N_VPWR_c_912_n 0.0143191f $X=2.955 $Y=1.54 $X2=0
+ $Y2=0
cc_715 N_A_27_297#_c_846_p N_VPWR_c_913_n 0.0149311f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_716 N_A_27_297#_c_794_n N_VPWR_c_914_n 0.0143191f $X=3.895 $Y=1.54 $X2=0
+ $Y2=0
cc_717 N_A_27_297#_c_789_n N_VPWR_c_915_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_718 N_A_27_297#_c_849_p N_VPWR_c_916_n 0.015002f $X=4.02 $Y=2.295 $X2=0 $Y2=0
cc_719 N_A_27_297#_c_829_n N_VPWR_c_916_n 0.0386815f $X=4.835 $Y=2.38 $X2=0
+ $Y2=0
cc_720 N_A_27_297#_c_831_n N_VPWR_c_916_n 0.0386815f $X=5.775 $Y=2.38 $X2=0
+ $Y2=0
cc_721 N_A_27_297#_c_833_n N_VPWR_c_916_n 0.0386815f $X=6.715 $Y=2.38 $X2=0
+ $Y2=0
cc_722 N_A_27_297#_c_796_n N_VPWR_c_916_n 0.057821f $X=7.655 $Y=2.38 $X2=0 $Y2=0
cc_723 N_A_27_297#_c_854_p N_VPWR_c_916_n 0.0149886f $X=4.96 $Y=2.38 $X2=0 $Y2=0
cc_724 N_A_27_297#_c_855_p N_VPWR_c_916_n 0.0149886f $X=5.9 $Y=2.38 $X2=0 $Y2=0
cc_725 N_A_27_297#_c_856_p N_VPWR_c_916_n 0.0149886f $X=6.84 $Y=2.38 $X2=0 $Y2=0
cc_726 N_A_27_297#_M1000_d N_VPWR_c_907_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_727 N_A_27_297#_M1003_d N_VPWR_c_907_n 0.00370124f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_728 N_A_27_297#_M1016_d N_VPWR_c_907_n 0.00370124f $X=1.995 $Y=1.485 $X2=0
+ $Y2=0
cc_729 N_A_27_297#_M1032_d N_VPWR_c_907_n 0.00370124f $X=2.935 $Y=1.485 $X2=0
+ $Y2=0
cc_730 N_A_27_297#_M1056_d N_VPWR_c_907_n 0.00297222f $X=3.875 $Y=1.485 $X2=0
+ $Y2=0
cc_731 N_A_27_297#_M1009_d N_VPWR_c_907_n 0.00231264f $X=4.815 $Y=1.485 $X2=0
+ $Y2=0
cc_732 N_A_27_297#_M1035_d N_VPWR_c_907_n 0.00231264f $X=5.755 $Y=1.485 $X2=0
+ $Y2=0
cc_733 N_A_27_297#_M1047_d N_VPWR_c_907_n 0.00231264f $X=6.695 $Y=1.485 $X2=0
+ $Y2=0
cc_734 N_A_27_297#_M1058_d N_VPWR_c_907_n 0.00217519f $X=7.635 $Y=1.485 $X2=0
+ $Y2=0
cc_735 N_A_27_297#_c_789_n N_VPWR_c_907_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_736 N_A_27_297#_c_842_p N_VPWR_c_907_n 0.00955092f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_737 N_A_27_297#_c_844_p N_VPWR_c_907_n 0.00955092f $X=2.14 $Y=2.3 $X2=0 $Y2=0
cc_738 N_A_27_297#_c_846_p N_VPWR_c_907_n 0.00955092f $X=3.08 $Y=2.3 $X2=0 $Y2=0
cc_739 N_A_27_297#_c_849_p N_VPWR_c_907_n 0.00962794f $X=4.02 $Y=2.295 $X2=0
+ $Y2=0
cc_740 N_A_27_297#_c_829_n N_VPWR_c_907_n 0.0239144f $X=4.835 $Y=2.38 $X2=0
+ $Y2=0
cc_741 N_A_27_297#_c_831_n N_VPWR_c_907_n 0.0239144f $X=5.775 $Y=2.38 $X2=0
+ $Y2=0
cc_742 N_A_27_297#_c_833_n N_VPWR_c_907_n 0.0239144f $X=6.715 $Y=2.38 $X2=0
+ $Y2=0
cc_743 N_A_27_297#_c_796_n N_VPWR_c_907_n 0.0350785f $X=7.655 $Y=2.38 $X2=0
+ $Y2=0
cc_744 N_A_27_297#_c_854_p N_VPWR_c_907_n 0.00962421f $X=4.96 $Y=2.38 $X2=0
+ $Y2=0
cc_745 N_A_27_297#_c_855_p N_VPWR_c_907_n 0.00962421f $X=5.9 $Y=2.38 $X2=0 $Y2=0
cc_746 N_A_27_297#_c_856_p N_VPWR_c_907_n 0.00962421f $X=6.84 $Y=2.38 $X2=0
+ $Y2=0
cc_747 N_A_27_297#_c_829_n N_A_869_297#_M1005_s 0.00352392f $X=4.835 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_748 N_A_27_297#_c_831_n N_A_869_297#_M1014_s 0.00352392f $X=5.775 $Y=2.38
+ $X2=0 $Y2=0
cc_749 N_A_27_297#_c_833_n N_A_869_297#_M1043_s 0.00352392f $X=6.715 $Y=2.38
+ $X2=0 $Y2=0
cc_750 N_A_27_297#_c_796_n N_A_869_297#_M1053_s 0.00352392f $X=7.655 $Y=2.38
+ $X2=0 $Y2=0
cc_751 N_A_27_297#_M1009_d N_A_869_297#_c_1090_n 0.00187091f $X=4.815 $Y=1.485
+ $X2=0 $Y2=0
cc_752 N_A_27_297#_c_829_n N_A_869_297#_c_1090_n 0.00385532f $X=4.835 $Y=2.38
+ $X2=0 $Y2=0
cc_753 N_A_27_297#_c_884_p N_A_869_297#_c_1090_n 0.0143018f $X=4.96 $Y=1.96
+ $X2=0 $Y2=0
cc_754 N_A_27_297#_c_831_n N_A_869_297#_c_1090_n 0.00385532f $X=5.775 $Y=2.38
+ $X2=0 $Y2=0
cc_755 N_A_27_297#_M1035_d N_A_869_297#_c_1091_n 0.00187091f $X=5.755 $Y=1.485
+ $X2=0 $Y2=0
cc_756 N_A_27_297#_c_831_n N_A_869_297#_c_1091_n 0.00385532f $X=5.775 $Y=2.38
+ $X2=0 $Y2=0
cc_757 N_A_27_297#_c_888_p N_A_869_297#_c_1091_n 0.0143018f $X=5.9 $Y=1.96 $X2=0
+ $Y2=0
cc_758 N_A_27_297#_c_833_n N_A_869_297#_c_1091_n 0.00385532f $X=6.715 $Y=2.38
+ $X2=0 $Y2=0
cc_759 N_A_27_297#_M1047_d N_A_869_297#_c_1092_n 0.00187091f $X=6.695 $Y=1.485
+ $X2=0 $Y2=0
cc_760 N_A_27_297#_c_833_n N_A_869_297#_c_1092_n 0.00385532f $X=6.715 $Y=2.38
+ $X2=0 $Y2=0
cc_761 N_A_27_297#_c_892_p N_A_869_297#_c_1092_n 0.0143018f $X=6.84 $Y=1.96
+ $X2=0 $Y2=0
cc_762 N_A_27_297#_c_796_n N_A_869_297#_c_1092_n 0.00385532f $X=7.655 $Y=2.38
+ $X2=0 $Y2=0
cc_763 N_A_27_297#_M1058_d N_A_869_297#_c_1093_n 0.00295666f $X=7.635 $Y=1.485
+ $X2=0 $Y2=0
cc_764 N_A_27_297#_c_796_n N_A_869_297#_c_1093_n 0.00385532f $X=7.655 $Y=2.38
+ $X2=0 $Y2=0
cc_765 N_A_27_297#_c_797_n N_A_869_297#_c_1093_n 0.0205983f $X=7.78 $Y=1.96
+ $X2=0 $Y2=0
cc_766 N_A_27_297#_c_795_n N_A_869_297#_c_1097_n 0.00226124f $X=4.02 $Y=1.625
+ $X2=0 $Y2=0
cc_767 N_A_27_297#_c_829_n N_A_869_297#_c_1097_n 0.013395f $X=4.835 $Y=2.38
+ $X2=0 $Y2=0
cc_768 N_A_27_297#_c_831_n N_A_869_297#_c_1098_n 0.013395f $X=5.775 $Y=2.38
+ $X2=0 $Y2=0
cc_769 N_A_27_297#_c_833_n N_A_869_297#_c_1099_n 0.013395f $X=6.715 $Y=2.38
+ $X2=0 $Y2=0
cc_770 N_A_27_297#_c_796_n N_A_869_297#_c_1100_n 0.013395f $X=7.655 $Y=2.38
+ $X2=0 $Y2=0
cc_771 N_A_27_297#_c_797_n N_A_1635_297#_c_1210_n 0.0376802f $X=7.78 $Y=1.96
+ $X2=0 $Y2=0
cc_772 N_A_27_297#_c_796_n N_A_1635_297#_c_1211_n 0.0147157f $X=7.655 $Y=2.38
+ $X2=0 $Y2=0
cc_773 N_A_27_297#_c_794_n N_Y_c_1334_n 0.00286947f $X=3.895 $Y=1.54 $X2=0 $Y2=0
cc_774 N_A_27_297#_c_795_n N_Y_c_1334_n 0.00936521f $X=4.02 $Y=1.625 $X2=0 $Y2=0
cc_775 N_A_27_297#_c_791_n N_VGND_c_1739_n 0.0106493f $X=0.425 $Y=1.54 $X2=0
+ $Y2=0
cc_776 N_VPWR_c_907_n N_A_869_297#_M1005_s 0.00232895f $X=15.87 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_777 N_VPWR_c_907_n N_A_869_297#_M1014_s 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_778 N_VPWR_c_907_n N_A_869_297#_M1043_s 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_779 N_VPWR_c_907_n N_A_869_297#_M1053_s 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_780 N_VPWR_c_907_n N_A_869_297#_M1001_d 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_781 N_VPWR_c_907_n N_A_869_297#_M1017_d 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_782 N_VPWR_c_907_n N_A_869_297#_M1025_d 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_783 N_VPWR_c_907_n N_A_869_297#_M1050_d 0.00232895f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_784 N_VPWR_c_907_n N_A_1635_297#_M1001_s 0.00217519f $X=15.87 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_785 N_VPWR_c_907_n N_A_1635_297#_M1013_s 0.00231263f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_786 N_VPWR_c_907_n N_A_1635_297#_M1021_s 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_787 N_VPWR_c_907_n N_A_1635_297#_M1034_s 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_788 N_VPWR_c_907_n N_A_1635_297#_M1059_s 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_789 N_VPWR_c_907_n N_A_1635_297#_M1011_d 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_790 N_VPWR_c_907_n N_A_1635_297#_M1029_d 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_791 N_VPWR_c_907_n N_A_1635_297#_M1037_d 0.00231264f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_792 N_VPWR_c_907_n N_A_1635_297#_M1060_d 0.00225717f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_793 N_VPWR_c_916_n N_A_1635_297#_c_1215_n 0.0367458f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_794 N_VPWR_c_907_n N_A_1635_297#_c_1215_n 0.0225861f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_795 N_VPWR_c_916_n N_A_1635_297#_c_1211_n 0.0191395f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_796 N_VPWR_c_907_n N_A_1635_297#_c_1211_n 0.0111641f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_797 N_VPWR_c_916_n N_A_1635_297#_c_1219_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_798 N_VPWR_c_907_n N_A_1635_297#_c_1219_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_799 N_VPWR_c_916_n N_A_1635_297#_c_1221_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_800 N_VPWR_c_907_n N_A_1635_297#_c_1221_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_801 N_VPWR_c_916_n N_A_1635_297#_c_1223_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_802 N_VPWR_c_907_n N_A_1635_297#_c_1223_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_803 N_VPWR_c_916_n N_A_1635_297#_c_1228_n 0.0386553f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_804 N_VPWR_c_907_n N_A_1635_297#_c_1228_n 0.023911f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_805 N_VPWR_c_916_n N_A_1635_297#_c_1230_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_806 N_VPWR_c_907_n N_A_1635_297#_c_1230_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_807 N_VPWR_c_916_n N_A_1635_297#_c_1232_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_808 N_VPWR_c_907_n N_A_1635_297#_c_1232_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_809 N_VPWR_c_916_n N_A_1635_297#_c_1234_n 0.0386815f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_810 N_VPWR_c_907_n N_A_1635_297#_c_1234_n 0.0239144f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_811 N_VPWR_c_916_n N_A_1635_297#_c_1213_n 0.0198621f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_812 N_VPWR_c_907_n N_A_1635_297#_c_1213_n 0.0115483f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_813 N_VPWR_c_916_n N_A_1635_297#_c_1226_n 0.0170278f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_814 N_VPWR_c_907_n N_A_1635_297#_c_1226_n 0.0110002f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_815 N_VPWR_c_916_n N_A_1635_297#_c_1270_n 0.0149886f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_816 N_VPWR_c_907_n N_A_1635_297#_c_1270_n 0.00962421f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_817 N_VPWR_c_916_n N_A_1635_297#_c_1272_n 0.0149886f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_818 N_VPWR_c_907_n N_A_1635_297#_c_1272_n 0.00962421f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_819 N_VPWR_c_916_n N_A_1635_297#_c_1274_n 0.015002f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_820 N_VPWR_c_907_n N_A_1635_297#_c_1274_n 0.00961749f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_821 N_VPWR_c_916_n N_A_1635_297#_c_1276_n 0.0149886f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_822 N_VPWR_c_907_n N_A_1635_297#_c_1276_n 0.00962421f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_823 N_VPWR_c_916_n N_A_1635_297#_c_1278_n 0.0149886f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_824 N_VPWR_c_907_n N_A_1635_297#_c_1278_n 0.00962421f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_825 N_VPWR_c_916_n N_A_1635_297#_c_1280_n 0.0149886f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_826 N_VPWR_c_907_n N_A_1635_297#_c_1280_n 0.00962421f $X=15.87 $Y=2.72 $X2=0
+ $Y2=0
cc_827 N_VPWR_c_907_n N_Y_M1006_s 0.00232895f $X=15.87 $Y=2.72 $X2=0 $Y2=0
cc_828 N_VPWR_c_907_n N_Y_M1023_s 0.00232895f $X=15.87 $Y=2.72 $X2=0 $Y2=0
cc_829 N_VPWR_c_907_n N_Y_M1036_s 0.00232895f $X=15.87 $Y=2.72 $X2=0 $Y2=0
cc_830 N_VPWR_c_907_n N_Y_M1044_s 0.00232895f $X=15.87 $Y=2.72 $X2=0 $Y2=0
cc_831 N_A_869_297#_c_1093_n N_A_1635_297#_M1001_s 0.00295666f $X=8.645 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_832 N_A_869_297#_c_1094_n N_A_1635_297#_M1013_s 0.00187091f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_833 N_A_869_297#_c_1095_n N_A_1635_297#_M1021_s 0.00187091f $X=10.525 $Y=1.54
+ $X2=0 $Y2=0
cc_834 N_A_869_297#_c_1096_n N_A_1635_297#_M1034_s 0.00187091f $X=11.465 $Y=1.54
+ $X2=0 $Y2=0
cc_835 N_A_869_297#_c_1093_n N_A_1635_297#_c_1210_n 0.0205983f $X=8.645 $Y=1.54
+ $X2=0 $Y2=0
cc_836 N_A_869_297#_M1001_d N_A_1635_297#_c_1215_n 0.00352392f $X=8.625 $Y=1.485
+ $X2=0 $Y2=0
cc_837 N_A_869_297#_c_1093_n N_A_1635_297#_c_1215_n 0.00385532f $X=8.645 $Y=1.54
+ $X2=0 $Y2=0
cc_838 N_A_869_297#_c_1094_n N_A_1635_297#_c_1215_n 0.00342456f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_839 N_A_869_297#_c_1101_n N_A_1635_297#_c_1215_n 0.013395f $X=8.77 $Y=1.62
+ $X2=0 $Y2=0
cc_840 N_A_869_297#_c_1094_n N_A_1635_297#_c_1217_n 0.0157053f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_841 N_A_869_297#_M1017_d N_A_1635_297#_c_1219_n 0.00352392f $X=9.565 $Y=1.485
+ $X2=0 $Y2=0
cc_842 N_A_869_297#_c_1094_n N_A_1635_297#_c_1219_n 0.00385532f $X=9.585 $Y=1.54
+ $X2=0 $Y2=0
cc_843 N_A_869_297#_c_1095_n N_A_1635_297#_c_1219_n 0.00385532f $X=10.525
+ $Y=1.54 $X2=0 $Y2=0
cc_844 N_A_869_297#_c_1102_n N_A_1635_297#_c_1219_n 0.013395f $X=9.71 $Y=1.62
+ $X2=0 $Y2=0
cc_845 N_A_869_297#_c_1095_n N_A_1635_297#_c_1296_n 0.0143018f $X=10.525 $Y=1.54
+ $X2=0 $Y2=0
cc_846 N_A_869_297#_M1025_d N_A_1635_297#_c_1221_n 0.00352392f $X=10.505
+ $Y=1.485 $X2=0 $Y2=0
cc_847 N_A_869_297#_c_1095_n N_A_1635_297#_c_1221_n 0.00385532f $X=10.525
+ $Y=1.54 $X2=0 $Y2=0
cc_848 N_A_869_297#_c_1096_n N_A_1635_297#_c_1221_n 0.00385532f $X=11.465
+ $Y=1.54 $X2=0 $Y2=0
cc_849 N_A_869_297#_c_1103_n N_A_1635_297#_c_1221_n 0.013395f $X=10.65 $Y=1.62
+ $X2=0 $Y2=0
cc_850 N_A_869_297#_c_1096_n N_A_1635_297#_c_1301_n 0.0143018f $X=11.465 $Y=1.54
+ $X2=0 $Y2=0
cc_851 N_A_869_297#_M1050_d N_A_1635_297#_c_1223_n 0.00352392f $X=11.445
+ $Y=1.485 $X2=0 $Y2=0
cc_852 N_A_869_297#_c_1096_n N_A_1635_297#_c_1223_n 0.00385532f $X=11.465
+ $Y=1.54 $X2=0 $Y2=0
cc_853 N_A_869_297#_c_1104_n N_A_1635_297#_c_1223_n 0.013395f $X=11.59 $Y=1.62
+ $X2=0 $Y2=0
cc_854 N_A_869_297#_c_1104_n N_A_1635_297#_c_1212_n 0.00209545f $X=11.59 $Y=1.62
+ $X2=0 $Y2=0
cc_855 N_A_869_297#_c_1093_n N_Y_c_1338_n 0.0271341f $X=8.645 $Y=1.54 $X2=0
+ $Y2=0
cc_856 N_A_1635_297#_c_1228_n N_Y_M1006_s 0.00352392f $X=12.875 $Y=2.38 $X2=0
+ $Y2=0
cc_857 N_A_1635_297#_c_1230_n N_Y_M1023_s 0.00352392f $X=13.815 $Y=2.38 $X2=0
+ $Y2=0
cc_858 N_A_1635_297#_c_1232_n N_Y_M1036_s 0.00352392f $X=14.755 $Y=2.38 $X2=0
+ $Y2=0
cc_859 N_A_1635_297#_c_1234_n N_Y_M1044_s 0.00352392f $X=15.695 $Y=2.38 $X2=0
+ $Y2=0
cc_860 N_A_1635_297#_c_1212_n N_Y_c_1342_n 0.00929029f $X=12.06 $Y=1.62 $X2=0
+ $Y2=0
cc_861 N_A_1635_297#_M1011_d N_Y_c_1361_n 0.00187091f $X=12.855 $Y=1.485 $X2=0
+ $Y2=0
cc_862 N_A_1635_297#_c_1228_n N_Y_c_1361_n 8.39986e-19 $X=12.875 $Y=2.38 $X2=0
+ $Y2=0
cc_863 N_A_1635_297#_c_1313_p N_Y_c_1361_n 0.0143018f $X=13 $Y=1.96 $X2=0 $Y2=0
cc_864 N_A_1635_297#_c_1230_n N_Y_c_1361_n 0.00385532f $X=13.815 $Y=2.38 $X2=0
+ $Y2=0
cc_865 N_A_1635_297#_M1029_d N_Y_c_1362_n 0.00187091f $X=13.795 $Y=1.485 $X2=0
+ $Y2=0
cc_866 N_A_1635_297#_c_1230_n N_Y_c_1362_n 0.00385532f $X=13.815 $Y=2.38 $X2=0
+ $Y2=0
cc_867 N_A_1635_297#_c_1317_p N_Y_c_1362_n 0.0143018f $X=13.94 $Y=1.96 $X2=0
+ $Y2=0
cc_868 N_A_1635_297#_c_1232_n N_Y_c_1362_n 0.00385532f $X=14.755 $Y=2.38 $X2=0
+ $Y2=0
cc_869 N_A_1635_297#_M1037_d N_Y_c_1363_n 0.00187091f $X=14.735 $Y=1.485 $X2=0
+ $Y2=0
cc_870 N_A_1635_297#_c_1232_n N_Y_c_1363_n 0.00385532f $X=14.755 $Y=2.38 $X2=0
+ $Y2=0
cc_871 N_A_1635_297#_c_1321_p N_Y_c_1363_n 0.0143018f $X=14.89 $Y=1.96 $X2=0
+ $Y2=0
cc_872 N_A_1635_297#_c_1234_n N_Y_c_1363_n 0.00385532f $X=15.695 $Y=2.38 $X2=0
+ $Y2=0
cc_873 N_A_1635_297#_c_1212_n N_Y_c_1557_n 0.00209545f $X=12.06 $Y=1.62 $X2=0
+ $Y2=0
cc_874 N_A_1635_297#_c_1228_n N_Y_c_1557_n 0.0167505f $X=12.875 $Y=2.38 $X2=0
+ $Y2=0
cc_875 N_A_1635_297#_c_1230_n N_Y_c_1364_n 0.013395f $X=13.815 $Y=2.38 $X2=0
+ $Y2=0
cc_876 N_A_1635_297#_c_1232_n N_Y_c_1365_n 0.013395f $X=14.755 $Y=2.38 $X2=0
+ $Y2=0
cc_877 N_A_1635_297#_c_1234_n N_Y_c_1366_n 0.013395f $X=15.695 $Y=2.38 $X2=0
+ $Y2=0
cc_878 N_A_1635_297#_c_1214_n N_Y_c_1366_n 0.00139065f $X=15.83 $Y=1.63 $X2=0
+ $Y2=0
cc_879 N_A_1635_297#_c_1214_n N_VGND_c_1759_n 0.0109198f $X=15.83 $Y=1.63 $X2=0
+ $Y2=0
cc_880 N_Y_c_1330_n N_VGND_M1019_d 0.00274794f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_881 N_Y_c_1332_n N_VGND_M1038_d 0.00274794f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_882 N_Y_c_1333_n N_VGND_M1051_d 0.00274794f $X=3.385 $Y=0.815 $X2=0 $Y2=0
cc_883 N_Y_c_1334_n N_VGND_M1062_d 0.00274794f $X=4.325 $Y=0.815 $X2=0 $Y2=0
cc_884 N_Y_c_1335_n N_VGND_M1012_s 0.00274794f $X=5.265 $Y=0.815 $X2=0 $Y2=0
cc_885 N_Y_c_1336_n N_VGND_M1024_s 0.00274794f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_886 N_Y_c_1337_n N_VGND_M1041_s 0.00274794f $X=7.145 $Y=0.815 $X2=0 $Y2=0
cc_887 N_Y_c_1338_n N_VGND_M1061_s 0.0127463f $X=8.605 $Y=0.815 $X2=0 $Y2=0
cc_888 N_Y_c_1339_n N_VGND_M1007_s 0.00274794f $X=9.545 $Y=0.815 $X2=0 $Y2=0
cc_889 N_Y_c_1340_n N_VGND_M1028_s 0.00274794f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_890 N_Y_c_1341_n N_VGND_M1054_s 0.00274794f $X=11.425 $Y=0.815 $X2=0 $Y2=0
cc_891 N_Y_c_1342_n N_VGND_M1063_s 0.00274794f $X=12.365 $Y=0.815 $X2=0 $Y2=0
cc_892 N_Y_c_1343_n N_VGND_M1022_s 0.00274794f $X=13.305 $Y=0.815 $X2=0 $Y2=0
cc_893 N_Y_c_1344_n N_VGND_M1030_s 0.00274794f $X=14.245 $Y=0.815 $X2=0 $Y2=0
cc_894 N_Y_c_1345_n N_VGND_M1042_s 0.00274794f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_895 N_Y_c_1331_n N_VGND_c_1739_n 0.00834802f $X=0.895 $Y=0.815 $X2=0 $Y2=0
cc_896 N_Y_c_1330_n N_VGND_c_1740_n 0.0201123f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_897 N_Y_c_1330_n N_VGND_c_1741_n 0.00198695f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_898 N_Y_c_1379_n N_VGND_c_1741_n 0.0188551f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_899 N_Y_c_1332_n N_VGND_c_1741_n 0.00198695f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_900 N_Y_c_1332_n N_VGND_c_1742_n 0.0201123f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_901 N_Y_c_1332_n N_VGND_c_1743_n 0.00198695f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_902 N_Y_c_1387_n N_VGND_c_1743_n 0.0188551f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_903 N_Y_c_1333_n N_VGND_c_1743_n 0.00198695f $X=3.385 $Y=0.815 $X2=0 $Y2=0
cc_904 N_Y_c_1333_n N_VGND_c_1744_n 0.0201123f $X=3.385 $Y=0.815 $X2=0 $Y2=0
cc_905 N_Y_c_1333_n N_VGND_c_1745_n 0.00198695f $X=3.385 $Y=0.815 $X2=0 $Y2=0
cc_906 N_Y_c_1395_n N_VGND_c_1745_n 0.0188551f $X=3.55 $Y=0.39 $X2=0 $Y2=0
cc_907 N_Y_c_1334_n N_VGND_c_1745_n 0.00198695f $X=4.325 $Y=0.815 $X2=0 $Y2=0
cc_908 N_Y_c_1334_n N_VGND_c_1746_n 0.0201123f $X=4.325 $Y=0.815 $X2=0 $Y2=0
cc_909 N_Y_c_1334_n N_VGND_c_1747_n 0.00198695f $X=4.325 $Y=0.815 $X2=0 $Y2=0
cc_910 N_Y_c_1401_n N_VGND_c_1747_n 0.0188551f $X=4.49 $Y=0.39 $X2=0 $Y2=0
cc_911 N_Y_c_1335_n N_VGND_c_1747_n 0.00198695f $X=5.265 $Y=0.815 $X2=0 $Y2=0
cc_912 N_Y_c_1335_n N_VGND_c_1748_n 0.0201123f $X=5.265 $Y=0.815 $X2=0 $Y2=0
cc_913 N_Y_c_1336_n N_VGND_c_1749_n 0.0201123f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_914 N_Y_c_1337_n N_VGND_c_1750_n 0.0201123f $X=7.145 $Y=0.815 $X2=0 $Y2=0
cc_915 N_Y_c_1339_n N_VGND_c_1751_n 0.0201123f $X=9.545 $Y=0.815 $X2=0 $Y2=0
cc_916 N_Y_c_1340_n N_VGND_c_1752_n 0.0201123f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_917 N_Y_c_1341_n N_VGND_c_1753_n 0.0201123f $X=11.425 $Y=0.815 $X2=0 $Y2=0
cc_918 N_Y_c_1342_n N_VGND_c_1754_n 0.0201123f $X=12.365 $Y=0.815 $X2=0 $Y2=0
cc_919 N_Y_c_1343_n N_VGND_c_1755_n 0.0201123f $X=13.305 $Y=0.815 $X2=0 $Y2=0
cc_920 N_Y_c_1344_n N_VGND_c_1756_n 0.0201123f $X=14.245 $Y=0.815 $X2=0 $Y2=0
cc_921 N_Y_c_1345_n N_VGND_c_1757_n 0.0201123f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_922 N_Y_c_1345_n N_VGND_c_1759_n 0.00835667f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_923 N_Y_c_1335_n N_VGND_c_1760_n 0.00198695f $X=5.265 $Y=0.815 $X2=0 $Y2=0
cc_924 N_Y_c_1425_n N_VGND_c_1760_n 0.0188551f $X=5.43 $Y=0.39 $X2=0 $Y2=0
cc_925 N_Y_c_1336_n N_VGND_c_1760_n 0.00198695f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_926 N_Y_c_1336_n N_VGND_c_1762_n 0.00198695f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_927 N_Y_c_1433_n N_VGND_c_1762_n 0.0188551f $X=6.37 $Y=0.39 $X2=0 $Y2=0
cc_928 N_Y_c_1337_n N_VGND_c_1762_n 0.00198695f $X=7.145 $Y=0.815 $X2=0 $Y2=0
cc_929 N_Y_c_1338_n N_VGND_c_1764_n 0.00198695f $X=8.605 $Y=0.815 $X2=0 $Y2=0
cc_930 N_Y_c_1466_n N_VGND_c_1764_n 0.0188551f $X=8.77 $Y=0.39 $X2=0 $Y2=0
cc_931 N_Y_c_1339_n N_VGND_c_1764_n 0.00198695f $X=9.545 $Y=0.815 $X2=0 $Y2=0
cc_932 N_Y_c_1339_n N_VGND_c_1766_n 0.00198695f $X=9.545 $Y=0.815 $X2=0 $Y2=0
cc_933 N_Y_c_1473_n N_VGND_c_1766_n 0.0188551f $X=9.71 $Y=0.39 $X2=0 $Y2=0
cc_934 N_Y_c_1340_n N_VGND_c_1766_n 0.00198695f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_935 N_Y_c_1340_n N_VGND_c_1768_n 0.00198695f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_936 N_Y_c_1481_n N_VGND_c_1768_n 0.0188551f $X=10.65 $Y=0.39 $X2=0 $Y2=0
cc_937 N_Y_c_1341_n N_VGND_c_1768_n 0.00198695f $X=11.425 $Y=0.815 $X2=0 $Y2=0
cc_938 N_Y_c_1341_n N_VGND_c_1770_n 0.00198695f $X=11.425 $Y=0.815 $X2=0 $Y2=0
cc_939 N_Y_c_1489_n N_VGND_c_1770_n 0.0188551f $X=11.59 $Y=0.39 $X2=0 $Y2=0
cc_940 N_Y_c_1342_n N_VGND_c_1770_n 0.00198695f $X=12.365 $Y=0.815 $X2=0 $Y2=0
cc_941 N_Y_c_1342_n N_VGND_c_1772_n 0.00198695f $X=12.365 $Y=0.815 $X2=0 $Y2=0
cc_942 N_Y_c_1495_n N_VGND_c_1772_n 0.0188977f $X=12.53 $Y=0.39 $X2=0 $Y2=0
cc_943 N_Y_c_1357_n N_VGND_c_1772_n 0.00177065f $X=12.59 $Y=0.815 $X2=0 $Y2=0
cc_944 N_Y_c_1343_n N_VGND_c_1774_n 0.00198695f $X=13.305 $Y=0.815 $X2=0 $Y2=0
cc_945 N_Y_c_1527_n N_VGND_c_1774_n 0.0188551f $X=13.47 $Y=0.39 $X2=0 $Y2=0
cc_946 N_Y_c_1344_n N_VGND_c_1774_n 0.00198695f $X=14.245 $Y=0.815 $X2=0 $Y2=0
cc_947 N_Y_c_1344_n N_VGND_c_1776_n 0.00198695f $X=14.245 $Y=0.815 $X2=0 $Y2=0
cc_948 N_Y_c_1539_n N_VGND_c_1776_n 0.0188551f $X=14.41 $Y=0.39 $X2=0 $Y2=0
cc_949 N_Y_c_1345_n N_VGND_c_1776_n 0.00198695f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_950 N_Y_c_1368_n N_VGND_c_1778_n 0.0188551f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_951 N_Y_c_1330_n N_VGND_c_1778_n 0.00198695f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_952 N_Y_c_1345_n N_VGND_c_1779_n 0.00198695f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_953 N_Y_c_1552_n N_VGND_c_1779_n 0.0188551f $X=15.35 $Y=0.39 $X2=0 $Y2=0
cc_954 N_Y_c_1337_n N_VGND_c_1785_n 0.00198695f $X=7.145 $Y=0.815 $X2=0 $Y2=0
cc_955 N_Y_c_1441_n N_VGND_c_1785_n 0.0188551f $X=7.31 $Y=0.39 $X2=0 $Y2=0
cc_956 N_Y_c_1338_n N_VGND_c_1785_n 0.00198695f $X=8.605 $Y=0.815 $X2=0 $Y2=0
cc_957 N_Y_c_1338_n N_VGND_c_1786_n 0.0606502f $X=8.605 $Y=0.815 $X2=0 $Y2=0
cc_958 N_Y_M1018_s N_VGND_c_1787_n 0.00215201f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_959 N_Y_M1031_s N_VGND_c_1787_n 0.00215201f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_960 N_Y_M1045_s N_VGND_c_1787_n 0.00215201f $X=2.475 $Y=0.235 $X2=0 $Y2=0
cc_961 N_Y_M1057_s N_VGND_c_1787_n 0.00215201f $X=3.415 $Y=0.235 $X2=0 $Y2=0
cc_962 N_Y_M1002_d N_VGND_c_1787_n 0.00215201f $X=4.355 $Y=0.235 $X2=0 $Y2=0
cc_963 N_Y_M1020_d N_VGND_c_1787_n 0.00215201f $X=5.295 $Y=0.235 $X2=0 $Y2=0
cc_964 N_Y_M1039_d N_VGND_c_1787_n 0.00215201f $X=6.235 $Y=0.235 $X2=0 $Y2=0
cc_965 N_Y_M1052_d N_VGND_c_1787_n 0.00215201f $X=7.175 $Y=0.235 $X2=0 $Y2=0
cc_966 N_Y_M1004_d N_VGND_c_1787_n 0.00215201f $X=8.635 $Y=0.235 $X2=0 $Y2=0
cc_967 N_Y_M1015_d N_VGND_c_1787_n 0.00215201f $X=9.575 $Y=0.235 $X2=0 $Y2=0
cc_968 N_Y_M1046_d N_VGND_c_1787_n 0.00215201f $X=10.515 $Y=0.235 $X2=0 $Y2=0
cc_969 N_Y_M1055_d N_VGND_c_1787_n 0.00215201f $X=11.455 $Y=0.235 $X2=0 $Y2=0
cc_970 N_Y_M1010_d N_VGND_c_1787_n 0.00215201f $X=12.395 $Y=0.235 $X2=0 $Y2=0
cc_971 N_Y_M1027_d N_VGND_c_1787_n 0.00215201f $X=13.335 $Y=0.235 $X2=0 $Y2=0
cc_972 N_Y_M1033_d N_VGND_c_1787_n 0.00215201f $X=14.275 $Y=0.235 $X2=0 $Y2=0
cc_973 N_Y_M1048_d N_VGND_c_1787_n 0.00215201f $X=15.215 $Y=0.235 $X2=0 $Y2=0
cc_974 N_Y_c_1368_n N_VGND_c_1787_n 0.0122069f $X=0.73 $Y=0.39 $X2=0 $Y2=0
cc_975 N_Y_c_1330_n N_VGND_c_1787_n 0.00874058f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_976 N_Y_c_1379_n N_VGND_c_1787_n 0.0122069f $X=1.67 $Y=0.39 $X2=0 $Y2=0
cc_977 N_Y_c_1332_n N_VGND_c_1787_n 0.00874058f $X=2.445 $Y=0.815 $X2=0 $Y2=0
cc_978 N_Y_c_1387_n N_VGND_c_1787_n 0.0122069f $X=2.61 $Y=0.39 $X2=0 $Y2=0
cc_979 N_Y_c_1333_n N_VGND_c_1787_n 0.00874058f $X=3.385 $Y=0.815 $X2=0 $Y2=0
cc_980 N_Y_c_1395_n N_VGND_c_1787_n 0.0122069f $X=3.55 $Y=0.39 $X2=0 $Y2=0
cc_981 N_Y_c_1334_n N_VGND_c_1787_n 0.00874058f $X=4.325 $Y=0.815 $X2=0 $Y2=0
cc_982 N_Y_c_1401_n N_VGND_c_1787_n 0.0122069f $X=4.49 $Y=0.39 $X2=0 $Y2=0
cc_983 N_Y_c_1335_n N_VGND_c_1787_n 0.00874058f $X=5.265 $Y=0.815 $X2=0 $Y2=0
cc_984 N_Y_c_1425_n N_VGND_c_1787_n 0.0122069f $X=5.43 $Y=0.39 $X2=0 $Y2=0
cc_985 N_Y_c_1336_n N_VGND_c_1787_n 0.00874058f $X=6.205 $Y=0.815 $X2=0 $Y2=0
cc_986 N_Y_c_1433_n N_VGND_c_1787_n 0.0122069f $X=6.37 $Y=0.39 $X2=0 $Y2=0
cc_987 N_Y_c_1337_n N_VGND_c_1787_n 0.00874058f $X=7.145 $Y=0.815 $X2=0 $Y2=0
cc_988 N_Y_c_1441_n N_VGND_c_1787_n 0.0122069f $X=7.31 $Y=0.39 $X2=0 $Y2=0
cc_989 N_Y_c_1338_n N_VGND_c_1787_n 0.0107088f $X=8.605 $Y=0.815 $X2=0 $Y2=0
cc_990 N_Y_c_1466_n N_VGND_c_1787_n 0.0122069f $X=8.77 $Y=0.39 $X2=0 $Y2=0
cc_991 N_Y_c_1339_n N_VGND_c_1787_n 0.00874058f $X=9.545 $Y=0.815 $X2=0 $Y2=0
cc_992 N_Y_c_1473_n N_VGND_c_1787_n 0.0122069f $X=9.71 $Y=0.39 $X2=0 $Y2=0
cc_993 N_Y_c_1340_n N_VGND_c_1787_n 0.00874058f $X=10.485 $Y=0.815 $X2=0 $Y2=0
cc_994 N_Y_c_1481_n N_VGND_c_1787_n 0.0122069f $X=10.65 $Y=0.39 $X2=0 $Y2=0
cc_995 N_Y_c_1341_n N_VGND_c_1787_n 0.00874058f $X=11.425 $Y=0.815 $X2=0 $Y2=0
cc_996 N_Y_c_1489_n N_VGND_c_1787_n 0.0122069f $X=11.59 $Y=0.39 $X2=0 $Y2=0
cc_997 N_Y_c_1342_n N_VGND_c_1787_n 0.00874058f $X=12.365 $Y=0.815 $X2=0 $Y2=0
cc_998 N_Y_c_1495_n N_VGND_c_1787_n 0.01222f $X=12.53 $Y=0.39 $X2=0 $Y2=0
cc_999 N_Y_c_1343_n N_VGND_c_1787_n 0.00617665f $X=13.305 $Y=0.815 $X2=0 $Y2=0
cc_1000 N_Y_c_1527_n N_VGND_c_1787_n 0.0122069f $X=13.47 $Y=0.39 $X2=0 $Y2=0
cc_1001 N_Y_c_1344_n N_VGND_c_1787_n 0.00874058f $X=14.245 $Y=0.815 $X2=0 $Y2=0
cc_1002 N_Y_c_1539_n N_VGND_c_1787_n 0.0122069f $X=14.41 $Y=0.39 $X2=0 $Y2=0
cc_1003 N_Y_c_1345_n N_VGND_c_1787_n 0.00874058f $X=15.185 $Y=0.815 $X2=0 $Y2=0
cc_1004 N_Y_c_1552_n N_VGND_c_1787_n 0.0122069f $X=15.35 $Y=0.39 $X2=0 $Y2=0
cc_1005 N_Y_c_1357_n N_VGND_c_1787_n 0.00274439f $X=12.59 $Y=0.815 $X2=0 $Y2=0
