* File: sky130_fd_sc_hdll__dlrtp_1.pex.spice
* Created: Thu Aug 27 19:05:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%GATE 4 5 7 8 10 13 19 20 24 26
c42 19 0 5.20423e-20 $X=0.23 $Y=1.19
c43 13 0 3.98209e-20 $X=0.52 $Y=0.805
r44 24 27 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.4
r45 24 26 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.07
r46 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.26 $Y=1.19
+ $X2=0.26 $Y2=1.53
r47 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.235 $X2=0.3 $Y2=1.235
r48 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r49 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r51 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.33 $Y=1.665
+ $X2=0.495 $Y2=1.665
r52 4 27 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=1.59 $X2=0.33
+ $Y2=1.4
r53 1 13 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.805
+ $X2=0.52 $Y2=0.805
r54 1 26 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.88 $X2=0.33
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%A_27_363# 1 2 9 13 15 17 18 20 21 25 27 32
+ 34 35 36 41 44 46 49 50 53 56 61 63 67
c155 67 0 3.47682e-19 $X=2.87 $Y=1.44
c156 27 0 2.60212e-20 $X=0.965 $Y=1.59
c157 18 0 1.43299e-19 $X=2.95 $Y=1.99
c158 9 0 2.60212e-20 $X=0.94 $Y=0.445
r159 66 68 43.3814 $w=3.15e-07 $l=1.95e-07 $layer=POLY_cond $X=2.892 $Y=1.44
+ $X2=2.892 $Y2=1.635
r160 66 67 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.44 $X2=2.87 $Y2=1.44
r161 63 66 21.9826 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=2.892 $Y=1.32
+ $X2=2.892 $Y2=1.44
r162 56 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.81 $Y=1.53
+ $X2=2.81 $Y2=1.53
r163 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=1.53
+ $X2=0.69 $Y2=1.53
r164 50 52 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.835 $Y=1.53
+ $X2=0.69 $Y2=1.53
r165 49 56 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=2.81 $Y2=1.53
r166 49 50 2.26485 $w=1.4e-07 $l=1.83e-06 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=0.835 $Y2=1.53
r167 48 53 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=1.795
+ $X2=0.69 $Y2=1.53
r168 47 53 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=0.69 $Y=1.4
+ $X2=0.69 $Y2=1.53
r169 45 61 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r170 44 47 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.235
+ $X2=0.75 $Y2=1.4
r171 44 46 8.51388 $w=2.88e-07 $l=1.65e-07 $layer=LI1_cond $X=0.75 $Y=1.235
+ $X2=0.75 $Y2=1.07
r172 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r173 38 46 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=0.805
+ $X2=0.69 $Y2=1.07
r174 37 41 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.88
+ $X2=0.24 $Y2=1.88
r175 36 48 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.69 $Y2=1.795
r176 36 37 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.395 $Y2=1.88
r177 34 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.69 $Y2=0.805
r178 34 35 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.395 $Y2=0.72
r179 30 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.395 $Y2=0.72
r180 30 32 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.31 $Y2=0.445
r181 23 25 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.465 $Y=1.245
+ $X2=3.465 $Y2=0.445
r182 22 63 20.1192 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=3.05 $Y=1.32
+ $X2=2.892 $Y2=1.32
r183 21 23 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.465 $Y2=1.245
r184 21 22 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.05 $Y2=1.32
r185 18 20 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99
+ $X2=2.95 $Y2=2.275
r186 17 18 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r187 17 68 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=2.95 $Y=1.89
+ $X2=2.95 $Y2=1.635
r188 13 27 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=1.59
r189 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r190 11 61 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.235
r191 11 27 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.59
r192 7 61 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r193 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r194 2 41 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r195 1 32 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%D 2 3 5 8 10 11 12
c43 12 0 5.01492e-20 $X=1.61 $Y=1.19
c44 2 0 1.74491e-19 $X=1.955 $Y=1.67
r45 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r46 10 15 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.6 $Y2=1.16
r47 10 11 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.955 $Y2=1.16
r48 6 11 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.955 $Y2=1.16
r49 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.445
r50 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r52 1 11 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.16
r53 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%A_319_369# 1 2 8 9 11 14 17 20 23 27 30 32
c78 32 0 1.14507e-19 $X=2.4 $Y=0.765
c79 30 0 1.2579e-19 $X=2.4 $Y=0.93
c80 17 0 1.74491e-19 $X=1.72 $Y=1.99
r81 30 33 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=1.095
r82 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=0.765
r83 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=0.93 $X2=2.4 $Y2=0.93
r84 27 29 12.2997 $w=3.67e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.03 $Y=0.72
+ $X2=2.4 $Y2=0.93
r85 26 27 8.64305 $w=3.67e-07 $l=2.6e-07 $layer=LI1_cond $X=1.77 $Y=0.72
+ $X2=2.03 $Y2=0.72
r86 20 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.58
r87 19 27 5.25812 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=2.03 $Y2=0.72
r88 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.03 $Y=1.095 $X2=2.03
+ $Y2=1.495
r89 15 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.72 $Y=1.58
+ $X2=2.03 $Y2=1.58
r90 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r91 14 32 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=0.445
+ $X2=2.425 $Y2=0.765
r92 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r93 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r94 8 33 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r95 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r96 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.77 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%A_203_47# 1 2 9 11 13 16 19 20 24 26 28 29
+ 32 35 36
c118 35 0 1.0603e-19 $X=3.365 $Y=1.87
c119 26 0 1.14507e-19 $X=3.21 $Y=0.915
c120 24 0 2.17725e-19 $X=2.945 $Y=0.9
c121 19 0 1.26282e-19 $X=3.21 $Y=1.575
c122 11 0 8.68433e-20 $X=3.42 $Y=1.99
r123 36 46 4.25306 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=3.365 $Y=1.785
+ $X2=3.21 $Y2=1.785
r124 36 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r125 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.365 $Y=1.87
+ $X2=3.365 $Y2=1.87
r126 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.2 $Y=1.87 $X2=1.2
+ $Y2=1.87
r127 29 31 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.345 $Y=1.87
+ $X2=1.2 $Y2=1.87
r128 28 35 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=3.365 $Y2=1.87
r129 28 29 2.32054 $w=1.4e-07 $l=1.875e-06 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=1.345 $Y2=1.87
r130 23 26 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.945 $Y=0.915
+ $X2=3.21 $Y2=0.915
r131 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.945
+ $Y=0.9 $X2=2.945 $Y2=0.9
r132 20 32 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.82 $X2=1.2
+ $Y2=1.87
r133 20 21 7.33542 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=1.82
+ $X2=1.2 $Y2=1.685
r134 19 46 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.21 $Y=1.575
+ $X2=3.21 $Y2=1.785
r135 18 26 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=0.915
r136 18 19 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=1.575
r137 16 21 80.8984 $w=1.68e-07 $l=1.24e-06 $layer=LI1_cond $X=1.15 $Y=0.445
+ $X2=1.15 $Y2=1.685
r138 11 41 48.3784 $w=2.91e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.425 $Y2=1.74
r139 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.42 $Y2=2.275
r140 7 24 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.9
r141 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.415
r142 2 32 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r143 1 16 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.15 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%A_750_21# 1 2 9 11 13 14 16 17 19 20 27 30
+ 33 35 38 39 44 48
c100 9 0 1.26282e-19 $X=3.825 $Y=0.445
r101 48 49 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.16 $X2=5.73 $Y2=1.16
r102 45 48 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.64 $Y=1.19 $X2=5.73
+ $Y2=1.19
r103 43 44 7.23989 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=1.7
+ $X2=5.17 $Y2=1.7
r104 41 43 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=5.027 $Y=1.7
+ $X2=5.04 $Y2=1.7
r105 40 41 13.6896 $w=3.28e-07 $l=3.92e-07 $layer=LI1_cond $X=4.635 $Y=1.7
+ $X2=5.027 $Y2=1.7
r106 37 45 3.44395 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.64 $Y2=1.19
r107 37 38 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.64 $Y2=1.535
r108 35 38 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.64 $Y2=1.535
r109 35 44 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.17 $Y2=1.62
r110 31 41 1.61437 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=5.027 $Y=1.865
+ $X2=5.027 $Y2=1.7
r111 31 33 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=5.027 $Y=1.865
+ $X2=5.027 $Y2=1.96
r112 30 40 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=1.7
r113 30 39 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=0.825
r114 25 39 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.825
r115 25 27 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.38
r116 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.7 $X2=4.105 $Y2=1.7
r117 20 40 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.635 $Y2=1.7
r118 20 22 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.105 $Y2=1.7
r119 17 49 51.486 $w=2.55e-07 $l=2.57391e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.73 $Y2=1.16
r120 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.985
r121 14 49 39.2931 $w=2.55e-07 $l=1.69926e-07 $layer=POLY_cond $X=5.72 $Y=0.995
+ $X2=5.73 $Y2=1.16
r122 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.72 $Y=0.995
+ $X2=5.72 $Y2=0.56
r123 11 23 53.3563 $w=3.12e-07 $l=3.38452e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=4.005 $Y2=1.7
r124 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=3.9 $Y2=2.275
r125 7 23 78.6992 $w=3.12e-07 $l=5.07075e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=4.005 $Y2=1.7
r126 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=3.825 $Y2=0.445
r127 2 43 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=1.62
r128 2 33 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=1.96
r129 1 27 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.495
+ $Y=0.235 $X2=4.62 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%A_604_47# 1 2 7 9 11 14 16 18 22 27 29 30
+ 32 33
c93 30 0 2.92347e-19 $X=3.85 $Y=1.16
c94 29 0 1.43299e-19 $X=3.765 $Y=2.165
r95 35 36 9.46122 $w=2.45e-07 $l=1.9e-07 $layer=LI1_cond $X=3.575 $Y=1.16
+ $X2=3.765 $Y2=1.16
r96 33 39 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.295 $Y=1.16
+ $X2=4.295 $Y2=1.25
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.16 $X2=4.295 $Y2=1.16
r98 30 36 3.97745 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=3.765 $Y2=1.16
r99 30 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=4.295 $Y2=1.16
r100 28 36 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=1.16
r101 28 29 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=2.165
r102 27 35 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r103 26 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.575 $Y=0.565
+ $X2=3.575 $Y2=0.995
r104 22 26 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.575 $Y2=0.565
r105 22 24 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.205 $Y2=0.422
r106 18 29 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.765 $Y2=2.165
r107 18 20 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.185 $Y2=2.275
r108 16 17 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=4.805 $Y=1.25
+ $X2=4.805 $Y2=1.175
r109 14 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.83 $Y=0.56
+ $X2=4.83 $Y2=1.175
r110 9 16 53.8601 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.25
r111 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.985
r112 8 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.43 $Y=1.25
+ $X2=4.295 $Y2=1.25
r113 7 16 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.805 $Y2=1.25
r114 7 8 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.43 $Y2=1.25
r115 2 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.185 $Y2=2.275
r116 1 24 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.235 $X2=3.205 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%RESET_B 1 3 4 6 7
r32 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r33 4 10 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.25 $Y2=1.16
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.275 $Y2=1.985
r35 1 10 39.2931 $w=2.55e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.25 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%VPWR 1 2 3 4 15 19 24 26 30 31 32 34 39 44
+ 57 58 61 64 67
r92 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r93 61 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r95 55 58 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r96 55 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r97 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 52 54 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.635 $Y=2.72
+ $X2=5.29 $Y2=2.72
r99 51 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r100 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r101 48 51 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r102 48 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r103 47 50 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r105 45 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.19 $Y2=2.72
r106 45 47 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 44 52 8.15384 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=4.342 $Y=2.72
+ $X2=4.635 $Y2=2.72
r108 44 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r109 44 67 8.58723 $w=5.83e-07 $l=4.2e-07 $layer=LI1_cond $X=4.342 $Y=2.72
+ $X2=4.342 $Y2=2.3
r110 44 50 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.05 $Y=2.72
+ $X2=3.91 $Y2=2.72
r111 43 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 43 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r113 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 40 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.73 $Y2=2.72
r115 40 42 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 39 64 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.19 $Y2=2.72
r117 39 42 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 34 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.73 $Y2=2.72
r119 34 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r120 32 62 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 32 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 30 54 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r123 30 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.495 $Y2=2.72
r124 29 57 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=6.21 $Y2=2.72
r125 29 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.495 $Y2=2.72
r126 26 28 6.40424 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.51 $Y=1.97
+ $X2=5.51 $Y2=2.15
r127 24 28 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=5.495 $Y=2.34
+ $X2=5.495 $Y2=2.15
r128 22 31 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.72
r129 22 24 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.34
r130 17 64 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r131 17 19 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r132 13 61 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r133 13 15 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.22
r134 4 26 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=1.97
r135 4 24 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=2.34
r136 3 67 300 $w=1.7e-07 $l=6.62156e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.065 $X2=4.545 $Y2=2.3
r137 2 19 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r138 1 15 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%Q 1 2 9 15 16 20 22
r23 21 22 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.18 $Y=1.495
+ $X2=6.18 $Y2=1.19
r24 20 21 6.81796 $w=3.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.095 $Y=1.66
+ $X2=6.095 $Y2=1.495
r25 15 16 2.48556 $w=4.78e-07 $l=8.5e-08 $layer=LI1_cond $X=6.055 $Y=2.34
+ $X2=6.055 $Y2=2.255
r26 11 13 8.3798 $w=4.95e-07 $l=3.4e-07 $layer=LI1_cond $X=6.03 $Y=0.38 $X2=6.03
+ $Y2=0.72
r27 9 22 15.2824 $w=2.28e-07 $l=3.05e-07 $layer=LI1_cond $X=6.18 $Y=0.885
+ $X2=6.18 $Y2=1.19
r28 9 13 7.59129 $w=4.95e-07 $l=2.2798e-07 $layer=LI1_cond $X=6.18 $Y=0.885
+ $X2=6.03 $Y2=0.72
r29 7 20 1.00839 $w=3.98e-07 $l=3.5e-08 $layer=LI1_cond $X=6.095 $Y=1.695
+ $X2=6.095 $Y2=1.66
r30 7 16 16.1342 $w=3.98e-07 $l=5.6e-07 $layer=LI1_cond $X=6.095 $Y=1.695
+ $X2=6.095 $Y2=2.255
r31 2 20 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=1.66
r32 2 15 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=2.34
r33 1 13 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.93 $Y2=0.72
r34 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.795
+ $Y=0.235 $X2=5.93 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTP_1%VGND 1 2 3 4 15 19 23 28 30 31 33 36 38 43
+ 48 61 62 65 68 71
c89 62 0 3.98209e-20 $X=6.21 $Y=0
r90 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r91 68 69 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r92 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r93 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r94 59 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r95 58 59 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r96 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r97 56 72 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r98 55 58 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r99 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r100 53 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.035
+ $Y2=0
r101 53 55 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.37
+ $Y2=0
r102 52 72 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r103 52 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r104 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r105 49 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.19
+ $Y2=0
r106 49 51 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r107 48 71 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.035
+ $Y2=0
r108 48 51 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.87 $Y=0 $X2=2.53
+ $Y2=0
r109 47 69 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r110 47 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r111 46 47 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r112 44 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r113 44 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r114 43 68 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.19
+ $Y2=0
r115 43 46 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=1.15 $Y2=0
r116 38 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r117 38 40 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.23 $Y2=0
r118 36 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r119 36 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r120 33 34 4.37018 $w=3.28e-07 $l=1.15e-07 $layer=LI1_cond $X=5.485 $Y=0.74
+ $X2=5.485 $Y2=0.625
r121 30 58 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.29
+ $Y2=0
r122 30 31 7.54988 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=5.32 $Y=0 $X2=5.457
+ $Y2=0
r123 29 61 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=5.595 $Y=0 $X2=6.21
+ $Y2=0
r124 29 31 7.54988 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=5.595 $Y=0
+ $X2=5.457 $Y2=0
r125 28 34 10.2672 $w=2.73e-07 $l=2.45e-07 $layer=LI1_cond $X=5.457 $Y=0.38
+ $X2=5.457 $Y2=0.625
r126 25 31 0.316938 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=5.457 $Y=0.085
+ $X2=5.457 $Y2=0
r127 25 28 12.3626 $w=2.73e-07 $l=2.95e-07 $layer=LI1_cond $X=5.457 $Y=0.085
+ $X2=5.457 $Y2=0.38
r128 21 71 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0
r129 21 23 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0.445
r130 17 68 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r131 17 19 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.36
r132 13 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r133 13 15 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r134 4 33 182 $w=1.7e-07 $l=5.86003e-07 $layer=licon1_NDIFF $count=1 $X=5.31
+ $Y=0.235 $X2=5.485 $Y2=0.74
r135 4 28 182 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=1 $X=5.31
+ $Y=0.235 $X2=5.485 $Y2=0.38
r136 3 23 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.035 $Y2=0.445
r137 2 19 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r138 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

