* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xor3_4 A B C VGND VNB VPB VPWR X
X0 VGND a_80_207# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_1225_365# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 a_658_49# a_1109_297# a_1225_365# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X3 a_80_207# a_528_297# a_652_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X4 VPWR a_80_207# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_80_207# a_528_297# a_658_49# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X6 a_652_325# a_1109_297# a_1225_365# VNB sky130_fd_pr__nfet_01v8 w=600000u l=150000u
X7 X a_80_207# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR a_1225_365# a_1510_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_1510_297# B a_652_325# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X10 X a_80_207# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_652_325# a_1109_297# a_1510_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X12 VPWR B a_1109_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_1225_365# B a_652_325# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X14 X a_80_207# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 VGND B a_1109_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VGND a_80_207# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_652_325# C a_80_207# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X18 a_1510_297# B a_658_49# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X19 VGND C a_528_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_658_49# C a_80_207# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X21 a_1225_365# A VGND VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X22 VPWR C a_528_297# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X23 VGND a_1225_365# a_1510_297# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X24 X a_80_207# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_658_49# a_1109_297# a_1510_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VPWR a_80_207# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_1225_365# B a_658_49# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
.ends
