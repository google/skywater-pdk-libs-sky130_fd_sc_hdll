# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a31oi_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a31oi_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.060000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.330000 0.995000 3.090000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.150000 0.995000 1.905000 1.615000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.145000 0.995000 0.870000 1.615000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.220000 1.075000 4.940000 1.275000 ;
        RECT 4.715000 1.275000 4.940000 1.625000 ;
    END
  END B1
  PIN VGND
    ANTENNADIFFAREA  0.468000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.060000 0.085000 ;
        RECT 0.515000  0.085000 0.895000 0.465000 ;
        RECT 4.025000  0.085000 4.405000 0.465000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.060000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.470000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.060000 2.805000 ;
        RECT 0.515000 2.125000 0.895000 2.635000 ;
        RECT 1.455000 2.125000 1.835000 2.635000 ;
        RECT 2.560000 2.125000 3.280000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.060000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.007000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.545000 0.655000 4.955000 0.825000 ;
        RECT 3.330000 0.825000 4.955000 0.845000 ;
        RECT 3.330000 0.845000 3.645000 1.445000 ;
        RECT 3.330000 1.445000 4.485000 1.615000 ;
        RECT 3.605000 0.255000 3.775000 0.655000 ;
        RECT 4.155000 1.615000 4.485000 2.115000 ;
        RECT 4.575000 0.295000 4.955000 0.655000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.095000 0.655000 2.305000 0.825000 ;
      RECT 0.175000 1.785000 3.855000 1.955000 ;
      RECT 0.175000 1.955000 0.345000 2.465000 ;
      RECT 1.115000 1.955000 1.285000 2.465000 ;
      RECT 1.455000 0.295000 3.375000 0.465000 ;
      RECT 2.055000 1.955000 2.225000 2.465000 ;
      RECT 3.685000 1.955000 3.855000 2.295000 ;
      RECT 3.685000 2.295000 4.875000 2.465000 ;
      RECT 4.705000 1.795000 4.875000 2.295000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a31oi_2
