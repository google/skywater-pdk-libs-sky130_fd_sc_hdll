* File: sky130_fd_sc_hdll__inv_12.pex.spice
* Created: Thu Aug 27 19:08:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__INV_12%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22 24
+ 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 58 60 61 63
+ 64 66 67 69 70 72 73 74 75 76 77 78 79 80 81 118 119 124 127 132 135 138 142
+ 144 147
r236 142 144 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.29 $Y=1.2
+ $X2=4.67 $Y2=1.2
r237 119 120 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.83 $Y=1.202
+ $X2=5.855 $Y2=1.202
r238 117 119 30.8638 $w=3.67e-07 $l=2.35e-07 $layer=POLY_cond $X=5.595 $Y=1.202
+ $X2=5.83 $Y2=1.202
r239 117 118 26.4145 $w=1.7e-07 $l=9.35e-07 $layer=licon1_POLY $count=5 $X=5.595
+ $Y=1.16 $X2=5.595 $Y2=1.16
r240 115 117 30.8638 $w=3.67e-07 $l=2.35e-07 $layer=POLY_cond $X=5.36 $Y=1.202
+ $X2=5.595 $Y2=1.202
r241 114 115 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=5.335 $Y=1.202
+ $X2=5.36 $Y2=1.202
r242 113 114 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=4.89 $Y=1.202
+ $X2=5.335 $Y2=1.202
r243 112 113 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.865 $Y=1.202
+ $X2=4.89 $Y2=1.202
r244 111 112 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=4.42 $Y=1.202
+ $X2=4.865 $Y2=1.202
r245 110 111 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.395 $Y=1.202
+ $X2=4.42 $Y2=1.202
r246 109 110 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=3.95 $Y=1.202
+ $X2=4.395 $Y2=1.202
r247 108 109 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.925 $Y=1.202
+ $X2=3.95 $Y2=1.202
r248 107 108 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=3.48 $Y=1.202
+ $X2=3.925 $Y2=1.202
r249 106 107 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=3.455 $Y=1.202
+ $X2=3.48 $Y2=1.202
r250 105 106 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=3.01 $Y=1.202
+ $X2=3.455 $Y2=1.202
r251 104 105 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.985 $Y=1.202
+ $X2=3.01 $Y2=1.202
r252 103 104 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=2.54 $Y=1.202
+ $X2=2.985 $Y2=1.202
r253 102 103 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.515 $Y=1.202
+ $X2=2.54 $Y2=1.202
r254 101 102 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=2.07 $Y=1.202
+ $X2=2.515 $Y2=1.202
r255 100 101 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.045 $Y=1.202
+ $X2=2.07 $Y2=1.202
r256 99 100 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=1.6 $Y=1.202
+ $X2=2.045 $Y2=1.202
r257 98 99 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.575 $Y=1.202
+ $X2=1.6 $Y2=1.202
r258 97 98 58.4441 $w=3.67e-07 $l=4.45e-07 $layer=POLY_cond $X=1.13 $Y=1.202
+ $X2=1.575 $Y2=1.202
r259 96 97 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=1.105 $Y=1.202
+ $X2=1.13 $Y2=1.202
r260 95 124 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=1.2
+ $X2=1.15 $Y2=1.2
r261 94 96 27.5804 $w=3.67e-07 $l=2.1e-07 $layer=POLY_cond $X=0.895 $Y=1.202
+ $X2=1.105 $Y2=1.202
r262 94 95 26.4145 $w=1.7e-07 $l=9.35e-07 $layer=licon1_POLY $count=5 $X=0.895
+ $Y=1.16 $X2=0.895 $Y2=1.16
r263 92 94 30.8638 $w=3.67e-07 $l=2.35e-07 $layer=POLY_cond $X=0.66 $Y=1.202
+ $X2=0.895 $Y2=1.202
r264 91 92 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.635 $Y=1.202
+ $X2=0.66 $Y2=1.202
r265 81 118 19.5915 $w=2.48e-07 $l=4.25e-07 $layer=LI1_cond $X=5.17 $Y=1.2
+ $X2=5.595 $Y2=1.2
r266 81 147 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.17 $Y=1.2 $X2=5.09
+ $Y2=1.2
r267 80 147 16.1342 $w=2.48e-07 $l=3.5e-07 $layer=LI1_cond $X=4.74 $Y=1.2
+ $X2=5.09 $Y2=1.2
r268 80 144 3.22684 $w=2.48e-07 $l=7e-08 $layer=LI1_cond $X=4.74 $Y=1.2 $X2=4.67
+ $Y2=1.2
r269 79 142 2.76586 $w=2.48e-07 $l=6e-08 $layer=LI1_cond $X=4.23 $Y=1.2 $X2=4.29
+ $Y2=1.2
r270 78 79 35.2648 $w=2.48e-07 $l=7.65e-07 $layer=LI1_cond $X=3.465 $Y=1.2
+ $X2=4.23 $Y2=1.2
r271 78 138 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.465 $Y=1.2
+ $X2=3.45 $Y2=1.2
r272 77 138 20.5135 $w=2.48e-07 $l=4.45e-07 $layer=LI1_cond $X=3.005 $Y=1.2
+ $X2=3.45 $Y2=1.2
r273 77 135 0.691466 $w=2.48e-07 $l=1.5e-08 $layer=LI1_cond $X=3.005 $Y=1.2
+ $X2=2.99 $Y2=1.2
r274 76 135 20.9745 $w=2.48e-07 $l=4.55e-07 $layer=LI1_cond $X=2.535 $Y=1.2
+ $X2=2.99 $Y2=1.2
r275 76 132 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=2.535 $Y=1.2
+ $X2=2.53 $Y2=1.2
r276 75 132 21.205 $w=2.48e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=1.2
+ $X2=2.53 $Y2=1.2
r277 74 75 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=1.635 $Y=1.2
+ $X2=2.07 $Y2=1.2
r278 74 127 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=1.635 $Y=1.2
+ $X2=1.61 $Y2=1.2
r279 73 127 20.0525 $w=2.48e-07 $l=4.35e-07 $layer=LI1_cond $X=1.175 $Y=1.2
+ $X2=1.61 $Y2=1.2
r280 73 124 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=1.2
+ $X2=1.15 $Y2=1.2
r281 70 120 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.855 $Y=0.995
+ $X2=5.855 $Y2=1.202
r282 70 72 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.855 $Y=0.995
+ $X2=5.855 $Y2=0.56
r283 67 119 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.83 $Y=1.41
+ $X2=5.83 $Y2=1.202
r284 67 69 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.83 $Y=1.41
+ $X2=5.83 $Y2=1.985
r285 64 115 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.36 $Y=1.41
+ $X2=5.36 $Y2=1.202
r286 64 66 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.36 $Y=1.41
+ $X2=5.36 $Y2=1.985
r287 61 114 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.335 $Y=0.995
+ $X2=5.335 $Y2=1.202
r288 61 63 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.335 $Y=0.995
+ $X2=5.335 $Y2=0.56
r289 58 113 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.89 $Y=1.41
+ $X2=4.89 $Y2=1.202
r290 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.89 $Y=1.41
+ $X2=4.89 $Y2=1.985
r291 55 112 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.865 $Y=0.995
+ $X2=4.865 $Y2=1.202
r292 55 57 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.865 $Y=0.995
+ $X2=4.865 $Y2=0.56
r293 52 111 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.42 $Y=1.41
+ $X2=4.42 $Y2=1.202
r294 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.42 $Y=1.41
+ $X2=4.42 $Y2=1.985
r295 49 110 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.395 $Y=0.995
+ $X2=4.395 $Y2=1.202
r296 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.395 $Y=0.995
+ $X2=4.395 $Y2=0.56
r297 46 109 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.202
r298 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.985
r299 43 108 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.925 $Y=0.995
+ $X2=3.925 $Y2=1.202
r300 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.925 $Y=0.995
+ $X2=3.925 $Y2=0.56
r301 40 107 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.48 $Y2=1.202
r302 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.48 $Y=1.41
+ $X2=3.48 $Y2=1.985
r303 37 106 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=1.202
r304 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.455 $Y=0.995
+ $X2=3.455 $Y2=0.56
r305 34 105 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.01 $Y=1.41
+ $X2=3.01 $Y2=1.202
r306 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.01 $Y=1.41
+ $X2=3.01 $Y2=1.985
r307 31 104 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.985 $Y2=1.202
r308 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.985 $Y2=0.56
r309 28 103 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.54 $Y=1.41
+ $X2=2.54 $Y2=1.202
r310 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.54 $Y=1.41
+ $X2=2.54 $Y2=1.985
r311 25 102 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=1.202
r312 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.515 $Y=0.995
+ $X2=2.515 $Y2=0.56
r313 22 101 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.07 $Y=1.41
+ $X2=2.07 $Y2=1.202
r314 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.07 $Y=1.41
+ $X2=2.07 $Y2=1.985
r315 19 100 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.045 $Y2=1.202
r316 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.045 $Y=0.995
+ $X2=2.045 $Y2=0.56
r317 16 99 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.6 $Y=1.41
+ $X2=1.6 $Y2=1.202
r318 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.6 $Y=1.41
+ $X2=1.6 $Y2=1.985
r319 13 98 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.575 $Y=0.995
+ $X2=1.575 $Y2=1.202
r320 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.575 $Y=0.995
+ $X2=1.575 $Y2=0.56
r321 10 97 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.202
r322 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.13 $Y=1.41
+ $X2=1.13 $Y2=1.985
r323 7 96 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=1.202
r324 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.105 $Y=0.995
+ $X2=1.105 $Y2=0.56
r325 4 92 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.66 $Y=1.41
+ $X2=0.66 $Y2=1.202
r326 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.66 $Y=1.41
+ $X2=0.66 $Y2=1.985
r327 1 91 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=1.202
r328 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.635 $Y=0.995
+ $X2=0.635 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_12%VPWR 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46
+ 48 51 52 54 55 57 58 60 61 63 64 65 83 92
c102 7 0 4.98153e-20 $X=5.92 $Y=1.485
r103 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r104 86 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.21 $Y2=2.72
r105 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r106 83 91 3.94577 $w=1.7e-07 $l=2.32e-07 $layer=LI1_cond $X=5.975 $Y=2.72
+ $X2=6.207 $Y2=2.72
r107 83 85 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=5.975 $Y=2.72
+ $X2=5.75 $Y2=2.72
r108 82 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r110 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r112 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r114 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r115 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r116 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 67 88 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=0.255 $Y2=2.72
r119 67 69 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 65 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r121 65 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 63 81 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.04 $Y=2.72
+ $X2=4.83 $Y2=2.72
r123 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=2.72
+ $X2=5.125 $Y2=2.72
r124 62 85 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r125 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=2.72
+ $X2=5.125 $Y2=2.72
r126 60 78 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=2.72
+ $X2=4.185 $Y2=2.72
r128 59 81 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.27 $Y=2.72
+ $X2=4.83 $Y2=2.72
r129 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=2.72
+ $X2=4.185 $Y2=2.72
r130 57 75 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=2.99 $Y2=2.72
r131 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=2.72
+ $X2=3.245 $Y2=2.72
r132 56 78 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.91 $Y2=2.72
r133 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=2.72
+ $X2=3.245 $Y2=2.72
r134 54 72 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.07 $Y2=2.72
r135 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=2.72
+ $X2=2.305 $Y2=2.72
r136 53 75 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.39 $Y=2.72 $X2=2.99
+ $Y2=2.72
r137 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=2.72
+ $X2=2.305 $Y2=2.72
r138 51 69 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.15 $Y2=2.72
r139 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=2.72
+ $X2=1.365 $Y2=2.72
r140 50 72 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r141 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=2.72
+ $X2=1.365 $Y2=2.72
r142 46 91 3.23145 $w=2.55e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.102 $Y=2.635
+ $X2=6.207 $Y2=2.72
r143 46 48 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=6.102 $Y=2.635
+ $X2=6.102 $Y2=2
r144 42 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=2.635
+ $X2=5.125 $Y2=2.72
r145 42 44 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.125 $Y=2.635
+ $X2=5.125 $Y2=2
r146 38 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=2.635
+ $X2=4.185 $Y2=2.72
r147 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.185 $Y=2.635
+ $X2=4.185 $Y2=2
r148 34 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=2.635
+ $X2=3.245 $Y2=2.72
r149 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.245 $Y=2.635
+ $X2=3.245 $Y2=2
r150 30 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=2.635
+ $X2=2.305 $Y2=2.72
r151 30 32 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.305 $Y=2.635
+ $X2=2.305 $Y2=2
r152 26 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2.72
r153 26 28 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.365 $Y=2.635
+ $X2=1.365 $Y2=2
r154 22 88 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.255 $Y2=2.72
r155 22 24 28.6981 $w=2.53e-07 $l=6.35e-07 $layer=LI1_cond $X=0.382 $Y=2.635
+ $X2=0.382 $Y2=2
r156 7 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.92
+ $Y=1.485 $X2=6.065 $Y2=2
r157 6 44 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.98
+ $Y=1.485 $X2=5.125 $Y2=2
r158 5 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.04
+ $Y=1.485 $X2=4.185 $Y2=2
r159 4 36 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.1
+ $Y=1.485 $X2=3.245 $Y2=2
r160 3 32 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.16
+ $Y=1.485 $X2=2.305 $Y2=2
r161 2 28 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.22
+ $Y=1.485 $X2=1.365 $Y2=2
r162 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.3
+ $Y=1.485 $X2=0.425 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_12%Y 1 2 3 4 5 6 7 8 9 10 11 12 39 43 45 46 47
+ 48 51 55 57 59 63 67 69 71 75 79 81 83 87 91 93 95 99 103 105 107 118 120 121
+ 123 124 126 127 129 130 132 135 136
c257 136 0 4.98153e-20 $X=6.18 $Y=1.19
r258 134 136 10.0427 $w=3.48e-07 $l=3.05e-07 $layer=LI1_cond $X=6.145 $Y=1.495
+ $X2=6.145 $Y2=1.19
r259 133 136 9.38418 $w=3.48e-07 $l=2.85e-07 $layer=LI1_cond $X=6.145 $Y=0.905
+ $X2=6.145 $Y2=1.19
r260 114 135 8.27047 $w=4.23e-07 $l=3.05e-07 $layer=LI1_cond $X=0.297 $Y=1.495
+ $X2=0.297 $Y2=1.19
r261 110 135 7.72815 $w=4.23e-07 $l=2.85e-07 $layer=LI1_cond $X=0.297 $Y=0.905
+ $X2=0.297 $Y2=1.19
r262 108 132 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.76 $Y=1.58
+ $X2=5.57 $Y2=1.58
r263 107 134 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=6.145 $Y2=1.495
r264 107 108 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.97 $Y=1.58
+ $X2=5.76 $Y2=1.58
r265 106 130 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.76 $Y=0.81
+ $X2=5.57 $Y2=0.81
r266 105 133 7.62524 $w=1.9e-07 $l=2.17371e-07 $layer=LI1_cond $X=5.97 $Y=0.81
+ $X2=6.145 $Y2=0.905
r267 105 106 12.2584 $w=1.88e-07 $l=2.1e-07 $layer=LI1_cond $X=5.97 $Y=0.81
+ $X2=5.76 $Y2=0.81
r268 101 132 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.57 $Y=1.665
+ $X2=5.57 $Y2=1.58
r269 101 103 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.57 $Y=1.665
+ $X2=5.57 $Y2=2.34
r270 97 130 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.57 $Y=0.715
+ $X2=5.57 $Y2=0.81
r271 97 99 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.57 $Y=0.715
+ $X2=5.57 $Y2=0.38
r272 96 129 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.82 $Y=1.58
+ $X2=4.63 $Y2=1.58
r273 95 132 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.38 $Y=1.58
+ $X2=5.57 $Y2=1.58
r274 95 96 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.38 $Y=1.58
+ $X2=4.82 $Y2=1.58
r275 94 127 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.82 $Y=0.81
+ $X2=4.63 $Y2=0.81
r276 93 130 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.38 $Y=0.81
+ $X2=5.57 $Y2=0.81
r277 93 94 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=5.38 $Y=0.81
+ $X2=4.82 $Y2=0.81
r278 89 129 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.63 $Y=1.665
+ $X2=4.63 $Y2=1.58
r279 89 91 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.63 $Y=1.665
+ $X2=4.63 $Y2=2.34
r280 85 127 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=4.63 $Y=0.715
+ $X2=4.63 $Y2=0.81
r281 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.63 $Y=0.715
+ $X2=4.63 $Y2=0.38
r282 84 126 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.88 $Y=1.58
+ $X2=3.69 $Y2=1.58
r283 83 129 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.44 $Y=1.58
+ $X2=4.63 $Y2=1.58
r284 83 84 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.44 $Y=1.58
+ $X2=3.88 $Y2=1.58
r285 82 124 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.88 $Y=0.81
+ $X2=3.69 $Y2=0.81
r286 81 127 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=4.44 $Y=0.81
+ $X2=4.63 $Y2=0.81
r287 81 82 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=4.44 $Y=0.81
+ $X2=3.88 $Y2=0.81
r288 77 126 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=1.58
r289 77 79 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=3.69 $Y=1.665
+ $X2=3.69 $Y2=2.34
r290 73 124 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=3.69 $Y=0.715
+ $X2=3.69 $Y2=0.81
r291 73 75 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.69 $Y=0.715
+ $X2=3.69 $Y2=0.38
r292 72 123 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.94 $Y=1.58
+ $X2=2.75 $Y2=1.58
r293 71 126 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.5 $Y=1.58
+ $X2=3.69 $Y2=1.58
r294 71 72 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.5 $Y=1.58
+ $X2=2.94 $Y2=1.58
r295 70 121 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.94 $Y=0.81
+ $X2=2.75 $Y2=0.81
r296 69 124 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=3.5 $Y=0.81
+ $X2=3.69 $Y2=0.81
r297 69 70 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=3.5 $Y=0.81 $X2=2.94
+ $Y2=0.81
r298 65 123 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=1.665
+ $X2=2.75 $Y2=1.58
r299 65 67 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=2.75 $Y=1.665
+ $X2=2.75 $Y2=2.34
r300 61 121 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=2.75 $Y=0.715
+ $X2=2.75 $Y2=0.81
r301 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.75 $Y=0.715
+ $X2=2.75 $Y2=0.38
r302 60 120 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2 $Y=1.58 $X2=1.81
+ $Y2=1.58
r303 59 123 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=1.58
+ $X2=2.75 $Y2=1.58
r304 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.56 $Y=1.58 $X2=2
+ $Y2=1.58
r305 58 118 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2 $Y=0.81 $X2=1.81
+ $Y2=0.81
r306 57 121 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=0.81
+ $X2=2.75 $Y2=0.81
r307 57 58 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=2.56 $Y=0.81 $X2=2
+ $Y2=0.81
r308 53 120 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.81 $Y=1.665
+ $X2=1.81 $Y2=1.58
r309 53 55 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.81 $Y=1.665
+ $X2=1.81 $Y2=2.34
r310 49 118 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=1.81 $Y=0.715
+ $X2=1.81 $Y2=0.81
r311 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.81 $Y=0.715
+ $X2=1.81 $Y2=0.38
r312 47 120 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=1.58
+ $X2=1.81 $Y2=1.58
r313 47 48 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.62 $Y=1.58
+ $X2=1.06 $Y2=1.58
r314 45 118 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=1.62 $Y=0.81
+ $X2=1.81 $Y2=0.81
r315 45 46 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=1.62 $Y=0.81
+ $X2=1.06 $Y2=0.81
r316 41 48 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.87 $Y=1.58
+ $X2=1.06 $Y2=1.58
r317 41 114 37.3829 $w=1.68e-07 $l=5.73e-07 $layer=LI1_cond $X=0.87 $Y=1.58
+ $X2=0.297 $Y2=1.58
r318 41 43 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=0.87 $Y=1.665
+ $X2=0.87 $Y2=2.34
r319 37 46 11.0909 $w=1.88e-07 $l=1.9e-07 $layer=LI1_cond $X=0.87 $Y=0.81
+ $X2=1.06 $Y2=0.81
r320 37 110 33.4478 $w=1.88e-07 $l=5.73e-07 $layer=LI1_cond $X=0.87 $Y=0.81
+ $X2=0.297 $Y2=0.81
r321 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.87 $Y=0.715
+ $X2=0.87 $Y2=0.38
r322 12 132 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.45
+ $Y=1.485 $X2=5.595 $Y2=1.66
r323 12 103 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.45
+ $Y=1.485 $X2=5.595 $Y2=2.34
r324 11 129 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.485 $X2=4.655 $Y2=1.66
r325 11 91 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.51
+ $Y=1.485 $X2=4.655 $Y2=2.34
r326 10 126 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.485 $X2=3.715 $Y2=1.66
r327 10 79 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.57
+ $Y=1.485 $X2=3.715 $Y2=2.34
r328 9 123 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.775 $Y2=1.66
r329 9 67 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.775 $Y2=2.34
r330 8 120 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.835 $Y2=1.66
r331 8 55 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.69
+ $Y=1.485 $X2=1.835 $Y2=2.34
r332 7 41 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.895 $Y2=1.66
r333 7 43 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.75
+ $Y=1.485 $X2=0.895 $Y2=2.34
r334 6 99 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=5.41
+ $Y=0.235 $X2=5.595 $Y2=0.38
r335 5 87 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.47
+ $Y=0.235 $X2=4.655 $Y2=0.38
r336 4 75 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=3.53
+ $Y=0.235 $X2=3.715 $Y2=0.38
r337 3 63 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=2.59
+ $Y=0.235 $X2=2.775 $Y2=0.38
r338 2 51 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=1.65
+ $Y=0.235 $X2=1.835 $Y2=0.38
r339 1 39 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=0.71
+ $Y=0.235 $X2=0.895 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__INV_12%VGND 1 2 3 4 5 6 7 22 24 28 32 36 40 44 46
+ 48 51 52 54 55 57 58 60 61 63 64 65 83 92
r114 91 92 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r115 86 92 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r116 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r117 83 91 4.06587 $w=1.7e-07 $l=2.4e-07 $layer=LI1_cond $X=5.96 $Y=0 $X2=6.2
+ $Y2=0
r118 83 85 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.96 $Y=0 $X2=5.75
+ $Y2=0
r119 82 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r120 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r121 79 82 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r122 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r123 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r124 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r125 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r126 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r127 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r128 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r129 67 88 3.91904 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=0.255
+ $Y2=0
r130 67 69 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=0.51 $Y=0 $X2=1.15
+ $Y2=0
r131 65 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r132 65 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r133 63 81 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.04 $Y=0 $X2=4.83
+ $Y2=0
r134 63 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.04 $Y=0 $X2=5.125
+ $Y2=0
r135 62 85 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.75
+ $Y2=0
r136 62 64 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.21 $Y=0 $X2=5.125
+ $Y2=0
r137 60 78 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=4.1 $Y=0 $X2=3.91
+ $Y2=0
r138 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0 $X2=4.185
+ $Y2=0
r139 59 81 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.83
+ $Y2=0
r140 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.27 $Y=0 $X2=4.185
+ $Y2=0
r141 57 75 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.16 $Y=0 $X2=2.99
+ $Y2=0
r142 57 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.16 $Y=0 $X2=3.245
+ $Y2=0
r143 56 78 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.91
+ $Y2=0
r144 56 58 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.33 $Y=0 $X2=3.245
+ $Y2=0
r145 54 72 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.07
+ $Y2=0
r146 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.22 $Y=0 $X2=2.305
+ $Y2=0
r147 53 75 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.99
+ $Y2=0
r148 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.39 $Y=0 $X2=2.305
+ $Y2=0
r149 51 69 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.15
+ $Y2=0
r150 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.28 $Y=0 $X2=1.365
+ $Y2=0
r151 50 72 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.45 $Y=0 $X2=2.07
+ $Y2=0
r152 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.45 $Y=0 $X2=1.365
+ $Y2=0
r153 46 91 3.21882 $w=2.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.095 $Y=0.085
+ $X2=6.2 $Y2=0
r154 46 48 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.095 $Y=0.085
+ $X2=6.095 $Y2=0.38
r155 42 64 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0
r156 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.125 $Y=0.085
+ $X2=5.125 $Y2=0.38
r157 38 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.185 $Y=0.085
+ $X2=4.185 $Y2=0
r158 38 40 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.185 $Y=0.085
+ $X2=4.185 $Y2=0.38
r159 34 58 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0
r160 34 36 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.245 $Y=0.085
+ $X2=3.245 $Y2=0.38
r161 30 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0
r162 30 32 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.305 $Y=0.085
+ $X2=2.305 $Y2=0.38
r163 26 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0
r164 26 28 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.365 $Y=0.085
+ $X2=1.365 $Y2=0.38
r165 22 88 3.25818 $w=2.55e-07 $l=1.64085e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.255 $Y2=0
r166 22 24 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.382 $Y=0.085
+ $X2=0.382 $Y2=0.38
r167 7 48 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.93
+ $Y=0.235 $X2=6.065 $Y2=0.38
r168 6 44 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.94
+ $Y=0.235 $X2=5.125 $Y2=0.38
r169 5 40 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.185 $Y2=0.38
r170 4 36 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.235 $X2=3.245 $Y2=0.38
r171 3 32 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.235 $X2=2.305 $Y2=0.38
r172 2 28 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=1.18
+ $Y=0.235 $X2=1.365 $Y2=0.38
r173 1 24 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.38
.ends

