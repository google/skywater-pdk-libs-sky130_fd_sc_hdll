* File: sky130_fd_sc_hdll__clkbuf_4.pxi.spice
* Created: Thu Aug 27 19:01:49 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_4%A N_A_c_61_n N_A_M1003_g N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__CLKBUF_4%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_4%A_27_47# N_A_27_47#_M1000_s N_A_27_47#_M1003_s
+ N_A_27_47#_M1001_g N_A_27_47#_c_107_n N_A_27_47#_M1004_g N_A_27_47#_M1002_g
+ N_A_27_47#_c_108_n N_A_27_47#_M1006_g N_A_27_47#_c_96_n N_A_27_47#_M1005_g
+ N_A_27_47#_c_109_n N_A_27_47#_M1007_g N_A_27_47#_c_98_n N_A_27_47#_c_110_n
+ N_A_27_47#_M1008_g N_A_27_47#_M1009_g N_A_27_47#_c_100_n N_A_27_47#_c_101_n
+ N_A_27_47#_c_102_n N_A_27_47#_c_103_n N_A_27_47#_c_104_n N_A_27_47#_c_115_n
+ N_A_27_47#_c_127_n N_A_27_47#_c_116_n N_A_27_47#_c_131_n N_A_27_47#_c_159_p
+ N_A_27_47#_c_105_n N_A_27_47#_c_106_n N_A_27_47#_c_118_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_4%VPWR N_VPWR_M1003_d N_VPWR_M1006_d
+ N_VPWR_M1008_d N_VPWR_c_201_n N_VPWR_c_202_n N_VPWR_c_203_n N_VPWR_c_204_n
+ N_VPWR_c_205_n N_VPWR_c_206_n N_VPWR_c_207_n VPWR N_VPWR_c_208_n
+ N_VPWR_c_200_n N_VPWR_c_210_n PM_SKY130_FD_SC_HDLL__CLKBUF_4%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_4%X N_X_M1001_d N_X_M1005_d N_X_M1004_s
+ N_X_M1007_s N_X_c_245_n N_X_c_290_n N_X_c_246_n N_X_c_247_n N_X_c_267_n
+ N_X_c_271_n N_X_c_248_n N_X_c_297_n X X X N_X_c_251_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_4%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_4%VGND N_VGND_M1000_d N_VGND_M1002_s
+ N_VGND_M1009_s N_VGND_c_315_n N_VGND_c_316_n N_VGND_c_317_n N_VGND_c_318_n
+ N_VGND_c_319_n N_VGND_c_320_n N_VGND_c_321_n VGND N_VGND_c_322_n
+ N_VGND_c_323_n N_VGND_c_324_n N_VGND_c_325_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_4%VGND
cc_1 VNB N_A_c_61_n 0.0290211f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_2 VNB N_A_M1000_g 0.0338609f $X=-0.19 $Y=-0.24 $X2=0.525 $Y2=0.445
cc_3 VNB A 0.00882584f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=0.765
cc_4 VNB N_A_27_47#_M1001_g 0.0305549f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.105
cc_5 VNB N_A_27_47#_M1002_g 0.0297352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_c_96_n 0.0205679f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1005_g 0.030394f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_98_n 0.0193336f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1009_g 0.0378445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_100_n 0.0112911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_101_n 0.0202094f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_102_n 0.00639652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_103_n 0.0143585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_104_n 0.0331263f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_105_n 0.0063974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_106_n 0.0131987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VPWR_c_200_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_X_c_245_n 7.7005e-19 $X=-0.19 $Y=-0.24 $X2=0.625 $Y2=0.85
cc_19 VNB N_X_c_246_n 0.00738088f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_X_c_247_n 0.0025078f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_X_c_248_n 0.00154712f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB X 0.0341382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_315_n 0.00528656f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_24 VNB N_VGND_c_316_n 0.00520797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_317_n 0.0053486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_318_n 0.0200491f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_319_n 0.0048778f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_320_n 0.018696f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_321_n 0.00535855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_322_n 0.0179145f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_323_n 0.0132796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_324_n 0.189653f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_325_n 0.0052624f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_c_61_n 0.0313201f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_35 VPB A 0.00221606f $X=-0.19 $Y=1.305 $X2=0.655 $Y2=0.765
cc_36 VPB N_A_27_47#_c_107_n 0.0166394f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A_27_47#_c_108_n 0.0164072f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_38 VPB N_A_27_47#_c_109_n 0.0163105f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_A_27_47#_c_110_n 0.01843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_A_27_47#_c_100_n 0.00630734f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_47#_c_102_n 0.00650179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_47#_c_103_n 0.0076017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_43 VPB N_A_27_47#_c_104_n 0.00911296f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_47#_c_115_n 0.0313553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_A_27_47#_c_116_n 0.00182082f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_105_n 0.00651103f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_27_47#_c_118_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_201_n 0.00550303f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.16
cc_49 VPB N_VPWR_c_202_n 0.00466331f $X=-0.19 $Y=1.305 $X2=0.625 $Y2=1.16
cc_50 VPB N_VPWR_c_203_n 0.026657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_204_n 0.0189422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_VPWR_c_205_n 0.00487698f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_VPWR_c_206_n 0.0167627f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_VPWR_c_207_n 0.00516759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_VPWR_c_208_n 0.0131219f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_VPWR_c_200_n 0.0536295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_210_n 0.0247531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB X 0.00595667f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_X_c_251_n 0.0151804f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 N_A_c_61_n N_A_27_47#_M1001_g 0.0184312f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_M1000_g N_A_27_47#_M1001_g 0.0187281f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_62 A N_A_27_47#_M1001_g 0.00771044f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_63 N_A_c_61_n N_A_27_47#_c_107_n 0.0278268f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_61_n N_A_27_47#_c_100_n 0.00306202f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_61_n N_A_27_47#_c_104_n 0.0142883f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_M1000_g N_A_27_47#_c_104_n 0.00676678f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_67 A N_A_27_47#_c_104_n 0.0444892f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_68 N_A_c_61_n N_A_27_47#_c_127_n 0.0165266f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_69 A N_A_27_47#_c_127_n 0.0289325f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_70 N_A_c_61_n N_A_27_47#_c_116_n 0.00100022f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_71 A N_A_27_47#_c_116_n 0.00621264f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_72 A N_A_27_47#_c_131_n 0.014474f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_73 N_A_c_61_n N_A_27_47#_c_106_n 0.0012545f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_61_n N_A_27_47#_c_118_n 0.00120597f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_61_n N_VPWR_c_201_n 0.00313892f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_61_n N_VPWR_c_200_n 0.0134989f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_61_n N_VPWR_c_210_n 0.00702461f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_M1000_g N_X_c_245_n 7.69134e-19 $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_79 N_A_M1000_g N_X_c_247_n 2.13835e-19 $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_80 A N_X_c_247_n 0.0103401f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_81 N_A_c_61_n N_VGND_c_315_n 3.07485e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_M1000_g N_VGND_c_315_n 0.0031795f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_83 A N_VGND_c_315_n 0.0152693f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_84 N_A_M1000_g N_VGND_c_322_n 0.00441743f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_85 A N_VGND_c_322_n 0.00250701f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_86 N_A_M1000_g N_VGND_c_324_n 0.00701594f $X=0.525 $Y=0.445 $X2=0 $Y2=0
cc_87 A N_VGND_c_324_n 0.00497578f $X=0.655 $Y=0.765 $X2=0 $Y2=0
cc_88 N_A_27_47#_c_127_n N_VPWR_M1003_d 0.00653203f $X=0.995 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_27_47#_c_107_n N_VPWR_c_201_n 0.00695536f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_47#_c_127_n N_VPWR_c_201_n 0.0192006f $X=0.995 $Y=1.58 $X2=0 $Y2=0
cc_91 N_A_27_47#_c_108_n N_VPWR_c_202_n 0.0030005f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_27_47#_c_109_n N_VPWR_c_202_n 0.00169564f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_93 N_A_27_47#_c_109_n N_VPWR_c_203_n 5.61462e-19 $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_27_47#_c_110_n N_VPWR_c_203_n 0.0122616f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_95 N_A_27_47#_c_107_n N_VPWR_c_204_n 0.00702461f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_27_47#_c_108_n N_VPWR_c_204_n 0.00523784f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_27_47#_c_109_n N_VPWR_c_206_n 0.00523784f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_27_47#_c_110_n N_VPWR_c_206_n 0.00642146f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_99 N_A_27_47#_M1003_s N_VPWR_c_200_n 0.00273689f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_100 N_A_27_47#_c_107_n N_VPWR_c_200_n 0.0127458f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_27_47#_c_108_n N_VPWR_c_200_n 0.00689717f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_27_47#_c_109_n N_VPWR_c_200_n 0.00683736f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_27_47#_c_110_n N_VPWR_c_200_n 0.0107337f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_27_47#_c_115_n N_VPWR_c_200_n 0.0118616f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_105 N_A_27_47#_c_115_n N_VPWR_c_210_n 0.0202977f $X=0.26 $Y=1.69 $X2=0 $Y2=0
cc_106 N_A_27_47#_c_127_n N_X_M1004_s 0.00279542f $X=0.995 $Y=1.58 $X2=0 $Y2=0
cc_107 N_A_27_47#_M1001_g N_X_c_245_n 0.00691963f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_108 N_A_27_47#_M1002_g N_X_c_245_n 0.00234073f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_109 N_A_27_47#_c_106_n N_X_c_245_n 4.97219e-19 $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_110 N_A_27_47#_M1002_g N_X_c_246_n 0.0128827f $X=1.49 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_27_47#_c_96_n N_X_c_246_n 0.00345722f $X=1.89 $Y=1.157 $X2=0 $Y2=0
cc_112 N_A_27_47#_M1005_g N_X_c_246_n 0.0130843f $X=1.97 $Y=0.445 $X2=0 $Y2=0
cc_113 N_A_27_47#_c_159_p N_X_c_246_n 0.0487363f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_27_47#_M1001_g N_X_c_247_n 0.00497832f $X=1.005 $Y=0.445 $X2=0 $Y2=0
cc_115 N_A_27_47#_c_101_n N_X_c_247_n 0.00369359f $X=1.41 $Y=1.157 $X2=0 $Y2=0
cc_116 N_A_27_47#_c_131_n N_X_c_247_n 0.0141685f $X=1.215 $Y=1.16 $X2=0 $Y2=0
cc_117 N_A_27_47#_c_159_p N_X_c_247_n 0.0150431f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_118 N_A_27_47#_c_108_n N_X_c_267_n 0.0157325f $X=1.51 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_27_47#_c_96_n N_X_c_267_n 0.00471411f $X=1.89 $Y=1.157 $X2=0 $Y2=0
cc_120 N_A_27_47#_c_109_n N_X_c_267_n 0.0142921f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_27_47#_c_159_p N_X_c_267_n 0.0154613f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_101_n N_X_c_271_n 0.00366589f $X=1.41 $Y=1.157 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_127_n N_X_c_271_n 0.00332702f $X=0.995 $Y=1.58 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_159_p N_X_c_271_n 0.00488011f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_125 N_A_27_47#_M1005_g N_X_c_248_n 0.00493215f $X=1.97 $Y=0.445 $X2=0 $Y2=0
cc_126 N_A_27_47#_M1009_g N_X_c_248_n 0.00212407f $X=2.495 $Y=0.445 $X2=0 $Y2=0
cc_127 N_A_27_47#_M1005_g X 0.00240256f $X=1.97 $Y=0.445 $X2=0 $Y2=0
cc_128 N_A_27_47#_c_98_n X 0.00511421f $X=2.37 $Y=1.157 $X2=0 $Y2=0
cc_129 N_A_27_47#_c_110_n X 5.25855e-19 $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_M1009_g X 0.0168311f $X=2.495 $Y=0.445 $X2=0 $Y2=0
cc_131 N_A_27_47#_c_103_n X 0.0235658f $X=2.47 $Y=1.215 $X2=0 $Y2=0
cc_132 N_A_27_47#_c_159_p X 0.0245385f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_133 N_A_27_47#_c_105_n X 6.77943e-19 $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_27_47#_c_109_n N_X_c_251_n 0.00227075f $X=1.99 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_27_47#_c_98_n N_X_c_251_n 0.00699157f $X=2.37 $Y=1.157 $X2=0 $Y2=0
cc_136 N_A_27_47#_c_110_n N_X_c_251_n 0.0184846f $X=2.47 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_27_47#_c_103_n N_X_c_251_n 6.12827e-19 $X=2.47 $Y=1.215 $X2=0 $Y2=0
cc_138 N_A_27_47#_c_159_p N_X_c_251_n 0.00991119f $X=2.07 $Y=1.16 $X2=0 $Y2=0
cc_139 N_A_27_47#_M1001_g N_VGND_c_315_n 0.00291251f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_140 N_A_27_47#_M1002_g N_VGND_c_316_n 0.00597974f $X=1.49 $Y=0.445 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_M1005_g N_VGND_c_316_n 0.00309457f $X=1.97 $Y=0.445 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_M1009_g N_VGND_c_317_n 0.00481644f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_143 N_A_27_47#_M1001_g N_VGND_c_318_n 0.00544863f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_144 N_A_27_47#_M1002_g N_VGND_c_318_n 0.00439206f $X=1.49 $Y=0.445 $X2=0
+ $Y2=0
cc_145 N_A_27_47#_M1005_g N_VGND_c_320_n 0.00439206f $X=1.97 $Y=0.445 $X2=0
+ $Y2=0
cc_146 N_A_27_47#_M1009_g N_VGND_c_320_n 0.00439071f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_106_n N_VGND_c_322_n 0.0199572f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_148 N_A_27_47#_M1000_s N_VGND_c_324_n 0.00409197f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_149 N_A_27_47#_M1001_g N_VGND_c_324_n 0.0098879f $X=1.005 $Y=0.445 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_M1002_g N_VGND_c_324_n 0.00630094f $X=1.49 $Y=0.445 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1005_g N_VGND_c_324_n 0.00628201f $X=1.97 $Y=0.445 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_M1009_g N_VGND_c_324_n 0.00725365f $X=2.495 $Y=0.445 $X2=0
+ $Y2=0
cc_153 N_A_27_47#_c_106_n N_VGND_c_324_n 0.0113402f $X=0.26 $Y=0.42 $X2=0 $Y2=0
cc_154 N_VPWR_c_200_n N_X_M1004_s 0.00337588f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_155 N_VPWR_c_200_n N_X_M1007_s 0.00302135f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_156 N_VPWR_c_204_n N_X_c_290_n 0.0155613f $X=1.625 $Y=2.72 $X2=0 $Y2=0
cc_157 N_VPWR_c_200_n N_X_c_290_n 0.00991615f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_M1006_d N_X_c_267_n 0.00502677f $X=1.6 $Y=1.485 $X2=0 $Y2=0
cc_159 N_VPWR_c_202_n N_X_c_267_n 0.0145212f $X=1.75 $Y=2.34 $X2=0 $Y2=0
cc_160 N_VPWR_c_204_n N_X_c_267_n 0.00276696f $X=1.625 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_206_n N_X_c_267_n 0.00280673f $X=2.545 $Y=2.72 $X2=0 $Y2=0
cc_162 N_VPWR_c_200_n N_X_c_267_n 0.0108807f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_163 N_VPWR_c_206_n N_X_c_297_n 0.0156343f $X=2.545 $Y=2.72 $X2=0 $Y2=0
cc_164 N_VPWR_c_200_n N_X_c_297_n 0.00993603f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_165 N_VPWR_M1008_d N_X_c_251_n 0.00400241f $X=2.56 $Y=1.485 $X2=0 $Y2=0
cc_166 N_VPWR_c_203_n N_X_c_251_n 0.0202479f $X=2.71 $Y=1.93 $X2=0 $Y2=0
cc_167 N_X_c_246_n N_VGND_c_316_n 0.018338f $X=2.105 $Y=0.82 $X2=0 $Y2=0
cc_168 X N_VGND_c_317_n 0.0227235f $X=2.695 $Y=0.765 $X2=0 $Y2=0
cc_169 N_X_c_245_n N_VGND_c_318_n 0.0132798f $X=1.275 $Y=0.51 $X2=0 $Y2=0
cc_170 N_X_c_246_n N_VGND_c_318_n 0.00299761f $X=2.105 $Y=0.82 $X2=0 $Y2=0
cc_171 N_X_c_246_n N_VGND_c_320_n 0.00307237f $X=2.105 $Y=0.82 $X2=0 $Y2=0
cc_172 N_X_c_248_n N_VGND_c_320_n 0.0112742f $X=2.235 $Y=0.51 $X2=0 $Y2=0
cc_173 X N_VGND_c_320_n 0.00325257f $X=2.695 $Y=0.765 $X2=0 $Y2=0
cc_174 X N_VGND_c_323_n 7.44471e-19 $X=2.695 $Y=0.765 $X2=0 $Y2=0
cc_175 N_X_M1001_d N_VGND_c_324_n 0.00283937f $X=1.08 $Y=0.235 $X2=0 $Y2=0
cc_176 N_X_M1005_d N_VGND_c_324_n 0.00366774f $X=2.045 $Y=0.235 $X2=0 $Y2=0
cc_177 N_X_c_245_n N_VGND_c_324_n 0.0127216f $X=1.275 $Y=0.51 $X2=0 $Y2=0
cc_178 N_X_c_246_n N_VGND_c_324_n 0.0110695f $X=2.105 $Y=0.82 $X2=0 $Y2=0
cc_179 N_X_c_248_n N_VGND_c_324_n 0.00940193f $X=2.235 $Y=0.51 $X2=0 $Y2=0
cc_180 X N_VGND_c_324_n 0.00772618f $X=2.695 $Y=0.765 $X2=0 $Y2=0
