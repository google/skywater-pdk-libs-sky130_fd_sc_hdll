* File: sky130_fd_sc_hdll__o221a_1.spice
* Created: Thu Aug 27 19:20:17 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o221a_1.pex.spice"
.subckt sky130_fd_sc_hdll__o221a_1  VNB VPB C1 B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1010 N_A_124_47#_M1010_d N_C1_M1010_g N_A_27_297#_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.1235 AS=0.169 PD=1.03 PS=1.82 NRD=19.38 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1008 N_A_230_47#_M1008_d N_B1_M1008_g N_A_124_47#_M1010_d VNB NSHORT L=0.15
+ W=0.65 AD=0.095875 AS=0.1235 PD=0.945 PS=1.03 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1000 N_A_124_47#_M1000_d N_B2_M1000_g N_A_230_47#_M1008_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.095875 PD=1.82 PS=0.945 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75001.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_230_47#_M1007_d N_A2_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=8.304 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1002_d N_A1_M1002_g N_A_230_47#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_27_297#_M1006_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2145 AS=0.08775 PD=1.96 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1011 N_VPWR_M1011_d N_C1_M1011_g N_A_27_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.295 PD=1.35 PS=2.59 NRD=4.9053 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1003 A_228_297# N_B1_M1003_g N_VPWR_M1011_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.175 PD=1.23 PS=1.35 NRD=11.8003 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1005 N_A_27_297#_M1005_d N_B2_M1005_g A_228_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.4225 AS=0.115 PD=1.845 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90001.1 SB=90002.2 A=0.18 P=2.36 MULT=1
MM1004 A_515_297# N_A2_M1004_g N_A_27_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.4225 PD=1.23 PS=1.845 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90002.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_515_297# VPB PHIGHVT L=0.18 W=1 AD=0.175
+ AS=0.115 PD=1.35 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90002.6
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1009 N_X_M1009_d N_A_27_297#_M1009_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.175 PD=2.58 PS=1.35 NRD=4.9053 NRS=12.7853 M=1 R=5.55556
+ SA=90003.1 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_16 A2 A2 PROBETYPE=1
pX14_noxref noxref_17 A2 A2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o221a_1.pxi.spice"
*
.ends
*
*
