* File: sky130_fd_sc_hdll__o211ai_1.pex.spice
* Created: Thu Aug 27 19:18:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%A1 1 3 4 6 7
c23 7 0 1.99521e-19 $X=0.23 $Y=1.19
r24 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.16 $X2=0.31 $Y2=1.16
r25 4 10 39.1844 $w=3.78e-07 $l=2.23596e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.387 $Y2=1.16
r26 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.525 $Y=0.995
+ $X2=0.525 $Y2=0.56
r27 1 10 45.167 $w=3.78e-07 $l=3.01247e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.387 $Y2=1.16
r28 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%A2 1 3 4 6 11 14
c36 1 0 1.99521e-19 $X=0.91 $Y=1.41
r37 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.945
+ $Y=1.16 $X2=0.945 $Y2=1.16
r38 8 14 9.61923 $w=2.6e-07 $l=2.05e-07 $layer=LI1_cond $X=0.695 $Y=1.325
+ $X2=0.695 $Y2=1.53
r39 7 11 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.945 $Y2=1.16
r40 7 8 2.13598 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=0.695 $Y=1.16
+ $X2=0.695 $Y2=1.325
r41 4 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=0.945 $Y2=1.16
r42 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.005 $Y=0.995
+ $X2=1.005 $Y2=0.56
r43 1 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.91 $Y=1.41
+ $X2=0.945 $Y2=1.16
r44 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.91 $Y=1.41 $X2=0.91
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%B1 1 3 4 6 7 8
r30 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.505
+ $Y=1.16 $X2=1.505 $Y2=1.16
r31 7 8 14.2055 $w=2.92e-07 $l=3.4e-07 $layer=LI1_cond $X=1.582 $Y=1.19
+ $X2=1.582 $Y2=1.53
r32 7 13 1.25342 $w=2.92e-07 $l=3e-08 $layer=LI1_cond $X=1.582 $Y=1.19 $X2=1.582
+ $Y2=1.16
r33 4 12 48.4451 $w=2.9e-07 $l=2.77038e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.527 $Y2=1.16
r34 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.41 $X2=1.47
+ $Y2=1.985
r35 1 12 38.6157 $w=2.9e-07 $l=2.01879e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.527 $Y2=1.16
r36 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.445 $Y=0.995
+ $X2=1.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%C1 1 3 4 6 7 11
r26 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.105
+ $Y=1.16 $X2=2.105 $Y2=1.16
r27 7 11 12.0114 $w=3.53e-07 $l=3.7e-07 $layer=LI1_cond $X=2.092 $Y=1.53
+ $X2=2.092 $Y2=1.16
r28 4 10 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=1.995 $Y=1.41
+ $X2=2.095 $Y2=1.16
r29 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.995 $Y=1.41
+ $X2=1.995 $Y2=1.985
r30 1 10 38.8967 $w=3.59e-07 $l=2.18746e-07 $layer=POLY_cond $X=1.97 $Y=0.995
+ $X2=2.095 $Y2=1.16
r31 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.97 $Y=0.995 $X2=1.97
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%VPWR 1 2 7 9 15 17 19 26 27 33
r36 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r37 27 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r38 26 27 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 24 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.87 $Y=2.72
+ $X2=1.705 $Y2=2.72
r40 24 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.87 $Y=2.72
+ $X2=2.53 $Y2=2.72
r41 23 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r42 22 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 20 30 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r44 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r45 19 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=1.705 $Y2=2.72
r46 19 22 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=0.69 $Y2=2.72
r47 17 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r48 17 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r49 13 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=2.635
+ $X2=1.705 $Y2=2.72
r50 13 15 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.705 $Y=2.635
+ $X2=1.705 $Y2=2.36
r51 9 12 26.122 $w=2.98e-07 $l=6.8e-07 $layer=LI1_cond $X=0.245 $Y=1.66
+ $X2=0.245 $Y2=2.34
r52 7 30 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.197 $Y2=2.72
r53 7 12 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2.34
r54 2 15 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.485 $X2=1.705 $Y2=2.36
r55 1 12 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r56 1 9 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%Y 1 2 3 12 14 17 21 22 23 27 30
r44 27 30 2.46759 $w=5.7e-07 $l=1.17e-07 $layer=LI1_cond $X=2.557 $Y=0.54
+ $X2=2.44 $Y2=0.54
r45 27 30 0.171228 $w=5.7e-07 $l=8e-09 $layer=LI1_cond $X=2.432 $Y=0.54 $X2=2.44
+ $Y2=0.54
r46 27 32 0.042807 $w=5.7e-07 $l=2e-09 $layer=LI1_cond $X=2.432 $Y=0.54 $X2=2.43
+ $Y2=0.54
r47 22 25 1.79412 $w=5.98e-07 $l=9e-08 $layer=LI1_cond $X=2.375 $Y=1.93
+ $X2=2.375 $Y2=2.02
r48 22 23 6.88405 $w=5.98e-07 $l=1.15e-07 $layer=LI1_cond $X=2.375 $Y=1.93
+ $X2=2.375 $Y2=1.815
r49 19 21 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=1.16 $Y=1.93 $X2=1.16
+ $Y2=2.02
r50 17 19 8.73063 $w=3.28e-07 $l=2.5e-07 $layer=LI1_cond $X=1.16 $Y=1.68
+ $X2=1.16 $Y2=1.93
r51 14 27 6.01081 $w=2.35e-07 $l=2.85e-07 $layer=LI1_cond $X=2.557 $Y=0.825
+ $X2=2.557 $Y2=0.54
r52 14 23 48.5497 $w=2.33e-07 $l=9.9e-07 $layer=LI1_cond $X=2.557 $Y=0.825
+ $X2=2.557 $Y2=1.815
r53 13 19 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=1.93
+ $X2=1.16 $Y2=1.93
r54 12 22 6.41018 $w=2.3e-07 $l=3e-07 $layer=LI1_cond $X=2.075 $Y=1.93 $X2=2.375
+ $Y2=1.93
r55 12 13 37.5797 $w=2.28e-07 $l=7.5e-07 $layer=LI1_cond $X=2.075 $Y=1.93
+ $X2=1.325 $Y2=1.93
r56 3 25 300 $w=1.7e-07 $l=6.90036e-07 $layer=licon1_PDIFF $count=2 $X=2.085
+ $Y=1.485 $X2=2.44 $Y2=2.02
r57 2 21 300 $w=1.7e-07 $l=6.09775e-07 $layer=licon1_PDIFF $count=2 $X=1
+ $Y=1.485 $X2=1.16 $Y2=2.02
r58 2 17 600 $w=1.7e-07 $l=2.63106e-07 $layer=licon1_PDIFF $count=1 $X=1
+ $Y=1.485 $X2=1.16 $Y2=1.68
r59 1 32 91 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_NDIFF $count=2 $X=2.045
+ $Y=0.235 $X2=2.43 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%A_27_47# 1 2 9 11 12 14
r26 14 16 10.3113 $w=3.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.26 $Y=0.38
+ $X2=1.26 $Y2=0.72
r27 11 16 4.20859 $w=2.1e-07 $l=1.9e-07 $layer=LI1_cond $X=1.07 $Y=0.72 $X2=1.26
+ $Y2=0.72
r28 11 12 35.3853 $w=2.08e-07 $l=6.7e-07 $layer=LI1_cond $X=1.07 $Y=0.72 $X2=0.4
+ $Y2=0.72
r29 7 12 7.12258 $w=2.1e-07 $l=1.98681e-07 $layer=LI1_cond $X=0.247 $Y=0.615
+ $X2=0.4 $Y2=0.72
r30 7 9 4.91205 $w=3.03e-07 $l=1.3e-07 $layer=LI1_cond $X=0.247 $Y=0.615
+ $X2=0.247 $Y2=0.485
r31 2 14 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=1.08
+ $Y=0.235 $X2=1.235 $Y2=0.38
r32 1 9 182 $w=1.7e-07 $l=3.06186e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.485
.ends

.subckt PM_SKY130_FD_SC_HDLL__O211AI_1%VGND 1 6 8 10 20 21 24
r32 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r33 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r34 18 21 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r35 18 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r36 17 20 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r37 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r38 15 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=0.735
+ $Y2=0
r39 15 17 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.9 $Y=0 $X2=1.15
+ $Y2=0
r40 10 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.735
+ $Y2=0
r41 10 12 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.57 $Y=0 $X2=0.23
+ $Y2=0
r42 8 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r43 8 12 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r44 4 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0
r45 4 6 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.735 $Y=0.085
+ $X2=0.735 $Y2=0.36
r46 1 6 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.735 $Y2=0.36
.ends

