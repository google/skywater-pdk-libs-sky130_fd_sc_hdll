# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__dlygate4sd1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__dlygate4sd1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.605000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.830000 0.255000 3.120000 0.825000 ;
        RECT 2.860000 1.495000 3.120000 2.465000 ;
        RECT 2.950000 0.825000 3.120000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.600000  0.085000 0.815000 0.545000 ;
        RECT 2.145000  0.085000 2.555000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.600000 2.175000 0.815000 2.635000 ;
        RECT 2.145000 1.915000 2.515000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 1.785000 0.945000 2.005000 ;
      RECT 0.085000 2.005000 0.380000 2.465000 ;
      RECT 0.095000 0.255000 0.380000 0.715000 ;
      RECT 0.095000 0.715000 0.945000 0.885000 ;
      RECT 0.775000 0.885000 0.945000 0.995000 ;
      RECT 0.775000 0.995000 1.080000 1.325000 ;
      RECT 0.775000 1.325000 0.945000 1.785000 ;
      RECT 0.985000 0.255000 1.420000 0.545000 ;
      RECT 0.985000 2.175000 1.420000 2.465000 ;
      RECT 1.250000 0.545000 1.420000 1.075000 ;
      RECT 1.250000 1.075000 2.000000 1.275000 ;
      RECT 1.250000 1.275000 1.420000 2.175000 ;
      RECT 1.615000 0.255000 1.840000 0.735000 ;
      RECT 1.615000 0.735000 2.610000 0.905000 ;
      RECT 1.615000 1.575000 2.610000 1.745000 ;
      RECT 1.615000 1.745000 1.840000 2.430000 ;
      RECT 2.400000 0.905000 2.610000 0.995000 ;
      RECT 2.400000 0.995000 2.730000 1.325000 ;
      RECT 2.400000 1.325000 2.610000 1.575000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__dlygate4sd1_1
