* File: sky130_fd_sc_hdll__and4b_1.pex.spice
* Created: Wed Sep  2 08:23:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%A_N 2 3 5 8 10 11 19
c37 19 0 1.66235e-19 $X=0.52 $Y=1.16
r38 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r39 15 18 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=1.16
+ $X2=0.495 $Y2=1.16
r40 10 11 11.6823 $w=3.63e-07 $l=3.7e-07 $layer=LI1_cond $X=0.267 $Y=1.16
+ $X2=0.267 $Y2=1.53
r41 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r42 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r43 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r44 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r45 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r46 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r47 1 2 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%A_27_47# 1 2 7 8 9 11 12 14 16 19 23 25 26
+ 27 28 30 32 36
c84 27 0 1.66235e-19 $X=0.68 $Y=1.93
r85 37 39 77.4253 $w=2.21e-07 $l=3.55e-07 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.94 $Y2=0.805
r86 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r87 33 36 6.11144 $w=3.28e-07 $l=1.75e-07 $layer=LI1_cond $X=0.765 $Y=1.16
+ $X2=0.94 $Y2=1.16
r88 31 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.16
r89 31 32 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=0.765 $Y=1.325
+ $X2=0.765 $Y2=1.845
r90 30 33 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.765 $Y=0.995
+ $X2=0.765 $Y2=1.16
r91 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.765 $Y=0.825
+ $X2=0.765 $Y2=0.995
r92 27 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=1.93
+ $X2=0.765 $Y2=1.845
r93 27 28 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=1.93
+ $X2=0.345 $Y2=1.93
r94 25 29 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.765 $Y2=0.825
r95 25 26 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.68 $Y=0.74
+ $X2=0.345 $Y2=0.74
r96 21 28 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=2.015
+ $X2=0.345 $Y2=1.93
r97 21 23 18.0623 $w=1.73e-07 $l=2.85e-07 $layer=LI1_cond $X=0.257 $Y=2.015
+ $X2=0.257 $Y2=2.3
r98 17 26 6.81835 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.257 $Y=0.655
+ $X2=0.345 $Y2=0.74
r99 17 19 14.8935 $w=1.73e-07 $l=2.35e-07 $layer=LI1_cond $X=0.257 $Y=0.655
+ $X2=0.257 $Y2=0.42
r100 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.46 $Y=0.73
+ $X2=1.46 $Y2=0.445
r101 13 39 11.8763 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.075 $Y=0.805
+ $X2=0.94 $Y2=0.805
r102 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.385 $Y=0.805
+ $X2=1.46 $Y2=0.73
r103 12 13 158.957 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=1.385 $Y=0.805
+ $X2=1.075 $Y2=0.805
r104 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.975 $Y=1.99
+ $X2=0.975 $Y2=2.275
r105 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.975 $Y=1.89 $X2=0.975
+ $Y2=1.99
r106 7 37 36.5218 $w=2.21e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.94 $Y2=1.16
r107 7 8 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.975 $Y=1.325
+ $X2=0.975 $Y2=1.89
r108 2 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r109 1 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%B 2 3 5 8 10 11 12 13 23
r44 21 23 10.4917 $w=3.3e-07 $l=6e-08 $layer=POLY_cond $X=1.76 $Y=1.3 $X2=1.82
+ $Y2=1.3
r45 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.76
+ $Y=1.3 $X2=1.76 $Y2=1.3
r46 18 21 30.6007 $w=3.3e-07 $l=1.75e-07 $layer=POLY_cond $X=1.585 $Y=1.3
+ $X2=1.76 $Y2=1.3
r47 13 22 5.73121 $w=4.78e-07 $l=2.3e-07 $layer=LI1_cond $X=1.915 $Y=1.53
+ $X2=1.915 $Y2=1.3
r48 12 22 2.74101 $w=4.78e-07 $l=1.1e-07 $layer=LI1_cond $X=1.915 $Y=1.19
+ $X2=1.915 $Y2=1.3
r49 11 12 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.915 $Y=0.85
+ $X2=1.915 $Y2=1.19
r50 10 11 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=1.915 $Y=0.51
+ $X2=1.915 $Y2=0.85
r51 6 23 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.82 $Y=1.135
+ $X2=1.82 $Y2=1.3
r52 6 8 353.809 $w=1.5e-07 $l=6.9e-07 $layer=POLY_cond $X=1.82 $Y=1.135 $X2=1.82
+ $Y2=0.445
r53 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.585 $Y=1.99
+ $X2=1.585 $Y2=2.275
r54 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.585 $Y=1.89 $X2=1.585
+ $Y2=1.99
r55 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.585 $Y=1.465
+ $X2=1.585 $Y2=1.3
r56 1 2 140.92 $w=2e-07 $l=4.25e-07 $layer=POLY_cond $X=1.585 $Y=1.465 $X2=1.585
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%C 2 3 5 8 10 11 12 13 19
r44 19 22 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.16
+ $X2=2.41 $Y2=1.325
r45 19 21 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.41 $Y=1.16
+ $X2=2.41 $Y2=0.995
r46 12 13 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.47 $Y=1.16
+ $X2=2.47 $Y2=1.53
r47 12 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.41
+ $Y=1.16 $X2=2.41 $Y2=1.16
r48 11 12 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.47 $Y=0.85
+ $X2=2.47 $Y2=1.16
r49 10 11 13.5114 $w=2.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.47 $Y=0.51
+ $X2=2.47 $Y2=0.85
r50 8 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.47 $Y=0.445
+ $X2=2.47 $Y2=0.995
r51 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.445 $Y=1.99
+ $X2=2.445 $Y2=2.275
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.445 $Y=1.89 $X2=2.445
+ $Y2=1.99
r53 2 22 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.445 $Y=1.89
+ $X2=2.445 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%D 2 3 5 8 10 11 12 17
c45 17 0 1.60968e-19 $X=2.915 $Y=1.16
r46 17 20 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.915 $Y2=1.325
r47 17 19 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.915 $Y=1.16
+ $X2=2.915 $Y2=0.995
r48 11 12 14.7036 $w=2.88e-07 $l=3.7e-07 $layer=LI1_cond $X=2.93 $Y=1.16
+ $X2=2.93 $Y2=1.53
r49 11 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.915
+ $Y=1.16 $X2=2.915 $Y2=1.16
r50 10 11 12.3192 $w=2.88e-07 $l=3.1e-07 $layer=LI1_cond $X=2.93 $Y=0.85
+ $X2=2.93 $Y2=1.16
r51 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.975 $Y=0.445
+ $X2=2.975 $Y2=0.995
r52 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99 $X2=2.95
+ $Y2=2.275
r53 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r54 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%A_213_413# 1 2 3 10 12 13 15 17 20 22 26
+ 28 31 33 36 37 41
c98 28 0 1.60968e-19 $X=3.245 $Y=1.96
r99 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.45
+ $Y=1.16 $X2=3.45 $Y2=1.16
r100 38 41 4.1907 $w=3.28e-07 $l=1.2e-07 $layer=LI1_cond $X=3.33 $Y=1.16
+ $X2=3.45 $Y2=1.16
r101 33 35 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=1.255 $Y=0.42
+ $X2=1.255 $Y2=0.585
r102 30 38 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.33 $Y=1.325
+ $X2=3.33 $Y2=1.16
r103 30 31 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=3.33 $Y=1.325
+ $X2=3.33 $Y2=1.875
r104 29 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.8 $Y=1.96
+ $X2=2.715 $Y2=1.96
r105 28 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.245 $Y=1.96
+ $X2=3.33 $Y2=1.875
r106 28 29 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=3.245 $Y=1.96
+ $X2=2.8 $Y2=1.96
r107 24 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.715 $Y=2.045
+ $X2=2.715 $Y2=1.96
r108 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.715 $Y=2.045
+ $X2=2.715 $Y2=2.3
r109 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=1.96
+ $X2=1.285 $Y2=1.96
r110 22 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.63 $Y=1.96
+ $X2=2.715 $Y2=1.96
r111 22 23 82.2032 $w=1.68e-07 $l=1.26e-06 $layer=LI1_cond $X=2.63 $Y=1.96
+ $X2=1.37 $Y2=1.96
r112 18 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.045
+ $X2=1.285 $Y2=1.96
r113 18 20 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.285 $Y=2.045
+ $X2=1.285 $Y2=2.3
r114 17 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=1.875
+ $X2=1.285 $Y2=1.96
r115 17 35 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=1.285 $Y=1.875
+ $X2=1.285 $Y2=0.585
r116 13 42 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.45 $Y2=1.16
r117 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.51 $Y=0.995
+ $X2=3.51 $Y2=0.56
r118 10 42 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.45 $Y2=1.16
r119 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.485 $Y=1.41
+ $X2=3.485 $Y2=1.985
r120 3 26 600 $w=1.7e-07 $l=3.1229e-07 $layer=licon1_PDIFF $count=1 $X=2.535
+ $Y=2.065 $X2=2.715 $Y2=2.3
r121 2 20 600 $w=1.7e-07 $l=3.26994e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=2.065 $X2=1.285 $Y2=2.3
r122 1 33 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%VPWR 1 2 3 12 16 19 20 21 23 38 39 42 47
+ 50
r61 49 50 10.0259 $w=5.78e-07 $l=1.65e-07 $layer=LI1_cond $X=2.21 $Y=2.515
+ $X2=2.375 $Y2=2.515
r62 45 49 2.88709 $w=5.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.07 $Y=2.515
+ $X2=2.21 $Y2=2.515
r63 45 47 15.1814 $w=5.78e-07 $l=4.15e-07 $layer=LI1_cond $X=2.07 $Y=2.515
+ $X2=1.655 $Y2=2.515
r64 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r65 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r67 36 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 36 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r69 35 50 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.375 $Y2=2.72
r70 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 32 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r72 32 43 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r73 31 47 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=1.655 $Y2=2.72
r74 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r75 29 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r76 29 31 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 23 42 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r78 23 25 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r79 21 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r80 21 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r81 19 35 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=3.06 $Y=2.72 $X2=2.99
+ $Y2=2.72
r82 19 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.06 $Y=2.72
+ $X2=3.225 $Y2=2.72
r83 18 38 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=3.91 $Y2=2.72
r84 18 20 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.39 $Y=2.72
+ $X2=3.225 $Y2=2.72
r85 14 20 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.225 $Y=2.635
+ $X2=3.225 $Y2=2.72
r86 14 16 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.225 $Y=2.635
+ $X2=3.225 $Y2=2.31
r87 10 42 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r88 10 12 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.34
r89 3 16 600 $w=1.7e-07 $l=3.24577e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.225 $Y2=2.31
r90 2 49 300 $w=1.7e-07 $l=6.45988e-07 $layer=licon1_PDIFF $count=2 $X=1.675
+ $Y=2.065 $X2=2.21 $Y2=2.31
r91 1 12 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%X 1 2 11 12 13 14 15 25
r24 14 15 10.8842 $w=3.58e-07 $l=3.4e-07 $layer=LI1_cond $X=3.815 $Y=1.87
+ $X2=3.815 $Y2=2.21
r25 13 29 9.63763 $w=4.73e-07 $l=2.95e-07 $layer=LI1_cond $X=3.757 $Y=0.51
+ $X2=3.757 $Y2=0.805
r26 13 25 3.27348 $w=4.73e-07 $l=1.3e-07 $layer=LI1_cond $X=3.757 $Y=0.51
+ $X2=3.757 $Y2=0.38
r27 12 29 29.4513 $w=2.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.86 $Y=1.495
+ $X2=3.86 $Y2=0.805
r28 11 12 6.02816 $w=3.58e-07 $l=1.65e-07 $layer=LI1_cond $X=3.815 $Y=1.66
+ $X2=3.815 $Y2=1.495
r29 9 14 6.2424 $w=3.58e-07 $l=1.95e-07 $layer=LI1_cond $X=3.815 $Y=1.675
+ $X2=3.815 $Y2=1.87
r30 9 11 0.480185 $w=3.58e-07 $l=1.5e-08 $layer=LI1_cond $X=3.815 $Y=1.675
+ $X2=3.815 $Y2=1.66
r31 2 11 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=3.575
+ $Y=1.485 $X2=3.72 $Y2=1.66
r32 1 25 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=3.585
+ $Y=0.235 $X2=3.72 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_1%VGND 1 2 7 9 14 21 22 26
r52 26 29 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.705
+ $Y2=0.38
r53 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r54 22 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r55 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r56 19 21 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.91
+ $Y2=0
r57 18 34 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.99
+ $Y2=0
r58 18 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r59 17 18 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r60 15 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r61 15 17 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=1.15
+ $Y2=0
r62 14 36 11.0868 $w=3.93e-07 $l=3.8e-07 $layer=LI1_cond $X=3.152 $Y=0 $X2=3.152
+ $Y2=0.38
r63 14 19 5.70203 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=3.152 $Y=0 $X2=3.35
+ $Y2=0
r64 14 34 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r65 14 17 117.759 $w=1.68e-07 $l=1.805e-06 $layer=LI1_cond $X=2.955 $Y=0
+ $X2=1.15 $Y2=0
r66 9 26 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r67 9 11 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r68 7 27 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r69 7 11 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r70 2 36 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.05
+ $Y=0.235 $X2=3.185 $Y2=0.38
r71 1 29 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

