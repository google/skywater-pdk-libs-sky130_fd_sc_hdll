* File: sky130_fd_sc_hdll__clkinv_4.spice
* Created: Wed Sep  2 08:26:29 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_4.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_4  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1001 N_Y_M1001_d N_A_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.1596 PD=0.75 PS=1.6 NRD=14.28 NRS=0 M=1 R=2.8 SA=75000.3 SB=75001.8
+ A=0.063 P=1.14 MULT=1
MM1002 N_Y_M1001_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=14.28 M=1 R=2.8 SA=75000.8 SB=75001.3
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1006_d N_A_M1006_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.0693 PD=0.75 PS=0.75 NRD=14.28 NRS=0 M=1 R=2.8 SA=75001.3 SB=75000.8
+ A=0.063 P=1.14 MULT=1
MM1008 N_Y_M1006_d N_A_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.42 AD=0.0693
+ AS=0.1869 PD=0.75 PS=1.73 NRD=0 NRS=14.28 M=1 R=2.8 SA=75001.7 SB=75000.4
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.315
+ AS=0.15 PD=2.63 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A_M1003_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1003_d N_A_M1004_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.2
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_M1005_g N_Y_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1005_d N_A_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_M1009_g N_Y_M1007_s VPB PHIGHVT L=0.18 W=1 AD=0.355
+ AS=0.15 PD=2.71 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.6
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_7 A A PROBETYPE=1
pX12_noxref noxref_8 A A PROBETYPE=1
pX13_noxref noxref_9 A A PROBETYPE=1
pX14_noxref noxref_10 A A PROBETYPE=1
*
.include "sky130_fd_sc_hdll__clkinv_4.pxi.spice"
*
.ends
*
*
