* File: sky130_fd_sc_hdll__muxb8to1_4.pex.spice
* Created: Thu Aug 27 19:12:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[0] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c112 30 0 1.3204e-19 $X=2.78 $Y=0.255
r113 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.23 $Y=1.16
+ $X2=0.58 $Y2=1.16
r114 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.62 $Y=0.255
+ $X2=3.62 $Y2=0.59
r115 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.275 $Y=0.18
+ $X2=3.2 $Y2=0.18
r116 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.545 $Y=0.18
+ $X2=3.62 $Y2=0.255
r117 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.545 $Y=0.18
+ $X2=3.275 $Y2=0.18
r118 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.2 $Y=0.255
+ $X2=3.2 $Y2=0.18
r119 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.2 $Y=0.255
+ $X2=3.2 $Y2=0.59
r120 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=0.18
+ $X2=2.78 $Y2=0.18
r121 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.125 $Y=0.18
+ $X2=3.2 $Y2=0.18
r122 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.125 $Y=0.18
+ $X2=2.855 $Y2=0.18
r123 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=0.255
+ $X2=2.78 $Y2=0.18
r124 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.78 $Y=0.255
+ $X2=2.78 $Y2=0.59
r125 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=0.18
+ $X2=2.36 $Y2=0.18
r126 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=0.18
+ $X2=2.78 $Y2=0.18
r127 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.705 $Y=0.18
+ $X2=2.435 $Y2=0.18
r128 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=0.255
+ $X2=2.36 $Y2=0.18
r129 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.36 $Y=0.255
+ $X2=2.36 $Y2=0.59
r130 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=0.18
+ $X2=2.36 $Y2=0.18
r131 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.285 $Y=0.18
+ $X2=1.675 $Y2=0.18
r132 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=0.255
+ $X2=1.675 $Y2=0.18
r133 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.6 $Y=0.255
+ $X2=1.6 $Y2=0.735
r134 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.19 $Y=0.81 $X2=1.09
+ $Y2=0.81
r135 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.525 $Y=0.81
+ $X2=1.6 $Y2=0.735
r136 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.525 $Y=0.81
+ $X2=1.19 $Y2=0.81
r137 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=1.09 $Y=1.55
+ $X2=1.09 $Y2=2.035
r138 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.09 $Y=1.45 $X2=1.09
+ $Y2=1.55
r139 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.09 $Y=0.885
+ $X2=1.09 $Y2=0.81
r140 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.09 $Y=0.885
+ $X2=1.09 $Y2=1.45
r141 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.065 $Y=0.735
+ $X2=1.09 $Y2=0.81
r142 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.065 $Y=0.735
+ $X2=1.065 $Y2=0.445
r143 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.72 $Y=0.81 $X2=0.62
+ $Y2=0.81
r144 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.99 $Y=0.81 $X2=1.09
+ $Y2=0.81
r145 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.99 $Y=0.81
+ $X2=0.72 $Y2=0.81
r146 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.645 $Y=0.735
+ $X2=0.62 $Y2=0.81
r147 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.645 $Y=0.735
+ $X2=0.645 $Y2=0.445
r148 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=0.62 $Y=1.55
+ $X2=0.62 $Y2=2.035
r149 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=0.62 $Y=1.16
+ $X2=0.62 $Y2=1.55
r150 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=1.16 $X2=0.58 $Y2=1.16
r151 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=0.62 $Y=1.16
+ $X2=0.62 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[1] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c118 30 0 1.3204e-19 $X=2.78 $Y=5.185
r119 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=0.23 $Y=4.28
+ $X2=0.58 $Y2=4.28
r120 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.62 $Y=5.185
+ $X2=3.62 $Y2=4.85
r121 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.275 $Y=5.26
+ $X2=3.2 $Y2=5.26
r122 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.545 $Y=5.26
+ $X2=3.62 $Y2=5.185
r123 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.545 $Y=5.26
+ $X2=3.275 $Y2=5.26
r124 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.2 $Y=5.185
+ $X2=3.2 $Y2=5.26
r125 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=3.2 $Y=5.185
+ $X2=3.2 $Y2=4.85
r126 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.855 $Y=5.26
+ $X2=2.78 $Y2=5.26
r127 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.125 $Y=5.26
+ $X2=3.2 $Y2=5.26
r128 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=3.125 $Y=5.26
+ $X2=2.855 $Y2=5.26
r129 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.78 $Y=5.185
+ $X2=2.78 $Y2=5.26
r130 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.78 $Y=5.185
+ $X2=2.78 $Y2=4.85
r131 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.435 $Y=5.26
+ $X2=2.36 $Y2=5.26
r132 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.705 $Y=5.26
+ $X2=2.78 $Y2=5.26
r133 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=2.705 $Y=5.26
+ $X2=2.435 $Y2=5.26
r134 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.36 $Y=5.185
+ $X2=2.36 $Y2=5.26
r135 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.36 $Y=5.185
+ $X2=2.36 $Y2=4.85
r136 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.285 $Y=5.26
+ $X2=2.36 $Y2=5.26
r137 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=2.285 $Y=5.26
+ $X2=1.675 $Y2=5.26
r138 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.6 $Y=5.185
+ $X2=1.675 $Y2=5.26
r139 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=1.6 $Y=4.705
+ $X2=1.6 $Y2=5.185
r140 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.19 $Y=4.63 $X2=1.09
+ $Y2=4.63
r141 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.525 $Y=4.63
+ $X2=1.6 $Y2=4.705
r142 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=1.525 $Y=4.63
+ $X2=1.19 $Y2=4.63
r143 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=1.09 $Y=3.89
+ $X2=1.09 $Y2=3.405
r144 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=1.065 $Y=4.705
+ $X2=1.09 $Y2=4.63
r145 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.065 $Y=4.705
+ $X2=1.065 $Y2=4.995
r146 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.09 $Y=4.555
+ $X2=1.09 $Y2=4.63
r147 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.09 $Y=3.99 $X2=1.09
+ $Y2=3.89
r148 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=1.09 $Y=3.99
+ $X2=1.09 $Y2=4.555
r149 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.72 $Y=4.63 $X2=0.62
+ $Y2=4.63
r150 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.99 $Y=4.63 $X2=1.09
+ $Y2=4.63
r151 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=0.99 $Y=4.63
+ $X2=0.72 $Y2=4.63
r152 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=0.645 $Y=4.705
+ $X2=0.62 $Y2=4.63
r153 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=0.645 $Y=4.705
+ $X2=0.645 $Y2=4.995
r154 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=0.62 $Y=3.89
+ $X2=0.62 $Y2=3.405
r155 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=0.62 $Y=4.28
+ $X2=0.62 $Y2=4.63
r156 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.58
+ $Y=4.28 $X2=0.58 $Y2=4.28
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=0.62 $Y=4.28
+ $X2=0.62 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_325# 1 2 7 9 10 11 12 14 15 17 19
+ 20 22 24 25 26 29 33 36 44 47 48 49 50
c112 22 0 9.37986e-20 $X=3.545 $Y=1.475
c113 20 0 1.74242e-19 $X=3.455 $Y=1.4
c114 17 0 9.37986e-20 $X=3.075 $Y=1.475
c115 12 0 9.37986e-20 $X=2.605 $Y=1.475
c116 7 0 9.37986e-20 $X=2.135 $Y=1.475
r117 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=1.905 $Y=1.285
+ $X2=1.815 $Y2=1.23
r118 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=1.23 $X2=1.905 $Y2=1.23
r119 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=1.565 $Y=1.23
+ $X2=1.815 $Y2=1.23
r120 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.565 $Y=1.23
+ $X2=1.905 $Y2=1.23
r121 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.23 $X2=1.565 $Y2=1.23
r122 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=1.23
+ $X2=0.935 $Y2=1.23
r123 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.02 $Y=1.23
+ $X2=1.565 $Y2=1.23
r124 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.395
+ $X2=0.935 $Y2=1.23
r125 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.935 $Y=1.395
+ $X2=0.935 $Y2=1.605
r126 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=1.065
+ $X2=0.935 $Y2=1.23
r127 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.935 $Y=1.065
+ $X2=0.935 $Y2=0.825
r128 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=0.7
+ $X2=0.895 $Y2=0.825
r129 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0.7
+ $X2=0.895 $Y2=0.445
r130 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=1.77
+ $X2=0.855 $Y2=1.605
r131 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.545 $Y=1.475
+ $X2=3.545 $Y2=1.965
r132 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.165 $Y=1.4
+ $X2=3.075 $Y2=1.4
r133 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.455 $Y=1.4
+ $X2=3.545 $Y2=1.475
r134 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.455 $Y=1.4
+ $X2=3.165 $Y2=1.4
r135 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=1.475
+ $X2=3.075 $Y2=1.4
r136 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.075 $Y=1.475
+ $X2=3.075 $Y2=1.965
r137 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.695 $Y=1.4
+ $X2=2.605 $Y2=1.4
r138 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.985 $Y=1.4
+ $X2=3.075 $Y2=1.4
r139 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.985 $Y=1.4
+ $X2=2.695 $Y2=1.4
r140 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=1.475
+ $X2=2.605 $Y2=1.4
r141 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.605 $Y=1.475
+ $X2=2.605 $Y2=1.965
r142 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.515 $Y=1.4
+ $X2=2.605 $Y2=1.4
r143 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.515 $Y=1.4
+ $X2=2.225 $Y2=1.4
r144 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.135 $Y=1.475
+ $X2=2.225 $Y2=1.4
r145 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=2.135 $Y=1.475
+ $X2=1.905 $Y2=1.285
r146 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.135 $Y=1.475
+ $X2=2.135 $Y2=1.965
r147 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.71
+ $Y=1.625 $X2=0.855 $Y2=1.77
r148 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.72
+ $Y=0.235 $X2=0.855 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_142_599# 1 2 7 9 10 11 12 14 15 17 19
+ 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c118 22 0 9.37986e-20 $X=3.545 $Y=3.965
c119 20 0 1.74242e-19 $X=3.455 $Y=4.04
c120 17 0 9.37986e-20 $X=3.075 $Y=3.965
c121 12 0 9.37986e-20 $X=2.605 $Y=3.965
c122 7 0 9.37986e-20 $X=2.135 $Y=3.965
r123 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=1.905 $Y=4.155
+ $X2=1.815 $Y2=4.21
r124 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.905
+ $Y=4.21 $X2=1.905 $Y2=4.21
r125 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=1.565 $Y=4.21
+ $X2=1.815 $Y2=4.21
r126 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.565 $Y=4.21
+ $X2=1.905 $Y2=4.21
r127 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=4.21 $X2=1.565 $Y2=4.21
r128 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.02 $Y=4.21
+ $X2=0.935 $Y2=4.21
r129 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=1.02 $Y=4.21
+ $X2=1.565 $Y2=4.21
r130 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=4.375
+ $X2=0.935 $Y2=4.21
r131 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=0.935 $Y=4.375
+ $X2=0.935 $Y2=4.615
r132 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.935 $Y=4.045
+ $X2=0.935 $Y2=4.21
r133 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.935 $Y=4.045
+ $X2=0.935 $Y2=3.835
r134 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=4.74
+ $X2=0.895 $Y2=4.615
r135 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=4.74
+ $X2=0.895 $Y2=4.995
r136 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.855 $Y=3.67
+ $X2=0.855 $Y2=3.835
r137 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=0.855 $Y=3.67
+ $X2=0.855 $Y2=3.14
r138 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.545 $Y=3.965
+ $X2=3.545 $Y2=3.475
r139 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=3.165 $Y=4.04
+ $X2=3.075 $Y2=4.04
r140 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=3.455 $Y=4.04
+ $X2=3.545 $Y2=3.965
r141 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=3.455 $Y=4.04
+ $X2=3.165 $Y2=4.04
r142 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=3.075 $Y=3.965
+ $X2=3.075 $Y2=4.04
r143 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=3.075 $Y=3.965
+ $X2=3.075 $Y2=3.475
r144 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.695 $Y=4.04
+ $X2=2.605 $Y2=4.04
r145 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.985 $Y=4.04
+ $X2=3.075 $Y2=4.04
r146 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.985 $Y=4.04
+ $X2=2.695 $Y2=4.04
r147 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=2.605 $Y=3.965
+ $X2=2.605 $Y2=4.04
r148 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.605 $Y=3.965
+ $X2=2.605 $Y2=3.475
r149 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.515 $Y=4.04
+ $X2=2.605 $Y2=4.04
r150 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.515 $Y=4.04
+ $X2=2.225 $Y2=4.04
r151 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.135 $Y=3.965
+ $X2=2.225 $Y2=4.04
r152 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=2.135 $Y=3.965
+ $X2=1.905 $Y2=4.155
r153 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=2.135 $Y=3.965
+ $X2=2.135 $Y2=3.475
r154 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=0.71
+ $Y=2.995 $X2=0.855 $Y2=3.14
r155 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.72
+ $Y=4.785 $X2=0.855 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[0] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
c99 52 0 1.35498e-19 $X=5.84 $Y=1.16
c100 31 0 1.35498e-19 $X=5.945 $Y=1.985
r101 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=1.16
+ $X2=5.945 $Y2=1.16
r102 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=5.84 $Y=1.16 $X2=5.92
+ $Y2=1.16
r103 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.84
+ $Y=1.16 $X2=5.84 $Y2=1.16
r104 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=5.5 $Y=1.16
+ $X2=5.84 $Y2=1.16
r105 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.5 $Y2=1.16
r106 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.98 $Y=1.16
+ $X2=5.005 $Y2=1.16
r107 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=4.82 $Y=1.16
+ $X2=4.98 $Y2=1.16
r108 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=1.16 $X2=4.82 $Y2=1.16
r109 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=4.56 $Y=1.16
+ $X2=4.82 $Y2=1.16
r110 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.535 $Y=1.16
+ $X2=4.56 $Y2=1.16
r111 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.16 $Y=1.19
+ $X2=4.82 $Y2=1.19
r112 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.16
+ $Y=1.16 $X2=5.16 $Y2=1.16
r113 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.095 $Y=1.16
+ $X2=5.005 $Y2=1.16
r114 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=5.095 $Y=1.16
+ $X2=5.16 $Y2=1.16
r115 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.385 $Y=1.16
+ $X2=5.475 $Y2=1.16
r116 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=5.385 $Y=1.16
+ $X2=5.16 $Y2=1.16
r117 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.75 $Y=1.19 $X2=5.84
+ $Y2=1.19
r118 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.75 $Y=1.19
+ $X2=5.16 $Y2=1.19
r119 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.16
r120 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.985
r121 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=1.16
r122 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=0.56
r123 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=1.025
+ $X2=5.5 $Y2=1.16
r124 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=1.025
+ $X2=5.5 $Y2=0.56
r125 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.16
r126 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.985
r127 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.005 $Y=1.295
+ $X2=5.005 $Y2=1.16
r128 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.005 $Y=1.295
+ $X2=5.005 $Y2=1.985
r129 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=1.025
+ $X2=4.98 $Y2=1.16
r130 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.98 $Y=1.025
+ $X2=4.98 $Y2=0.56
r131 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.56 $Y=1.025
+ $X2=4.56 $Y2=1.16
r132 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.56 $Y=1.025
+ $X2=4.56 $Y2=0.56
r133 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.535 $Y=1.295
+ $X2=4.535 $Y2=1.16
r134 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=4.535 $Y=1.295
+ $X2=4.535 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[1] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
c97 52 0 1.35498e-19 $X=5.84 $Y=4.28
c98 31 0 1.35498e-19 $X=5.945 $Y=3.455
r99 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=4.28
+ $X2=5.945 $Y2=4.28
r100 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=5.84 $Y=4.28 $X2=5.92
+ $Y2=4.28
r101 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.84
+ $Y=4.28 $X2=5.84 $Y2=4.28
r102 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=5.5 $Y=4.28
+ $X2=5.84 $Y2=4.28
r103 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=4.28
+ $X2=5.5 $Y2=4.28
r104 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.98 $Y=4.28
+ $X2=5.005 $Y2=4.28
r105 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=4.82 $Y=4.28
+ $X2=4.98 $Y2=4.28
r106 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.82
+ $Y=4.28 $X2=4.82 $Y2=4.28
r107 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=4.56 $Y=4.28
+ $X2=4.82 $Y2=4.28
r108 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=4.535 $Y=4.28
+ $X2=4.56 $Y2=4.28
r109 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.16 $Y=4.25
+ $X2=4.82 $Y2=4.25
r110 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.16
+ $Y=4.28 $X2=5.16 $Y2=4.28
r111 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.095 $Y=4.28
+ $X2=5.005 $Y2=4.28
r112 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=5.095 $Y=4.28
+ $X2=5.16 $Y2=4.28
r113 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=5.385 $Y=4.28
+ $X2=5.475 $Y2=4.28
r114 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=5.385 $Y=4.28
+ $X2=5.16 $Y2=4.28
r115 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=5.75 $Y=4.25 $X2=5.84
+ $Y2=4.25
r116 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=5.75 $Y=4.25
+ $X2=5.16 $Y2=4.25
r117 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=4.145
+ $X2=5.945 $Y2=4.28
r118 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=4.145
+ $X2=5.945 $Y2=3.455
r119 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=4.415
+ $X2=5.92 $Y2=4.28
r120 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=4.415
+ $X2=5.92 $Y2=4.88
r121 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=4.415
+ $X2=5.5 $Y2=4.28
r122 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=4.415
+ $X2=5.5 $Y2=4.88
r123 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=4.145
+ $X2=5.475 $Y2=4.28
r124 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=4.145
+ $X2=5.475 $Y2=3.455
r125 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.005 $Y=4.145
+ $X2=5.005 $Y2=4.28
r126 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.005 $Y=4.145
+ $X2=5.005 $Y2=3.455
r127 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.98 $Y=4.415
+ $X2=4.98 $Y2=4.28
r128 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.98 $Y=4.415
+ $X2=4.98 $Y2=4.88
r129 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.56 $Y=4.415
+ $X2=4.56 $Y2=4.28
r130 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.56 $Y=4.415
+ $X2=4.56 $Y2=4.88
r131 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.535 $Y=4.145
+ $X2=4.535 $Y2=4.28
r132 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=4.535 $Y=4.145
+ $X2=4.535 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[2] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
c101 51 0 1.35498e-19 $X=7.6 $Y=1.16
c102 3 0 1.35498e-19 $X=6.475 $Y=1.985
r103 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.86 $Y=1.16
+ $X2=7.885 $Y2=1.16
r104 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=7.6 $Y=1.16
+ $X2=7.86 $Y2=1.16
r105 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=1.16 $X2=7.6 $Y2=1.16
r106 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=7.44 $Y=1.16
+ $X2=7.6 $Y2=1.16
r107 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.415 $Y=1.16
+ $X2=7.44 $Y2=1.16
r108 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.92 $Y=1.16
+ $X2=6.945 $Y2=1.16
r109 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.92
+ $Y=1.16 $X2=6.92 $Y2=1.16
r110 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.5 $Y=1.16 $X2=6.92
+ $Y2=1.16
r111 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.475 $Y=1.16
+ $X2=6.5 $Y2=1.16
r112 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.26 $Y=1.19
+ $X2=7.6 $Y2=1.19
r113 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.26 $Y=1.19
+ $X2=6.92 $Y2=1.19
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=1.16 $X2=7.26 $Y2=1.16
r115 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.035 $Y=1.16
+ $X2=6.945 $Y2=1.16
r116 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=7.035 $Y=1.16
+ $X2=7.26 $Y2=1.16
r117 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.325 $Y=1.16
+ $X2=7.415 $Y2=1.16
r118 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=7.325 $Y=1.16
+ $X2=7.26 $Y2=1.16
r119 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.67 $Y=1.19
+ $X2=6.92 $Y2=1.19
r120 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.885 $Y=1.295
+ $X2=7.885 $Y2=1.16
r121 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.885 $Y=1.295
+ $X2=7.885 $Y2=1.985
r122 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.86 $Y=1.025
+ $X2=7.86 $Y2=1.16
r123 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.86 $Y=1.025
+ $X2=7.86 $Y2=0.56
r124 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.44 $Y=1.025
+ $X2=7.44 $Y2=1.16
r125 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.44 $Y=1.025
+ $X2=7.44 $Y2=0.56
r126 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.415 $Y=1.295
+ $X2=7.415 $Y2=1.16
r127 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.415 $Y=1.295
+ $X2=7.415 $Y2=1.985
r128 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.945 $Y=1.295
+ $X2=6.945 $Y2=1.16
r129 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.945 $Y=1.295
+ $X2=6.945 $Y2=1.985
r130 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.92 $Y=1.025
+ $X2=6.92 $Y2=1.16
r131 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.92 $Y=1.025
+ $X2=6.92 $Y2=0.56
r132 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.5 $Y=1.025
+ $X2=6.5 $Y2=1.16
r133 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.5 $Y=1.025 $X2=6.5
+ $Y2=0.56
r134 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.475 $Y=1.295
+ $X2=6.475 $Y2=1.16
r135 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.475 $Y=1.295
+ $X2=6.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[3] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
c97 51 0 1.35498e-19 $X=7.6 $Y=4.28
c98 3 0 1.35498e-19 $X=6.475 $Y=3.455
r99 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.86 $Y=4.28
+ $X2=7.885 $Y2=4.28
r100 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=7.6 $Y=4.28
+ $X2=7.86 $Y2=4.28
r101 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.6
+ $Y=4.28 $X2=7.6 $Y2=4.28
r102 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=7.44 $Y=4.28
+ $X2=7.6 $Y2=4.28
r103 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.415 $Y=4.28
+ $X2=7.44 $Y2=4.28
r104 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.92 $Y=4.28
+ $X2=6.945 $Y2=4.28
r105 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.92
+ $Y=4.28 $X2=6.92 $Y2=4.28
r106 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=6.5 $Y=4.28 $X2=6.92
+ $Y2=4.28
r107 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.475 $Y=4.28
+ $X2=6.5 $Y2=4.28
r108 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.26 $Y=4.25
+ $X2=7.6 $Y2=4.25
r109 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=7.26 $Y=4.25
+ $X2=6.92 $Y2=4.25
r110 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.26
+ $Y=4.28 $X2=7.26 $Y2=4.28
r111 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.035 $Y=4.28
+ $X2=6.945 $Y2=4.28
r112 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=7.035 $Y=4.28
+ $X2=7.26 $Y2=4.28
r113 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=7.325 $Y=4.28
+ $X2=7.415 $Y2=4.28
r114 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=7.325 $Y=4.28
+ $X2=7.26 $Y2=4.28
r115 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=6.67 $Y=4.25
+ $X2=6.92 $Y2=4.25
r116 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.885 $Y=4.145
+ $X2=7.885 $Y2=4.28
r117 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.885 $Y=4.145
+ $X2=7.885 $Y2=3.455
r118 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.86 $Y=4.415
+ $X2=7.86 $Y2=4.28
r119 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.86 $Y=4.415
+ $X2=7.86 $Y2=4.88
r120 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.44 $Y=4.415
+ $X2=7.44 $Y2=4.28
r121 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.44 $Y=4.415
+ $X2=7.44 $Y2=4.88
r122 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.415 $Y=4.145
+ $X2=7.415 $Y2=4.28
r123 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.415 $Y=4.145
+ $X2=7.415 $Y2=3.455
r124 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.945 $Y=4.145
+ $X2=6.945 $Y2=4.28
r125 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.945 $Y=4.145
+ $X2=6.945 $Y2=3.455
r126 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.92 $Y=4.415
+ $X2=6.92 $Y2=4.28
r127 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.92 $Y=4.415
+ $X2=6.92 $Y2=4.88
r128 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.5 $Y=4.415
+ $X2=6.5 $Y2=4.28
r129 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.5 $Y=4.415 $X2=6.5
+ $Y2=4.88
r130 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.475 $Y=4.145
+ $X2=6.475 $Y2=4.28
r131 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.475 $Y=4.145
+ $X2=6.475 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c119 22 0 9.37986e-20 $X=10.285 $Y=1.475
c120 20 0 1.10627e-19 $X=10.195 $Y=1.4
c121 17 0 9.37986e-20 $X=9.815 $Y=1.475
c122 12 0 9.37986e-20 $X=9.345 $Y=1.475
c123 11 0 1.74242e-19 $X=8.965 $Y=1.4
c124 7 0 9.37986e-20 $X=8.875 $Y=1.475
r125 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.565 $Y=1.77
+ $X2=11.565 $Y2=1.605
r126 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.485 $Y=1.395
+ $X2=11.485 $Y2=1.23
r127 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.485 $Y=1.395
+ $X2=11.485 $Y2=1.605
r128 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.485 $Y=1.065
+ $X2=11.485 $Y2=1.23
r129 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.485 $Y=1.065
+ $X2=11.485 $Y2=0.825
r130 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.525 $Y=0.7
+ $X2=11.525 $Y2=0.825
r131 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.525 $Y=0.7
+ $X2=11.525 $Y2=0.445
r132 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=10.855 $Y=1.23
+ $X2=10.605 $Y2=1.23
r133 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.855
+ $Y=1.23 $X2=10.855 $Y2=1.23
r134 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=10.515
+ $Y=1.285 $X2=10.605 $Y2=1.23
r135 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.515 $Y=1.23
+ $X2=10.855 $Y2=1.23
r136 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.515
+ $Y=1.23 $X2=10.515 $Y2=1.23
r137 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.4 $Y=1.23
+ $X2=11.485 $Y2=1.23
r138 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=11.4 $Y=1.23
+ $X2=10.855 $Y2=1.23
r139 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=10.285
+ $Y=1.475 $X2=10.515 $Y2=1.285
r140 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=10.285 $Y=1.475
+ $X2=10.285 $Y2=1.965
r141 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.905 $Y=1.4
+ $X2=9.815 $Y2=1.4
r142 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.195 $Y=1.4
+ $X2=10.285 $Y2=1.475
r143 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.195 $Y=1.4
+ $X2=9.905 $Y2=1.4
r144 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.815 $Y=1.475
+ $X2=9.815 $Y2=1.4
r145 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.815 $Y=1.475
+ $X2=9.815 $Y2=1.965
r146 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.435 $Y=1.4
+ $X2=9.345 $Y2=1.4
r147 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.725 $Y=1.4
+ $X2=9.815 $Y2=1.4
r148 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.725 $Y=1.4
+ $X2=9.435 $Y2=1.4
r149 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.345 $Y=1.475
+ $X2=9.345 $Y2=1.4
r150 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.345 $Y=1.475
+ $X2=9.345 $Y2=1.965
r151 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.255 $Y=1.4
+ $X2=9.345 $Y2=1.4
r152 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.255 $Y=1.4
+ $X2=8.965 $Y2=1.4
r153 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.875 $Y=1.475
+ $X2=8.965 $Y2=1.4
r154 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=8.875 $Y=1.475
+ $X2=8.875 $Y2=1.965
r155 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.42
+ $Y=1.625 $X2=11.565 $Y2=1.77
r156 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=11.43
+ $Y=0.235 $X2=11.565 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1755_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c125 22 0 9.37986e-20 $X=10.285 $Y=3.965
c126 20 0 1.10627e-19 $X=10.195 $Y=4.04
c127 17 0 9.37986e-20 $X=9.815 $Y=3.965
c128 12 0 9.37986e-20 $X=9.345 $Y=3.965
c129 11 0 1.74242e-19 $X=8.965 $Y=4.04
c130 7 0 9.37986e-20 $X=8.875 $Y=3.965
r131 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=11.525 $Y=4.74
+ $X2=11.525 $Y2=4.615
r132 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=11.525 $Y=4.74
+ $X2=11.525 $Y2=4.995
r133 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.485 $Y=4.375
+ $X2=11.485 $Y2=4.21
r134 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=11.485 $Y=4.375
+ $X2=11.485 $Y2=4.615
r135 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=11.485 $Y=4.045
+ $X2=11.485 $Y2=4.21
r136 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=11.485 $Y=4.045
+ $X2=11.485 $Y2=3.835
r137 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=11.565 $Y=3.67
+ $X2=11.565 $Y2=3.835
r138 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=11.565 $Y=3.67
+ $X2=11.565 $Y2=3.14
r139 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=10.855 $Y=4.21
+ $X2=10.605 $Y2=4.21
r140 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.855
+ $Y=4.21 $X2=10.855 $Y2=4.21
r141 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=10.515
+ $Y=4.155 $X2=10.605 $Y2=4.21
r142 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=10.515 $Y=4.21
+ $X2=10.855 $Y2=4.21
r143 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.515
+ $Y=4.21 $X2=10.515 $Y2=4.21
r144 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=11.4 $Y=4.21
+ $X2=11.485 $Y2=4.21
r145 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=11.4 $Y=4.21
+ $X2=10.855 $Y2=4.21
r146 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=10.285
+ $Y=3.965 $X2=10.515 $Y2=4.155
r147 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=10.285 $Y=3.965
+ $X2=10.285 $Y2=3.475
r148 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.905 $Y=4.04
+ $X2=9.815 $Y2=4.04
r149 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=10.195 $Y=4.04
+ $X2=10.285 $Y2=3.965
r150 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=10.195 $Y=4.04
+ $X2=9.905 $Y2=4.04
r151 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.815 $Y=3.965
+ $X2=9.815 $Y2=4.04
r152 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.815 $Y=3.965
+ $X2=9.815 $Y2=3.475
r153 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.435 $Y=4.04
+ $X2=9.345 $Y2=4.04
r154 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.725 $Y=4.04
+ $X2=9.815 $Y2=4.04
r155 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.725 $Y=4.04
+ $X2=9.435 $Y2=4.04
r156 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=9.345 $Y=3.965
+ $X2=9.345 $Y2=4.04
r157 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=9.345 $Y=3.965
+ $X2=9.345 $Y2=3.475
r158 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=9.255 $Y=4.04
+ $X2=9.345 $Y2=4.04
r159 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=9.255 $Y=4.04
+ $X2=8.965 $Y2=4.04
r160 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=8.875 $Y=3.965
+ $X2=8.965 $Y2=4.04
r161 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=8.875 $Y=3.965
+ $X2=8.875 $Y2=3.475
r162 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.42
+ $Y=2.995 $X2=11.565 $Y2=3.14
r163 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=11.43
+ $Y=4.785 $X2=11.565 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[2] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c117 11 0 1.3204e-19 $X=9.64 $Y=0.255
r118 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.18
+ $Y=1.16 $X2=12.18 $Y2=1.16
r119 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=11.8 $Y=1.55
+ $X2=12.007 $Y2=1.16
r120 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=11.8 $Y=1.55
+ $X2=11.8 $Y2=2.035
r121 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.775 $Y=0.735
+ $X2=11.775 $Y2=0.445
r122 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=11.43 $Y=0.81
+ $X2=11.33 $Y2=0.81
r123 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=11.7 $Y=0.81
+ $X2=12.007 $Y2=1.16
r124 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.7 $Y=0.81
+ $X2=11.775 $Y2=0.735
r125 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.7 $Y=0.81
+ $X2=11.43 $Y2=0.81
r126 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=11.355 $Y=0.735
+ $X2=11.33 $Y2=0.81
r127 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.355 $Y=0.735
+ $X2=11.355 $Y2=0.445
r128 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=11.33 $Y=1.55
+ $X2=11.33 $Y2=2.035
r129 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=11.33 $Y=1.45 $X2=11.33
+ $Y2=1.55
r130 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=11.33 $Y=0.885
+ $X2=11.33 $Y2=0.81
r131 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=11.33 $Y=0.885
+ $X2=11.33 $Y2=1.45
r132 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=11.23 $Y=0.81
+ $X2=11.33 $Y2=0.81
r133 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.23 $Y=0.81
+ $X2=10.895 $Y2=0.81
r134 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.82 $Y=0.735
+ $X2=10.895 $Y2=0.81
r135 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.82 $Y=0.255
+ $X2=10.82 $Y2=0.735
r136 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.135 $Y=0.18
+ $X2=10.06 $Y2=0.18
r137 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.745 $Y=0.18
+ $X2=10.82 $Y2=0.255
r138 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.745 $Y=0.18
+ $X2=10.135 $Y2=0.18
r139 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.06 $Y=0.255
+ $X2=10.06 $Y2=0.18
r140 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.06 $Y=0.255
+ $X2=10.06 $Y2=0.59
r141 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.715 $Y=0.18
+ $X2=9.64 $Y2=0.18
r142 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=10.06 $Y2=0.18
r143 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.985 $Y=0.18
+ $X2=9.715 $Y2=0.18
r144 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.18
r145 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.64 $Y=0.255
+ $X2=9.64 $Y2=0.59
r146 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.295 $Y=0.18
+ $X2=9.22 $Y2=0.18
r147 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.64 $Y2=0.18
r148 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.565 $Y=0.18
+ $X2=9.295 $Y2=0.18
r149 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.18
r150 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.22 $Y=0.255
+ $X2=9.22 $Y2=0.59
r151 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=9.22 $Y2=0.18
r152 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.145 $Y=0.18
+ $X2=8.875 $Y2=0.18
r153 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.8 $Y=0.255
+ $X2=8.875 $Y2=0.18
r154 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.8 $Y=0.255 $X2=8.8
+ $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[3] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c125 11 0 1.3204e-19 $X=9.64 $Y=5.185
r126 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=12.18
+ $Y=4.28 $X2=12.18 $Y2=4.28
r127 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=11.8 $Y=3.89
+ $X2=12.007 $Y2=4.28
r128 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=11.8 $Y=3.89
+ $X2=11.8 $Y2=3.405
r129 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.775 $Y=4.705
+ $X2=11.775 $Y2=4.995
r130 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=11.43 $Y=4.63
+ $X2=11.33 $Y2=4.63
r131 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.7 $Y=4.63
+ $X2=11.775 $Y2=4.705
r132 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=11.7 $Y=4.63
+ $X2=12.007 $Y2=4.28
r133 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.7 $Y=4.63
+ $X2=11.43 $Y2=4.63
r134 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=11.355 $Y=4.705
+ $X2=11.33 $Y2=4.63
r135 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.355 $Y=4.705
+ $X2=11.355 $Y2=4.995
r136 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=11.33 $Y=3.89
+ $X2=11.33 $Y2=3.405
r137 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=11.33 $Y=4.555
+ $X2=11.33 $Y2=4.63
r138 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=11.33 $Y=3.99 $X2=11.33
+ $Y2=3.89
r139 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=11.33 $Y=3.99
+ $X2=11.33 $Y2=4.555
r140 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=11.23 $Y=4.63
+ $X2=11.33 $Y2=4.63
r141 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=11.23 $Y=4.63
+ $X2=10.895 $Y2=4.63
r142 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.82 $Y=4.705
+ $X2=10.895 $Y2=4.63
r143 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=10.82 $Y=4.705
+ $X2=10.82 $Y2=5.185
r144 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.135 $Y=5.26
+ $X2=10.06 $Y2=5.26
r145 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.745 $Y=5.26
+ $X2=10.82 $Y2=5.185
r146 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=10.745 $Y=5.26
+ $X2=10.135 $Y2=5.26
r147 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.06 $Y=5.185
+ $X2=10.06 $Y2=5.26
r148 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.06 $Y=5.185
+ $X2=10.06 $Y2=4.85
r149 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.715 $Y=5.26
+ $X2=9.64 $Y2=5.26
r150 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.985 $Y=5.26
+ $X2=10.06 $Y2=5.26
r151 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.985 $Y=5.26
+ $X2=9.715 $Y2=5.26
r152 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.64 $Y=5.185
+ $X2=9.64 $Y2=5.26
r153 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.64 $Y=5.185
+ $X2=9.64 $Y2=4.85
r154 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.295 $Y=5.26
+ $X2=9.22 $Y2=5.26
r155 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.565 $Y=5.26
+ $X2=9.64 $Y2=5.26
r156 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.565 $Y=5.26
+ $X2=9.295 $Y2=5.26
r157 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.22 $Y=5.185
+ $X2=9.22 $Y2=5.26
r158 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=9.22 $Y=5.185
+ $X2=9.22 $Y2=4.85
r159 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=9.145 $Y=5.26
+ $X2=9.22 $Y2=5.26
r160 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=9.145 $Y=5.26
+ $X2=8.875 $Y2=5.26
r161 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.8 $Y=5.185
+ $X2=8.875 $Y2=5.26
r162 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.8 $Y=5.185 $X2=8.8
+ $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[4] 1 3 5 6 8 9 11 13 15 16 18 19 22
+ 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 52
c120 30 0 1.3204e-19 $X=15.2 $Y=0.255
r121 47 52 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.65 $Y=1.16
+ $X2=13 $Y2=1.16
r122 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.04 $Y=0.255
+ $X2=16.04 $Y2=0.59
r123 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.695 $Y=0.18
+ $X2=15.62 $Y2=0.18
r124 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.965 $Y=0.18
+ $X2=16.04 $Y2=0.255
r125 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.965 $Y=0.18
+ $X2=15.695 $Y2=0.18
r126 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.62 $Y=0.255
+ $X2=15.62 $Y2=0.18
r127 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.62 $Y=0.255
+ $X2=15.62 $Y2=0.59
r128 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.275 $Y=0.18
+ $X2=15.2 $Y2=0.18
r129 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.545 $Y=0.18
+ $X2=15.62 $Y2=0.18
r130 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.545 $Y=0.18
+ $X2=15.275 $Y2=0.18
r131 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.2 $Y=0.255
+ $X2=15.2 $Y2=0.18
r132 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.2 $Y=0.255
+ $X2=15.2 $Y2=0.59
r133 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.855 $Y=0.18
+ $X2=14.78 $Y2=0.18
r134 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.125 $Y=0.18
+ $X2=15.2 $Y2=0.18
r135 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.125 $Y=0.18
+ $X2=14.855 $Y2=0.18
r136 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.78 $Y=0.255
+ $X2=14.78 $Y2=0.18
r137 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=14.78 $Y=0.255
+ $X2=14.78 $Y2=0.59
r138 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.705 $Y=0.18
+ $X2=14.78 $Y2=0.18
r139 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=14.705 $Y=0.18
+ $X2=14.095 $Y2=0.18
r140 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.02 $Y=0.255
+ $X2=14.095 $Y2=0.18
r141 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.02 $Y=0.255
+ $X2=14.02 $Y2=0.735
r142 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.61 $Y=0.81
+ $X2=13.51 $Y2=0.81
r143 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.945 $Y=0.81
+ $X2=14.02 $Y2=0.735
r144 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=13.945 $Y=0.81
+ $X2=13.61 $Y2=0.81
r145 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=13.51 $Y=1.55
+ $X2=13.51 $Y2=2.035
r146 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=13.51 $Y=1.45 $X2=13.51
+ $Y2=1.55
r147 14 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=13.51 $Y=0.885
+ $X2=13.51 $Y2=0.81
r148 14 15 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=13.51 $Y=0.885
+ $X2=13.51 $Y2=1.45
r149 11 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=13.485 $Y=0.735
+ $X2=13.51 $Y2=0.81
r150 11 13 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=13.485 $Y=0.735
+ $X2=13.485 $Y2=0.445
r151 10 49 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.14 $Y=0.81
+ $X2=13.04 $Y2=0.81
r152 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.41 $Y=0.81
+ $X2=13.51 $Y2=0.81
r153 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.41 $Y=0.81
+ $X2=13.14 $Y2=0.81
r154 6 49 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=13.065 $Y=0.735
+ $X2=13.04 $Y2=0.81
r155 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=13.065 $Y=0.735
+ $X2=13.065 $Y2=0.445
r156 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=13.04 $Y=1.55
+ $X2=13.04 $Y2=2.035
r157 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=13.04 $Y=1.16
+ $X2=13.04 $Y2=1.55
r158 1 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13 $Y=1.16
+ $X2=13 $Y2=1.16
r159 1 49 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=13.04 $Y=1.16
+ $X2=13.04 $Y2=0.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[5] 1 3 5 6 8 9 11 12 13 15 16 18 19
+ 22 23 24 25 27 28 30 32 33 35 37 38 40 42 43 44 45 46 47 51
c128 30 0 1.3204e-19 $X=15.2 $Y=5.185
r129 47 51 12.2229 $w=3.28e-07 $l=3.5e-07 $layer=LI1_cond $X=12.65 $Y=4.28
+ $X2=13 $Y2=4.28
r130 40 42 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=16.04 $Y=5.185
+ $X2=16.04 $Y2=4.85
r131 39 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.695 $Y=5.26
+ $X2=15.62 $Y2=5.26
r132 38 40 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.965 $Y=5.26
+ $X2=16.04 $Y2=5.185
r133 38 39 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.965 $Y=5.26
+ $X2=15.695 $Y2=5.26
r134 35 46 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.62 $Y=5.185
+ $X2=15.62 $Y2=5.26
r135 35 37 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.62 $Y=5.185
+ $X2=15.62 $Y2=4.85
r136 34 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.275 $Y=5.26
+ $X2=15.2 $Y2=5.26
r137 33 46 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.545 $Y=5.26
+ $X2=15.62 $Y2=5.26
r138 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.545 $Y=5.26
+ $X2=15.275 $Y2=5.26
r139 30 45 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.2 $Y=5.185
+ $X2=15.2 $Y2=5.26
r140 30 32 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.2 $Y=5.185
+ $X2=15.2 $Y2=4.85
r141 29 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.855 $Y=5.26
+ $X2=14.78 $Y2=5.26
r142 28 45 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=15.125 $Y=5.26
+ $X2=15.2 $Y2=5.26
r143 28 29 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=15.125 $Y=5.26
+ $X2=14.855 $Y2=5.26
r144 25 44 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.78 $Y=5.185
+ $X2=14.78 $Y2=5.26
r145 25 27 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=14.78 $Y=5.185
+ $X2=14.78 $Y2=4.85
r146 23 44 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.705 $Y=5.26
+ $X2=14.78 $Y2=5.26
r147 23 24 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=14.705 $Y=5.26
+ $X2=14.095 $Y2=5.26
r148 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.02 $Y=5.185
+ $X2=14.095 $Y2=5.26
r149 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=14.02 $Y=4.705
+ $X2=14.02 $Y2=5.185
r150 20 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.61 $Y=4.63
+ $X2=13.51 $Y2=4.63
r151 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=13.945 $Y=4.63
+ $X2=14.02 $Y2=4.705
r152 19 20 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=13.945 $Y=4.63
+ $X2=13.61 $Y2=4.63
r153 16 18 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=13.51 $Y=3.89
+ $X2=13.51 $Y2=3.405
r154 13 43 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=13.485 $Y=4.705
+ $X2=13.51 $Y2=4.63
r155 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=13.485 $Y=4.705
+ $X2=13.485 $Y2=4.995
r156 12 43 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=13.51 $Y=4.555
+ $X2=13.51 $Y2=4.63
r157 11 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=13.51 $Y=3.99 $X2=13.51
+ $Y2=3.89
r158 11 12 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=13.51 $Y=3.99
+ $X2=13.51 $Y2=4.555
r159 10 52 7.64856 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.14 $Y=4.63
+ $X2=13.04 $Y2=4.63
r160 9 43 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=13.41 $Y=4.63
+ $X2=13.51 $Y2=4.63
r161 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=13.41 $Y=4.63
+ $X2=13.14 $Y2=4.63
r162 6 52 21.4346 $w=1.84e-07 $l=8.66025e-08 $layer=POLY_cond $X=13.065 $Y=4.705
+ $X2=13.04 $Y2=4.63
r163 6 8 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=13.065 $Y=4.705
+ $X2=13.065 $Y2=4.995
r164 3 5 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=13.04 $Y=3.89
+ $X2=13.04 $Y2=3.405
r165 1 52 91.6848 $w=1.84e-07 $l=3.5e-07 $layer=POLY_cond $X=13.04 $Y=4.28
+ $X2=13.04 $Y2=4.63
r166 1 51 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=13 $Y=4.28
+ $X2=13 $Y2=4.28
r167 1 3 102.163 $w=1.84e-07 $l=3.9e-07 $layer=POLY_cond $X=13.04 $Y=4.28
+ $X2=13.04 $Y2=3.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_325# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 33 36 44 47 48 49 50
c116 22 0 9.37986e-20 $X=15.965 $Y=1.475
c117 20 0 1.74242e-19 $X=15.875 $Y=1.4
c118 17 0 9.37986e-20 $X=15.495 $Y=1.475
c119 12 0 9.37986e-20 $X=15.025 $Y=1.475
c120 7 0 9.37986e-20 $X=14.555 $Y=1.475
r121 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=14.325
+ $Y=1.285 $X2=14.235 $Y2=1.23
r122 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.325
+ $Y=1.23 $X2=14.325 $Y2=1.23
r123 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=13.985 $Y=1.23
+ $X2=14.235 $Y2=1.23
r124 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=13.985 $Y=1.23
+ $X2=14.325 $Y2=1.23
r125 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.985
+ $Y=1.23 $X2=13.985 $Y2=1.23
r126 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.44 $Y=1.23
+ $X2=13.355 $Y2=1.23
r127 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=13.44 $Y=1.23
+ $X2=13.985 $Y2=1.23
r128 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.355 $Y=1.395
+ $X2=13.355 $Y2=1.23
r129 37 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=13.355 $Y=1.395
+ $X2=13.355 $Y2=1.605
r130 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.355 $Y=1.065
+ $X2=13.355 $Y2=1.23
r131 36 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=13.355 $Y=1.065
+ $X2=13.355 $Y2=0.825
r132 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=13.315 $Y=0.7
+ $X2=13.315 $Y2=0.825
r133 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=13.315 $Y=0.7
+ $X2=13.315 $Y2=0.445
r134 29 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.275 $Y=1.77
+ $X2=13.275 $Y2=1.605
r135 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.965 $Y=1.475
+ $X2=15.965 $Y2=1.965
r136 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.585 $Y=1.4
+ $X2=15.495 $Y2=1.4
r137 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=15.875 $Y=1.4
+ $X2=15.965 $Y2=1.475
r138 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=15.875 $Y=1.4
+ $X2=15.585 $Y2=1.4
r139 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=15.495 $Y=1.475
+ $X2=15.495 $Y2=1.4
r140 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.495 $Y=1.475
+ $X2=15.495 $Y2=1.965
r141 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.115 $Y=1.4
+ $X2=15.025 $Y2=1.4
r142 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.405 $Y=1.4
+ $X2=15.495 $Y2=1.4
r143 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=15.405 $Y=1.4
+ $X2=15.115 $Y2=1.4
r144 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=15.025 $Y=1.475
+ $X2=15.025 $Y2=1.4
r145 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.025 $Y=1.475
+ $X2=15.025 $Y2=1.965
r146 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.935 $Y=1.4
+ $X2=15.025 $Y2=1.4
r147 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.935 $Y=1.4
+ $X2=14.645 $Y2=1.4
r148 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=14.555 $Y=1.475
+ $X2=14.645 $Y2=1.4
r149 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=14.555 $Y=1.475
+ $X2=14.325 $Y2=1.285
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=14.555 $Y=1.475
+ $X2=14.555 $Y2=1.965
r151 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.13
+ $Y=1.625 $X2=13.275 $Y2=1.77
r152 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=13.14
+ $Y=0.235 $X2=13.275 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2626_599# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 29 31 33 36 44 47 48 49 50
c122 22 0 9.37986e-20 $X=15.965 $Y=3.965
c123 20 0 1.74242e-19 $X=15.875 $Y=4.04
c124 17 0 9.37986e-20 $X=15.495 $Y=3.965
c125 12 0 9.37986e-20 $X=15.025 $Y=3.965
c126 7 0 9.37986e-20 $X=14.555 $Y=3.965
r127 45 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=14.325
+ $Y=4.155 $X2=14.235 $Y2=4.21
r128 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=14.325
+ $Y=4.21 $X2=14.325 $Y2=4.21
r129 42 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=13.985 $Y=4.21
+ $X2=14.235 $Y2=4.21
r130 41 44 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=13.985 $Y=4.21
+ $X2=14.325 $Y2=4.21
r131 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.985
+ $Y=4.21 $X2=13.985 $Y2=4.21
r132 39 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.44 $Y=4.21
+ $X2=13.355 $Y2=4.21
r133 39 41 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=13.44 $Y=4.21
+ $X2=13.985 $Y2=4.21
r134 37 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.355 $Y=4.375
+ $X2=13.355 $Y2=4.21
r135 37 48 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=13.355 $Y=4.375
+ $X2=13.355 $Y2=4.615
r136 36 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=13.355 $Y=4.045
+ $X2=13.355 $Y2=4.21
r137 36 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=13.355 $Y=4.045
+ $X2=13.355 $Y2=3.835
r138 31 48 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=13.315 $Y=4.74
+ $X2=13.315 $Y2=4.615
r139 31 33 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=13.315 $Y=4.74
+ $X2=13.315 $Y2=4.995
r140 27 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.275 $Y=3.67
+ $X2=13.275 $Y2=3.835
r141 27 29 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=13.275 $Y=3.67
+ $X2=13.275 $Y2=3.14
r142 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.965 $Y=3.965
+ $X2=15.965 $Y2=3.475
r143 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.585 $Y=4.04
+ $X2=15.495 $Y2=4.04
r144 20 22 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=15.875 $Y=4.04
+ $X2=15.965 $Y2=3.965
r145 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=15.875 $Y=4.04
+ $X2=15.585 $Y2=4.04
r146 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=15.495 $Y=3.965
+ $X2=15.495 $Y2=4.04
r147 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.495 $Y=3.965
+ $X2=15.495 $Y2=3.475
r148 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.115 $Y=4.04
+ $X2=15.025 $Y2=4.04
r149 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=15.405 $Y=4.04
+ $X2=15.495 $Y2=4.04
r150 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=15.405 $Y=4.04
+ $X2=15.115 $Y2=4.04
r151 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=15.025 $Y=3.965
+ $X2=15.025 $Y2=4.04
r152 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=15.025 $Y=3.965
+ $X2=15.025 $Y2=3.475
r153 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=14.935 $Y=4.04
+ $X2=15.025 $Y2=4.04
r154 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.935 $Y=4.04
+ $X2=14.645 $Y2=4.04
r155 7 11 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=14.555 $Y=3.965
+ $X2=14.645 $Y2=4.04
r156 7 45 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=14.555 $Y=3.965
+ $X2=14.325 $Y2=4.155
r157 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=14.555 $Y=3.965
+ $X2=14.555 $Y2=3.475
r158 2 29 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.13
+ $Y=2.995 $X2=13.275 $Y2=3.14
r159 1 33 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=13.14
+ $Y=4.785 $X2=13.275 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[4] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
c99 52 0 1.35498e-19 $X=18.26 $Y=1.16
c100 31 0 1.35498e-19 $X=18.365 $Y=1.985
r101 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.34 $Y=1.16
+ $X2=18.365 $Y2=1.16
r102 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=18.26 $Y=1.16
+ $X2=18.34 $Y2=1.16
r103 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=18.26
+ $Y=1.16 $X2=18.26 $Y2=1.16
r104 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=17.92 $Y=1.16
+ $X2=18.26 $Y2=1.16
r105 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=17.895 $Y=1.16
+ $X2=17.92 $Y2=1.16
r106 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=17.4 $Y=1.16
+ $X2=17.425 $Y2=1.16
r107 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=17.24 $Y=1.16
+ $X2=17.4 $Y2=1.16
r108 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.24
+ $Y=1.16 $X2=17.24 $Y2=1.16
r109 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=16.98 $Y=1.16
+ $X2=17.24 $Y2=1.16
r110 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=16.955 $Y=1.16
+ $X2=16.98 $Y2=1.16
r111 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=17.58 $Y=1.19
+ $X2=17.24 $Y2=1.19
r112 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.58
+ $Y=1.16 $X2=17.58 $Y2=1.16
r113 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=17.515 $Y=1.16
+ $X2=17.425 $Y2=1.16
r114 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=17.515 $Y=1.16
+ $X2=17.58 $Y2=1.16
r115 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=17.805 $Y=1.16
+ $X2=17.895 $Y2=1.16
r116 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=17.805 $Y=1.16
+ $X2=17.58 $Y2=1.16
r117 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=18.17 $Y=1.19
+ $X2=18.26 $Y2=1.19
r118 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=18.17 $Y=1.19
+ $X2=17.58 $Y2=1.19
r119 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.365 $Y=1.295
+ $X2=18.365 $Y2=1.16
r120 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.365 $Y=1.295
+ $X2=18.365 $Y2=1.985
r121 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.34 $Y=1.025
+ $X2=18.34 $Y2=1.16
r122 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.34 $Y=1.025
+ $X2=18.34 $Y2=0.56
r123 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=17.92 $Y=1.025
+ $X2=17.92 $Y2=1.16
r124 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=17.92 $Y=1.025
+ $X2=17.92 $Y2=0.56
r125 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.895 $Y=1.295
+ $X2=17.895 $Y2=1.16
r126 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=17.895 $Y=1.295
+ $X2=17.895 $Y2=1.985
r127 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.425 $Y=1.295
+ $X2=17.425 $Y2=1.16
r128 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=17.425 $Y=1.295
+ $X2=17.425 $Y2=1.985
r129 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=17.4 $Y=1.025
+ $X2=17.4 $Y2=1.16
r130 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=17.4 $Y=1.025
+ $X2=17.4 $Y2=0.56
r131 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=16.98 $Y=1.025
+ $X2=16.98 $Y2=1.16
r132 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=16.98 $Y=1.025
+ $X2=16.98 $Y2=0.56
r133 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=16.955 $Y=1.295
+ $X2=16.955 $Y2=1.16
r134 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=16.955 $Y=1.295
+ $X2=16.955 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[5] 3 7 11 15 19 23 27 31 33 35 36 52
+ 54
c97 52 0 1.35498e-19 $X=18.26 $Y=4.28
c98 31 0 1.35498e-19 $X=18.365 $Y=3.455
r99 53 54 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.34 $Y=4.28
+ $X2=18.365 $Y2=4.28
r100 51 53 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=18.26 $Y=4.28
+ $X2=18.34 $Y2=4.28
r101 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=18.26
+ $Y=4.28 $X2=18.26 $Y2=4.28
r102 49 51 75.5391 $w=2.7e-07 $l=3.4e-07 $layer=POLY_cond $X=17.92 $Y=4.28
+ $X2=18.26 $Y2=4.28
r103 48 49 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=17.895 $Y=4.28
+ $X2=17.92 $Y2=4.28
r104 46 47 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=17.4 $Y=4.28
+ $X2=17.425 $Y2=4.28
r105 44 46 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=17.24 $Y=4.28
+ $X2=17.4 $Y2=4.28
r106 44 45 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.24
+ $Y=4.28 $X2=17.24 $Y2=4.28
r107 42 44 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=16.98 $Y=4.28
+ $X2=17.24 $Y2=4.28
r108 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=16.955 $Y=4.28
+ $X2=16.98 $Y2=4.28
r109 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=17.58 $Y=4.25
+ $X2=17.24 $Y2=4.25
r110 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.58
+ $Y=4.28 $X2=17.58 $Y2=4.28
r111 36 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=17.515 $Y=4.28
+ $X2=17.425 $Y2=4.28
r112 36 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=17.515 $Y=4.28
+ $X2=17.58 $Y2=4.28
r113 35 48 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=17.805 $Y=4.28
+ $X2=17.895 $Y2=4.28
r114 35 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=17.805 $Y=4.28
+ $X2=17.58 $Y2=4.28
r115 33 52 3.84148 $w=2.68e-07 $l=9e-08 $layer=LI1_cond $X=18.17 $Y=4.25
+ $X2=18.26 $Y2=4.25
r116 33 39 25.183 $w=2.68e-07 $l=5.9e-07 $layer=LI1_cond $X=18.17 $Y=4.25
+ $X2=17.58 $Y2=4.25
r117 29 54 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.365 $Y=4.145
+ $X2=18.365 $Y2=4.28
r118 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.365 $Y=4.145
+ $X2=18.365 $Y2=3.455
r119 25 53 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.34 $Y=4.415
+ $X2=18.34 $Y2=4.28
r120 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.34 $Y=4.415
+ $X2=18.34 $Y2=4.88
r121 21 49 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=17.92 $Y=4.415
+ $X2=17.92 $Y2=4.28
r122 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=17.92 $Y=4.415
+ $X2=17.92 $Y2=4.88
r123 17 48 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.895 $Y=4.145
+ $X2=17.895 $Y2=4.28
r124 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=17.895 $Y=4.145
+ $X2=17.895 $Y2=3.455
r125 13 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.425 $Y=4.145
+ $X2=17.425 $Y2=4.28
r126 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=17.425 $Y=4.145
+ $X2=17.425 $Y2=3.455
r127 9 46 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=17.4 $Y=4.415
+ $X2=17.4 $Y2=4.28
r128 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=17.4 $Y=4.415
+ $X2=17.4 $Y2=4.88
r129 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=16.98 $Y=4.415
+ $X2=16.98 $Y2=4.28
r130 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=16.98 $Y=4.415
+ $X2=16.98 $Y2=4.88
r131 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=16.955 $Y=4.145
+ $X2=16.955 $Y2=4.28
r132 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=16.955 $Y=4.145
+ $X2=16.955 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[6] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
c101 51 0 1.35498e-19 $X=20.02 $Y=1.16
c102 3 0 1.35498e-19 $X=18.895 $Y=1.985
r103 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=20.28 $Y=1.16
+ $X2=20.305 $Y2=1.16
r104 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=20.02 $Y=1.16
+ $X2=20.28 $Y2=1.16
r105 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.02
+ $Y=1.16 $X2=20.02 $Y2=1.16
r106 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=19.86 $Y=1.16
+ $X2=20.02 $Y2=1.16
r107 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.835 $Y=1.16
+ $X2=19.86 $Y2=1.16
r108 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.34 $Y=1.16
+ $X2=19.365 $Y2=1.16
r109 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.34
+ $Y=1.16 $X2=19.34 $Y2=1.16
r110 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=18.92 $Y=1.16
+ $X2=19.34 $Y2=1.16
r111 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.895 $Y=1.16
+ $X2=18.92 $Y2=1.16
r112 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.68 $Y=1.19
+ $X2=20.02 $Y2=1.19
r113 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.68 $Y=1.19
+ $X2=19.34 $Y2=1.19
r114 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.68
+ $Y=1.16 $X2=19.68 $Y2=1.16
r115 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=19.455 $Y=1.16
+ $X2=19.365 $Y2=1.16
r116 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=19.455 $Y=1.16
+ $X2=19.68 $Y2=1.16
r117 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=19.745 $Y=1.16
+ $X2=19.835 $Y2=1.16
r118 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=19.745 $Y=1.16
+ $X2=19.68 $Y2=1.16
r119 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=19.09 $Y=1.19
+ $X2=19.34 $Y2=1.19
r120 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=20.305 $Y=1.295
+ $X2=20.305 $Y2=1.16
r121 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=20.305 $Y=1.295
+ $X2=20.305 $Y2=1.985
r122 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=20.28 $Y=1.025
+ $X2=20.28 $Y2=1.16
r123 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=20.28 $Y=1.025
+ $X2=20.28 $Y2=0.56
r124 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.86 $Y=1.025
+ $X2=19.86 $Y2=1.16
r125 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.86 $Y=1.025
+ $X2=19.86 $Y2=0.56
r126 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.835 $Y=1.295
+ $X2=19.835 $Y2=1.16
r127 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.835 $Y=1.295
+ $X2=19.835 $Y2=1.985
r128 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.365 $Y=1.295
+ $X2=19.365 $Y2=1.16
r129 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.365 $Y=1.295
+ $X2=19.365 $Y2=1.985
r130 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.34 $Y=1.025
+ $X2=19.34 $Y2=1.16
r131 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.34 $Y=1.025
+ $X2=19.34 $Y2=0.56
r132 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.92 $Y=1.025
+ $X2=18.92 $Y2=1.16
r133 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.92 $Y=1.025
+ $X2=18.92 $Y2=0.56
r134 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.895 $Y=1.295
+ $X2=18.895 $Y2=1.16
r135 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.895 $Y=1.295
+ $X2=18.895 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%D[7] 3 7 11 15 19 23 27 31 33 35 36 51
+ 53
c97 51 0 1.35498e-19 $X=20.02 $Y=4.28
c98 3 0 1.35498e-19 $X=18.895 $Y=3.455
r99 52 53 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=20.28 $Y=4.28
+ $X2=20.305 $Y2=4.28
r100 50 52 57.7652 $w=2.7e-07 $l=2.6e-07 $layer=POLY_cond $X=20.02 $Y=4.28
+ $X2=20.28 $Y2=4.28
r101 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.02
+ $Y=4.28 $X2=20.02 $Y2=4.28
r102 48 50 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=19.86 $Y=4.28
+ $X2=20.02 $Y2=4.28
r103 47 48 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.835 $Y=4.28
+ $X2=19.86 $Y2=4.28
r104 44 46 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.34 $Y=4.28
+ $X2=19.365 $Y2=4.28
r105 44 45 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=19.34
+ $Y=4.28 $X2=19.34 $Y2=4.28
r106 42 44 93.313 $w=2.7e-07 $l=4.2e-07 $layer=POLY_cond $X=18.92 $Y=4.28
+ $X2=19.34 $Y2=4.28
r107 40 42 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.895 $Y=4.28
+ $X2=18.92 $Y2=4.28
r108 39 51 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.68 $Y=4.25
+ $X2=20.02 $Y2=4.25
r109 39 45 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.68 $Y=4.25
+ $X2=19.34 $Y2=4.25
r110 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.68
+ $Y=4.28 $X2=19.68 $Y2=4.28
r111 36 46 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=19.455 $Y=4.28
+ $X2=19.365 $Y2=4.28
r112 36 38 49.9891 $w=2.7e-07 $l=2.25e-07 $layer=POLY_cond $X=19.455 $Y=4.28
+ $X2=19.68 $Y2=4.28
r113 35 47 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=19.745 $Y=4.28
+ $X2=19.835 $Y2=4.28
r114 35 38 14.4413 $w=2.7e-07 $l=6.5e-08 $layer=POLY_cond $X=19.745 $Y=4.28
+ $X2=19.68 $Y2=4.28
r115 33 45 10.6708 $w=2.68e-07 $l=2.5e-07 $layer=LI1_cond $X=19.09 $Y=4.25
+ $X2=19.34 $Y2=4.25
r116 29 53 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=20.305 $Y=4.145
+ $X2=20.305 $Y2=4.28
r117 29 31 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=20.305 $Y=4.145
+ $X2=20.305 $Y2=3.455
r118 25 52 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=20.28 $Y=4.415
+ $X2=20.28 $Y2=4.28
r119 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=20.28 $Y=4.415
+ $X2=20.28 $Y2=4.88
r120 21 48 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.86 $Y=4.415
+ $X2=19.86 $Y2=4.28
r121 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.86 $Y=4.415
+ $X2=19.86 $Y2=4.88
r122 17 47 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.835 $Y=4.145
+ $X2=19.835 $Y2=4.28
r123 17 19 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.835 $Y=4.145
+ $X2=19.835 $Y2=3.455
r124 13 46 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.365 $Y=4.145
+ $X2=19.365 $Y2=4.28
r125 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.365 $Y=4.145
+ $X2=19.365 $Y2=3.455
r126 9 44 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.34 $Y=4.415
+ $X2=19.34 $Y2=4.28
r127 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.34 $Y=4.415
+ $X2=19.34 $Y2=4.88
r128 5 42 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.92 $Y=4.415
+ $X2=18.92 $Y2=4.28
r129 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.92 $Y=4.415
+ $X2=18.92 $Y2=4.88
r130 1 40 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.895 $Y=4.145
+ $X2=18.895 $Y2=4.28
r131 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.895 $Y=4.145
+ $X2=18.895 $Y2=3.455
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_265# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 45 47 48 49 50
c115 22 0 9.37986e-20 $X=22.705 $Y=1.475
c116 20 0 1.10627e-19 $X=22.615 $Y=1.4
c117 17 0 9.37986e-20 $X=22.235 $Y=1.475
c118 12 0 9.37986e-20 $X=21.765 $Y=1.475
c119 11 0 1.74242e-19 $X=21.385 $Y=1.4
c120 7 0 9.37986e-20 $X=21.295 $Y=1.475
r121 45 49 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=23.985 $Y=1.77
+ $X2=23.985 $Y2=1.605
r122 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.905 $Y=1.395
+ $X2=23.905 $Y2=1.23
r123 41 49 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=23.905 $Y=1.395
+ $X2=23.905 $Y2=1.605
r124 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.905 $Y=1.065
+ $X2=23.905 $Y2=1.23
r125 40 47 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=23.905 $Y=1.065
+ $X2=23.905 $Y2=0.825
r126 35 47 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=23.945 $Y=0.7
+ $X2=23.945 $Y2=0.825
r127 35 37 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=23.945 $Y=0.7
+ $X2=23.945 $Y2=0.445
r128 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=23.275 $Y=1.23
+ $X2=23.025 $Y2=1.23
r129 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=23.275
+ $Y=1.23 $X2=23.275 $Y2=1.23
r130 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=22.935
+ $Y=1.285 $X2=23.025 $Y2=1.23
r131 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=22.935 $Y=1.23
+ $X2=23.275 $Y2=1.23
r132 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.935
+ $Y=1.23 $X2=22.935 $Y2=1.23
r133 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=23.82 $Y=1.23
+ $X2=23.905 $Y2=1.23
r134 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=23.82 $Y=1.23
+ $X2=23.275 $Y2=1.23
r135 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=22.705
+ $Y=1.475 $X2=22.935 $Y2=1.285
r136 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.705 $Y=1.475
+ $X2=22.705 $Y2=1.965
r137 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.325 $Y=1.4
+ $X2=22.235 $Y2=1.4
r138 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=22.615 $Y=1.4
+ $X2=22.705 $Y2=1.475
r139 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.615 $Y=1.4
+ $X2=22.325 $Y2=1.4
r140 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=22.235 $Y=1.475
+ $X2=22.235 $Y2=1.4
r141 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.235 $Y=1.475
+ $X2=22.235 $Y2=1.965
r142 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.855 $Y=1.4
+ $X2=21.765 $Y2=1.4
r143 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.145 $Y=1.4
+ $X2=22.235 $Y2=1.4
r144 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.145 $Y=1.4
+ $X2=21.855 $Y2=1.4
r145 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=21.765 $Y=1.475
+ $X2=21.765 $Y2=1.4
r146 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.765 $Y=1.475
+ $X2=21.765 $Y2=1.965
r147 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.675 $Y=1.4
+ $X2=21.765 $Y2=1.4
r148 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.675 $Y=1.4
+ $X2=21.385 $Y2=1.4
r149 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=21.295 $Y=1.475
+ $X2=21.385 $Y2=1.4
r150 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.295 $Y=1.475
+ $X2=21.295 $Y2=1.965
r151 2 45 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=23.84
+ $Y=1.625 $X2=23.985 $Y2=1.77
r152 1 37 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=23.85
+ $Y=0.235 $X2=23.985 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_4239_793# 1 2 7 9 10 11 12 14 15 17
+ 19 20 22 24 25 26 27 34 37 40 43 45 47 48 49 50
c121 22 0 9.37986e-20 $X=22.705 $Y=3.965
c122 20 0 1.10627e-19 $X=22.615 $Y=4.04
c123 17 0 9.37986e-20 $X=22.235 $Y=3.965
c124 12 0 9.37986e-20 $X=21.765 $Y=3.965
c125 11 0 1.74242e-19 $X=21.385 $Y=4.04
c126 7 0 9.37986e-20 $X=21.295 $Y=3.965
r127 43 49 6.94937 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=23.945 $Y=4.74
+ $X2=23.945 $Y2=4.615
r128 43 45 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=23.945 $Y=4.74
+ $X2=23.945 $Y2=4.995
r129 41 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.905 $Y=4.375
+ $X2=23.905 $Y2=4.21
r130 41 49 15.6578 $w=1.68e-07 $l=2.4e-07 $layer=LI1_cond $X=23.905 $Y=4.375
+ $X2=23.905 $Y2=4.615
r131 40 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=23.905 $Y=4.045
+ $X2=23.905 $Y2=4.21
r132 40 47 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=23.905 $Y=4.045
+ $X2=23.905 $Y2=3.835
r133 35 47 8.46218 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=23.985 $Y=3.67
+ $X2=23.985 $Y2=3.835
r134 35 37 18.5089 $w=3.28e-07 $l=5.3e-07 $layer=LI1_cond $X=23.985 $Y=3.67
+ $X2=23.985 $Y2=3.14
r135 34 50 55.5434 $w=2.7e-07 $l=2.5e-07 $layer=POLY_cond $X=23.275 $Y=4.21
+ $X2=23.025 $Y2=4.21
r136 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=23.275
+ $Y=4.21 $X2=23.275 $Y2=4.21
r137 30 50 15.1848 $w=2.93e-07 $l=1.14237e-07 $layer=POLY_cond $X=22.935
+ $Y=4.155 $X2=23.025 $Y2=4.21
r138 29 33 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=22.935 $Y=4.21
+ $X2=23.275 $Y2=4.21
r139 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.935
+ $Y=4.21 $X2=22.935 $Y2=4.21
r140 27 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=23.82 $Y=4.21
+ $X2=23.905 $Y2=4.21
r141 27 33 19.0328 $w=3.28e-07 $l=5.45e-07 $layer=LI1_cond $X=23.82 $Y=4.21
+ $X2=23.275 $Y2=4.21
r142 22 30 37.8362 $w=2.93e-07 $l=3.10805e-07 $layer=POLY_cond $X=22.705
+ $Y=3.965 $X2=22.935 $Y2=4.155
r143 22 24 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.705 $Y=3.965
+ $X2=22.705 $Y2=3.475
r144 21 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.325 $Y=4.04
+ $X2=22.235 $Y2=4.04
r145 20 22 26.2537 $w=2.93e-07 $l=1.21861e-07 $layer=POLY_cond $X=22.615 $Y=4.04
+ $X2=22.705 $Y2=3.965
r146 20 21 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.615 $Y=4.04
+ $X2=22.325 $Y2=4.04
r147 17 26 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=22.235 $Y=3.965
+ $X2=22.235 $Y2=4.04
r148 17 19 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=22.235 $Y=3.965
+ $X2=22.235 $Y2=3.475
r149 16 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.855 $Y=4.04
+ $X2=21.765 $Y2=4.04
r150 15 26 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=22.145 $Y=4.04
+ $X2=22.235 $Y2=4.04
r151 15 16 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=22.145 $Y=4.04
+ $X2=21.855 $Y2=4.04
r152 12 25 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=21.765 $Y=3.965
+ $X2=21.765 $Y2=4.04
r153 12 14 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.765 $Y=3.965
+ $X2=21.765 $Y2=3.475
r154 10 25 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=21.675 $Y=4.04
+ $X2=21.765 $Y2=4.04
r155 10 11 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.675 $Y=4.04
+ $X2=21.385 $Y2=4.04
r156 7 11 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=21.295 $Y=3.965
+ $X2=21.385 $Y2=4.04
r157 7 9 131.211 $w=1.8e-07 $l=4.9e-07 $layer=POLY_cond $X=21.295 $Y=3.965
+ $X2=21.295 $Y2=3.475
r158 2 37 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=23.84
+ $Y=2.995 $X2=23.985 $Y2=3.14
r159 1 45 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=23.85
+ $Y=4.785 $X2=23.985 $Y2=4.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[6] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c110 11 0 1.3204e-19 $X=22.06 $Y=0.255
r111 45 49 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=24.6
+ $Y=1.16 $X2=24.6 $Y2=1.16
r112 38 49 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=24.22 $Y=1.55
+ $X2=24.427 $Y2=1.16
r113 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=24.22 $Y=1.55
+ $X2=24.22 $Y2=2.035
r114 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=24.195 $Y=0.735
+ $X2=24.195 $Y2=0.445
r115 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=23.85 $Y=0.81
+ $X2=23.75 $Y2=0.81
r116 33 49 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=24.12 $Y=0.81
+ $X2=24.427 $Y2=1.16
r117 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=24.12 $Y=0.81
+ $X2=24.195 $Y2=0.735
r118 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=24.12 $Y=0.81
+ $X2=23.85 $Y2=0.81
r119 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=23.775 $Y=0.735
+ $X2=23.75 $Y2=0.81
r120 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=23.775 $Y=0.735
+ $X2=23.775 $Y2=0.445
r121 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=23.75 $Y=1.55
+ $X2=23.75 $Y2=2.035
r122 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=23.75 $Y=1.45 $X2=23.75
+ $Y2=1.55
r123 25 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=23.75 $Y=0.885
+ $X2=23.75 $Y2=0.81
r124 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=23.75 $Y=0.885
+ $X2=23.75 $Y2=1.45
r125 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=23.65 $Y=0.81
+ $X2=23.75 $Y2=0.81
r126 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=23.65 $Y=0.81
+ $X2=23.315 $Y2=0.81
r127 22 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.24 $Y=0.735
+ $X2=23.315 $Y2=0.81
r128 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=23.24 $Y=0.255
+ $X2=23.24 $Y2=0.735
r129 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.555 $Y=0.18
+ $X2=22.48 $Y2=0.18
r130 19 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.165 $Y=0.18
+ $X2=23.24 $Y2=0.255
r131 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=23.165 $Y=0.18
+ $X2=22.555 $Y2=0.18
r132 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.48 $Y=0.255
+ $X2=22.48 $Y2=0.18
r133 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.48 $Y=0.255
+ $X2=22.48 $Y2=0.59
r134 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.135 $Y=0.18
+ $X2=22.06 $Y2=0.18
r135 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.405 $Y=0.18
+ $X2=22.48 $Y2=0.18
r136 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.405 $Y=0.18
+ $X2=22.135 $Y2=0.18
r137 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.06 $Y=0.255
+ $X2=22.06 $Y2=0.18
r138 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.06 $Y=0.255
+ $X2=22.06 $Y2=0.59
r139 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.715 $Y=0.18
+ $X2=21.64 $Y2=0.18
r140 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.985 $Y=0.18
+ $X2=22.06 $Y2=0.18
r141 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.985 $Y=0.18
+ $X2=21.715 $Y2=0.18
r142 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.64 $Y=0.255
+ $X2=21.64 $Y2=0.18
r143 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.64 $Y=0.255
+ $X2=21.64 $Y2=0.59
r144 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.565 $Y=0.18
+ $X2=21.64 $Y2=0.18
r145 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.565 $Y=0.18
+ $X2=21.295 $Y2=0.18
r146 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.22 $Y=0.255
+ $X2=21.295 $Y2=0.18
r147 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.22 $Y=0.255
+ $X2=21.22 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%S[7] 1 3 4 5 6 8 9 11 13 14 16 18 19 22
+ 23 24 25 26 27 29 30 32 33 35 37 38 40 41 42 43 44 45
c116 11 0 1.3204e-19 $X=22.06 $Y=5.185
r117 45 48 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=24.6
+ $Y=4.28 $X2=24.6 $Y2=4.28
r118 38 48 64.8801 $w=3.52e-07 $l=4.82525e-07 $layer=POLY_cond $X=24.22 $Y=3.89
+ $X2=24.427 $Y2=4.28
r119 38 40 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=24.22 $Y=3.89
+ $X2=24.22 $Y2=3.405
r120 35 37 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=24.195 $Y=4.705
+ $X2=24.195 $Y2=4.995
r121 34 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=23.85 $Y=4.63
+ $X2=23.75 $Y2=4.63
r122 33 35 26.4837 $w=3.52e-07 $l=1.06066e-07 $layer=POLY_cond $X=24.12 $Y=4.63
+ $X2=24.195 $Y2=4.705
r123 33 48 47.9261 $w=3.52e-07 $l=4.79531e-07 $layer=POLY_cond $X=24.12 $Y=4.63
+ $X2=24.427 $Y2=4.28
r124 33 34 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=24.12 $Y=4.63
+ $X2=23.85 $Y2=4.63
r125 30 44 10.2464 $w=1.5e-07 $l=8.66025e-08 $layer=POLY_cond $X=23.775 $Y=4.705
+ $X2=23.75 $Y2=4.63
r126 30 32 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=23.775 $Y=4.705
+ $X2=23.775 $Y2=4.995
r127 27 29 129.872 $w=1.8e-07 $l=4.85e-07 $layer=POLY_cond $X=23.75 $Y=3.89
+ $X2=23.75 $Y2=3.405
r128 26 44 10.2464 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=23.75 $Y=4.555
+ $X2=23.75 $Y2=4.63
r129 25 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=23.75 $Y=3.99 $X2=23.75
+ $Y2=3.89
r130 25 26 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=23.75 $Y=3.99
+ $X2=23.75 $Y2=4.555
r131 23 44 13.9575 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=23.65 $Y=4.63
+ $X2=23.75 $Y2=4.63
r132 23 24 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=23.65 $Y=4.63
+ $X2=23.315 $Y2=4.63
r133 21 24 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.24 $Y=4.705
+ $X2=23.315 $Y2=4.63
r134 21 22 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=23.24 $Y=4.705
+ $X2=23.24 $Y2=5.185
r135 20 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.555 $Y=5.26
+ $X2=22.48 $Y2=5.26
r136 19 22 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.165 $Y=5.26
+ $X2=23.24 $Y2=5.185
r137 19 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=23.165 $Y=5.26
+ $X2=22.555 $Y2=5.26
r138 16 43 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.48 $Y=5.185
+ $X2=22.48 $Y2=5.26
r139 16 18 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.48 $Y=5.185
+ $X2=22.48 $Y2=4.85
r140 15 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.135 $Y=5.26
+ $X2=22.06 $Y2=5.26
r141 14 43 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.405 $Y=5.26
+ $X2=22.48 $Y2=5.26
r142 14 15 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=22.405 $Y=5.26
+ $X2=22.135 $Y2=5.26
r143 11 42 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=22.06 $Y=5.185
+ $X2=22.06 $Y2=5.26
r144 11 13 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=22.06 $Y=5.185
+ $X2=22.06 $Y2=4.85
r145 10 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.715 $Y=5.26
+ $X2=21.64 $Y2=5.26
r146 9 42 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.985 $Y=5.26
+ $X2=22.06 $Y2=5.26
r147 9 10 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.985 $Y=5.26
+ $X2=21.715 $Y2=5.26
r148 6 41 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.64 $Y=5.185
+ $X2=21.64 $Y2=5.26
r149 6 8 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.64 $Y=5.185
+ $X2=21.64 $Y2=4.85
r150 4 41 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.565 $Y=5.26
+ $X2=21.64 $Y2=5.26
r151 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.565 $Y=5.26
+ $X2=21.295 $Y2=5.26
r152 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.22 $Y=5.185
+ $X2=21.295 $Y2=5.26
r153 1 3 107.647 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.22 $Y=5.185
+ $X2=21.22 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 111 115 119
+ 123 127 131 135 139 143 149 155 159 161 165 169 173 177 181 185 187 191 195
+ 199 203 207 211 215 219 223 229 235 239 241 245 249 253 257 261 265 267 268
+ 269 271 272 274 275 276 277 278 279 280 282 283 285 286 287 288 289 304 308
+ 313 320 340 344 349 356 362 367 370 373 376 379 382 385 388 391 394 397 398
c748 356 0 3.94334e-19 $X=20.93 $Y=2.72
c749 349 0 3.95698e-19 $X=19.465 $Y=2.72
c750 344 0 3.95698e-19 $X=18.465 $Y=2.72
c751 340 0 3.95698e-19 $X=17.525 $Y=2.72
c752 320 0 3.94334e-19 $X=8.51 $Y=2.72
c753 313 0 3.95698e-19 $X=7.045 $Y=2.72
c754 308 0 3.95698e-19 $X=6.045 $Y=2.72
c755 304 0 3.95698e-19 $X=5.105 $Y=2.72
c756 285 0 3.94334e-19 $X=23.35 $Y=2.72
c757 282 0 3.94334e-19 $X=16.585 $Y=2.72
c758 278 0 3.94334e-19 $X=13.91 $Y=2.72
c759 274 0 3.94334e-19 $X=10.93 $Y=2.72
c760 271 0 3.94334e-19 $X=4.165 $Y=2.72
c761 267 0 3.94334e-19 $X=1.49 $Y=2.72
c762 241 0 3.95698e-19 $X=20.405 $Y=2.72
c763 161 0 3.95698e-19 $X=7.985 $Y=2.72
c764 32 0 9.57576e-20 $X=20.395 $Y=2.955
c765 31 0 9.57576e-20 $X=20.395 $Y=1.485
c766 30 0 1.91515e-19 $X=19.455 $Y=2.955
c767 29 0 1.91515e-19 $X=19.455 $Y=1.485
c768 26 0 1.91515e-19 $X=17.515 $Y=2.955
c769 25 0 1.91515e-19 $X=17.515 $Y=1.485
c770 24 0 9.57576e-20 $X=16.595 $Y=2.955
c771 23 0 9.57576e-20 $X=16.595 $Y=1.485
c772 14 0 9.57576e-20 $X=7.975 $Y=2.955
c773 13 0 9.57576e-20 $X=7.975 $Y=1.485
c774 12 0 1.91515e-19 $X=7.035 $Y=2.955
c775 11 0 1.91515e-19 $X=7.035 $Y=1.485
c776 8 0 1.91515e-19 $X=5.095 $Y=2.955
c777 7 0 1.91515e-19 $X=5.095 $Y=1.485
c778 6 0 9.57576e-20 $X=4.175 $Y=2.955
c779 5 0 9.57576e-20 $X=4.175 $Y=1.485
r780 397 398 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=2.72
+ $X2=24.61 $Y2=2.72
r781 394 395 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=2.72
+ $X2=20.47 $Y2=2.72
r782 392 395 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=2.72
+ $X2=20.47 $Y2=2.72
r783 391 392 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.55 $Y=2.72
+ $X2=19.55 $Y2=2.72
r784 385 386 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=2.72
+ $X2=17.71 $Y2=2.72
r785 382 383 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r786 379 380 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r787 377 380 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=8.05 $Y2=2.72
r788 376 377 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r789 370 371 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r790 365 398 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=2.72
+ $X2=24.61 $Y2=2.72
r791 364 365 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=2.72
+ $X2=24.15 $Y2=2.72
r792 362 397 3.44808 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=24.32 $Y=2.72
+ $X2=24.58 $Y2=2.72
r793 362 364 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=24.32 $Y=2.72
+ $X2=24.15 $Y2=2.72
r794 361 365 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=2.72
+ $X2=24.15 $Y2=2.72
r795 360 361 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=23.23 $Y=2.72
+ $X2=23.23 $Y2=2.72
r796 357 361 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=2.72
+ $X2=23.23 $Y2=2.72
r797 357 395 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.93 $Y=2.72
+ $X2=20.47 $Y2=2.72
r798 356 357 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.93 $Y=2.72
+ $X2=20.93 $Y2=2.72
r799 354 394 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=20.675 $Y=2.72
+ $X2=20.54 $Y2=2.72
r800 354 356 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=20.675 $Y=2.72
+ $X2=20.93 $Y2=2.72
r801 353 392 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=2.72
+ $X2=19.55 $Y2=2.72
r802 352 353 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.09 $Y=2.72
+ $X2=19.09 $Y2=2.72
r803 350 388 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.795 $Y=2.72
+ $X2=18.63 $Y2=2.72
r804 350 352 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.795 $Y=2.72
+ $X2=19.09 $Y2=2.72
r805 349 391 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.465 $Y=2.72
+ $X2=19.6 $Y2=2.72
r806 349 352 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=19.465 $Y=2.72
+ $X2=19.09 $Y2=2.72
r807 348 386 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=2.72
+ $X2=17.71 $Y2=2.72
r808 347 348 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=2.72
+ $X2=18.17 $Y2=2.72
r809 345 385 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.795 $Y=2.72
+ $X2=17.66 $Y2=2.72
r810 345 347 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=17.795 $Y=2.72
+ $X2=18.17 $Y2=2.72
r811 344 388 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=2.72
+ $X2=18.63 $Y2=2.72
r812 344 347 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.465 $Y=2.72
+ $X2=18.17 $Y2=2.72
r813 343 386 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=17.25 $Y=2.72
+ $X2=17.71 $Y2=2.72
r814 342 343 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.25 $Y=2.72
+ $X2=17.25 $Y2=2.72
r815 340 385 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.525 $Y=2.72
+ $X2=17.66 $Y2=2.72
r816 340 342 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=17.525 $Y=2.72
+ $X2=17.25 $Y2=2.72
r817 338 343 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.33 $Y=2.72
+ $X2=17.25 $Y2=2.72
r818 337 338 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r819 335 338 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=16.33 $Y2=2.72
r820 334 335 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r821 332 335 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.03 $Y2=2.72
r822 332 383 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=12.65 $Y2=2.72
r823 331 332 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r824 329 382 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.94 $Y=2.72
+ $X2=12.79 $Y2=2.72
r825 329 331 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=12.94 $Y=2.72
+ $X2=13.57 $Y2=2.72
r826 328 383 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.65 $Y2=2.72
r827 327 328 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r828 325 328 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.73 $Y2=2.72
r829 324 325 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r830 321 325 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=10.81 $Y2=2.72
r831 321 380 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=8.05 $Y2=2.72
r832 320 321 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r833 318 379 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.12 $Y2=2.72
r834 318 320 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.255 $Y=2.72
+ $X2=8.51 $Y2=2.72
r835 317 377 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r836 316 317 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r837 314 373 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=2.72
+ $X2=6.21 $Y2=2.72
r838 314 316 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.375 $Y=2.72
+ $X2=6.67 $Y2=2.72
r839 313 376 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.045 $Y=2.72
+ $X2=7.18 $Y2=2.72
r840 313 316 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.045 $Y=2.72
+ $X2=6.67 $Y2=2.72
r841 312 371 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=5.29 $Y2=2.72
r842 311 312 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r843 309 370 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.375 $Y=2.72
+ $X2=5.24 $Y2=2.72
r844 309 311 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=2.72
+ $X2=5.75 $Y2=2.72
r845 308 373 11.8412 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=6.21 $Y2=2.72
r846 308 311 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.045 $Y=2.72
+ $X2=5.75 $Y2=2.72
r847 307 371 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r848 306 307 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r849 304 370 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=5.24 $Y2=2.72
r850 304 306 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.105 $Y=2.72
+ $X2=4.83 $Y2=2.72
r851 302 307 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r852 301 302 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r853 299 302 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=3.91 $Y2=2.72
r854 298 299 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r855 296 299 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r856 295 296 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r857 293 367 3.44808 $w=1.7e-07 $l=2.6e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.26 $Y2=2.72
r858 293 295 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=1.15 $Y2=2.72
r859 289 353 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=2.72
+ $X2=19.09 $Y2=2.72
r860 289 348 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=2.72
+ $X2=18.17 $Y2=2.72
r861 289 388 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.63 $Y=2.72
+ $X2=18.63 $Y2=2.72
r862 288 317 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r863 288 312 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r864 288 373 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r865 287 296 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r866 287 367 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r867 285 360 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=23.35 $Y=2.72
+ $X2=23.23 $Y2=2.72
r868 285 286 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=23.35 $Y=2.72
+ $X2=23.487 $Y2=2.72
r869 284 364 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=23.625 $Y=2.72
+ $X2=24.15 $Y2=2.72
r870 284 286 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=23.625 $Y=2.72
+ $X2=23.487 $Y2=2.72
r871 282 337 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=16.585 $Y=2.72
+ $X2=16.33 $Y2=2.72
r872 282 283 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.585 $Y=2.72
+ $X2=16.72 $Y2=2.72
r873 281 342 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=16.855 $Y=2.72
+ $X2=17.25 $Y2=2.72
r874 281 283 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=16.855 $Y=2.72
+ $X2=16.72 $Y2=2.72
r875 279 331 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=13.635 $Y=2.72
+ $X2=13.57 $Y2=2.72
r876 279 280 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=13.635 $Y=2.72
+ $X2=13.772 $Y2=2.72
r877 278 334 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=13.91 $Y=2.72
+ $X2=14.03 $Y2=2.72
r878 278 280 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=13.91 $Y=2.72
+ $X2=13.772 $Y2=2.72
r879 276 327 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=11.9 $Y=2.72
+ $X2=11.73 $Y2=2.72
r880 276 277 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.9 $Y=2.72
+ $X2=12.05 $Y2=2.72
r881 274 324 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=10.93 $Y=2.72
+ $X2=10.81 $Y2=2.72
r882 274 275 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=10.93 $Y=2.72
+ $X2=11.067 $Y2=2.72
r883 273 327 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=11.73 $Y2=2.72
r884 273 275 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=11.067 $Y2=2.72
r885 271 301 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r886 271 272 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.165 $Y=2.72
+ $X2=4.3 $Y2=2.72
r887 270 306 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.83 $Y2=2.72
r888 270 272 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.435 $Y=2.72
+ $X2=4.3 $Y2=2.72
r889 268 295 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.215 $Y=2.72
+ $X2=1.15 $Y2=2.72
r890 268 269 9.83177 $w=1.7e-07 $l=1.37e-07 $layer=LI1_cond $X=1.215 $Y=2.72
+ $X2=1.352 $Y2=2.72
r891 267 298 8.61176 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=1.49 $Y=2.72
+ $X2=1.61 $Y2=2.72
r892 267 269 9.83177 $w=1.7e-07 $l=1.38e-07 $layer=LI1_cond $X=1.49 $Y=2.72
+ $X2=1.352 $Y2=2.72
r893 263 397 3.14896 $w=3e-07 $l=1.46458e-07 $layer=LI1_cond $X=24.47 $Y=2.805
+ $X2=24.58 $Y2=2.72
r894 263 265 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=24.47 $Y=2.805
+ $X2=24.47 $Y2=3.14
r895 259 397 3.14896 $w=3e-07 $l=1.46458e-07 $layer=LI1_cond $X=24.47 $Y=2.635
+ $X2=24.58 $Y2=2.72
r896 259 261 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=24.47 $Y=2.635
+ $X2=24.47 $Y2=1.77
r897 255 286 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=23.487 $Y=2.805
+ $X2=23.487 $Y2=2.72
r898 255 257 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=23.487 $Y=2.805
+ $X2=23.487 $Y2=3.14
r899 251 286 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=23.487 $Y=2.635
+ $X2=23.487 $Y2=2.72
r900 251 253 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=23.487 $Y=2.635
+ $X2=23.487 $Y2=1.77
r901 247 394 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.54 $Y=2.805
+ $X2=20.54 $Y2=2.72
r902 247 249 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=20.54 $Y=2.805
+ $X2=20.54 $Y2=3.1
r903 243 394 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=20.54 $Y=2.635
+ $X2=20.54 $Y2=2.72
r904 243 245 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=20.54 $Y=2.635
+ $X2=20.54 $Y2=2
r905 242 391 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.735 $Y=2.72
+ $X2=19.6 $Y2=2.72
r906 241 394 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=20.405 $Y=2.72
+ $X2=20.54 $Y2=2.72
r907 241 242 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=20.405 $Y=2.72
+ $X2=19.735 $Y2=2.72
r908 237 391 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.6 $Y=2.805
+ $X2=19.6 $Y2=2.72
r909 237 239 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=19.6 $Y=2.805
+ $X2=19.6 $Y2=3.1
r910 233 391 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.6 $Y=2.635
+ $X2=19.6 $Y2=2.72
r911 233 235 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=19.6 $Y=2.635
+ $X2=19.6 $Y2=2
r912 229 231 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=18.63 $Y=3.1
+ $X2=18.63 $Y2=3.78
r913 227 388 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.63 $Y=2.805
+ $X2=18.63 $Y2=2.72
r914 227 229 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=18.63 $Y=2.805
+ $X2=18.63 $Y2=3.1
r915 223 226 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=18.63 $Y=1.66
+ $X2=18.63 $Y2=2.34
r916 221 388 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.63 $Y=2.635
+ $X2=18.63 $Y2=2.72
r917 221 226 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=18.63 $Y=2.635
+ $X2=18.63 $Y2=2.34
r918 217 385 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.66 $Y=2.805
+ $X2=17.66 $Y2=2.72
r919 217 219 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.66 $Y=2.805
+ $X2=17.66 $Y2=3.1
r920 213 385 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.66 $Y=2.635
+ $X2=17.66 $Y2=2.72
r921 213 215 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=17.66 $Y=2.635
+ $X2=17.66 $Y2=2
r922 209 283 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.72 $Y=2.805
+ $X2=16.72 $Y2=2.72
r923 209 211 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=16.72 $Y=2.805
+ $X2=16.72 $Y2=3.1
r924 205 283 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=16.72 $Y=2.635
+ $X2=16.72 $Y2=2.72
r925 205 207 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=16.72 $Y=2.635
+ $X2=16.72 $Y2=2
r926 201 280 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=13.772 $Y=2.805
+ $X2=13.772 $Y2=2.72
r927 201 203 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=13.772 $Y=2.805
+ $X2=13.772 $Y2=3.14
r928 197 280 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=13.772 $Y=2.635
+ $X2=13.772 $Y2=2.72
r929 197 199 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=13.772 $Y=2.635
+ $X2=13.772 $Y2=1.77
r930 193 382 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.79 $Y=2.805
+ $X2=12.79 $Y2=2.72
r931 193 195 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.79 $Y=2.805
+ $X2=12.79 $Y2=3.14
r932 189 382 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.79 $Y=2.635
+ $X2=12.79 $Y2=2.72
r933 189 191 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=12.79 $Y=2.635
+ $X2=12.79 $Y2=1.77
r934 188 277 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.2 $Y=2.72
+ $X2=12.05 $Y2=2.72
r935 187 382 10.7647 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.64 $Y=2.72
+ $X2=12.79 $Y2=2.72
r936 187 188 28.7059 $w=1.68e-07 $l=4.4e-07 $layer=LI1_cond $X=12.64 $Y=2.72
+ $X2=12.2 $Y2=2.72
r937 183 277 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.05 $Y=2.805
+ $X2=12.05 $Y2=2.72
r938 183 185 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=12.05 $Y=2.805
+ $X2=12.05 $Y2=3.14
r939 179 277 3.45667 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.05 $Y=2.635
+ $X2=12.05 $Y2=2.72
r940 179 181 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=12.05 $Y=2.635
+ $X2=12.05 $Y2=1.77
r941 175 275 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.067 $Y=2.805
+ $X2=11.067 $Y2=2.72
r942 175 177 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=11.067 $Y=2.805
+ $X2=11.067 $Y2=3.14
r943 171 275 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=11.067 $Y=2.635
+ $X2=11.067 $Y2=2.72
r944 171 173 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=11.067 $Y=2.635
+ $X2=11.067 $Y2=1.77
r945 167 379 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=2.805
+ $X2=8.12 $Y2=2.72
r946 167 169 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=8.12 $Y=2.805
+ $X2=8.12 $Y2=3.1
r947 163 379 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.12 $Y=2.635
+ $X2=8.12 $Y2=2.72
r948 163 165 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.12 $Y=2.635
+ $X2=8.12 $Y2=2
r949 162 376 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.315 $Y=2.72
+ $X2=7.18 $Y2=2.72
r950 161 379 9.68824 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.985 $Y=2.72
+ $X2=8.12 $Y2=2.72
r951 161 162 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.985 $Y=2.72
+ $X2=7.315 $Y2=2.72
r952 157 376 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=2.805
+ $X2=7.18 $Y2=2.72
r953 157 159 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.18 $Y=2.805
+ $X2=7.18 $Y2=3.1
r954 153 376 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=2.635
+ $X2=7.18 $Y2=2.72
r955 153 155 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.18 $Y=2.635
+ $X2=7.18 $Y2=2
r956 149 151 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.21 $Y=3.1
+ $X2=6.21 $Y2=3.78
r957 147 373 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.805
+ $X2=6.21 $Y2=2.72
r958 147 149 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.21 $Y=2.805
+ $X2=6.21 $Y2=3.1
r959 143 146 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=6.21 $Y=1.66
+ $X2=6.21 $Y2=2.34
r960 141 373 3.14242 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=2.635
+ $X2=6.21 $Y2=2.72
r961 141 146 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.21 $Y=2.635
+ $X2=6.21 $Y2=2.34
r962 137 370 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=2.805
+ $X2=5.24 $Y2=2.72
r963 137 139 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.24 $Y=2.805
+ $X2=5.24 $Y2=3.1
r964 133 370 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2.72
r965 133 135 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.24 $Y=2.635
+ $X2=5.24 $Y2=2
r966 129 272 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=2.805
+ $X2=4.3 $Y2=2.72
r967 129 131 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.3 $Y=2.805
+ $X2=4.3 $Y2=3.1
r968 125 272 3.84074 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=2.635
+ $X2=4.3 $Y2=2.72
r969 125 127 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.3 $Y=2.635
+ $X2=4.3 $Y2=2
r970 121 269 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.352 $Y=2.805
+ $X2=1.352 $Y2=2.72
r971 121 123 14.0389 $w=2.73e-07 $l=3.35e-07 $layer=LI1_cond $X=1.352 $Y=2.805
+ $X2=1.352 $Y2=3.14
r972 117 269 3.77091 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=1.352 $Y=2.635
+ $X2=1.352 $Y2=2.72
r973 117 119 36.2496 $w=2.73e-07 $l=8.65e-07 $layer=LI1_cond $X=1.352 $Y=2.635
+ $X2=1.352 $Y2=1.77
r974 113 367 3.14896 $w=3e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.37 $Y=2.805
+ $X2=0.26 $Y2=2.72
r975 113 115 12.8689 $w=2.98e-07 $l=3.35e-07 $layer=LI1_cond $X=0.37 $Y=2.805
+ $X2=0.37 $Y2=3.14
r976 109 367 3.14896 $w=3e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.37 $Y=2.635
+ $X2=0.26 $Y2=2.72
r977 109 111 33.2288 $w=2.98e-07 $l=8.65e-07 $layer=LI1_cond $X=0.37 $Y=2.635
+ $X2=0.37 $Y2=1.77
r978 36 265 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=24.31
+ $Y=2.995 $X2=24.455 $Y2=3.14
r979 35 261 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=24.31
+ $Y=1.625 $X2=24.455 $Y2=1.77
r980 34 257 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=23.39
+ $Y=2.995 $X2=23.515 $Y2=3.14
r981 33 253 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=23.39
+ $Y=1.625 $X2=23.515 $Y2=1.77
r982 32 249 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=20.395
+ $Y=2.955 $X2=20.54 $Y2=3.1
r983 31 245 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=20.395
+ $Y=1.485 $X2=20.54 $Y2=2
r984 30 239 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=19.455
+ $Y=2.955 $X2=19.6 $Y2=3.1
r985 29 235 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=19.455
+ $Y=1.485 $X2=19.6 $Y2=2
r986 28 231 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=18.455
+ $Y=2.955 $X2=18.63 $Y2=3.78
r987 28 229 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=18.455
+ $Y=2.955 $X2=18.63 $Y2=3.1
r988 27 226 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=18.455
+ $Y=1.485 $X2=18.63 $Y2=2.34
r989 27 223 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=18.455
+ $Y=1.485 $X2=18.63 $Y2=1.66
r990 26 219 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=17.515
+ $Y=2.955 $X2=17.66 $Y2=3.1
r991 25 215 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=17.515
+ $Y=1.485 $X2=17.66 $Y2=2
r992 24 211 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=16.595
+ $Y=2.955 $X2=16.72 $Y2=3.1
r993 23 207 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=16.595
+ $Y=1.485 $X2=16.72 $Y2=2
r994 22 203 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.6
+ $Y=2.995 $X2=13.745 $Y2=3.14
r995 21 199 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=13.6
+ $Y=1.625 $X2=13.745 $Y2=1.77
r996 20 195 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.68
+ $Y=2.995 $X2=12.805 $Y2=3.14
r997 19 191 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=12.68
+ $Y=1.625 $X2=12.805 $Y2=1.77
r998 18 185 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.89
+ $Y=2.995 $X2=12.035 $Y2=3.14
r999 17 181 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=11.89
+ $Y=1.625 $X2=12.035 $Y2=1.77
r1000 16 177 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.97
+ $Y=2.995 $X2=11.095 $Y2=3.14
r1001 15 173 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.97
+ $Y=1.625 $X2=11.095 $Y2=1.77
r1002 14 169 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.975
+ $Y=2.955 $X2=8.12 $Y2=3.1
r1003 13 165 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.975
+ $Y=1.485 $X2=8.12 $Y2=2
r1004 12 159 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=7.035
+ $Y=2.955 $X2=7.18 $Y2=3.1
r1005 11 155 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.035
+ $Y=1.485 $X2=7.18 $Y2=2
r1006 10 151 400 $w=1.7e-07 $l=9.08295e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=2.955 $X2=6.21 $Y2=3.78
r1007 10 149 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=2.955 $X2=6.21 $Y2=3.1
r1008 9 146 400 $w=1.7e-07 $l=9.3843e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.21 $Y2=2.34
r1009 9 143 400 $w=1.7e-07 $l=2.47487e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.21 $Y2=1.66
r1010 8 139 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=2.955 $X2=5.24 $Y2=3.1
r1011 7 135 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.095
+ $Y=1.485 $X2=5.24 $Y2=2
r1012 6 131 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=2.955 $X2=4.3 $Y2=3.1
r1013 5 127 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=4.175
+ $Y=1.485 $X2=4.3 $Y2=2
r1014 4 123 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=2.995 $X2=1.325 $Y2=3.14
r1015 3 119 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.18
+ $Y=1.625 $X2=1.325 $Y2=1.77
r1016 2 115 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.26
+ $Y=2.995 $X2=0.385 $Y2=3.14
r1017 1 111 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.26
+ $Y=1.625 $X2=0.385 $Y2=1.77
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_311# 1 2 3 4 5 16 17 18 23 24 27
+ 28 29 30 31 32 33 34 47 49 50 53 58 63
c127 58 0 1.3204e-19 $X=2.84 $Y=1.7
c128 49 0 1.97849e-19 $X=5.71 $Y=2.225
c129 34 0 1.97849e-19 $X=4.915 $Y=2.225
c130 33 0 1.91515e-19 $X=5.565 $Y=2.225
c131 32 0 1.97167e-19 $X=3.935 $Y=2.225
c132 31 0 9.57576e-20 $X=4.625 $Y=2.225
c133 29 0 1.87597e-19 $X=3.645 $Y=2.225
c134 28 0 1.97167e-19 $X=2.035 $Y=2.225
c135 27 0 1.87597e-19 $X=2.695 $Y=2.225
r136 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.71 $Y=2.225
+ $X2=5.71 $Y2=2.225
r137 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.77 $Y=2.225
+ $X2=4.77 $Y2=2.225
r138 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=3.795 $Y=2.225
+ $X2=3.795 $Y2=1.7
r139 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.79 $Y=2.225
+ $X2=3.79 $Y2=2.225
r140 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.84 $Y=2.225
+ $X2=2.84 $Y2=1.7
r141 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=2.225
+ $X2=2.84 $Y2=2.225
r142 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=1.885 $Y=2.225
+ $X2=1.885 $Y2=1.73
r143 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.89 $Y=2.225
+ $X2=1.89 $Y2=2.225
r144 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.915 $Y=2.225
+ $X2=4.77 $Y2=2.225
r145 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.565 $Y=2.225
+ $X2=5.71 $Y2=2.225
r146 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=5.565 $Y=2.225
+ $X2=4.915 $Y2=2.225
r147 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=2.225
+ $X2=3.79 $Y2=2.225
r148 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.625 $Y=2.225
+ $X2=4.77 $Y2=2.225
r149 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=4.625 $Y=2.225
+ $X2=3.935 $Y2=2.225
r150 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=2.225
+ $X2=2.84 $Y2=2.225
r151 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.645 $Y=2.225
+ $X2=3.79 $Y2=2.225
r152 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=3.645 $Y=2.225
+ $X2=2.985 $Y2=2.225
r153 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.035 $Y=2.225
+ $X2=1.89 $Y2=2.225
r154 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=2.225
+ $X2=2.84 $Y2=2.225
r155 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=2.695 $Y=2.225
+ $X2=2.035 $Y2=2.225
r156 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=5.71 $Y=1.665
+ $X2=5.71 $Y2=2.225
r157 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=1.665
+ $X2=5.71 $Y2=1.58
r158 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=4.77 $Y=1.665
+ $X2=4.77 $Y2=2.225
r159 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=1.665
+ $X2=4.77 $Y2=1.58
r160 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=3.795 $Y=1.665
+ $X2=3.795 $Y2=1.7
r161 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=1.58
+ $X2=4.77 $Y2=1.58
r162 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=1.58
+ $X2=5.71 $Y2=1.58
r163 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.545 $Y=1.58
+ $X2=4.935 $Y2=1.58
r164 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.945 $Y=1.58
+ $X2=3.795 $Y2=1.665
r165 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=1.58
+ $X2=4.77 $Y2=1.58
r166 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.605 $Y=1.58
+ $X2=3.945 $Y2=1.58
r167 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.34
r168 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.66
r169 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=2.34
r170 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=1.485 $X2=4.77 $Y2=1.66
r171 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.635
+ $Y=1.555 $X2=3.78 $Y2=1.7
r172 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.695
+ $Y=1.555 $X2=2.84 $Y2=1.7
r173 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=1.775
+ $Y=1.555 $X2=1.9 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_355_613# 1 2 3 4 5 16 17 18 23 24 27
+ 28 29 30 31 32 33 34 49 53 57 61 64 67
c127 57 0 1.3204e-19 $X=2.84 $Y=3.21
c128 49 0 1.97849e-19 $X=5.71 $Y=3.215
c129 34 0 1.97849e-19 $X=4.915 $Y=3.215
c130 33 0 1.91515e-19 $X=5.565 $Y=3.215
c131 32 0 1.97167e-19 $X=3.935 $Y=3.215
c132 31 0 9.57576e-20 $X=4.625 $Y=3.215
c133 29 0 1.87597e-19 $X=3.645 $Y=3.215
c134 28 0 1.97167e-19 $X=2.035 $Y=3.215
c135 27 0 1.87597e-19 $X=2.695 $Y=3.215
r136 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.71 $Y=3.215
+ $X2=5.71 $Y2=3.215
r137 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.77 $Y=3.215
+ $X2=4.77 $Y2=3.215
r138 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.79 $Y=3.215
+ $X2=3.79 $Y2=3.215
r139 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.84 $Y=3.215
+ $X2=2.84 $Y2=3.215
r140 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.89 $Y=3.215
+ $X2=1.89 $Y2=3.215
r141 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.915 $Y=3.215
+ $X2=4.77 $Y2=3.215
r142 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.565 $Y=3.215
+ $X2=5.71 $Y2=3.215
r143 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=5.565 $Y=3.215
+ $X2=4.915 $Y2=3.215
r144 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.935 $Y=3.215
+ $X2=3.79 $Y2=3.215
r145 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.625 $Y=3.215
+ $X2=4.77 $Y2=3.215
r146 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=4.625 $Y=3.215
+ $X2=3.935 $Y2=3.215
r147 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.985 $Y=3.215
+ $X2=2.84 $Y2=3.215
r148 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.645 $Y=3.215
+ $X2=3.79 $Y2=3.215
r149 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=3.645 $Y=3.215
+ $X2=2.985 $Y2=3.215
r150 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.035 $Y=3.215
+ $X2=1.89 $Y2=3.215
r151 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.695 $Y=3.215
+ $X2=2.84 $Y2=3.215
r152 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=2.695 $Y=3.215
+ $X2=2.035 $Y2=3.215
r153 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=5.71 $Y=3.775
+ $X2=5.71 $Y2=3.1
r154 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.71 $Y=3.775
+ $X2=5.71 $Y2=3.86
r155 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=4.77 $Y=3.775
+ $X2=4.77 $Y2=3.1
r156 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=3.775
+ $X2=4.77 $Y2=3.86
r157 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=3.795 $Y=3.775
+ $X2=3.795 $Y2=3.21
r158 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=3.86
+ $X2=4.77 $Y2=3.86
r159 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=3.86
+ $X2=5.71 $Y2=3.86
r160 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.545 $Y=3.86
+ $X2=4.935 $Y2=3.86
r161 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=3.945 $Y=3.86
+ $X2=3.795 $Y2=3.775
r162 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=3.86
+ $X2=4.77 $Y2=3.86
r163 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.605 $Y=3.86
+ $X2=3.945 $Y2=3.86
r164 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.955 $X2=5.71 $Y2=3.1
r165 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=2.955 $X2=5.71 $Y2=3.78
r166 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=2.955 $X2=4.77 $Y2=3.1
r167 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.625
+ $Y=2.955 $X2=4.77 $Y2=3.78
r168 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.635
+ $Y=3.065 $X2=3.78 $Y2=3.21
r169 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.695
+ $Y=3.065 $X2=2.84 $Y2=3.21
r170 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.775
+ $Y=3.065 $X2=1.9 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 99 103 105 107 110 114 117
+ 119 123 127 131 135 137 139 142 146 149 151 155 159 162 164 166 168 170 174
+ 175 178 182 183 186 188 190 192 194 196 198 200 202 206 207 210 214 215 218
+ 220 222 224 225 226 227 228 229 230 231 232 233 234 235 236 237 241 245 249
+ 253 257 261 265 269 270 271 272 273 274 275 276 294 303 308 313 322 331 336
+ 341
c914 235 0 3.48484e-19 $X=21.385 $Y=3.57
c915 233 0 3.48484e-19 $X=21.385 $Y=1.87
c916 227 0 3.48484e-19 $X=8.965 $Y=3.57
c917 225 0 3.48484e-19 $X=8.965 $Y=1.87
c918 224 0 1.20815e-19 $X=22.37 $Y=4.225
c919 222 0 1.20815e-19 $X=22.37 $Y=1.215
c920 196 0 1.20815e-19 $X=14.89 $Y=4.225
c921 194 0 1.20815e-19 $X=14.89 $Y=1.215
c922 192 0 1.20815e-19 $X=9.95 $Y=4.225
c923 190 0 1.20815e-19 $X=9.95 $Y=1.215
c924 164 0 1.20815e-19 $X=2.47 $Y=4.225
c925 162 0 1.20815e-19 $X=2.47 $Y=1.215
r926 345 347 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=22.47 $Y=3.21
+ $X2=22.47 $Y2=3.57
r927 341 345 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=22.47 $Y=1.7
+ $X2=22.47 $Y2=3.21
r928 336 338 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=21.53 $Y=1.7
+ $X2=21.53 $Y2=3.21
r929 331 333 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=15.73 $Y=1.7
+ $X2=15.73 $Y2=3.21
r930 326 328 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=14.79 $Y=3.21
+ $X2=14.79 $Y2=3.57
r931 322 326 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=14.79 $Y=1.7
+ $X2=14.79 $Y2=3.21
r932 317 319 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=10.05 $Y=3.21
+ $X2=10.05 $Y2=3.57
r933 313 317 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=10.05 $Y=1.7
+ $X2=10.05 $Y2=3.21
r934 308 310 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=9.11 $Y=1.7
+ $X2=9.11 $Y2=3.21
r935 303 305 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=3.31 $Y=1.7
+ $X2=3.31 $Y2=3.21
r936 298 300 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=2.37 $Y=3.21
+ $X2=2.37 $Y2=3.57
r937 294 298 52.733 $w=3.28e-07 $l=1.51e-06 $layer=LI1_cond $X=2.37 $Y=1.7
+ $X2=2.37 $Y2=3.21
r938 276 347 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.47 $Y=3.57
+ $X2=22.47 $Y2=3.57
r939 275 341 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.47 $Y=1.87
+ $X2=22.47 $Y2=1.87
r940 274 328 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.79 $Y=3.57
+ $X2=14.79 $Y2=3.57
r941 273 322 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.79 $Y=1.87
+ $X2=14.79 $Y2=1.87
r942 272 319 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.05 $Y=3.57
+ $X2=10.05 $Y2=3.57
r943 271 313 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.05 $Y=1.87
+ $X2=10.05 $Y2=1.87
r944 270 300 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.37 $Y=3.57
+ $X2=2.37 $Y2=3.57
r945 269 294 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.37 $Y=1.87
+ $X2=2.37 $Y2=1.87
r946 268 338 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=21.53 $Y=3.57
+ $X2=21.53 $Y2=3.21
r947 267 268 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.53 $Y=3.57
+ $X2=21.53 $Y2=3.57
r948 265 276 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=21.675 $Y=3.57
+ $X2=22.325 $Y2=3.57
r949 265 267 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.675 $Y=3.57
+ $X2=21.53 $Y2=3.57
r950 263 336 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.53 $Y=1.87
+ $X2=21.53 $Y2=1.87
r951 261 275 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=21.675 $Y=1.87
+ $X2=22.325 $Y2=1.87
r952 261 263 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.675 $Y=1.87
+ $X2=21.53 $Y2=1.87
r953 260 333 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=15.73 $Y=3.57
+ $X2=15.73 $Y2=3.21
r954 259 260 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.73 $Y=3.57
+ $X2=15.73 $Y2=3.57
r955 257 274 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=15.585 $Y=3.57
+ $X2=14.935 $Y2=3.57
r956 257 259 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.585 $Y=3.57
+ $X2=15.73 $Y2=3.57
r957 255 331 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.73 $Y=1.87
+ $X2=15.73 $Y2=1.87
r958 253 273 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=15.585 $Y=1.87
+ $X2=14.935 $Y2=1.87
r959 253 255 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.585 $Y=1.87
+ $X2=15.73 $Y2=1.87
r960 252 310 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=9.11 $Y=3.57
+ $X2=9.11 $Y2=3.21
r961 251 252 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.11 $Y=3.57
+ $X2=9.11 $Y2=3.57
r962 249 272 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=9.255 $Y=3.57
+ $X2=9.905 $Y2=3.57
r963 249 251 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.255 $Y=3.57
+ $X2=9.11 $Y2=3.57
r964 247 308 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.11 $Y=1.87
+ $X2=9.11 $Y2=1.87
r965 245 271 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=9.255 $Y=1.87
+ $X2=9.905 $Y2=1.87
r966 245 247 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.255 $Y=1.87
+ $X2=9.11 $Y2=1.87
r967 244 305 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=3.31 $Y=3.57
+ $X2=3.31 $Y2=3.21
r968 243 244 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.31 $Y=3.57
+ $X2=3.31 $Y2=3.57
r969 241 270 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=3.165 $Y=3.57
+ $X2=2.515 $Y2=3.57
r970 241 243 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.165 $Y=3.57
+ $X2=3.31 $Y2=3.57
r971 239 303 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.31 $Y=1.87
+ $X2=3.31 $Y2=1.87
r972 237 269 0.361005 $w=2.8e-07 $l=6.5e-07 $layer=MET1_cond $X=3.165 $Y=1.87
+ $X2=2.515 $Y2=1.87
r973 237 239 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.165 $Y=1.87
+ $X2=3.31 $Y2=1.87
r974 236 259 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.875 $Y=3.57
+ $X2=15.73 $Y2=3.57
r975 235 267 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.385 $Y=3.57
+ $X2=21.53 $Y2=3.57
r976 235 236 6.81929 $w=1.4e-07 $l=5.51e-06 $layer=MET1_cond $X=21.385 $Y=3.57
+ $X2=15.875 $Y2=3.57
r977 234 255 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.875 $Y=1.87
+ $X2=15.73 $Y2=1.87
r978 233 263 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.385 $Y=1.87
+ $X2=21.53 $Y2=1.87
r979 233 234 6.81929 $w=1.4e-07 $l=5.51e-06 $layer=MET1_cond $X=21.385 $Y=1.87
+ $X2=15.875 $Y2=1.87
r980 232 272 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=10.195 $Y=3.57
+ $X2=9.99 $Y2=3.57
r981 231 274 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.645 $Y=3.57
+ $X2=14.79 $Y2=3.57
r982 231 232 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=14.645 $Y=3.57
+ $X2=10.195 $Y2=3.57
r983 230 271 0.153963 $w=2.3e-07 $l=2.05e-07 $layer=MET1_cond $X=10.195 $Y=1.87
+ $X2=9.99 $Y2=1.87
r984 229 273 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.645 $Y=1.87
+ $X2=14.79 $Y2=1.87
r985 229 230 5.50742 $w=1.4e-07 $l=4.45e-06 $layer=MET1_cond $X=14.645 $Y=1.87
+ $X2=10.195 $Y2=1.87
r986 228 243 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=3.57
+ $X2=3.31 $Y2=3.57
r987 227 251 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.965 $Y=3.57
+ $X2=9.11 $Y2=3.57
r988 227 228 6.81929 $w=1.4e-07 $l=5.51e-06 $layer=MET1_cond $X=8.965 $Y=3.57
+ $X2=3.455 $Y2=3.57
r989 226 239 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.455 $Y=1.87
+ $X2=3.31 $Y2=1.87
r990 225 247 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.965 $Y=1.87
+ $X2=9.11 $Y2=1.87
r991 225 226 6.81929 $w=1.4e-07 $l=5.51e-06 $layer=MET1_cond $X=8.965 $Y=1.87
+ $X2=3.455 $Y2=1.87
r992 223 347 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=22.47 $Y=4.075
+ $X2=22.47 $Y2=3.57
r993 223 224 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=22.47 $Y=4.075
+ $X2=22.37 $Y2=4.225
r994 221 341 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=22.47 $Y=1.365
+ $X2=22.47 $Y2=1.7
r995 221 222 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=22.47 $Y=1.365
+ $X2=22.37 $Y2=1.215
r996 219 268 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=21.53 $Y=4.075
+ $X2=21.53 $Y2=3.57
r997 219 220 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=21.53 $Y=4.075
+ $X2=21.53 $Y2=4.225
r998 217 336 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=21.53 $Y=1.365
+ $X2=21.53 $Y2=1.7
r999 217 218 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=21.53 $Y=1.365
+ $X2=21.53 $Y2=1.215
r1000 214 215 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=21.43 $Y=4.76
+ $X2=21.43 $Y2=4.555
r1001 210 212 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=21.43 $Y=0.68
+ $X2=21.43 $Y2=0.885
r1002 206 207 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.83 $Y=4.76
+ $X2=15.83 $Y2=4.555
r1003 202 204 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=15.83 $Y=0.68
+ $X2=15.83 $Y2=0.885
r1004 199 260 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=15.73 $Y=4.075
+ $X2=15.73 $Y2=3.57
r1005 199 200 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=15.73 $Y=4.075
+ $X2=15.73 $Y2=4.225
r1006 197 331 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=15.73 $Y=1.365
+ $X2=15.73 $Y2=1.7
r1007 197 198 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=15.73 $Y=1.365
+ $X2=15.73 $Y2=1.215
r1008 195 328 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=14.79 $Y=4.075
+ $X2=14.79 $Y2=3.57
r1009 195 196 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=14.79
+ $Y=4.075 $X2=14.89 $Y2=4.225
r1010 193 322 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=14.79 $Y=1.365
+ $X2=14.79 $Y2=1.7
r1011 193 194 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=14.79
+ $Y=1.365 $X2=14.89 $Y2=1.215
r1012 191 319 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=10.05 $Y=4.075
+ $X2=10.05 $Y2=3.57
r1013 191 192 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=10.05
+ $Y=4.075 $X2=9.95 $Y2=4.225
r1014 189 313 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=10.05 $Y=1.365
+ $X2=10.05 $Y2=1.7
r1015 189 190 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=10.05
+ $Y=1.365 $X2=9.95 $Y2=1.215
r1016 187 252 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=9.11 $Y=4.075
+ $X2=9.11 $Y2=3.57
r1017 187 188 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=9.11 $Y=4.075
+ $X2=9.11 $Y2=4.225
r1018 185 308 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=9.11 $Y=1.365
+ $X2=9.11 $Y2=1.7
r1019 185 186 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=9.11 $Y=1.365
+ $X2=9.11 $Y2=1.215
r1020 182 183 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.01 $Y=4.76
+ $X2=9.01 $Y2=4.555
r1021 178 180 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=9.01 $Y=0.68
+ $X2=9.01 $Y2=0.885
r1022 174 175 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.41 $Y=4.76
+ $X2=3.41 $Y2=4.555
r1023 170 172 8.22951 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=3.41 $Y=0.68
+ $X2=3.41 $Y2=0.885
r1024 167 244 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=3.31 $Y=4.075
+ $X2=3.31 $Y2=3.57
r1025 167 168 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.31 $Y=4.075
+ $X2=3.31 $Y2=4.225
r1026 165 303 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=3.31 $Y=1.365
+ $X2=3.31 $Y2=1.7
r1027 165 166 5.46921 $w=2.8e-07 $l=1.5e-07 $layer=LI1_cond $X=3.31 $Y=1.365
+ $X2=3.31 $Y2=1.215
r1028 163 300 17.6359 $w=3.28e-07 $l=5.05e-07 $layer=LI1_cond $X=2.37 $Y=4.075
+ $X2=2.37 $Y2=3.57
r1029 163 164 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=2.37 $Y=4.075
+ $X2=2.47 $Y2=4.225
r1030 161 294 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=2.37 $Y=1.365
+ $X2=2.37 $Y2=1.7
r1031 161 162 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=2.37 $Y=1.365
+ $X2=2.47 $Y2=1.215
r1032 157 224 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=22.27
+ $Y=4.375 $X2=22.37 $Y2=4.225
r1033 157 159 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=22.27 $Y=4.375
+ $X2=22.27 $Y2=4.76
r1034 153 222 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=22.27
+ $Y=1.065 $X2=22.37 $Y2=1.215
r1035 153 155 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=22.27 $Y=1.065
+ $X2=22.27 $Y2=0.68
r1036 152 220 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=21.695 $Y=4.225
+ $X2=21.53 $Y2=4.225
r1037 151 224 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=22.105 $Y=4.225
+ $X2=22.37 $Y2=4.225
r1038 151 152 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=22.105 $Y=4.225
+ $X2=21.695 $Y2=4.225
r1039 150 218 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=21.695 $Y=1.215
+ $X2=21.53 $Y2=1.215
r1040 149 222 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=22.105 $Y=1.215
+ $X2=22.37 $Y2=1.215
r1041 149 150 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=22.105 $Y=1.215
+ $X2=21.695 $Y2=1.215
r1042 147 220 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=21.48
+ $Y=4.375 $X2=21.53 $Y2=4.225
r1043 147 215 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=21.48 $Y=4.375
+ $X2=21.48 $Y2=4.555
r1044 146 218 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=21.48
+ $Y=1.065 $X2=21.53 $Y2=1.215
r1045 146 212 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=21.48 $Y=1.065
+ $X2=21.48 $Y2=0.885
r1046 143 200 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=15.78
+ $Y=4.375 $X2=15.73 $Y2=4.225
r1047 143 207 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=15.78 $Y=4.375
+ $X2=15.78 $Y2=4.555
r1048 142 198 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=15.78
+ $Y=1.065 $X2=15.73 $Y2=1.215
r1049 142 204 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=15.78 $Y=1.065
+ $X2=15.78 $Y2=0.885
r1050 140 196 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=15.155 $Y=4.225
+ $X2=14.89 $Y2=4.225
r1051 139 200 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=15.565 $Y=4.225
+ $X2=15.73 $Y2=4.225
r1052 139 140 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=15.565 $Y=4.225
+ $X2=15.155 $Y2=4.225
r1053 138 194 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=15.155 $Y=1.215
+ $X2=14.89 $Y2=1.215
r1054 137 198 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=15.565 $Y=1.215
+ $X2=15.73 $Y2=1.215
r1055 137 138 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=15.565 $Y=1.215
+ $X2=15.155 $Y2=1.215
r1056 133 196 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=14.99
+ $Y=4.375 $X2=14.89 $Y2=4.225
r1057 133 135 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=14.99 $Y=4.375
+ $X2=14.99 $Y2=4.76
r1058 129 194 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=14.99
+ $Y=1.065 $X2=14.89 $Y2=1.215
r1059 129 131 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=14.99 $Y=1.065
+ $X2=14.99 $Y2=0.68
r1060 125 192 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.85 $Y=4.375
+ $X2=9.95 $Y2=4.225
r1061 125 127 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.85 $Y=4.375
+ $X2=9.85 $Y2=4.76
r1062 121 190 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=9.85 $Y=1.065
+ $X2=9.95 $Y2=1.215
r1063 121 123 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=9.85 $Y=1.065
+ $X2=9.85 $Y2=0.68
r1064 120 188 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=4.225
+ $X2=9.11 $Y2=4.225
r1065 119 192 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=9.685 $Y=4.225
+ $X2=9.95 $Y2=4.225
r1066 119 120 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=9.685 $Y=4.225
+ $X2=9.275 $Y2=4.225
r1067 118 186 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=9.275 $Y=1.215
+ $X2=9.11 $Y2=1.215
r1068 117 190 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=9.685 $Y=1.215
+ $X2=9.95 $Y2=1.215
r1069 117 118 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=9.685 $Y=1.215
+ $X2=9.275 $Y2=1.215
r1070 115 188 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=9.06 $Y=4.375
+ $X2=9.11 $Y2=4.225
r1071 115 183 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.06 $Y=4.375
+ $X2=9.06 $Y2=4.555
r1072 114 186 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=9.06 $Y=1.065
+ $X2=9.11 $Y2=1.215
r1073 114 180 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=9.06 $Y=1.065
+ $X2=9.06 $Y2=0.885
r1074 111 168 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.36 $Y=4.375
+ $X2=3.31 $Y2=4.225
r1075 111 175 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.36 $Y=4.375
+ $X2=3.36 $Y2=4.555
r1076 110 166 5.46921 $w=2.8e-07 $l=1.73205e-07 $layer=LI1_cond $X=3.36 $Y=1.065
+ $X2=3.31 $Y2=1.215
r1077 110 172 9.01912 $w=2.28e-07 $l=1.8e-07 $layer=LI1_cond $X=3.36 $Y=1.065
+ $X2=3.36 $Y2=0.885
r1078 108 164 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=2.735 $Y=4.225
+ $X2=2.47 $Y2=4.225
r1079 107 168 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=4.225
+ $X2=3.31 $Y2=4.225
r1080 107 108 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.145 $Y=4.225
+ $X2=2.735 $Y2=4.225
r1081 106 162 1.68792 $w=3e-07 $l=2.65e-07 $layer=LI1_cond $X=2.735 $Y=1.215
+ $X2=2.47 $Y2=1.215
r1082 105 166 1.09533 $w=3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.145 $Y=1.215
+ $X2=3.31 $Y2=1.215
r1083 105 106 15.7501 $w=2.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.145 $Y=1.215
+ $X2=2.735 $Y2=1.215
r1084 101 164 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=2.57 $Y=4.375
+ $X2=2.47 $Y2=4.225
r1085 101 103 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.57 $Y=4.375
+ $X2=2.57 $Y2=4.76
r1086 97 162 4.76867 $w=3.3e-07 $l=1.93649e-07 $layer=LI1_cond $X=2.57 $Y=1.065
+ $X2=2.47 $Y2=1.215
r1087 97 99 13.4452 $w=3.28e-07 $l=3.85e-07 $layer=LI1_cond $X=2.57 $Y=1.065
+ $X2=2.57 $Y2=0.68
r1088 32 345 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=22.325 $Y=3.065 $X2=22.47 $Y2=3.21
r1089 31 341 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=22.325 $Y=1.555 $X2=22.47 $Y2=1.7
r1090 30 338 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=21.385 $Y=3.065 $X2=21.53 $Y2=3.21
r1091 29 336 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=21.385 $Y=1.555 $X2=21.53 $Y2=1.7
r1092 28 333 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=15.585 $Y=3.065 $X2=15.73 $Y2=3.21
r1093 27 331 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=15.585 $Y=1.555 $X2=15.73 $Y2=1.7
r1094 26 326 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=14.645 $Y=3.065 $X2=14.79 $Y2=3.21
r1095 25 322 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2
+ $X=14.645 $Y=1.555 $X2=14.79 $Y2=1.7
r1096 24 317 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.905
+ $Y=3.065 $X2=10.05 $Y2=3.21
r1097 23 313 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.905
+ $Y=1.555 $X2=10.05 $Y2=1.7
r1098 22 310 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.965
+ $Y=3.065 $X2=9.11 $Y2=3.21
r1099 21 308 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.965
+ $Y=1.555 $X2=9.11 $Y2=1.7
r1100 20 305 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=3.065 $X2=3.31 $Y2=3.21
r1101 19 303 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=3.165
+ $Y=1.555 $X2=3.31 $Y2=1.7
r1102 18 298 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=3.065 $X2=2.37 $Y2=3.21
r1103 17 294 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.225
+ $Y=1.555 $X2=2.37 $Y2=1.7
r1104 16 159 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=22.135 $Y=4.59 $X2=22.27 $Y2=4.76
r1105 15 155 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=22.135 $Y=0.33 $X2=22.27 $Y2=0.68
r1106 14 214 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=21.295 $Y=4.59 $X2=21.43 $Y2=4.76
r1107 13 210 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=21.295 $Y=0.33 $X2=21.43 $Y2=0.68
r1108 12 206 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=15.695 $Y=4.59 $X2=15.83 $Y2=4.76
r1109 11 202 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1
+ $X=15.695 $Y=0.33 $X2=15.83 $Y2=0.68
r1110 10 135 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1
+ $X=14.855 $Y=4.59 $X2=14.99 $Y2=4.76
r1111 9 131 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=14.855
+ $Y=0.33 $X2=14.99 $Y2=0.68
r1112 8 127 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=4.59 $X2=9.85 $Y2=4.76
r1113 7 123 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=0.33 $X2=9.85 $Y2=0.68
r1114 6 182 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=4.59 $X2=9.01 $Y2=4.76
r1115 5 178 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=8.875
+ $Y=0.33 $X2=9.01 $Y2=0.68
r1116 4 174 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=4.59 $X2=3.41 $Y2=4.76
r1117 3 170 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.33 $X2=3.41 $Y2=0.68
r1118 2 103 182 $w=1.7e-07 $l=2.27706e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=4.59 $X2=2.57 $Y2=4.76
r1119 1 99 182 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_NDIFF $count=1 $X=2.435
+ $Y=0.33 $X2=2.57 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_297# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 37 41 49 59 63 68
c128 63 0 1.3204e-19 $X=9.58 $Y=1.7
c129 49 0 1.97167e-19 $X=10.53 $Y=2.225
c130 33 0 1.87597e-19 $X=10.385 $Y=2.225
c131 32 0 1.97167e-19 $X=8.775 $Y=2.225
c132 31 0 1.87597e-19 $X=9.435 $Y=2.225
c133 30 0 1.97849e-19 $X=7.795 $Y=2.225
c134 29 0 9.57576e-20 $X=8.485 $Y=2.225
c135 28 0 1.97849e-19 $X=6.855 $Y=2.225
c136 27 0 1.91515e-19 $X=7.505 $Y=2.225
r137 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=10.535 $Y=2.225
+ $X2=10.535 $Y2=1.73
r138 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.53 $Y=2.225
+ $X2=10.53 $Y2=2.225
r139 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=9.58 $Y=2.225
+ $X2=9.58 $Y2=1.7
r140 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.58 $Y=2.225
+ $X2=9.58 $Y2=2.225
r141 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=8.625 $Y=2.225
+ $X2=8.625 $Y2=1.7
r142 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.63 $Y=2.225
+ $X2=8.63 $Y2=2.225
r143 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.65 $Y=2.225
+ $X2=7.65 $Y2=2.225
r144 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=2.225
+ $X2=6.71 $Y2=2.225
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.725 $Y=2.225
+ $X2=9.58 $Y2=2.225
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.385 $Y=2.225
+ $X2=10.53 $Y2=2.225
r147 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=10.385 $Y=2.225
+ $X2=9.725 $Y2=2.225
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.775 $Y=2.225
+ $X2=8.63 $Y2=2.225
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.435 $Y=2.225
+ $X2=9.58 $Y2=2.225
r150 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=9.435 $Y=2.225
+ $X2=8.775 $Y2=2.225
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.795 $Y=2.225
+ $X2=7.65 $Y2=2.225
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.485 $Y=2.225
+ $X2=8.63 $Y2=2.225
r153 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=8.485 $Y=2.225
+ $X2=7.795 $Y2=2.225
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.855 $Y=2.225
+ $X2=6.71 $Y2=2.225
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.505 $Y=2.225
+ $X2=7.65 $Y2=2.225
r156 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=7.505 $Y=2.225
+ $X2=6.855 $Y2=2.225
r157 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=8.625 $Y=1.665
+ $X2=8.625 $Y2=1.7
r158 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=7.65 $Y=1.665
+ $X2=7.65 $Y2=2.225
r159 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.65 $Y=1.665
+ $X2=7.65 $Y2=1.58
r160 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=6.71 $Y=1.665
+ $X2=6.71 $Y2=2.225
r161 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.71 $Y=1.665
+ $X2=6.71 $Y2=1.58
r162 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=1.58
+ $X2=7.65 $Y2=1.58
r163 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.475 $Y=1.58
+ $X2=8.625 $Y2=1.665
r164 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.475 $Y=1.58
+ $X2=7.815 $Y2=1.58
r165 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=1.58
+ $X2=6.71 $Y2=1.58
r166 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=1.58
+ $X2=7.65 $Y2=1.58
r167 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.485 $Y=1.58
+ $X2=6.875 $Y2=1.58
r168 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=10.375
+ $Y=1.555 $X2=10.52 $Y2=1.73
r169 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.435
+ $Y=1.555 $X2=9.58 $Y2=1.7
r170 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.515
+ $Y=1.555 $X2=8.64 $Y2=1.7
r171 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=1.485 $X2=7.65 $Y2=2.34
r172 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=1.485 $X2=7.65 $Y2=1.66
r173 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=1.485 $X2=6.71 $Y2=2.34
r174 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=1.485 $X2=6.71 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1313_591# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 49 53 56 59 62 66
c128 62 0 1.3204e-19 $X=9.58 $Y=3.21
c129 49 0 1.97167e-19 $X=10.53 $Y=3.215
c130 33 0 1.87597e-19 $X=10.385 $Y=3.215
c131 32 0 1.97167e-19 $X=8.775 $Y=3.215
c132 31 0 1.87597e-19 $X=9.435 $Y=3.215
c133 30 0 1.97849e-19 $X=7.795 $Y=3.215
c134 29 0 9.57576e-20 $X=8.485 $Y=3.215
c135 28 0 1.97849e-19 $X=6.855 $Y=3.215
c136 27 0 1.91515e-19 $X=7.505 $Y=3.215
r137 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.53 $Y=3.215
+ $X2=10.53 $Y2=3.215
r138 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.58 $Y=3.215
+ $X2=9.58 $Y2=3.215
r139 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.63 $Y=3.215
+ $X2=8.63 $Y2=3.215
r140 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.65 $Y=3.215
+ $X2=7.65 $Y2=3.215
r141 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.71 $Y=3.215
+ $X2=6.71 $Y2=3.215
r142 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.725 $Y=3.215
+ $X2=9.58 $Y2=3.215
r143 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=10.385 $Y=3.215
+ $X2=10.53 $Y2=3.215
r144 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=10.385 $Y=3.215
+ $X2=9.725 $Y2=3.215
r145 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.775 $Y=3.215
+ $X2=8.63 $Y2=3.215
r146 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.435 $Y=3.215
+ $X2=9.58 $Y2=3.215
r147 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=9.435 $Y=3.215
+ $X2=8.775 $Y2=3.215
r148 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.795 $Y=3.215
+ $X2=7.65 $Y2=3.215
r149 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.485 $Y=3.215
+ $X2=8.63 $Y2=3.215
r150 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=8.485 $Y=3.215
+ $X2=7.795 $Y2=3.215
r151 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.855 $Y=3.215
+ $X2=6.71 $Y2=3.215
r152 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.505 $Y=3.215
+ $X2=7.65 $Y2=3.215
r153 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=7.505 $Y=3.215
+ $X2=6.855 $Y2=3.215
r154 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=8.625 $Y=3.775
+ $X2=8.625 $Y2=3.21
r155 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=7.65 $Y=3.775
+ $X2=7.65 $Y2=3.1
r156 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.65 $Y=3.775
+ $X2=7.65 $Y2=3.86
r157 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=6.71 $Y=3.775
+ $X2=6.71 $Y2=3.1
r158 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.71 $Y=3.775
+ $X2=6.71 $Y2=3.86
r159 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=3.86
+ $X2=7.65 $Y2=3.86
r160 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=8.475 $Y=3.86
+ $X2=8.625 $Y2=3.775
r161 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=8.475 $Y=3.86
+ $X2=7.815 $Y2=3.86
r162 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=3.86
+ $X2=6.71 $Y2=3.86
r163 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=3.86
+ $X2=7.65 $Y2=3.86
r164 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.485 $Y=3.86
+ $X2=6.875 $Y2=3.86
r165 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=10.375
+ $Y=3.065 $X2=10.52 $Y2=3.21
r166 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=9.435
+ $Y=3.065 $X2=9.58 $Y2=3.21
r167 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=8.515
+ $Y=3.065 $X2=8.64 $Y2=3.21
r168 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=2.955 $X2=7.65 $Y2=3.1
r169 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.505
+ $Y=2.955 $X2=7.65 $Y2=3.78
r170 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=2.955 $X2=6.71 $Y2=3.1
r171 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.565
+ $Y=2.955 $X2=6.71 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_311# 1 2 3 4 5 16 17 18 23 24 27
+ 28 29 30 31 32 33 34 47 49 50 53 58 63
c131 58 0 1.3204e-19 $X=15.26 $Y=1.7
c132 49 0 1.97849e-19 $X=18.13 $Y=2.225
c133 34 0 1.97849e-19 $X=17.335 $Y=2.225
c134 33 0 1.91515e-19 $X=17.985 $Y=2.225
c135 32 0 1.97167e-19 $X=16.355 $Y=2.225
c136 31 0 9.57576e-20 $X=17.045 $Y=2.225
c137 29 0 1.87597e-19 $X=16.065 $Y=2.225
c138 28 0 1.97167e-19 $X=14.455 $Y=2.225
c139 27 0 1.87597e-19 $X=15.115 $Y=2.225
r140 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.13 $Y=2.225
+ $X2=18.13 $Y2=2.225
r141 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.19 $Y=2.225
+ $X2=17.19 $Y2=2.225
r142 44 63 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=16.215 $Y=2.225
+ $X2=16.215 $Y2=1.7
r143 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.21 $Y=2.225
+ $X2=16.21 $Y2=2.225
r144 41 58 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=15.26 $Y=2.225
+ $X2=15.26 $Y2=1.7
r145 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.26 $Y=2.225
+ $X2=15.26 $Y2=2.225
r146 37 53 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=14.305 $Y=2.225
+ $X2=14.305 $Y2=1.73
r147 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.31 $Y=2.225
+ $X2=14.31 $Y2=2.225
r148 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.335 $Y=2.225
+ $X2=17.19 $Y2=2.225
r149 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.985 $Y=2.225
+ $X2=18.13 $Y2=2.225
r150 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=17.985 $Y=2.225
+ $X2=17.335 $Y2=2.225
r151 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.355 $Y=2.225
+ $X2=16.21 $Y2=2.225
r152 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.045 $Y=2.225
+ $X2=17.19 $Y2=2.225
r153 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=17.045 $Y=2.225
+ $X2=16.355 $Y2=2.225
r154 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.405 $Y=2.225
+ $X2=15.26 $Y2=2.225
r155 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.065 $Y=2.225
+ $X2=16.21 $Y2=2.225
r156 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=16.065 $Y=2.225
+ $X2=15.405 $Y2=2.225
r157 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.455 $Y=2.225
+ $X2=14.31 $Y2=2.225
r158 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.115 $Y=2.225
+ $X2=15.26 $Y2=2.225
r159 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=15.115 $Y=2.225
+ $X2=14.455 $Y2=2.225
r160 24 50 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=18.13 $Y=1.665
+ $X2=18.13 $Y2=2.225
r161 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.13 $Y=1.665
+ $X2=18.13 $Y2=1.58
r162 21 47 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=17.19 $Y=1.665
+ $X2=17.19 $Y2=2.225
r163 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.19 $Y=1.665
+ $X2=17.19 $Y2=1.58
r164 20 63 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=16.215 $Y=1.665
+ $X2=16.215 $Y2=1.7
r165 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.355 $Y=1.58
+ $X2=17.19 $Y2=1.58
r166 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.965 $Y=1.58
+ $X2=18.13 $Y2=1.58
r167 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=17.965 $Y=1.58
+ $X2=17.355 $Y2=1.58
r168 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=16.365 $Y=1.58
+ $X2=16.215 $Y2=1.665
r169 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.025 $Y=1.58
+ $X2=17.19 $Y2=1.58
r170 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=17.025 $Y=1.58
+ $X2=16.365 $Y2=1.58
r171 5 50 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=17.985
+ $Y=1.485 $X2=18.13 $Y2=2.34
r172 5 26 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=17.985
+ $Y=1.485 $X2=18.13 $Y2=1.66
r173 4 47 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=17.045
+ $Y=1.485 $X2=17.19 $Y2=2.34
r174 4 23 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=17.045
+ $Y=1.485 $X2=17.19 $Y2=1.66
r175 3 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.055
+ $Y=1.555 $X2=16.2 $Y2=1.7
r176 2 58 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=15.115
+ $Y=1.555 $X2=15.26 $Y2=1.7
r177 1 53 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=14.195
+ $Y=1.555 $X2=14.32 $Y2=1.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2839_613# 1 2 3 4 5 16 17 18 23 24 27
+ 28 29 30 31 32 33 34 49 53 57 61 64 67
c131 57 0 1.3204e-19 $X=15.26 $Y=3.21
c132 49 0 1.97849e-19 $X=18.13 $Y=3.215
c133 34 0 1.97849e-19 $X=17.335 $Y=3.215
c134 33 0 1.91515e-19 $X=17.985 $Y=3.215
c135 32 0 1.97167e-19 $X=16.355 $Y=3.215
c136 31 0 9.57576e-20 $X=17.045 $Y=3.215
c137 29 0 1.87597e-19 $X=16.065 $Y=3.215
c138 28 0 1.97167e-19 $X=14.455 $Y=3.215
c139 27 0 1.87597e-19 $X=15.115 $Y=3.215
r140 49 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.13 $Y=3.215
+ $X2=18.13 $Y2=3.215
r141 46 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.19 $Y=3.215
+ $X2=17.19 $Y2=3.215
r142 43 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=16.21 $Y=3.215
+ $X2=16.21 $Y2=3.215
r143 40 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=15.26 $Y=3.215
+ $X2=15.26 $Y2=3.215
r144 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.31 $Y=3.215
+ $X2=14.31 $Y2=3.215
r145 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.335 $Y=3.215
+ $X2=17.19 $Y2=3.215
r146 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.985 $Y=3.215
+ $X2=18.13 $Y2=3.215
r147 33 34 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=17.985 $Y=3.215
+ $X2=17.335 $Y2=3.215
r148 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.355 $Y=3.215
+ $X2=16.21 $Y2=3.215
r149 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.045 $Y=3.215
+ $X2=17.19 $Y2=3.215
r150 31 32 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=17.045 $Y=3.215
+ $X2=16.355 $Y2=3.215
r151 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.405 $Y=3.215
+ $X2=15.26 $Y2=3.215
r152 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=16.065 $Y=3.215
+ $X2=16.21 $Y2=3.215
r153 29 30 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=16.065 $Y=3.215
+ $X2=15.405 $Y2=3.215
r154 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.455 $Y=3.215
+ $X2=14.31 $Y2=3.215
r155 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=15.115 $Y=3.215
+ $X2=15.26 $Y2=3.215
r156 27 28 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=15.115 $Y=3.215
+ $X2=14.455 $Y2=3.215
r157 24 67 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=18.13 $Y=3.775
+ $X2=18.13 $Y2=3.1
r158 24 26 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.13 $Y=3.775
+ $X2=18.13 $Y2=3.86
r159 21 64 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=17.19 $Y=3.775
+ $X2=17.19 $Y2=3.1
r160 21 23 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.19 $Y=3.775
+ $X2=17.19 $Y2=3.86
r161 20 61 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=16.215 $Y=3.775
+ $X2=16.215 $Y2=3.21
r162 19 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.355 $Y=3.86
+ $X2=17.19 $Y2=3.86
r163 18 26 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.965 $Y=3.86
+ $X2=18.13 $Y2=3.86
r164 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=17.965 $Y=3.86
+ $X2=17.355 $Y2=3.86
r165 17 20 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=16.365 $Y=3.86
+ $X2=16.215 $Y2=3.775
r166 16 23 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.025 $Y=3.86
+ $X2=17.19 $Y2=3.86
r167 16 17 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=17.025 $Y=3.86
+ $X2=16.365 $Y2=3.86
r168 5 67 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=17.985
+ $Y=2.955 $X2=18.13 $Y2=3.1
r169 5 26 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=17.985
+ $Y=2.955 $X2=18.13 $Y2=3.78
r170 4 64 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=17.045
+ $Y=2.955 $X2=17.19 $Y2=3.1
r171 4 23 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=17.045
+ $Y=2.955 $X2=17.19 $Y2=3.78
r172 3 61 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=16.055
+ $Y=3.065 $X2=16.2 $Y2=3.21
r173 2 57 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=15.115
+ $Y=3.065 $X2=15.26 $Y2=3.21
r174 1 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=14.195
+ $Y=3.065 $X2=14.32 $Y2=3.21
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_297# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 37 41 49 59 63 68
c122 63 0 1.3204e-19 $X=22 $Y=1.7
c123 49 0 1.97167e-19 $X=22.95 $Y=2.225
c124 33 0 1.87597e-19 $X=22.805 $Y=2.225
c125 32 0 1.97167e-19 $X=21.195 $Y=2.225
c126 31 0 1.87597e-19 $X=21.855 $Y=2.225
c127 30 0 1.97849e-19 $X=20.215 $Y=2.225
c128 29 0 9.57576e-20 $X=20.905 $Y=2.225
c129 28 0 1.97849e-19 $X=19.275 $Y=2.225
c130 27 0 1.91515e-19 $X=19.925 $Y=2.225
r131 50 68 19.0153 $w=2.98e-07 $l=4.95e-07 $layer=LI1_cond $X=22.955 $Y=2.225
+ $X2=22.955 $Y2=1.73
r132 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.95 $Y=2.225
+ $X2=22.95 $Y2=2.225
r133 47 63 22.4086 $w=2.68e-07 $l=5.25e-07 $layer=LI1_cond $X=22 $Y=2.225 $X2=22
+ $Y2=1.7
r134 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22 $Y=2.225 $X2=22
+ $Y2=2.225
r135 44 59 20.1678 $w=2.98e-07 $l=5.25e-07 $layer=LI1_cond $X=21.045 $Y=2.225
+ $X2=21.045 $Y2=1.7
r136 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.05 $Y=2.225
+ $X2=21.05 $Y2=2.225
r137 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.07 $Y=2.225
+ $X2=20.07 $Y2=2.225
r138 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.13 $Y=2.225
+ $X2=19.13 $Y2=2.225
r139 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.145 $Y=2.225
+ $X2=22 $Y2=2.225
r140 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.805 $Y=2.225
+ $X2=22.95 $Y2=2.225
r141 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.805 $Y=2.225
+ $X2=22.145 $Y2=2.225
r142 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.195 $Y=2.225
+ $X2=21.05 $Y2=2.225
r143 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.855 $Y=2.225
+ $X2=22 $Y2=2.225
r144 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=21.855 $Y=2.225
+ $X2=21.195 $Y2=2.225
r145 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.215 $Y=2.225
+ $X2=20.07 $Y2=2.225
r146 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.905 $Y=2.225
+ $X2=21.05 $Y2=2.225
r147 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=20.905 $Y=2.225
+ $X2=20.215 $Y2=2.225
r148 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.275 $Y=2.225
+ $X2=19.13 $Y2=2.225
r149 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.925 $Y=2.225
+ $X2=20.07 $Y2=2.225
r150 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=19.925 $Y=2.225
+ $X2=19.275 $Y2=2.225
r151 26 59 1.34452 $w=2.98e-07 $l=3.5e-08 $layer=LI1_cond $X=21.045 $Y=1.665
+ $X2=21.045 $Y2=1.7
r152 23 41 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=20.07 $Y=1.665
+ $X2=20.07 $Y2=2.225
r153 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.07 $Y=1.665
+ $X2=20.07 $Y2=1.58
r154 20 37 19.5566 $w=3.28e-07 $l=5.6e-07 $layer=LI1_cond $X=19.13 $Y=1.665
+ $X2=19.13 $Y2=2.225
r155 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.13 $Y=1.665
+ $X2=19.13 $Y2=1.58
r156 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.235 $Y=1.58
+ $X2=20.07 $Y2=1.58
r157 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=20.895 $Y=1.58
+ $X2=21.045 $Y2=1.665
r158 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=20.895 $Y=1.58
+ $X2=20.235 $Y2=1.58
r159 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.295 $Y=1.58
+ $X2=19.13 $Y2=1.58
r160 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.905 $Y=1.58
+ $X2=20.07 $Y2=1.58
r161 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=19.905 $Y=1.58
+ $X2=19.295 $Y2=1.58
r162 5 68 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=22.795
+ $Y=1.555 $X2=22.94 $Y2=1.73
r163 4 63 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=21.855
+ $Y=1.555 $X2=22 $Y2=1.7
r164 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=20.935
+ $Y=1.555 $X2=21.06 $Y2=1.7
r165 2 41 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=19.925
+ $Y=1.485 $X2=20.07 $Y2=2.34
r166 2 25 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=19.925
+ $Y=1.485 $X2=20.07 $Y2=1.66
r167 1 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=18.985
+ $Y=1.485 $X2=19.13 $Y2=2.34
r168 1 22 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=18.985
+ $Y=1.485 $X2=19.13 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3797_591# 1 2 3 4 5 16 18 20 25 27 28
+ 29 30 31 32 33 34 49 53 56 59 62 66
c122 62 0 1.3204e-19 $X=22 $Y=3.21
c123 49 0 1.97167e-19 $X=22.95 $Y=3.215
c124 33 0 1.87597e-19 $X=22.805 $Y=3.215
c125 32 0 1.97167e-19 $X=21.195 $Y=3.215
c126 31 0 1.87597e-19 $X=21.855 $Y=3.215
c127 30 0 1.97849e-19 $X=20.215 $Y=3.215
c128 29 0 9.57576e-20 $X=20.905 $Y=3.215
c129 28 0 1.97849e-19 $X=19.275 $Y=3.215
c130 27 0 1.91515e-19 $X=19.925 $Y=3.215
r131 49 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22.95 $Y=3.215
+ $X2=22.95 $Y2=3.215
r132 46 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=22 $Y=3.215 $X2=22
+ $Y2=3.215
r133 43 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=21.05 $Y=3.215
+ $X2=21.05 $Y2=3.215
r134 40 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.07 $Y=3.215
+ $X2=20.07 $Y2=3.215
r135 36 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.13 $Y=3.215
+ $X2=19.13 $Y2=3.215
r136 34 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.145 $Y=3.215
+ $X2=22 $Y2=3.215
r137 33 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=22.805 $Y=3.215
+ $X2=22.95 $Y2=3.215
r138 33 34 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=22.805 $Y=3.215
+ $X2=22.145 $Y2=3.215
r139 32 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.195 $Y=3.215
+ $X2=21.05 $Y2=3.215
r140 31 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.855 $Y=3.215
+ $X2=22 $Y2=3.215
r141 31 32 0.81683 $w=1.4e-07 $l=6.6e-07 $layer=MET1_cond $X=21.855 $Y=3.215
+ $X2=21.195 $Y2=3.215
r142 30 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.215 $Y=3.215
+ $X2=20.07 $Y2=3.215
r143 29 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.905 $Y=3.215
+ $X2=21.05 $Y2=3.215
r144 29 30 0.853959 $w=1.4e-07 $l=6.9e-07 $layer=MET1_cond $X=20.905 $Y=3.215
+ $X2=20.215 $Y2=3.215
r145 28 36 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.275 $Y=3.215
+ $X2=19.13 $Y2=3.215
r146 27 40 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=19.925 $Y=3.215
+ $X2=20.07 $Y2=3.215
r147 27 28 0.804454 $w=1.4e-07 $l=6.5e-07 $layer=MET1_cond $X=19.925 $Y=3.215
+ $X2=19.275 $Y2=3.215
r148 26 59 21.7043 $w=2.98e-07 $l=5.65e-07 $layer=LI1_cond $X=21.045 $Y=3.775
+ $X2=21.045 $Y2=3.21
r149 23 56 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=20.07 $Y=3.775
+ $X2=20.07 $Y2=3.1
r150 23 25 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.07 $Y=3.775
+ $X2=20.07 $Y2=3.86
r151 20 53 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=19.13 $Y=3.775
+ $X2=19.13 $Y2=3.1
r152 20 22 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.13 $Y=3.775
+ $X2=19.13 $Y2=3.86
r153 19 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.235 $Y=3.86
+ $X2=20.07 $Y2=3.86
r154 18 26 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=20.895 $Y=3.86
+ $X2=21.045 $Y2=3.775
r155 18 19 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=20.895 $Y=3.86
+ $X2=20.235 $Y2=3.86
r156 17 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.295 $Y=3.86
+ $X2=19.13 $Y2=3.86
r157 16 25 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.905 $Y=3.86
+ $X2=20.07 $Y2=3.86
r158 16 17 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=19.905 $Y=3.86
+ $X2=19.295 $Y2=3.86
r159 5 66 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=22.795
+ $Y=3.065 $X2=22.94 $Y2=3.21
r160 4 62 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=21.855
+ $Y=3.065 $X2=22 $Y2=3.21
r161 3 59 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=20.935
+ $Y=3.065 $X2=21.06 $Y2=3.21
r162 2 56 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=19.925
+ $Y=2.955 $X2=20.07 $Y2=3.1
r163 2 25 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=19.925
+ $Y=2.955 $X2=20.07 $Y2=3.78
r164 1 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=18.985
+ $Y=2.955 $X2=19.13 $Y2=3.1
r165 1 22 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=18.985
+ $Y=2.955 $X2=19.13 $Y2=3.78
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%VGND 1 2 3 4 5 6 7 8 9 10 11 12 13 14
+ 15 16 17 18 19 20 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 109 111 113
+ 115 119 123 127 131 135 139 143 147 151 155 157 159 163 167 171 175 179 183
+ 187 191 195 199 203 207 211 215 219 223 227 231 233 235 239 243 247 251 253
+ 255 257 259 262 263 265 266 268 269 271 272 274 275 277 278 280 281 283 284
+ 286 287 289 290 292 293 295 296 298 299 301 302 304 305 307 308 309 310 311
+ 312 313 314 341 345 349 354 359 364 413 417 421 426 431 436 455 459 470 473
+ 476 479 482 485 488 491 494 497 500 503 506 509 512 515 519 522
r662 521 522 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=5.44
+ $X2=24.61 $Y2=5.44
r663 518 519 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.61 $Y=0
+ $X2=24.61 $Y2=0
r664 515 516 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=5.44
+ $X2=20.47 $Y2=5.44
r665 512 513 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.47 $Y=0
+ $X2=20.47 $Y2=0
r666 510 516 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=5.44
+ $X2=20.47 $Y2=5.44
r667 509 510 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.55 $Y=5.44
+ $X2=19.55 $Y2=5.44
r668 507 513 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=19.55 $Y=0
+ $X2=20.47 $Y2=0
r669 506 507 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.55 $Y=0
+ $X2=19.55 $Y2=0
r670 497 498 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=5.44
+ $X2=17.71 $Y2=5.44
r671 494 495 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=0
+ $X2=17.71 $Y2=0
r672 491 492 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=5.44
+ $X2=8.05 $Y2=5.44
r673 488 489 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r674 486 492 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=5.44
+ $X2=8.05 $Y2=5.44
r675 485 486 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=5.44
+ $X2=7.13 $Y2=5.44
r676 483 489 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r677 482 483 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r678 473 474 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=5.44
+ $X2=5.29 $Y2=5.44
r679 470 471 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r680 462 522 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=5.44
+ $X2=24.61 $Y2=5.44
r681 461 462 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=5.44
+ $X2=24.15 $Y2=5.44
r682 459 521 4.16519 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=24.28 $Y=5.44
+ $X2=24.56 $Y2=5.44
r683 459 461 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=24.28 $Y=5.44
+ $X2=24.15 $Y2=5.44
r684 458 519 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.15 $Y=0
+ $X2=24.61 $Y2=0
r685 457 458 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=24.15 $Y=0
+ $X2=24.15 $Y2=0
r686 455 518 4.16519 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=24.28 $Y=0
+ $X2=24.56 $Y2=0
r687 455 457 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=24.28 $Y=0
+ $X2=24.15 $Y2=0
r688 454 462 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=5.44
+ $X2=24.15 $Y2=5.44
r689 453 454 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=5.44
+ $X2=23.23 $Y2=5.44
r690 451 454 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=5.44
+ $X2=23.23 $Y2=5.44
r691 451 516 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.93 $Y=5.44
+ $X2=20.47 $Y2=5.44
r692 450 453 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=5.44
+ $X2=23.23 $Y2=5.44
r693 450 451 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=5.44
+ $X2=20.93 $Y2=5.44
r694 448 515 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=20.655 $Y=5.44
+ $X2=20.53 $Y2=5.44
r695 448 450 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=20.655 $Y=5.44
+ $X2=20.93 $Y2=5.44
r696 447 458 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=23.23 $Y=0
+ $X2=24.15 $Y2=0
r697 446 447 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=23.23 $Y=0
+ $X2=23.23 $Y2=0
r698 444 447 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r699 444 513 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.93 $Y=0
+ $X2=20.47 $Y2=0
r700 443 446 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=20.93 $Y=0
+ $X2=23.23 $Y2=0
r701 443 444 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=20.93 $Y=0
+ $X2=20.93 $Y2=0
r702 441 512 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=20.655 $Y=0
+ $X2=20.53 $Y2=0
r703 441 443 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=20.655 $Y=0
+ $X2=20.93 $Y2=0
r704 440 510 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=5.44
+ $X2=19.55 $Y2=5.44
r705 439 440 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.09 $Y=5.44
+ $X2=19.09 $Y2=5.44
r706 437 503 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.795 $Y=5.44
+ $X2=18.63 $Y2=5.44
r707 437 439 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.795 $Y=5.44
+ $X2=19.09 $Y2=5.44
r708 436 509 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.465 $Y=5.44
+ $X2=19.6 $Y2=5.44
r709 436 439 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=19.465 $Y=5.44
+ $X2=19.09 $Y2=5.44
r710 435 507 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=0
+ $X2=19.55 $Y2=0
r711 434 435 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=19.09 $Y=0
+ $X2=19.09 $Y2=0
r712 432 500 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.795 $Y=0
+ $X2=18.63 $Y2=0
r713 432 434 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.795 $Y=0
+ $X2=19.09 $Y2=0
r714 431 506 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.465 $Y=0
+ $X2=19.6 $Y2=0
r715 431 434 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=19.465 $Y=0
+ $X2=19.09 $Y2=0
r716 430 498 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=5.44
+ $X2=17.71 $Y2=5.44
r717 429 430 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=5.44
+ $X2=18.17 $Y2=5.44
r718 427 497 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.795 $Y=5.44
+ $X2=17.66 $Y2=5.44
r719 427 429 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=17.795 $Y=5.44
+ $X2=18.17 $Y2=5.44
r720 426 503 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=5.44
+ $X2=18.63 $Y2=5.44
r721 426 429 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.465 $Y=5.44
+ $X2=18.17 $Y2=5.44
r722 425 495 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=0
+ $X2=17.71 $Y2=0
r723 424 425 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.17 $Y=0
+ $X2=18.17 $Y2=0
r724 422 494 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.795 $Y=0
+ $X2=17.66 $Y2=0
r725 422 424 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=17.795 $Y=0
+ $X2=18.17 $Y2=0
r726 421 500 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=18.465 $Y=0
+ $X2=18.63 $Y2=0
r727 421 424 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=18.465 $Y=0
+ $X2=18.17 $Y2=0
r728 420 498 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=17.25 $Y=5.44
+ $X2=17.71 $Y2=5.44
r729 419 420 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.25 $Y=5.44
+ $X2=17.25 $Y2=5.44
r730 417 497 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.525 $Y=5.44
+ $X2=17.66 $Y2=5.44
r731 417 419 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=17.525 $Y=5.44
+ $X2=17.25 $Y2=5.44
r732 416 495 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=17.25 $Y=0
+ $X2=17.71 $Y2=0
r733 415 416 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=17.25 $Y=0
+ $X2=17.25 $Y2=0
r734 413 494 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=17.525 $Y=0
+ $X2=17.66 $Y2=0
r735 413 415 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=17.525 $Y=0
+ $X2=17.25 $Y2=0
r736 412 420 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.33 $Y=5.44
+ $X2=17.25 $Y2=5.44
r737 411 412 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=16.33 $Y=5.44
+ $X2=16.33 $Y2=5.44
r738 409 412 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=14.03 $Y=5.44
+ $X2=16.33 $Y2=5.44
r739 408 411 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=14.03 $Y=5.44
+ $X2=16.33 $Y2=5.44
r740 408 409 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.03 $Y=5.44
+ $X2=14.03 $Y2=5.44
r741 406 416 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=16.33 $Y=0
+ $X2=17.25 $Y2=0
r742 405 406 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r743 403 406 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=16.33 $Y2=0
r744 402 405 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=14.03 $Y=0
+ $X2=16.33 $Y2=0
r745 402 403 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r746 400 409 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=5.44
+ $X2=14.03 $Y2=5.44
r747 399 400 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=5.44
+ $X2=13.57 $Y2=5.44
r748 397 403 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.03 $Y2=0
r749 396 397 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r750 394 400 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=5.44
+ $X2=13.57 $Y2=5.44
r751 393 394 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=5.44
+ $X2=12.65 $Y2=5.44
r752 391 397 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.57 $Y2=0
r753 390 391 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r754 388 394 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=5.44
+ $X2=12.65 $Y2=5.44
r755 387 388 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=5.44
+ $X2=11.73 $Y2=5.44
r756 385 391 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.65 $Y2=0
r757 384 385 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r758 382 388 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=5.44
+ $X2=11.73 $Y2=5.44
r759 381 382 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=5.44
+ $X2=10.81 $Y2=5.44
r760 379 382 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=5.44
+ $X2=10.81 $Y2=5.44
r761 379 492 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=5.44
+ $X2=8.05 $Y2=5.44
r762 378 381 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.51 $Y=5.44
+ $X2=10.81 $Y2=5.44
r763 378 379 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=5.44
+ $X2=8.51 $Y2=5.44
r764 376 491 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=5.44
+ $X2=8.11 $Y2=5.44
r765 376 378 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.235 $Y=5.44
+ $X2=8.51 $Y2=5.44
r766 375 385 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.73 $Y2=0
r767 374 375 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r768 372 375 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r769 372 489 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r770 371 374 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r771 371 372 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r772 369 488 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.235 $Y=0
+ $X2=8.11 $Y2=0
r773 369 371 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=8.235 $Y=0
+ $X2=8.51 $Y2=0
r774 368 486 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=5.44
+ $X2=7.13 $Y2=5.44
r775 367 368 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=5.44
+ $X2=6.67 $Y2=5.44
r776 365 479 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=5.44
+ $X2=6.21 $Y2=5.44
r777 365 367 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.375 $Y=5.44
+ $X2=6.67 $Y2=5.44
r778 364 485 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.045 $Y=5.44
+ $X2=7.18 $Y2=5.44
r779 364 367 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.045 $Y=5.44
+ $X2=6.67 $Y2=5.44
r780 363 483 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r781 362 363 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r782 360 476 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=0
+ $X2=6.21 $Y2=0
r783 360 362 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.375 $Y=0
+ $X2=6.67 $Y2=0
r784 359 482 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=7.18 $Y2=0
r785 359 362 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=7.045 $Y=0
+ $X2=6.67 $Y2=0
r786 358 474 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=5.44
+ $X2=5.29 $Y2=5.44
r787 357 358 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=5.44
+ $X2=5.75 $Y2=5.44
r788 355 473 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.375 $Y=5.44
+ $X2=5.24 $Y2=5.44
r789 355 357 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=5.44
+ $X2=5.75 $Y2=5.44
r790 354 479 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=5.44
+ $X2=6.21 $Y2=5.44
r791 354 357 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.045 $Y=5.44
+ $X2=5.75 $Y2=5.44
r792 353 471 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r793 352 353 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r794 350 470 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.24 $Y2=0
r795 350 352 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=5.375 $Y=0
+ $X2=5.75 $Y2=0
r796 349 476 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.045 $Y=0
+ $X2=6.21 $Y2=0
r797 349 352 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.045 $Y=0
+ $X2=5.75 $Y2=0
r798 348 474 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=5.44
+ $X2=5.29 $Y2=5.44
r799 347 348 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=5.44
+ $X2=4.83 $Y2=5.44
r800 345 473 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.105 $Y=5.44
+ $X2=5.24 $Y2=5.44
r801 345 347 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.105 $Y=5.44
+ $X2=4.83 $Y2=5.44
r802 344 471 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r803 343 344 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r804 341 470 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=5.105 $Y=0
+ $X2=5.24 $Y2=0
r805 341 343 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=5.105 $Y=0
+ $X2=4.83 $Y2=0
r806 340 348 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=5.44
+ $X2=4.83 $Y2=5.44
r807 339 340 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=5.44
+ $X2=3.91 $Y2=5.44
r808 337 340 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=5.44
+ $X2=3.91 $Y2=5.44
r809 336 339 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=5.44
+ $X2=3.91 $Y2=5.44
r810 336 337 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=5.44
+ $X2=1.61 $Y2=5.44
r811 334 344 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r812 333 334 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r813 331 334 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=1.61 $Y=0
+ $X2=3.91 $Y2=0
r814 330 333 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=1.61 $Y=0
+ $X2=3.91 $Y2=0
r815 330 331 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r816 328 337 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=5.44
+ $X2=1.61 $Y2=5.44
r817 327 328 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=5.44
+ $X2=1.15 $Y2=5.44
r818 325 467 4.16519 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=0.56 $Y=5.44
+ $X2=0.28 $Y2=5.44
r819 325 327 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.56 $Y=5.44
+ $X2=1.15 $Y2=5.44
r820 324 331 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r821 323 324 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r822 321 464 4.16519 $w=1.7e-07 $l=2.8e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=0.28
+ $Y2=0
r823 321 323 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=0.56 $Y=0 $X2=1.15
+ $Y2=0
r824 314 440 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=5.44
+ $X2=19.09 $Y2=5.44
r825 314 430 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=5.44
+ $X2=18.17 $Y2=5.44
r826 314 503 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.63 $Y=5.44
+ $X2=18.63 $Y2=5.44
r827 313 435 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=0
+ $X2=19.09 $Y2=0
r828 313 425 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.63 $Y=0
+ $X2=18.17 $Y2=0
r829 313 500 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.63 $Y=0
+ $X2=18.63 $Y2=0
r830 312 368 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=5.44
+ $X2=6.67 $Y2=5.44
r831 312 358 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=5.44
+ $X2=5.75 $Y2=5.44
r832 312 479 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=5.44
+ $X2=6.21 $Y2=5.44
r833 311 363 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r834 311 353 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r835 311 476 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r836 310 328 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=5.44
+ $X2=1.15 $Y2=5.44
r837 310 467 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=5.44
+ $X2=0.23 $Y2=5.44
r838 309 324 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r839 309 464 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r840 307 453 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=23.36 $Y=5.44
+ $X2=23.23 $Y2=5.44
r841 307 308 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=23.36 $Y=5.44
+ $X2=23.505 $Y2=5.44
r842 306 461 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=23.65 $Y=5.44
+ $X2=24.15 $Y2=5.44
r843 306 308 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=23.65 $Y=5.44
+ $X2=23.505 $Y2=5.44
r844 304 446 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=23.36 $Y=0
+ $X2=23.23 $Y2=0
r845 304 305 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=23.36 $Y=0
+ $X2=23.505 $Y2=0
r846 303 457 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=23.65 $Y=0
+ $X2=24.15 $Y2=0
r847 303 305 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=23.65 $Y=0
+ $X2=23.505 $Y2=0
r848 301 411 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.605 $Y=5.44
+ $X2=16.33 $Y2=5.44
r849 301 302 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.605 $Y=5.44
+ $X2=16.73 $Y2=5.44
r850 300 419 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=16.855 $Y=5.44
+ $X2=17.25 $Y2=5.44
r851 300 302 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.855 $Y=5.44
+ $X2=16.73 $Y2=5.44
r852 298 405 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=16.605 $Y=0
+ $X2=16.33 $Y2=0
r853 298 299 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.605 $Y=0
+ $X2=16.73 $Y2=0
r854 297 415 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=17.25 $Y2=0
r855 297 299 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.855 $Y=0
+ $X2=16.73 $Y2=0
r856 295 399 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=13.61 $Y=5.44
+ $X2=13.57 $Y2=5.44
r857 295 296 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.61 $Y=5.44
+ $X2=13.755 $Y2=5.44
r858 294 408 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=13.9 $Y=5.44
+ $X2=14.03 $Y2=5.44
r859 294 296 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.9 $Y=5.44
+ $X2=13.755 $Y2=5.44
r860 292 396 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=13.61 $Y=0
+ $X2=13.57 $Y2=0
r861 292 293 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.61 $Y=0
+ $X2=13.755 $Y2=0
r862 291 402 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=13.9 $Y=0
+ $X2=14.03 $Y2=0
r863 291 293 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=13.9 $Y=0
+ $X2=13.755 $Y2=0
r864 289 393 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=12.69 $Y=5.44
+ $X2=12.65 $Y2=5.44
r865 289 290 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.69 $Y=5.44
+ $X2=12.835 $Y2=5.44
r866 288 399 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.98 $Y=5.44
+ $X2=13.57 $Y2=5.44
r867 288 290 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.98 $Y=5.44
+ $X2=12.835 $Y2=5.44
r868 286 390 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=12.69 $Y=0
+ $X2=12.65 $Y2=0
r869 286 287 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.69 $Y=0
+ $X2=12.835 $Y2=0
r870 285 396 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=12.98 $Y=0
+ $X2=13.57 $Y2=0
r871 285 287 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.98 $Y=0
+ $X2=12.835 $Y2=0
r872 283 387 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.86 $Y=5.44
+ $X2=11.73 $Y2=5.44
r873 283 284 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.86 $Y=5.44
+ $X2=12.005 $Y2=5.44
r874 282 393 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=12.15 $Y=5.44
+ $X2=12.65 $Y2=5.44
r875 282 284 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.15 $Y=5.44
+ $X2=12.005 $Y2=5.44
r876 280 384 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=11.86 $Y=0
+ $X2=11.73 $Y2=0
r877 280 281 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.86 $Y=0
+ $X2=12.005 $Y2=0
r878 279 390 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=12.65 $Y2=0
r879 279 281 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=12.15 $Y=0
+ $X2=12.005 $Y2=0
r880 277 381 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=10.94 $Y=5.44
+ $X2=10.81 $Y2=5.44
r881 277 278 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.94 $Y=5.44
+ $X2=11.085 $Y2=5.44
r882 276 387 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.23 $Y=5.44
+ $X2=11.73 $Y2=5.44
r883 276 278 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.23 $Y=5.44
+ $X2=11.085 $Y2=5.44
r884 274 374 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=10.94 $Y=0
+ $X2=10.81 $Y2=0
r885 274 275 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=10.94 $Y=0
+ $X2=11.085 $Y2=0
r886 273 384 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=11.23 $Y=0
+ $X2=11.73 $Y2=0
r887 273 275 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=11.23 $Y=0
+ $X2=11.085 $Y2=0
r888 271 339 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=5.44
+ $X2=3.91 $Y2=5.44
r889 271 272 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=5.44
+ $X2=4.31 $Y2=5.44
r890 270 347 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=5.44
+ $X2=4.83 $Y2=5.44
r891 270 272 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=5.44
+ $X2=4.31 $Y2=5.44
r892 268 333 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=3.91 $Y2=0
r893 268 269 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.185 $Y=0
+ $X2=4.31 $Y2=0
r894 267 343 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.83 $Y2=0
r895 267 269 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.435 $Y=0
+ $X2=4.31 $Y2=0
r896 265 327 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.19 $Y=5.44
+ $X2=1.15 $Y2=5.44
r897 265 266 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.19 $Y=5.44
+ $X2=1.335 $Y2=5.44
r898 264 336 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.48 $Y=5.44
+ $X2=1.61 $Y2=5.44
r899 264 266 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.48 $Y=5.44
+ $X2=1.335 $Y2=5.44
r900 262 323 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=1.19 $Y=0 $X2=1.15
+ $Y2=0
r901 262 263 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.19 $Y=0
+ $X2=1.335 $Y2=0
r902 261 330 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=1.48 $Y=0
+ $X2=1.61 $Y2=0
r903 261 263 7.85057 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.48 $Y=0
+ $X2=1.335 $Y2=0
r904 257 521 3.27265 $w=2.9e-07 $l=1.72337e-07 $layer=LI1_cond $X=24.425
+ $Y=5.355 $X2=24.56 $Y2=5.44
r905 257 259 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=24.425 $Y=5.355
+ $X2=24.425 $Y2=4.995
r906 253 518 3.27265 $w=2.9e-07 $l=1.72337e-07 $layer=LI1_cond $X=24.425
+ $Y=0.085 $X2=24.56 $Y2=0
r907 253 255 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=24.425 $Y=0.085
+ $X2=24.425 $Y2=0.445
r908 249 308 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=23.505 $Y=5.355
+ $X2=23.505 $Y2=5.44
r909 249 251 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=23.505 $Y=5.355
+ $X2=23.505 $Y2=4.995
r910 245 305 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=23.505 $Y=0.085
+ $X2=23.505 $Y2=0
r911 245 247 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=23.505 $Y=0.085
+ $X2=23.505 $Y2=0.445
r912 241 515 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=20.53 $Y=5.355
+ $X2=20.53 $Y2=5.44
r913 241 243 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=20.53 $Y=5.355
+ $X2=20.53 $Y2=5.06
r914 237 512 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=20.53 $Y=0.085
+ $X2=20.53 $Y2=0
r915 237 239 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=20.53 $Y=0.085
+ $X2=20.53 $Y2=0.38
r916 236 509 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.735 $Y=5.44
+ $X2=19.6 $Y2=5.44
r917 235 515 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=20.405 $Y=5.44
+ $X2=20.53 $Y2=5.44
r918 235 236 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=20.405 $Y=5.44
+ $X2=19.735 $Y2=5.44
r919 234 506 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=19.735 $Y=0
+ $X2=19.6 $Y2=0
r920 233 512 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=20.405 $Y=0
+ $X2=20.53 $Y2=0
r921 233 234 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=20.405 $Y=0
+ $X2=19.735 $Y2=0
r922 229 509 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.6 $Y=5.355
+ $X2=19.6 $Y2=5.44
r923 229 231 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=19.6 $Y=5.355
+ $X2=19.6 $Y2=5.06
r924 225 506 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=19.6 $Y=0.085
+ $X2=19.6 $Y2=0
r925 225 227 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=19.6 $Y=0.085
+ $X2=19.6 $Y2=0.38
r926 221 503 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.63 $Y=5.355
+ $X2=18.63 $Y2=5.44
r927 221 223 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=18.63 $Y=5.355
+ $X2=18.63 $Y2=4.72
r928 217 500 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.63 $Y=0.085
+ $X2=18.63 $Y2=0
r929 217 219 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=18.63 $Y=0.085
+ $X2=18.63 $Y2=0.38
r930 213 497 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.66 $Y=5.355
+ $X2=17.66 $Y2=5.44
r931 213 215 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.66 $Y=5.355
+ $X2=17.66 $Y2=5.06
r932 209 494 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=17.66 $Y=0.085
+ $X2=17.66 $Y2=0
r933 209 211 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=17.66 $Y=0.085
+ $X2=17.66 $Y2=0.38
r934 205 302 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.73 $Y=5.355
+ $X2=16.73 $Y2=5.44
r935 205 207 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=16.73 $Y=5.355
+ $X2=16.73 $Y2=5.06
r936 201 299 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.73 $Y=0.085
+ $X2=16.73 $Y2=0
r937 201 203 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=16.73 $Y=0.085
+ $X2=16.73 $Y2=0.38
r938 197 296 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=5.355
+ $X2=13.755 $Y2=5.44
r939 197 199 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=13.755 $Y=5.355
+ $X2=13.755 $Y2=4.995
r940 193 293 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0
r941 193 195 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=13.755 $Y=0.085
+ $X2=13.755 $Y2=0.445
r942 189 290 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=5.355
+ $X2=12.835 $Y2=5.44
r943 189 191 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=12.835 $Y=5.355
+ $X2=12.835 $Y2=4.995
r944 185 287 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.835 $Y=0.085
+ $X2=12.835 $Y2=0
r945 185 187 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=12.835 $Y=0.085
+ $X2=12.835 $Y2=0.445
r946 181 284 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.005 $Y=5.355
+ $X2=12.005 $Y2=5.44
r947 181 183 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=12.005 $Y=5.355
+ $X2=12.005 $Y2=4.995
r948 177 281 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=12.005 $Y=0.085
+ $X2=12.005 $Y2=0
r949 177 179 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=12.005 $Y=0.085
+ $X2=12.005 $Y2=0.445
r950 173 278 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.085 $Y=5.355
+ $X2=11.085 $Y2=5.44
r951 173 175 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=11.085 $Y=5.355
+ $X2=11.085 $Y2=4.995
r952 169 275 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=11.085 $Y=0.085
+ $X2=11.085 $Y2=0
r953 169 171 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=11.085 $Y=0.085
+ $X2=11.085 $Y2=0.445
r954 165 491 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=5.355
+ $X2=8.11 $Y2=5.44
r955 165 167 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.11 $Y=5.355
+ $X2=8.11 $Y2=5.06
r956 161 488 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0
r957 161 163 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=8.11 $Y=0.085
+ $X2=8.11 $Y2=0.38
r958 160 485 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.315 $Y=5.44
+ $X2=7.18 $Y2=5.44
r959 159 491 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.985 $Y=5.44
+ $X2=8.11 $Y2=5.44
r960 159 160 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.985 $Y=5.44
+ $X2=7.315 $Y2=5.44
r961 158 482 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=7.315 $Y=0
+ $X2=7.18 $Y2=0
r962 157 488 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.985 $Y=0
+ $X2=8.11 $Y2=0
r963 157 158 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=7.985 $Y=0
+ $X2=7.315 $Y2=0
r964 153 485 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=5.355
+ $X2=7.18 $Y2=5.44
r965 153 155 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.18 $Y=5.355
+ $X2=7.18 $Y2=5.06
r966 149 482 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0
r967 149 151 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.18 $Y=0.085
+ $X2=7.18 $Y2=0.38
r968 145 479 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=5.355
+ $X2=6.21 $Y2=5.44
r969 145 147 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=6.21 $Y=5.355
+ $X2=6.21 $Y2=4.72
r970 141 476 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.21 $Y=0.085
+ $X2=6.21 $Y2=0
r971 141 143 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=6.21 $Y=0.085
+ $X2=6.21 $Y2=0.38
r972 137 473 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=5.355
+ $X2=5.24 $Y2=5.44
r973 137 139 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.24 $Y=5.355
+ $X2=5.24 $Y2=5.06
r974 133 470 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.24 $Y=0.085
+ $X2=5.24 $Y2=0
r975 133 135 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.24 $Y=0.085
+ $X2=5.24 $Y2=0.38
r976 129 272 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=5.355
+ $X2=4.31 $Y2=5.44
r977 129 131 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.31 $Y=5.355
+ $X2=4.31 $Y2=5.06
r978 125 269 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0
r979 125 127 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=4.31 $Y=0.085
+ $X2=4.31 $Y2=0.38
r980 121 266 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=5.355
+ $X2=1.335 $Y2=5.44
r981 121 123 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.335 $Y=5.355
+ $X2=1.335 $Y2=4.995
r982 117 263 0.489042 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.335 $Y=0.085
+ $X2=1.335 $Y2=0
r983 117 119 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=1.335 $Y=0.085
+ $X2=1.335 $Y2=0.445
r984 113 467 3.27265 $w=2.9e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.415 $Y=5.355
+ $X2=0.28 $Y2=5.44
r985 113 115 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.415 $Y=5.355
+ $X2=0.415 $Y2=4.995
r986 109 464 3.27265 $w=2.9e-07 $l=1.72337e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.28 $Y2=0
r987 109 111 14.3062 $w=2.88e-07 $l=3.6e-07 $layer=LI1_cond $X=0.415 $Y=0.085
+ $X2=0.415 $Y2=0.445
r988 36 259 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=24.27
+ $Y=4.785 $X2=24.405 $Y2=4.995
r989 35 255 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=24.27
+ $Y=0.235 $X2=24.405 $Y2=0.445
r990 34 251 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=23.44
+ $Y=4.785 $X2=23.565 $Y2=4.995
r991 33 247 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=23.44
+ $Y=0.235 $X2=23.565 $Y2=0.445
r992 32 243 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=20.355
+ $Y=4.555 $X2=20.49 $Y2=5.06
r993 31 239 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=20.355
+ $Y=0.235 $X2=20.49 $Y2=0.38
r994 30 231 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=19.415
+ $Y=4.555 $X2=19.6 $Y2=5.06
r995 29 227 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=19.415
+ $Y=0.235 $X2=19.6 $Y2=0.38
r996 28 223 91 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=2 $X=18.415
+ $Y=4.555 $X2=18.63 $Y2=4.72
r997 27 219 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=18.415
+ $Y=0.235 $X2=18.63 $Y2=0.38
r998 26 215 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=17.475
+ $Y=4.555 $X2=17.66 $Y2=5.06
r999 25 211 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=17.475
+ $Y=0.235 $X2=17.66 $Y2=0.38
r1000 24 207 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1
+ $X=16.645 $Y=4.555 $X2=16.77 $Y2=5.06
r1001 23 203 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1
+ $X=16.645 $Y=0.235 $X2=16.77 $Y2=0.38
r1002 22 199 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=13.56
+ $Y=4.785 $X2=13.695 $Y2=4.995
r1003 21 195 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=13.56
+ $Y=0.235 $X2=13.695 $Y2=0.445
r1004 20 191 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.73
+ $Y=4.785 $X2=12.855 $Y2=4.995
r1005 19 187 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=12.73
+ $Y=0.235 $X2=12.855 $Y2=0.445
r1006 18 183 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=11.85
+ $Y=4.785 $X2=11.985 $Y2=4.995
r1007 17 179 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=11.85
+ $Y=0.235 $X2=11.985 $Y2=0.445
r1008 16 175 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.02
+ $Y=4.785 $X2=11.145 $Y2=4.995
r1009 15 171 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=11.02
+ $Y=0.235 $X2=11.145 $Y2=0.445
r1010 14 167 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=7.935
+ $Y=4.555 $X2=8.07 $Y2=5.06
r1011 13 163 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.935
+ $Y=0.235 $X2=8.07 $Y2=0.38
r1012 12 155 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=4.555 $X2=7.18 $Y2=5.06
r1013 11 151 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.995
+ $Y=0.235 $X2=7.18 $Y2=0.38
r1014 10 147 91 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=4.555 $X2=6.21 $Y2=4.72
r1015 9 143 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.235 $X2=6.21 $Y2=0.38
r1016 8 139 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=4.555 $X2=5.24 $Y2=5.06
r1017 7 135 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.24 $Y2=0.38
r1018 6 131 182 $w=1.7e-07 $l=5.64048e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=4.555 $X2=4.35 $Y2=5.06
r1019 5 127 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.235 $X2=4.35 $Y2=0.38
r1020 4 123 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=4.785 $X2=1.275 $Y2=4.995
r1021 3 119 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.14
+ $Y=0.235 $X2=1.275 $Y2=0.445
r1022 2 115 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=4.785 $X2=0.435 $Y2=4.995
r1023 1 111 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.31
+ $Y=0.235 $X2=0.435 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=5.71 $Y=0.715
+ $X2=5.71 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=0.8
+ $X2=4.77 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.545 $Y=0.8
+ $X2=5.71 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.545 $Y=0.8
+ $X2=4.935 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.77 $Y=0.715
+ $X2=4.77 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.77 $Y=0.715
+ $X2=4.77 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=0.8
+ $X2=4.77 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.605 $Y=0.8
+ $X2=4.015 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.88 $Y=0.715
+ $X2=4.015 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.88 $Y=0.715
+ $X2=3.88 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=0.425
+ $X2=3.88 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=0.34
+ $X2=2.99 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.745 $Y=0.34
+ $X2=3.88 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.745 $Y=0.34
+ $X2=3.075 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=0.425
+ $X2=2.99 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=0.425
+ $X2=2.99 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.99 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.905 $Y=0.34
+ $X2=2.235 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.11 $Y=0.425
+ $X2=2.235 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=0.425
+ $X2=2.11 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=4.635
+ $Y=0.235 $X2=4.77 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=0.33 $X2=3.83 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=0.33 $X2=2.99 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.33 $X2=2.15 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_405_918# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.935 $Y=4.64
+ $X2=4.77 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.545 $Y=4.64
+ $X2=5.71 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.545 $Y=4.64
+ $X2=4.935 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.605 $Y=4.64
+ $X2=4.77 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=4.605 $Y=4.64
+ $X2=4.015 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.88 $Y=5.015
+ $X2=3.88 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.88 $Y=4.725
+ $X2=4.015 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=3.88 $Y=4.725
+ $X2=3.88 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.075 $Y=5.1 $X2=2.99
+ $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.745 $Y=5.1
+ $X2=3.88 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.745 $Y=5.1
+ $X2=3.075 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.99 $Y=5.015
+ $X2=2.99 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.99 $Y=5.015
+ $X2=2.99 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.905 $Y=5.1 $X2=2.99
+ $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.905 $Y=5.1
+ $X2=2.235 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.11 $Y=5.015
+ $X2=2.235 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=2.11 $Y=5.015
+ $X2=2.11 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=5.575
+ $Y=4.555 $X2=5.71 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=4.635
+ $Y=4.555 $X2=4.77 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.695
+ $Y=4.59 $X2=3.83 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=2.855
+ $Y=4.59 $X2=2.99 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=4.59 $X2=2.15 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=10.27 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=10.31 $Y=0.425
+ $X2=10.31 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=0.34
+ $X2=9.43 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=10.31 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.185 $Y=0.34
+ $X2=9.515 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.43 $Y=0.425
+ $X2=9.43 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=9.43 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.345 $Y=0.34
+ $X2=8.675 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.54 $Y=0.715
+ $X2=8.54 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.54 $Y=0.425
+ $X2=8.675 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.54 $Y=0.425
+ $X2=8.54 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=0.8
+ $X2=7.65 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.405 $Y=0.8
+ $X2=8.54 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.405 $Y=0.8
+ $X2=7.815 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.65 $Y=0.715
+ $X2=7.65 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=7.65 $Y=0.715
+ $X2=7.65 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=0.8
+ $X2=7.65 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.485 $Y=0.8
+ $X2=6.875 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.71 $Y=0.715
+ $X2=6.875 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.71 $Y=0.715
+ $X2=6.71 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=0.33 $X2=10.27 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=0.33 $X2=9.43 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=0.33 $X2=8.59 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=7.515
+ $Y=0.235 $X2=7.65 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=0.235 $X2=6.71 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_1315_911# 1 2 3 4 5 18 22 27 28 29 32
+ 34 38 41 43 44
c79 38 0 1.10627e-19 $X=10.27 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=10.31 $Y=5.015
+ $X2=10.31 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.515 $Y=5.1 $X2=9.43
+ $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=10.185 $Y=5.1
+ $X2=10.31 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.185 $Y=5.1
+ $X2=9.515 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.43 $Y=5.015
+ $X2=9.43 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=9.43 $Y=5.015
+ $X2=9.43 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.345 $Y=5.1 $X2=9.43
+ $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=9.345 $Y=5.1
+ $X2=8.675 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.54 $Y=5.015
+ $X2=8.675 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=8.54 $Y=5.015
+ $X2=8.54 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.54 $Y=4.725
+ $X2=8.54 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.815 $Y=4.64
+ $X2=7.65 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=8.405 $Y=4.64
+ $X2=8.54 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=8.405 $Y=4.64
+ $X2=7.815 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.875 $Y=4.64
+ $X2=6.71 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.485 $Y=4.64
+ $X2=7.65 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=7.485 $Y=4.64
+ $X2=6.875 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=10.135
+ $Y=4.59 $X2=10.27 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.295
+ $Y=4.59 $X2=9.43 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=8.465
+ $Y=4.59 $X2=8.59 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=7.515
+ $Y=4.555 $X2=7.65 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=4.555 $X2=6.71 $Y2=4.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_66# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
r84 40 42 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=18.13 $Y=0.715
+ $X2=18.13 $Y2=0.38
r85 39 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.355 $Y=0.8
+ $X2=17.19 $Y2=0.8
r86 38 40 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=17.965 $Y=0.8
+ $X2=18.13 $Y2=0.715
r87 38 39 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=17.965 $Y=0.8
+ $X2=17.355 $Y2=0.8
r88 34 45 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=17.19 $Y=0.715
+ $X2=17.19 $Y2=0.8
r89 34 36 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=17.19 $Y=0.715
+ $X2=17.19 $Y2=0.38
r90 32 45 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.025 $Y=0.8
+ $X2=17.19 $Y2=0.8
r91 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=17.025 $Y=0.8
+ $X2=16.435 $Y2=0.8
r92 29 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.3 $Y=0.715
+ $X2=16.435 $Y2=0.8
r93 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=16.3 $Y=0.715
+ $X2=16.3 $Y2=0.59
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.3 $Y=0.425
+ $X2=16.3 $Y2=0.59
r95 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.495 $Y=0.34
+ $X2=15.41 $Y2=0.34
r96 26 28 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.165 $Y=0.34
+ $X2=16.3 $Y2=0.425
r97 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.165 $Y=0.34
+ $X2=15.495 $Y2=0.34
r98 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.41 $Y=0.425
+ $X2=15.41 $Y2=0.34
r99 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.41 $Y=0.425
+ $X2=15.41 $Y2=0.59
r100 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.325 $Y=0.34
+ $X2=15.41 $Y2=0.34
r101 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=15.325 $Y=0.34
+ $X2=14.655 $Y2=0.34
r102 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=14.53 $Y=0.425
+ $X2=14.655 $Y2=0.34
r103 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=14.53 $Y=0.425
+ $X2=14.53 $Y2=0.59
r104 5 42 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=17.995
+ $Y=0.235 $X2=18.13 $Y2=0.38
r105 4 36 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=17.055
+ $Y=0.235 $X2=17.19 $Y2=0.38
r106 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.115
+ $Y=0.33 $X2=16.25 $Y2=0.59
r107 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=15.275
+ $Y=0.33 $X2=15.41 $Y2=0.59
r108 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=14.445
+ $Y=0.33 $X2=14.57 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_2889_918# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 40 42 44
r82 37 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.355 $Y=4.64
+ $X2=17.19 $Y2=4.64
r83 36 44 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.965 $Y=4.64
+ $X2=18.13 $Y2=4.64
r84 36 37 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=17.965 $Y=4.64
+ $X2=17.355 $Y2=4.64
r85 32 42 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=17.025 $Y=4.64
+ $X2=17.19 $Y2=4.64
r86 32 33 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=17.025 $Y=4.64
+ $X2=16.435 $Y2=4.64
r87 29 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=16.3 $Y=5.015
+ $X2=16.3 $Y2=4.85
r88 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.3 $Y=4.725
+ $X2=16.435 $Y2=4.64
r89 28 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=16.3 $Y=4.725
+ $X2=16.3 $Y2=4.85
r90 27 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.495 $Y=5.1
+ $X2=15.41 $Y2=5.1
r91 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=16.165 $Y=5.1
+ $X2=16.3 $Y2=5.015
r92 26 27 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=16.165 $Y=5.1
+ $X2=15.495 $Y2=5.1
r93 22 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.41 $Y=5.015
+ $X2=15.41 $Y2=5.1
r94 22 24 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=15.41 $Y=5.015
+ $X2=15.41 $Y2=4.85
r95 20 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=15.325 $Y=5.1
+ $X2=15.41 $Y2=5.1
r96 20 21 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=15.325 $Y=5.1
+ $X2=14.655 $Y2=5.1
r97 16 21 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=14.53 $Y=5.015
+ $X2=14.655 $Y2=5.1
r98 16 18 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=14.53 $Y=5.015
+ $X2=14.53 $Y2=4.85
r99 5 44 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=17.995
+ $Y=4.555 $X2=18.13 $Y2=4.72
r100 4 42 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=17.055
+ $Y=4.555 $X2=17.19 $Y2=4.72
r101 3 31 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.115
+ $Y=4.59 $X2=16.25 $Y2=4.85
r102 2 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=15.275
+ $Y=4.59 $X2=15.41 $Y2=4.85
r103 1 18 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=14.445
+ $Y=4.59 $X2=14.57 $Y2=4.85
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_47# 1 2 3 4 5 18 20 21 24 26 31
+ 32 33 36 38 42 44 45
c83 42 0 1.10627e-19 $X=22.69 $Y=0.59
r84 40 42 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=22.73 $Y=0.425
+ $X2=22.73 $Y2=0.59
r85 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.935 $Y=0.34
+ $X2=21.85 $Y2=0.34
r86 38 40 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=22.605 $Y=0.34
+ $X2=22.73 $Y2=0.425
r87 38 39 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.605 $Y=0.34
+ $X2=21.935 $Y2=0.34
r88 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.85 $Y=0.425
+ $X2=21.85 $Y2=0.34
r89 34 36 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=21.85 $Y=0.425
+ $X2=21.85 $Y2=0.59
r90 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.765 $Y=0.34
+ $X2=21.85 $Y2=0.34
r91 32 33 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=21.765 $Y=0.34
+ $X2=21.095 $Y2=0.34
r92 29 31 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=20.96 $Y=0.715
+ $X2=20.96 $Y2=0.59
r93 28 33 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=20.96 $Y=0.425
+ $X2=21.095 $Y2=0.34
r94 28 31 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=20.96 $Y=0.425
+ $X2=20.96 $Y2=0.59
r95 27 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.235 $Y=0.8
+ $X2=20.07 $Y2=0.8
r96 26 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=20.825 $Y=0.8
+ $X2=20.96 $Y2=0.715
r97 26 27 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=20.825 $Y=0.8
+ $X2=20.235 $Y2=0.8
r98 22 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.07 $Y=0.715
+ $X2=20.07 $Y2=0.8
r99 22 24 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=20.07 $Y=0.715
+ $X2=20.07 $Y2=0.38
r100 20 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.905 $Y=0.8
+ $X2=20.07 $Y2=0.8
r101 20 21 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=19.905 $Y=0.8
+ $X2=19.295 $Y2=0.8
r102 16 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=19.13 $Y=0.715
+ $X2=19.295 $Y2=0.8
r103 16 18 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=19.13 $Y=0.715
+ $X2=19.13 $Y2=0.38
r104 5 42 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.555
+ $Y=0.33 $X2=22.69 $Y2=0.59
r105 4 36 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=21.715
+ $Y=0.33 $X2=21.85 $Y2=0.59
r106 3 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=20.885
+ $Y=0.33 $X2=21.01 $Y2=0.59
r107 2 24 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=19.935
+ $Y=0.235 $X2=20.07 $Y2=0.38
r108 1 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=18.995
+ $Y=0.235 $X2=19.13 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_4%A_3799_911# 1 2 3 4 5 18 22 27 28 29 32
+ 34 38 41 43 44
c79 38 0 1.10627e-19 $X=22.69 $Y=4.85
r80 36 38 7.60612 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=22.73 $Y=5.015
+ $X2=22.73 $Y2=4.85
r81 35 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.935 $Y=5.1
+ $X2=21.85 $Y2=5.1
r82 34 36 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=22.605 $Y=5.1
+ $X2=22.73 $Y2=5.015
r83 34 35 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=22.605 $Y=5.1
+ $X2=21.935 $Y2=5.1
r84 30 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.85 $Y=5.015
+ $X2=21.85 $Y2=5.1
r85 30 32 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=21.85 $Y=5.015
+ $X2=21.85 $Y2=4.85
r86 28 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=21.765 $Y=5.1
+ $X2=21.85 $Y2=5.1
r87 28 29 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=21.765 $Y=5.1
+ $X2=21.095 $Y2=5.1
r88 25 29 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=20.96 $Y=5.015
+ $X2=21.095 $Y2=5.1
r89 25 27 7.04271 $w=2.68e-07 $l=1.65e-07 $layer=LI1_cond $X=20.96 $Y=5.015
+ $X2=20.96 $Y2=4.85
r90 24 27 5.33538 $w=2.68e-07 $l=1.25e-07 $layer=LI1_cond $X=20.96 $Y=4.725
+ $X2=20.96 $Y2=4.85
r91 23 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=20.235 $Y=4.64
+ $X2=20.07 $Y2=4.64
r92 22 24 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=20.825 $Y=4.64
+ $X2=20.96 $Y2=4.725
r93 22 23 38.492 $w=1.68e-07 $l=5.9e-07 $layer=LI1_cond $X=20.825 $Y=4.64
+ $X2=20.235 $Y2=4.64
r94 19 41 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.295 $Y=4.64
+ $X2=19.13 $Y2=4.64
r95 18 43 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=19.905 $Y=4.64
+ $X2=20.07 $Y2=4.64
r96 18 19 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=19.905 $Y=4.64
+ $X2=19.295 $Y2=4.64
r97 5 38 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.555
+ $Y=4.59 $X2=22.69 $Y2=4.85
r98 4 32 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=21.715
+ $Y=4.59 $X2=21.85 $Y2=4.85
r99 3 27 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=20.885
+ $Y=4.59 $X2=21.01 $Y2=4.85
r100 2 43 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=19.935
+ $Y=4.555 $X2=20.07 $Y2=4.72
r101 1 41 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=18.995
+ $Y=4.555 $X2=19.13 $Y2=4.72
.ends

