# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o21a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.760000 0.990000 4.115000 1.495000 ;
        RECT 3.760000 1.495000 5.880000 1.705000 ;
        RECT 5.410000 0.995000 5.880000 1.495000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.420000 0.995000 5.070000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.735000 1.075000 3.485000 1.615000 ;
    END
  END B1
  PIN X
    ANTENNADIFFAREA  1.029000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.635000 1.865000 0.805000 ;
        RECT 0.090000 0.805000 0.350000 1.530000 ;
        RECT 0.090000 1.530000 2.155000 1.700000 ;
        RECT 0.645000 0.615000 1.865000 0.635000 ;
        RECT 1.015000 1.700000 1.205000 2.465000 ;
        RECT 1.975000 1.700000 2.155000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  0.085000 0.425000 0.465000 ;
      RECT 0.415000  1.870000 0.795000 2.635000 ;
      RECT 0.520000  0.995000 2.565000 1.335000 ;
      RECT 1.055000  0.085000 1.385000 0.445000 ;
      RECT 1.375000  1.870000 1.755000 2.635000 ;
      RECT 2.015000  0.085000 2.345000 0.465000 ;
      RECT 2.315000  0.655000 3.385000 0.870000 ;
      RECT 2.315000  0.870000 2.565000 0.995000 ;
      RECT 2.325000  1.335000 2.565000 1.830000 ;
      RECT 2.325000  1.830000 3.195000 1.875000 ;
      RECT 2.325000  1.875000 4.875000 2.085000 ;
      RECT 2.335000  2.255000 2.735000 2.635000 ;
      RECT 2.585000  0.255000 3.885000 0.485000 ;
      RECT 2.955000  2.085000 4.875000 2.105000 ;
      RECT 2.955000  2.105000 3.195000 2.465000 ;
      RECT 3.515000  2.275000 3.845000 2.635000 ;
      RECT 3.555000  0.485000 3.885000 0.615000 ;
      RECT 3.555000  0.615000 5.835000 0.785000 ;
      RECT 4.055000  0.085000 4.395000 0.445000 ;
      RECT 4.495000  2.105000 4.875000 2.445000 ;
      RECT 4.975000  0.085000 5.355000 0.445000 ;
      RECT 5.455000  1.935000 5.865000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21a_4
END LIBRARY
