* NGSPICE file created from sky130_fd_sc_hdll__and3_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__and3_2 A B C VGND VNB VPB VPWR X
M1000 VGND a_29_311# X VNB nshort w=650000u l=150000u
+  ad=5.093e+11p pd=4.31e+06u as=2.21e+11p ps=1.98e+06u
M1001 VGND C a_194_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.281e+11p ps=1.45e+06u
M1002 VPWR C a_29_311# VPB phighvt w=420000u l=180000u
+  ad=8.325e+11p pd=6.94e+06u as=2.7055e+11p ps=3.05e+06u
M1003 a_29_311# B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_194_53# B a_122_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=8.82e+10p ps=1.26e+06u
M1005 VPWR a_29_311# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 X a_29_311# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1007 X a_29_311# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_122_53# A a_29_311# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1009 VPWR A a_29_311# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

