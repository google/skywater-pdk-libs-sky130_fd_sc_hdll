* File: sky130_fd_sc_hdll__isobufsrc_8.spice
* Created: Wed Sep  2 08:34:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__isobufsrc_8.pex.spice"
.subckt sky130_fd_sc_hdll__isobufsrc_8  VNB VPB A SLEEP VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* SLEEP	SLEEP
* A	A
* VPB	VPB
* VNB	VNB
MM1018 N_VGND_M1018_d N_A_M1018_g N_A_117_297#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.234 AS=0.104 PD=2.02 PS=0.97 NRD=4.608 NRS=2.76 M=1 R=4.33333 SA=75000.3
+ SB=75008.6 A=0.0975 P=1.6 MULT=1
MM1027 N_VGND_M1027_d N_A_M1027_g N_A_117_297#_M1018_s VNB NSHORT L=0.15 W=0.65
+ AD=0.21125 AS=0.104 PD=1.3 PS=0.97 NRD=6.456 NRS=4.608 M=1 R=4.33333
+ SA=75000.8 SB=75008.1 A=0.0975 P=1.6 MULT=1
MM1006 N_X_M1006_d N_A_117_297#_M1006_g N_VGND_M1027_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.21125 PD=0.97 PS=1.3 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1008 N_X_M1006_d N_A_117_297#_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1011 N_X_M1011_d N_A_117_297#_M1011_g N_VGND_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1019 N_X_M1011_d N_A_117_297#_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1020 N_X_M1020_d N_A_117_297#_M1020_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.4
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1026 N_X_M1020_d N_A_117_297#_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.9
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1029 N_X_M1029_d N_A_117_297#_M1029_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.4
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1032 N_X_M1029_d N_A_117_297#_M1032_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1009_d N_SLEEP_M1009_g N_VGND_M1032_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.3
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1009_d N_SLEEP_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.8
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1012 N_X_M1012_d N_SLEEP_M1012_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.3
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1013 N_X_M1012_d N_SLEEP_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75006.7
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1022 N_X_M1022_d N_SLEEP_M1022_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1024 N_X_M1022_d N_SLEEP_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75007.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1030 N_X_M1030_d N_SLEEP_M1030_g N_VGND_M1024_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1033 N_X_M1030_d N_SLEEP_M1033_g N_VGND_M1033_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75008.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.17 PD=2.54 PS=1.34 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1014_d N_A_M1014_g N_A_117_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.33 AS=0.17 PD=2.66 PS=1.34 NRD=0.9653 NRS=10.8153 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_A_117_297#_M1000_g N_A_345_297#_M1000_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90007.2 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1000_d N_A_117_297#_M1002_g N_A_345_297#_M1002_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.7 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_117_297#_M1004_g N_A_345_297#_M1002_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.1 SB=90006.3 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1004_d N_A_117_297#_M1005_g N_A_345_297#_M1005_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001.6 SB=90005.8 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_117_297#_M1015_g N_A_345_297#_M1005_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.1 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1015_d N_A_117_297#_M1017_g N_A_345_297#_M1017_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90002.5 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1023_d N_A_117_297#_M1023_g N_A_345_297#_M1017_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1031 N_VPWR_M1023_d N_A_117_297#_M1031_g N_A_345_297#_M1031_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90003.5 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1003 N_A_345_297#_M1031_s N_SLEEP_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1007 N_A_345_297#_M1007_d N_SLEEP_M1007_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.4 SB=90003 A=0.18 P=2.36 MULT=1
MM1016 N_A_345_297#_M1007_d N_SLEEP_M1016_g N_X_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.9 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1021 N_A_345_297#_M1021_d N_SLEEP_M1021_g N_X_M1016_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1025 N_A_345_297#_M1021_d N_SLEEP_M1025_g N_X_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.8 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1028 N_A_345_297#_M1028_d N_SLEEP_M1028_g N_X_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.3 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1034 N_A_345_297#_M1028_d N_SLEEP_M1034_g N_X_M1034_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.8 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1035 N_A_345_297#_M1035_d N_SLEEP_M1035_g N_X_M1034_s VPB PHIGHVT L=0.18 W=1
+ AD=0.28 AS=0.145 PD=2.56 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX36_noxref VNB VPB NWDIODE A=16.1142 P=23.29
pX37_noxref noxref_10 SLEEP SLEEP PROBETYPE=1
*
.include "sky130_fd_sc_hdll__isobufsrc_8.pxi.spice"
*
.ends
*
*
