# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdfsbp_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfsbp_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.64000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.855000 1.720000 3.335000 1.970000 ;
        RECT 3.155000 1.055000 3.815000 1.590000 ;
        RECT 3.155000 1.590000 3.335000 1.720000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.765000 1.425000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 14.700000 0.275000 15.080000 0.825000 ;
        RECT 14.700000 1.495000 15.080000 2.450000 ;
        RECT 14.805000 0.825000 15.080000 1.495000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.555000 0.255000 13.000000 2.465000 ;
    END
  END Q_N
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.365000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.570000 1.075000 0.860000 1.120000 ;
        RECT 0.570000 1.120000 2.875000 1.260000 ;
        RECT 0.570000 1.260000 0.860000 1.305000 ;
        RECT 2.585000 1.075000 2.875000 1.120000 ;
        RECT 2.585000 1.260000 2.875000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 7.385000 1.415000 7.725000 1.460000 ;
        RECT 7.385000 1.460000 9.965000 1.600000 ;
        RECT 7.385000 1.600000 7.725000 1.645000 ;
        RECT 9.675000 1.415000 9.965000 1.460000 ;
        RECT 9.675000 1.600000 9.965000 1.645000 ;
    END
  END SET_B
  PIN VGND
    ANTENNADIFFAREA  1.905350 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.625500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 15.640000 0.085000 ;
      RECT  0.000000  2.635000 15.640000 2.805000 ;
      RECT  0.085000  0.085000  0.430000 0.595000 ;
      RECT  0.085000  1.845000  1.205000 2.025000 ;
      RECT  0.085000  2.025000  0.345000 2.465000 ;
      RECT  0.515000  2.195000  0.815000 2.635000 ;
      RECT  0.550000  0.765000  0.860000 1.675000 ;
      RECT  0.975000  0.280000  1.845000 0.560000 ;
      RECT  1.035000  2.025000  1.205000 2.255000 ;
      RECT  1.035000  2.255000  2.245000 2.465000 ;
      RECT  1.395000  1.870000  1.845000 2.075000 ;
      RECT  1.655000  0.560000  1.845000 1.870000 ;
      RECT  2.025000  0.085000  2.205000 0.545000 ;
      RECT  2.065000  0.715000  2.715000 0.905000 ;
      RECT  2.065000  0.905000  2.400000 1.770000 ;
      RECT  2.065000  1.770000  2.685000 2.085000 ;
      RECT  2.460000  0.255000  2.715000 0.715000 ;
      RECT  2.470000  2.085000  2.685000 2.465000 ;
      RECT  2.570000  1.075000  2.950000 1.550000 ;
      RECT  2.940000  0.085000  3.280000 0.555000 ;
      RECT  2.940000  2.140000  3.280000 2.635000 ;
      RECT  3.505000  1.775000  4.295000 1.955000 ;
      RECT  3.505000  1.955000  3.675000 2.325000 ;
      RECT  3.520000  0.255000  3.705000 0.715000 ;
      RECT  3.520000  0.715000  4.295000 0.885000 ;
      RECT  3.845000  2.275000  4.225000 2.635000 ;
      RECT  3.930000  0.085000  4.240000 0.545000 ;
      RECT  4.035000  0.885000  4.295000 1.775000 ;
      RECT  4.445000  2.135000  4.790000 2.465000 ;
      RECT  4.460000  0.255000  4.685000 0.585000 ;
      RECT  4.515000  0.585000  4.685000 1.090000 ;
      RECT  4.515000  1.090000  4.840000 1.420000 ;
      RECT  4.515000  1.420000  4.790000 2.135000 ;
      RECT  4.855000  0.255000  5.180000 0.920000 ;
      RECT  4.960000  1.590000  5.180000 2.465000 ;
      RECT  5.010000  0.920000  5.180000 1.590000 ;
      RECT  5.400000  0.255000  5.890000 1.225000 ;
      RECT  5.400000  1.225000  8.360000 1.275000 ;
      RECT  5.430000  2.135000  6.205000 2.465000 ;
      RECT  5.485000  1.275000  6.935000 1.395000 ;
      RECT  5.605000  1.575000  5.865000 1.955000 ;
      RECT  6.035000  1.395000  6.205000 2.135000 ;
      RECT  6.060000  0.085000  6.595000 0.465000 ;
      RECT  6.060000  0.635000  7.085000 0.805000 ;
      RECT  6.060000  0.805000  6.475000 1.015000 ;
      RECT  6.425000  1.575000  6.595000 1.935000 ;
      RECT  6.425000  1.935000  7.365000 2.105000 ;
      RECT  6.445000  2.275000  6.775000 2.635000 ;
      RECT  6.750000  0.975000  8.360000 1.225000 ;
      RECT  6.775000  0.255000  7.085000 0.635000 ;
      RECT  7.100000  2.105000  7.365000 2.450000 ;
      RECT  7.190000  1.445000  7.725000 1.765000 ;
      RECT  7.540000  0.085000  8.275000 0.690000 ;
      RECT  7.655000  2.125000  8.710000 2.635000 ;
      RECT  7.910000  1.495000  8.755000 1.955000 ;
      RECT  7.950000  1.275000  8.360000 1.325000 ;
      RECT  8.535000  0.695000  9.890000 0.895000 ;
      RECT  8.535000  0.895000  8.755000 1.495000 ;
      RECT  8.880000  2.125000  9.735000 2.460000 ;
      RECT  9.115000  1.075000  9.395000 1.905000 ;
      RECT  9.160000  0.275000 10.775000 0.445000 ;
      RECT  9.565000  1.895000 11.465000 2.065000 ;
      RECT  9.565000  2.065000  9.735000 2.125000 ;
      RECT  9.610000  0.895000  9.890000 1.245000 ;
      RECT  9.685000  1.415000  9.960000 1.525000 ;
      RECT  9.685000  1.525000 11.075000 1.725000 ;
      RECT 10.045000  2.235000 10.425000 2.635000 ;
      RECT 10.140000  0.855000 10.365000 1.185000 ;
      RECT 10.140000  1.185000 11.945000 1.355000 ;
      RECT 10.605000  0.445000 10.775000 0.845000 ;
      RECT 10.605000  0.845000 11.545000 1.015000 ;
      RECT 10.645000  2.065000 10.860000 2.450000 ;
      RECT 11.135000  2.235000 11.465000 2.635000 ;
      RECT 11.220000  0.085000 11.390000 0.545000 ;
      RECT 11.245000  1.525000 11.465000 1.895000 ;
      RECT 11.560000  0.255000 11.945000 0.540000 ;
      RECT 11.685000  1.355000 11.945000 2.465000 ;
      RECT 11.765000  0.540000 11.945000 1.185000 ;
      RECT 12.170000  0.085000 12.380000 0.885000 ;
      RECT 12.170000  1.485000 12.380000 2.635000 ;
      RECT 13.215000  0.085000 13.505000 0.885000 ;
      RECT 13.215000  1.485000 13.505000 2.635000 ;
      RECT 13.720000  0.255000 13.905000 0.995000 ;
      RECT 13.720000  0.995000 14.585000 1.325000 ;
      RECT 13.720000  1.325000 13.905000 2.465000 ;
      RECT 14.075000  0.085000 14.480000 0.825000 ;
      RECT 14.075000  1.635000 14.480000 2.635000 ;
      RECT 15.250000  0.085000 15.515000 0.885000 ;
      RECT 15.250000  1.485000 15.515000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.630000  1.105000  0.800000 1.275000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.675000  1.445000  1.845000 1.615000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.645000  1.105000  2.815000 1.275000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.125000  1.785000  4.295000 1.955000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.585000  1.105000  4.755000 1.275000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.010000  1.445000  5.180000 1.615000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.605000  1.785000  5.775000 1.955000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.445000  1.445000  7.615000 1.615000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.205000  1.785000  8.375000 1.955000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.225000  1.105000  9.395000 1.275000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.735000  1.445000  9.905000 1.615000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
      RECT 12.105000 -0.085000 12.275000 0.085000 ;
      RECT 12.105000  2.635000 12.275000 2.805000 ;
      RECT 12.565000 -0.085000 12.735000 0.085000 ;
      RECT 12.565000  2.635000 12.735000 2.805000 ;
      RECT 13.025000 -0.085000 13.195000 0.085000 ;
      RECT 13.025000  2.635000 13.195000 2.805000 ;
      RECT 13.485000 -0.085000 13.655000 0.085000 ;
      RECT 13.485000  2.635000 13.655000 2.805000 ;
      RECT 13.945000 -0.085000 14.115000 0.085000 ;
      RECT 13.945000  2.635000 14.115000 2.805000 ;
      RECT 14.405000 -0.085000 14.575000 0.085000 ;
      RECT 14.405000  2.635000 14.575000 2.805000 ;
      RECT 14.865000 -0.085000 15.035000 0.085000 ;
      RECT 14.865000  2.635000 15.035000 2.805000 ;
      RECT 15.325000 -0.085000 15.495000 0.085000 ;
      RECT 15.325000  2.635000 15.495000 2.805000 ;
    LAYER met1 ;
      RECT 1.615000 1.415000 1.955000 1.460000 ;
      RECT 1.615000 1.460000 5.240000 1.600000 ;
      RECT 1.615000 1.600000 1.955000 1.645000 ;
      RECT 4.065000 1.755000 4.405000 1.800000 ;
      RECT 4.065000 1.800000 8.435000 1.940000 ;
      RECT 4.065000 1.940000 4.405000 1.985000 ;
      RECT 4.525000 1.075000 4.815000 1.120000 ;
      RECT 4.525000 1.120000 9.455000 1.260000 ;
      RECT 4.525000 1.260000 4.815000 1.305000 ;
      RECT 4.950000 1.415000 5.240000 1.460000 ;
      RECT 4.950000 1.600000 5.240000 1.645000 ;
      RECT 5.545000 1.755000 5.885000 1.800000 ;
      RECT 5.545000 1.940000 5.885000 1.985000 ;
      RECT 8.145000 1.755000 8.435000 1.800000 ;
      RECT 8.145000 1.940000 8.435000 1.985000 ;
      RECT 9.115000 1.075000 9.455000 1.120000 ;
      RECT 9.115000 1.260000 9.455000 1.305000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfsbp_2
