* File: sky130_fd_sc_hdll__a22o_2.pex.spice
* Created: Thu Aug 27 18:54:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22O_2%B2 1 3 4 6 7 11
c24 1 0 1.14637e-19 $X=0.495 $Y=1.41
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r26 7 11 9.70455 $w=1.98e-07 $l=1.75e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.41 $Y2=1.175
r27 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.435 $Y2=1.16
r28 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r29 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.435 $Y2=1.16
r30 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%B1 1 3 4 6 7 8 14 22
r36 14 22 2.48225 $w=2.08e-07 $l=4.7e-08 $layer=LI1_cond $X=1.202 $Y=1.18
+ $X2=1.155 $Y2=1.18
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.16 $X2=0.98 $Y2=1.16
r38 8 14 9.42908 $w=2.73e-07 $l=2.25e-07 $layer=LI1_cond $X=1.202 $Y=0.85
+ $X2=1.202 $Y2=1.075
r39 7 22 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=1.15 $Y=1.18 $X2=1.155
+ $Y2=1.18
r40 7 13 8.97835 $w=2.08e-07 $l=1.7e-07 $layer=LI1_cond $X=1.15 $Y=1.18 $X2=0.98
+ $Y2=1.18
r41 4 12 47.2262 $w=3.11e-07 $l=2.64575e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.995 $Y2=1.16
r42 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r43 1 12 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.9 $Y=0.995
+ $X2=0.995 $Y2=1.16
r44 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.9 $Y=0.995 $X2=0.9
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%A1 1 3 4 6 7 8 13
r36 13 19 3.34013 $w=4.13e-07 $l=8.5e-08 $layer=LI1_cond $X=1.732 $Y=1.16
+ $X2=1.732 $Y2=1.075
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.775
+ $Y=1.16 $X2=1.775 $Y2=1.16
r38 8 13 0.833091 $w=4.13e-07 $l=3e-08 $layer=LI1_cond $X=1.732 $Y=1.19
+ $X2=1.732 $Y2=1.16
r39 7 19 8.78982 $w=2.93e-07 $l=2.25e-07 $layer=LI1_cond $X=1.672 $Y=0.85
+ $X2=1.672 $Y2=1.075
r40 4 12 39.0558 $w=3.7e-07 $l=2.21743e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.847 $Y2=1.16
r41 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.56
r42 1 12 45.3064 $w=3.7e-07 $l=2.99165e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.847 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%A2 1 3 4 6 7
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=1.16 $X2=2.4 $Y2=1.16
r34 7 11 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=2.505 $Y=1.175
+ $X2=2.4 $Y2=1.175
r35 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.51 $Y=0.995
+ $X2=2.425 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.51 $Y=0.995 $X2=2.51
+ $Y2=0.56
r37 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.425 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.485 $Y=1.41
+ $X2=2.485 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%A_27_297# 1 2 3 4 13 15 16 18 19 21 22 24
+ 26 28 29 30 33 40 41 42 46 51 52 57
c125 51 0 1.14637e-19 $X=1.2 $Y=2.34
r126 57 58 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3.47 $Y=1.202
+ $X2=3.495 $Y2=1.202
r127 56 57 57.504 $w=3.73e-07 $l=4.45e-07 $layer=POLY_cond $X=3.025 $Y=1.202
+ $X2=3.47 $Y2=1.202
r128 55 56 3.23056 $w=3.73e-07 $l=2.5e-08 $layer=POLY_cond $X=3 $Y=1.202
+ $X2=3.025 $Y2=1.202
r129 51 52 9.14916 $w=2.08e-07 $l=1.65e-07 $layer=LI1_cond $X=1.2 $Y=2.36
+ $X2=1.035 $Y2=2.36
r130 47 55 9.04558 $w=3.73e-07 $l=7e-08 $layer=POLY_cond $X=2.93 $Y=1.202 $X2=3
+ $Y2=1.202
r131 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.93
+ $Y=1.16 $X2=2.93 $Y2=1.16
r132 44 46 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.93 $Y=1.455
+ $X2=2.93 $Y2=1.16
r133 43 46 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.93 $Y=0.905
+ $X2=2.93 $Y2=1.16
r134 41 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.845 $Y=0.82
+ $X2=2.93 $Y2=0.905
r135 41 42 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.845 $Y=0.82
+ $X2=2.295 $Y2=0.82
r136 40 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.21 $Y=0.735
+ $X2=2.295 $Y2=0.82
r137 39 40 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.21 $Y=0.505
+ $X2=2.21 $Y2=0.735
r138 35 38 25.8147 $w=2.48e-07 $l=5.6e-07 $layer=LI1_cond $X=1.16 $Y=0.38
+ $X2=1.72 $Y2=0.38
r139 33 39 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=2.125 $Y=0.38
+ $X2=2.21 $Y2=0.505
r140 33 38 18.6696 $w=2.48e-07 $l=4.05e-07 $layer=LI1_cond $X=2.125 $Y=0.38
+ $X2=1.72 $Y2=0.38
r141 32 49 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=0.26 $Y2=2.38
r142 32 52 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=0.425 $Y=2.38
+ $X2=1.035 $Y2=2.38
r143 29 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.845 $Y=1.54
+ $X2=2.93 $Y2=1.455
r144 29 30 157.882 $w=1.68e-07 $l=2.42e-06 $layer=LI1_cond $X=2.845 $Y=1.54
+ $X2=0.425 $Y2=1.54
r145 26 49 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=2.38
r146 26 28 22.1758 $w=3.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.66
r147 25 30 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.425 $Y2=1.54
r148 25 28 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=0.26 $Y=1.625
+ $X2=0.26 $Y2=1.66
r149 22 58 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.495 $Y2=1.202
r150 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.495 $Y2=0.56
r151 19 57 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.202
r152 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.985
r153 16 56 24.162 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=1.202
r154 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.025 $Y=0.995
+ $X2=3.025 $Y2=0.56
r155 13 55 19.8045 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3 $Y=1.41 $X2=3
+ $Y2=1.202
r156 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3 $Y=1.41 $X2=3
+ $Y2=1.985
r157 4 51 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r158 3 49 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r159 3 28 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r160 2 38 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.42
r161 1 35 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=0.975
+ $Y=0.235 $X2=1.16 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%A_117_297# 1 2 7 9 11 16
r23 14 16 5.94149 $w=3.28e-07 $l=1.45e-07 $layer=LI1_cond $X=0.73 $Y=1.96
+ $X2=0.875 $Y2=1.96
r24 9 18 3.3405 $w=2.5e-07 $l=1.2e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.255 $Y2=1.915
r25 9 11 12.2159 $w=2.48e-07 $l=2.65e-07 $layer=LI1_cond $X=2.255 $Y=2.035
+ $X2=2.255 $Y2=2.3
r26 7 18 3.47969 $w=2.4e-07 $l=1.25e-07 $layer=LI1_cond $X=2.13 $Y=1.915
+ $X2=2.255 $Y2=1.915
r27 7 16 60.2632 $w=2.38e-07 $l=1.255e-06 $layer=LI1_cond $X=2.13 $Y=1.915
+ $X2=0.875 $Y2=1.915
r28 2 18 600 $w=1.7e-07 $l=5.43392e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.215 $Y2=1.95
r29 2 11 600 $w=1.7e-07 $l=8.95977e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.215 $Y2=2.3
r30 1 14 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%VPWR 1 2 3 12 16 18 20 25 26 27 29 38 43 47
r57 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r58 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r59 41 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r60 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r61 38 46 3.40825 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.947 $Y2=2.72
r62 38 40 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=2.72
+ $X2=3.45 $Y2=2.72
r63 37 41 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r64 37 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r65 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r66 34 43 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=1.732 $Y2=2.72
r67 34 36 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=1.91 $Y=2.72
+ $X2=2.53 $Y2=2.72
r68 29 43 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.732 $Y2=2.72
r69 29 31 86.4438 $w=1.68e-07 $l=1.325e-06 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 27 44 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r71 27 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 25 36 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.6 $Y=2.72 $X2=2.53
+ $Y2=2.72
r73 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.6 $Y=2.72
+ $X2=2.765 $Y2=2.72
r74 24 40 33.9251 $w=1.68e-07 $l=5.2e-07 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=3.45 $Y2=2.72
r75 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.93 $Y=2.72
+ $X2=2.765 $Y2=2.72
r76 20 23 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.84 $Y=1.63
+ $X2=3.84 $Y2=2.31
r77 18 46 3.40825 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.947 $Y2=2.72
r78 18 23 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.84 $Y=2.635
+ $X2=3.84 $Y2=2.31
r79 14 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.765 $Y2=2.72
r80 14 16 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.765 $Y2=1.96
r81 10 43 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=2.72
r82 10 12 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=1.732 $Y=2.635
+ $X2=1.732 $Y2=2.3
r83 3 23 400 $w=1.7e-07 $l=9.54791e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.84 $Y2=2.31
r84 3 20 400 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=3.56
+ $Y=1.485 $X2=3.84 $Y2=1.63
r85 2 16 300 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_PDIFF $count=2 $X=2.575
+ $Y=1.485 $X2=2.765 $Y2=1.96
r86 1 12 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%X 1 2 7 8 9 10 11 12 36 40
r24 40 41 2.69457 $w=4.08e-07 $l=7.5e-08 $layer=LI1_cond $X=3.355 $Y=0.51
+ $X2=3.355 $Y2=0.585
r25 31 46 0.843251 $w=4.08e-07 $l=3e-08 $layer=LI1_cond $X=3.355 $Y=1.99
+ $X2=3.355 $Y2=1.96
r26 12 31 6.18384 $w=4.08e-07 $l=2.2e-07 $layer=LI1_cond $X=3.355 $Y=2.21
+ $X2=3.355 $Y2=1.99
r27 9 46 2.52975 $w=4.08e-07 $l=9e-08 $layer=LI1_cond $X=3.355 $Y=1.87 $X2=3.355
+ $Y2=1.96
r28 9 11 7.66305 $w=4.88e-07 $l=2.55e-07 $layer=LI1_cond $X=3.4 $Y=1.785 $X2=3.4
+ $Y2=1.53
r29 8 11 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.4 $Y=1.19 $X2=3.4
+ $Y2=1.53
r30 8 10 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=3.4 $Y=1.19 $X2=3.4
+ $Y2=0.85
r31 7 40 0.140542 $w=4.08e-07 $l=5e-09 $layer=LI1_cond $X=3.355 $Y=0.505
+ $X2=3.355 $Y2=0.51
r32 7 36 2.38921 $w=4.08e-07 $l=8.5e-08 $layer=LI1_cond $X=3.355 $Y=0.505
+ $X2=3.355 $Y2=0.42
r33 7 10 9.3636 $w=3.18e-07 $l=2.6e-07 $layer=LI1_cond $X=3.4 $Y=0.59 $X2=3.4
+ $Y2=0.85
r34 7 41 0.180069 $w=3.18e-07 $l=5e-09 $layer=LI1_cond $X=3.4 $Y=0.59 $X2=3.4
+ $Y2=0.585
r35 2 46 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.09
+ $Y=1.485 $X2=3.235 $Y2=1.96
r36 1 36 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.1
+ $Y=0.235 $X2=3.235 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_2%VGND 1 2 3 10 12 16 18 20 22 24 29 38 42
r49 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r50 38 39 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r51 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r52 33 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r53 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 30 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=2.695
+ $Y2=0
r55 30 32 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.885 $Y=0 $X2=3.45
+ $Y2=0
r56 29 41 3.40825 $w=1.7e-07 $l=1.92e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.947
+ $Y2=0
r57 29 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.755 $Y=0 $X2=3.45
+ $Y2=0
r58 28 39 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r59 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r60 25 35 6.38223 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.297
+ $Y2=0
r61 25 27 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.69
+ $Y2=0
r62 24 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.505 $Y=0 $X2=2.695
+ $Y2=0
r63 24 27 118.412 $w=1.68e-07 $l=1.815e-06 $layer=LI1_cond $X=2.505 $Y=0
+ $X2=0.69 $Y2=0
r64 22 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r65 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r66 18 41 3.40825 $w=1.7e-07 $l=1.43332e-07 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.947 $Y2=0
r67 18 20 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.84 $Y=0.085
+ $X2=3.84 $Y2=0.4
r68 14 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0
r69 14 16 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=2.695 $Y=0.085
+ $X2=2.695 $Y2=0.4
r70 10 35 2.84844 $w=5e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.297 $Y2=0
r71 10 12 7.53529 $w=4.98e-07 $l=3.15e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.4
r72 3 20 91 $w=1.7e-07 $l=3.4271e-07 $layer=licon1_NDIFF $count=2 $X=3.57
+ $Y=0.235 $X2=3.84 $Y2=0.4
r73 2 16 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.585
+ $Y=0.235 $X2=2.72 $Y2=0.4
r74 1 12 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

