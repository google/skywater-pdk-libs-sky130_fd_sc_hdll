* File: sky130_fd_sc_hdll__nand4bb_4.pxi.spice
* Created: Thu Aug 27 19:15:15 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_N N_A_N_c_136_n N_A_N_M1014_g N_A_N_c_133_n
+ N_A_N_M1021_g A_N A_N N_A_N_c_135_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%B_N N_B_N_c_161_n N_B_N_M1001_g N_B_N_c_162_n
+ N_B_N_M1013_g B_N B_N N_B_N_c_163_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%B_N
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_27_47# N_A_27_47#_M1021_s N_A_27_47#_M1014_s
+ N_A_27_47#_c_203_n N_A_27_47#_M1004_g N_A_27_47#_c_194_n N_A_27_47#_M1007_g
+ N_A_27_47#_c_204_n N_A_27_47#_M1010_g N_A_27_47#_M1032_g N_A_27_47#_c_205_n
+ N_A_27_47#_M1022_g N_A_27_47#_M1033_g N_A_27_47#_c_206_n N_A_27_47#_M1034_g
+ N_A_27_47#_M1035_g N_A_27_47#_c_198_n N_A_27_47#_c_207_n N_A_27_47#_c_214_n
+ N_A_27_47#_c_199_n N_A_27_47#_c_218_n N_A_27_47#_c_208_n N_A_27_47#_c_200_n
+ N_A_27_47#_c_250_p N_A_27_47#_c_201_n N_A_27_47#_c_202_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_206_47# N_A_206_47#_M1013_d
+ N_A_206_47#_M1001_d N_A_206_47#_M1002_g N_A_206_47#_c_344_n
+ N_A_206_47#_M1003_g N_A_206_47#_M1008_g N_A_206_47#_c_345_n
+ N_A_206_47#_M1015_g N_A_206_47#_M1025_g N_A_206_47#_c_346_n
+ N_A_206_47#_M1019_g N_A_206_47#_c_347_n N_A_206_47#_M1031_g
+ N_A_206_47#_M1028_g N_A_206_47#_c_348_n N_A_206_47#_c_340_n
+ N_A_206_47#_c_341_n N_A_206_47#_c_349_n N_A_206_47#_c_342_n
+ N_A_206_47#_c_378_n N_A_206_47#_c_381_n N_A_206_47#_c_350_n
+ N_A_206_47#_c_384_n N_A_206_47#_c_343_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_206_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%C N_C_c_479_n N_C_M1005_g N_C_M1000_g
+ N_C_c_480_n N_C_M1023_g N_C_M1009_g N_C_c_481_n N_C_M1027_g N_C_M1011_g
+ N_C_c_482_n N_C_M1029_g N_C_M1020_g C C C C N_C_c_476_n N_C_c_477_n
+ N_C_c_478_n C C C C PM_SKY130_FD_SC_HDLL__NAND4BB_4%C
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%D N_D_M1016_g N_D_c_555_n N_D_M1006_g
+ N_D_M1018_g N_D_c_556_n N_D_M1012_g N_D_M1026_g N_D_c_557_n N_D_M1017_g
+ N_D_M1030_g N_D_c_558_n N_D_M1024_g D D D D N_D_c_553_n N_D_c_554_n D D D
+ PM_SKY130_FD_SC_HDLL__NAND4BB_4%D
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%VPWR N_VPWR_M1014_d N_VPWR_M1004_d
+ N_VPWR_M1010_d N_VPWR_M1034_d N_VPWR_M1015_s N_VPWR_M1031_s N_VPWR_M1023_s
+ N_VPWR_M1029_s N_VPWR_M1012_d N_VPWR_M1024_d N_VPWR_c_623_n N_VPWR_c_624_n
+ N_VPWR_c_625_n N_VPWR_c_626_n N_VPWR_c_627_n N_VPWR_c_628_n N_VPWR_c_629_n
+ N_VPWR_c_630_n N_VPWR_c_631_n N_VPWR_c_632_n N_VPWR_c_633_n N_VPWR_c_634_n
+ N_VPWR_c_635_n N_VPWR_c_636_n N_VPWR_c_637_n N_VPWR_c_638_n N_VPWR_c_639_n
+ N_VPWR_c_640_n N_VPWR_c_641_n N_VPWR_c_642_n VPWR N_VPWR_c_643_n
+ N_VPWR_c_644_n N_VPWR_c_645_n N_VPWR_c_646_n N_VPWR_c_647_n N_VPWR_c_648_n
+ N_VPWR_c_649_n N_VPWR_c_650_n N_VPWR_c_651_n N_VPWR_c_652_n N_VPWR_c_622_n
+ PM_SKY130_FD_SC_HDLL__NAND4BB_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%Y N_Y_M1007_d N_Y_M1033_d N_Y_M1004_s
+ N_Y_M1022_s N_Y_M1003_d N_Y_M1019_d N_Y_M1005_d N_Y_M1027_d N_Y_M1006_s
+ N_Y_M1017_s N_Y_c_787_n N_Y_c_808_n N_Y_c_789_n N_Y_c_790_n N_Y_c_817_n
+ N_Y_c_820_n N_Y_c_791_n N_Y_c_792_n N_Y_c_848_n N_Y_c_793_n N_Y_c_867_n
+ N_Y_c_794_n N_Y_c_874_n N_Y_c_795_n N_Y_c_879_n N_Y_c_796_n N_Y_c_797_n
+ N_Y_c_903_n N_Y_c_798_n N_Y_c_799_n N_Y_c_800_n N_Y_c_801_n Y Y N_Y_c_830_n Y
+ PM_SKY130_FD_SC_HDLL__NAND4BB_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%VGND N_VGND_M1021_d N_VGND_M1016_s
+ N_VGND_M1026_s N_VGND_c_979_n N_VGND_c_980_n N_VGND_c_981_n N_VGND_c_982_n
+ N_VGND_c_983_n N_VGND_c_984_n VGND N_VGND_c_985_n N_VGND_c_986_n
+ N_VGND_c_987_n N_VGND_c_988_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_395_47# N_A_395_47#_M1007_s
+ N_A_395_47#_M1032_s N_A_395_47#_M1035_s N_A_395_47#_M1008_d
+ N_A_395_47#_M1028_d N_A_395_47#_c_1077_n N_A_395_47#_c_1090_n
+ N_A_395_47#_c_1078_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_395_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_853_47# N_A_853_47#_M1002_s
+ N_A_853_47#_M1025_s N_A_853_47#_M1000_s N_A_853_47#_M1011_s
+ N_A_853_47#_c_1120_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_853_47#
x_PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_1251_47# N_A_1251_47#_M1000_d
+ N_A_1251_47#_M1009_d N_A_1251_47#_M1020_d N_A_1251_47#_M1018_d
+ N_A_1251_47#_M1030_d N_A_1251_47#_c_1156_n N_A_1251_47#_c_1166_n
+ N_A_1251_47#_c_1160_n PM_SKY130_FD_SC_HDLL__NAND4BB_4%A_1251_47#
cc_1 VNB N_A_N_c_133_n 0.0218146f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB A_N 0.0132315f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_135_n 0.0374535f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_N_c_161_n 0.0204084f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_N_c_162_n 0.019471f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B_N_c_163_n 0.00277699f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_7 VNB N_A_27_47#_c_194_n 0.0200672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_M1032_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_M1033_g 0.0183474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_M1035_g 0.016866f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_198_n 0.0147604f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_199_n 0.00802475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_200_n 0.00399837f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_201_n 0.0649753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_202_n 0.084068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_206_47#_M1002_g 0.0182068f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_206_47#_M1008_g 0.0183665f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_18 VNB N_A_206_47#_M1025_g 0.0188863f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_206_47#_M1028_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_206_47#_c_340_n 0.00869179f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_206_47#_c_341_n 0.0114847f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_206_47#_c_342_n 0.00428644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_206_47#_c_343_n 0.0934346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C_M1000_g 0.0244378f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_25 VNB N_C_M1009_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_26 VNB N_C_M1011_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_C_M1020_g 0.0182512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_C_c_476_n 0.0306494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_C_c_477_n 0.00507666f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_C_c_478_n 0.0848272f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_D_M1016_g 0.0183452f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_32 VNB N_D_M1018_g 0.0183651f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_D_M1026_g 0.018595f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_D_M1030_g 0.0246977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB D 0.0103832f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_D_c_553_n 0.0835282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_D_c_554_n 0.0279824f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VPWR_c_622_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_787_n 0.00655553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB Y 0.00395553f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_979_n 0.00272748f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_42 VNB N_VGND_c_980_n 0.00220692f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.16
cc_43 VNB N_VGND_c_981_n 0.174993f $X=-0.19 $Y=-0.24 $X2=0.215 $Y2=1.53
cc_44 VNB N_VGND_c_982_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_983_n 0.015705f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_984_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_985_n 0.0143107f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_986_n 0.0220602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_987_n 0.504903f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_988_n 0.0055668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_395_47#_c_1077_n 0.00153527f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_395_47#_c_1078_n 0.00292796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_853_47#_c_1120_n 0.0296652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VPB N_A_N_c_136_n 0.0189297f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB A_N 0.0125739f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_56 VPB N_A_N_c_135_n 0.0154933f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_57 VPB N_B_N_c_161_n 0.027413f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_58 VPB N_B_N_c_163_n 4.94236e-19 $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_59 VPB N_A_27_47#_c_203_n 0.0193285f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_60 VPB N_A_27_47#_c_204_n 0.0154404f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_61 VPB N_A_27_47#_c_205_n 0.0158682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_206_n 0.0157857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_207_n 0.0180063f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_208_n 0.00912537f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_200_n 0.00256132f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_201_n 0.0374474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_202_n 0.025583f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_206_47#_c_344_n 0.0159745f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.202
cc_69 VPB N_A_206_47#_c_345_n 0.0158724f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_206_47#_c_346_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_206_47#_c_347_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_206_47#_c_348_n 0.0145641f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_206_47#_c_349_n 0.0176916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_206_47#_c_350_n 0.0018159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_206_47#_c_343_n 0.0286944f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_C_c_479_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_77 VPB N_C_c_480_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_78 VPB N_C_c_481_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.202
cc_79 VPB N_C_c_482_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_C_c_478_n 0.0287129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_D_c_555_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_82 VPB N_D_c_556_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_83 VPB N_D_c_557_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.215 $Y2=1.53
cc_84 VPB N_D_c_558_n 0.0198539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_D_c_553_n 0.028998f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_D_c_554_n 0.00844673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_623_n 0.00237984f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_624_n 0.00414143f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_625_n 0.00231485f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_626_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_627_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_628_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_629_n 0.00737229f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_630_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_631_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_632_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_633_n 0.0144823f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_634_n 0.047812f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_635_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_636_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_637_n 0.0215922f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_638_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_639_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_640_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_641_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_642_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_643_n 0.0151232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_644_n 0.0293088f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_645_n 0.016313f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_646_n 0.022232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_647_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_648_n 0.00392577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_649_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_650_n 0.00426174f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_651_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_652_n 0.0122844f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_622_n 0.0579871f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_789_n 0.00177751f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_790_n 0.00119387f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_Y_c_791_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_Y_c_792_n 0.00476286f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_Y_c_793_n 0.00912739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_Y_c_794_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_Y_c_795_n 0.0052852f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_Y_c_796_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_Y_c_797_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_Y_c_798_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Y_c_799_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Y_c_800_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_Y_c_801_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB Y 0.00192405f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 N_A_N_c_136_n N_B_N_c_161_n 0.0386899f $X=0.495 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_133 A_N N_B_N_c_161_n 2.08799e-19 $X=0.15 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_134 N_A_N_c_135_n N_B_N_c_161_n 0.0254519f $X=0.495 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_135 N_A_N_c_133_n N_B_N_c_162_n 0.0247499f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_N_c_136_n N_B_N_c_163_n 0.00144992f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_137 A_N N_B_N_c_163_n 0.0310761f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_N_c_135_n N_B_N_c_163_n 0.0115234f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_139 A_N N_A_27_47#_M1014_s 0.00452798f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A_N_c_133_n N_A_27_47#_c_198_n 0.00425507f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_N_c_133_n N_A_27_47#_c_214_n 0.0164992f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_N_c_135_n N_A_27_47#_c_214_n 0.00285708f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_143 A_N N_A_27_47#_c_199_n 0.0179334f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_144 N_A_N_c_135_n N_A_27_47#_c_199_n 0.00237938f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_145 N_A_N_c_136_n N_A_27_47#_c_218_n 0.0217802f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_146 A_N N_A_27_47#_c_208_n 0.0204787f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A_N_c_135_n N_A_27_47#_c_208_n 0.00187944f $X=0.495 $Y=1.202 $X2=0
+ $Y2=0
cc_148 N_A_N_c_136_n N_VPWR_c_623_n 0.010811f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_N_c_136_n N_VPWR_c_643_n 0.00395083f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_N_c_136_n N_VPWR_c_622_n 0.00565038f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_N_c_133_n N_VGND_c_985_n 0.00198377f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_N_c_133_n N_VGND_c_987_n 0.00367064f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_N_c_133_n N_VGND_c_988_n 0.0112861f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B_N_c_161_n N_A_27_47#_c_214_n 3.82953e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B_N_c_162_n N_A_27_47#_c_214_n 0.0137333f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B_N_c_163_n N_A_27_47#_c_214_n 0.0280928f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B_N_c_161_n N_A_27_47#_c_218_n 0.0172423f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_158 N_B_N_c_163_n N_A_27_47#_c_218_n 0.0257158f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_159 N_B_N_c_161_n N_A_27_47#_c_200_n 0.0146565f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_160 N_B_N_c_162_n N_A_27_47#_c_200_n 0.0069944f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B_N_c_163_n N_A_27_47#_c_200_n 0.0496343f $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_162 N_B_N_c_161_n N_A_27_47#_c_201_n 0.0202849f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B_N_c_163_n N_A_27_47#_c_201_n 3.13741e-19 $X=0.94 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B_N_c_161_n N_A_206_47#_c_348_n 0.00633362f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_165 N_B_N_c_162_n N_A_206_47#_c_340_n 0.00481341f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_166 N_B_N_c_162_n N_A_206_47#_c_341_n 0.00421702f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_B_N_c_161_n N_A_206_47#_c_349_n 0.00449466f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_B_N_c_163_n N_VPWR_M1014_d 0.00194964f $X=0.94 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_169 N_B_N_c_161_n N_VPWR_c_623_n 0.00403433f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_N_c_161_n N_VPWR_c_644_n 0.00489587f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B_N_c_161_n N_VPWR_c_622_n 0.00786743f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_N_c_162_n N_VGND_c_981_n 0.00382585f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_N_c_162_n N_VGND_c_987_n 0.0057921f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B_N_c_162_n N_VGND_c_988_n 0.00780407f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_214_n N_A_206_47#_M1013_d 0.0133504f $X=1.195 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_176 N_A_27_47#_c_200_n N_A_206_47#_M1013_d 0.00198604f $X=1.42 $Y=1.16
+ $X2=-0.19 $Y2=-0.24
cc_177 N_A_27_47#_c_218_n N_A_206_47#_M1001_d 0.0124559f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_200_n N_A_206_47#_M1001_d 0.0107398f $X=1.42 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_M1035_g N_A_206_47#_M1002_g 0.0219184f $X=3.77 $Y=0.56 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_206_n N_A_206_47#_c_344_n 0.0227632f $X=3.745 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_218_n N_A_206_47#_c_348_n 0.0362102f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_194_n N_A_206_47#_c_340_n 9.24457e-19 $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_183 N_A_27_47#_c_214_n N_A_206_47#_c_340_n 0.0297553f $X=1.195 $Y=0.72 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_201_n N_A_206_47#_c_340_n 0.00521991f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_194_n N_A_206_47#_c_341_n 0.002948f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_214_n N_A_206_47#_c_341_n 0.0140572f $X=1.195 $Y=0.72 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_200_n N_A_206_47#_c_341_n 0.0205136f $X=1.42 $Y=1.16 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_201_n N_A_206_47#_c_341_n 0.0101291f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_c_203_n N_A_206_47#_c_349_n 0.00261716f $X=2.335 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_c_218_n N_A_206_47#_c_349_n 0.0161245f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_200_n N_A_206_47#_c_349_n 0.0372192f $X=1.42 $Y=1.16 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_c_201_n N_A_206_47#_c_349_n 0.00574989f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_202_n N_A_206_47#_c_349_n 0.00238213f $X=3.745 $Y=1.202
+ $X2=0 $Y2=0
cc_194 N_A_27_47#_c_250_p N_A_206_47#_c_342_n 0.0277024f $X=3.035 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_201_n N_A_206_47#_c_342_n 0.00685773f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_196 N_A_27_47#_c_202_n N_A_206_47#_c_342_n 0.0263606f $X=3.745 $Y=1.202 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_200_n N_A_206_47#_c_378_n 0.00140036f $X=1.42 $Y=1.16 $X2=0
+ $Y2=0
cc_198 N_A_27_47#_c_250_p N_A_206_47#_c_378_n 3.24364e-19 $X=3.035 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_201_n N_A_206_47#_c_378_n 0.0152355f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_200 N_A_27_47#_c_200_n N_A_206_47#_c_381_n 0.0157992f $X=1.42 $Y=1.16 $X2=0
+ $Y2=0
cc_201 N_A_27_47#_c_250_p N_A_206_47#_c_381_n 0.00514048f $X=3.035 $Y=1.16 $X2=0
+ $Y2=0
cc_202 N_A_27_47#_c_201_n N_A_206_47#_c_381_n 0.0208353f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_203 N_A_27_47#_c_202_n N_A_206_47#_c_384_n 2.35565e-19 $X=3.745 $Y=1.202
+ $X2=0 $Y2=0
cc_204 N_A_27_47#_c_202_n N_A_206_47#_c_343_n 0.0219184f $X=3.745 $Y=1.202 $X2=0
+ $Y2=0
cc_205 N_A_27_47#_c_218_n N_VPWR_M1014_d 0.00384337f $X=1.195 $Y=1.882 $X2=-0.19
+ $Y2=-0.24
cc_206 N_A_27_47#_c_218_n N_VPWR_c_623_n 0.0136926f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_207 N_A_27_47#_c_203_n N_VPWR_c_624_n 0.00592862f $X=2.335 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_27_47#_c_201_n N_VPWR_c_624_n 0.00486132f $X=2.235 $Y=1.16 $X2=0
+ $Y2=0
cc_209 N_A_27_47#_c_203_n N_VPWR_c_625_n 7.42159e-19 $X=2.335 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_27_47#_c_204_n N_VPWR_c_625_n 0.0151075f $X=2.805 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_205_n N_VPWR_c_625_n 0.00519708f $X=3.275 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_27_47#_c_205_n N_VPWR_c_626_n 0.00597712f $X=3.275 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_27_47#_c_206_n N_VPWR_c_626_n 0.00673617f $X=3.745 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_27_47#_c_206_n N_VPWR_c_627_n 0.0052072f $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_207_n N_VPWR_c_643_n 0.0165425f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_218_n N_VPWR_c_643_n 0.00202029f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_217 N_A_27_47#_c_218_n N_VPWR_c_644_n 0.00189996f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_218 N_A_27_47#_c_203_n N_VPWR_c_645_n 0.00597712f $X=2.335 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_27_47#_c_204_n N_VPWR_c_645_n 0.00427505f $X=2.805 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_27_47#_M1014_s N_VPWR_c_622_n 0.002367f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_221 N_A_27_47#_c_203_n N_VPWR_c_622_n 0.0112769f $X=2.335 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_204_n N_VPWR_c_622_n 0.00732977f $X=2.805 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_27_47#_c_205_n N_VPWR_c_622_n 0.00999457f $X=3.275 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_27_47#_c_206_n N_VPWR_c_622_n 0.011869f $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_27_47#_c_207_n N_VPWR_c_622_n 0.0107554f $X=0.26 $Y=2.275 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_218_n N_VPWR_c_622_n 0.00918143f $X=1.195 $Y=1.882 $X2=0
+ $Y2=0
cc_227 N_A_27_47#_c_194_n N_Y_c_787_n 0.00597217f $X=2.36 $Y=0.995 $X2=0 $Y2=0
cc_228 N_A_27_47#_M1032_g N_Y_c_787_n 0.0111034f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A_27_47#_M1033_g N_Y_c_787_n 0.0124988f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_250_p N_Y_c_787_n 0.0558172f $X=3.035 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_202_n N_Y_c_787_n 0.0103219f $X=3.745 $Y=1.202 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_203_n N_Y_c_808_n 0.0133529f $X=2.335 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_204_n N_Y_c_808_n 0.00416059f $X=2.805 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_204_n N_Y_c_789_n 0.0167108f $X=2.805 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_27_47#_c_205_n N_Y_c_789_n 0.0122386f $X=3.275 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_27_47#_c_250_p N_Y_c_789_n 0.0286833f $X=3.035 $Y=1.16 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_202_n N_Y_c_789_n 0.00900439f $X=3.745 $Y=1.202 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_203_n N_Y_c_790_n 0.00647857f $X=2.335 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_250_p N_Y_c_790_n 0.0174674f $X=3.035 $Y=1.16 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_202_n N_Y_c_790_n 0.00593229f $X=3.745 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_204_n N_Y_c_817_n 4.85405e-19 $X=2.805 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_205_n N_Y_c_817_n 0.0135107f $X=3.275 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_27_47#_c_206_n N_Y_c_817_n 0.0107001f $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_27_47#_c_206_n N_Y_c_820_n 6.49214e-19 $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_205_n N_Y_c_792_n 0.00369149f $X=3.275 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_206_n N_Y_c_792_n 0.0149171f $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_202_n N_Y_c_792_n 0.0085966f $X=3.745 $Y=1.202 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_205_n Y 2.107e-19 $X=3.275 $Y=1.41 $X2=0 $Y2=0
cc_249 N_A_27_47#_M1033_g Y 0.00249961f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_206_n Y 0.00183971f $X=3.745 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_27_47#_M1035_g Y 0.00312934f $X=3.77 $Y=0.56 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_250_p Y 0.00376631f $X=3.035 $Y=1.16 $X2=0 $Y2=0
cc_253 N_A_27_47#_c_202_n Y 0.0196048f $X=3.745 $Y=1.202 $X2=0 $Y2=0
cc_254 N_A_27_47#_M1035_g N_Y_c_830_n 0.00780112f $X=3.77 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_214_n N_VGND_M1021_d 0.00361179f $X=1.195 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_256 N_A_27_47#_c_194_n N_VGND_c_981_n 0.00357877f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_257 N_A_27_47#_M1032_g N_VGND_c_981_n 0.00357877f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A_27_47#_M1033_g N_VGND_c_981_n 0.00357877f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_27_47#_M1035_g N_VGND_c_981_n 0.00357877f $X=3.77 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_214_n N_VGND_c_981_n 0.00325692f $X=1.195 $Y=0.72 $X2=0
+ $Y2=0
cc_261 N_A_27_47#_c_198_n N_VGND_c_985_n 0.0179288f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_214_n N_VGND_c_985_n 0.00244154f $X=1.195 $Y=0.72 $X2=0
+ $Y2=0
cc_263 N_A_27_47#_M1021_s N_VGND_c_987_n 0.00289329f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_264 N_A_27_47#_c_194_n N_VGND_c_987_n 0.00677297f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_27_47#_M1032_g N_VGND_c_987_n 0.00548399f $X=2.83 $Y=0.56 $X2=0 $Y2=0
cc_266 N_A_27_47#_M1033_g N_VGND_c_987_n 0.00548399f $X=3.3 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_27_47#_M1035_g N_VGND_c_987_n 0.00538422f $X=3.77 $Y=0.56 $X2=0 $Y2=0
cc_268 N_A_27_47#_c_198_n N_VGND_c_987_n 0.00988152f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_269 N_A_27_47#_c_214_n N_VGND_c_987_n 0.0118754f $X=1.195 $Y=0.72 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_198_n N_VGND_c_988_n 0.0161786f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_214_n N_VGND_c_988_n 0.0196063f $X=1.195 $Y=0.72 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_194_n N_A_395_47#_c_1077_n 0.0052818f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_273 N_A_27_47#_c_201_n N_A_395_47#_c_1077_n 0.00536536f $X=2.235 $Y=1.16
+ $X2=0 $Y2=0
cc_274 N_A_27_47#_c_194_n N_A_395_47#_c_1078_n 0.0163476f $X=2.36 $Y=0.995 $X2=0
+ $Y2=0
cc_275 N_A_27_47#_M1032_g N_A_395_47#_c_1078_n 0.00958923f $X=2.83 $Y=0.56 $X2=0
+ $Y2=0
cc_276 N_A_27_47#_M1033_g N_A_395_47#_c_1078_n 0.00958923f $X=3.3 $Y=0.56 $X2=0
+ $Y2=0
cc_277 N_A_27_47#_M1035_g N_A_395_47#_c_1078_n 0.00958301f $X=3.77 $Y=0.56 $X2=0
+ $Y2=0
cc_278 N_A_27_47#_c_201_n N_A_395_47#_c_1078_n 0.00206727f $X=2.235 $Y=1.16
+ $X2=0 $Y2=0
cc_279 N_A_27_47#_M1035_g N_A_853_47#_c_1120_n 2.04286e-19 $X=3.77 $Y=0.56 $X2=0
+ $Y2=0
cc_280 N_A_206_47#_c_343_n N_C_c_476_n 0.00693702f $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_281 N_A_206_47#_c_384_n N_C_c_477_n 0.00793987f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_282 N_A_206_47#_c_343_n N_C_c_477_n 0.00233204f $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_283 N_A_206_47#_c_348_n N_VPWR_c_623_n 0.0218754f $X=1.675 $Y=2.307 $X2=0
+ $Y2=0
cc_284 N_A_206_47#_c_348_n N_VPWR_c_624_n 0.026185f $X=1.675 $Y=2.307 $X2=0
+ $Y2=0
cc_285 N_A_206_47#_c_349_n N_VPWR_c_624_n 0.0484095f $X=1.76 $Y=2.15 $X2=0 $Y2=0
cc_286 N_A_206_47#_c_342_n N_VPWR_c_624_n 0.00433199f $X=4.235 $Y=1.19 $X2=0
+ $Y2=0
cc_287 N_A_206_47#_c_378_n N_VPWR_c_624_n 2.19293e-19 $X=2.025 $Y=1.19 $X2=0
+ $Y2=0
cc_288 N_A_206_47#_c_381_n N_VPWR_c_624_n 5.51824e-19 $X=1.88 $Y=1.19 $X2=0
+ $Y2=0
cc_289 N_A_206_47#_c_344_n N_VPWR_c_627_n 0.004751f $X=4.215 $Y=1.41 $X2=0 $Y2=0
cc_290 N_A_206_47#_c_345_n N_VPWR_c_628_n 0.0052072f $X=4.685 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_206_47#_c_346_n N_VPWR_c_628_n 0.004751f $X=5.155 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_206_47#_c_347_n N_VPWR_c_629_n 0.00799044f $X=5.625 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_206_47#_c_344_n N_VPWR_c_635_n 0.00597712f $X=4.215 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_206_47#_c_345_n N_VPWR_c_635_n 0.00673617f $X=4.685 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_206_47#_c_348_n N_VPWR_c_644_n 0.0560407f $X=1.675 $Y=2.307 $X2=0
+ $Y2=0
cc_296 N_A_206_47#_c_346_n N_VPWR_c_646_n 0.00597712f $X=5.155 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_206_47#_c_347_n N_VPWR_c_646_n 0.00673617f $X=5.625 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_206_47#_M1001_d N_VPWR_c_622_n 0.00369224f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_299 N_A_206_47#_c_344_n N_VPWR_c_622_n 0.0100198f $X=4.215 $Y=1.41 $X2=0
+ $Y2=0
cc_300 N_A_206_47#_c_345_n N_VPWR_c_622_n 0.0118438f $X=4.685 $Y=1.41 $X2=0
+ $Y2=0
cc_301 N_A_206_47#_c_346_n N_VPWR_c_622_n 0.00999457f $X=5.155 $Y=1.41 $X2=0
+ $Y2=0
cc_302 N_A_206_47#_c_347_n N_VPWR_c_622_n 0.0132238f $X=5.625 $Y=1.41 $X2=0
+ $Y2=0
cc_303 N_A_206_47#_c_348_n N_VPWR_c_622_n 0.032206f $X=1.675 $Y=2.307 $X2=0
+ $Y2=0
cc_304 N_A_206_47#_c_342_n N_Y_c_787_n 0.017628f $X=4.235 $Y=1.19 $X2=0 $Y2=0
cc_305 N_A_206_47#_c_342_n N_Y_c_789_n 0.0238812f $X=4.235 $Y=1.19 $X2=0 $Y2=0
cc_306 N_A_206_47#_c_349_n N_Y_c_790_n 0.00173574f $X=1.76 $Y=2.15 $X2=0 $Y2=0
cc_307 N_A_206_47#_c_342_n N_Y_c_790_n 0.00674912f $X=4.235 $Y=1.19 $X2=0 $Y2=0
cc_308 N_A_206_47#_c_344_n N_Y_c_817_n 6.25403e-19 $X=4.215 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_206_47#_c_344_n N_Y_c_820_n 0.0133058f $X=4.215 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_206_47#_c_345_n N_Y_c_820_n 0.0107003f $X=4.685 $Y=1.41 $X2=0 $Y2=0
cc_311 N_A_206_47#_c_346_n N_Y_c_820_n 6.25403e-19 $X=5.155 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A_206_47#_c_345_n N_Y_c_791_n 0.0153933f $X=4.685 $Y=1.41 $X2=0 $Y2=0
cc_313 N_A_206_47#_c_346_n N_Y_c_791_n 0.0113962f $X=5.155 $Y=1.41 $X2=0 $Y2=0
cc_314 N_A_206_47#_c_343_n N_Y_c_791_n 0.00725062f $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_315 N_A_206_47#_c_344_n N_Y_c_792_n 0.0146193f $X=4.215 $Y=1.41 $X2=0 $Y2=0
cc_316 N_A_206_47#_c_345_n N_Y_c_792_n 0.00119493f $X=4.685 $Y=1.41 $X2=0 $Y2=0
cc_317 N_A_206_47#_c_342_n N_Y_c_792_n 0.00934565f $X=4.235 $Y=1.19 $X2=0 $Y2=0
cc_318 N_A_206_47#_c_350_n N_Y_c_792_n 0.00937583f $X=4.415 $Y=1.19 $X2=0 $Y2=0
cc_319 N_A_206_47#_c_384_n N_Y_c_792_n 0.0677883f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_320 N_A_206_47#_c_343_n N_Y_c_792_n 0.00614215f $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_321 N_A_206_47#_c_345_n N_Y_c_848_n 6.48386e-19 $X=4.685 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A_206_47#_c_346_n N_Y_c_848_n 0.0130707f $X=5.155 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A_206_47#_c_347_n N_Y_c_848_n 0.0161846f $X=5.625 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A_206_47#_c_347_n N_Y_c_793_n 0.0199408f $X=5.625 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A_206_47#_c_343_n N_Y_c_793_n 3.62813e-19 $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_326 N_A_206_47#_c_346_n N_Y_c_798_n 0.00292783f $X=5.155 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_206_47#_c_347_n N_Y_c_798_n 0.00116723f $X=5.625 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A_206_47#_c_384_n N_Y_c_798_n 0.0305808f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_206_47#_c_343_n N_Y_c_798_n 0.00723098f $X=5.625 $Y=1.217 $X2=0 $Y2=0
cc_330 N_A_206_47#_M1002_g Y 0.00936626f $X=4.19 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A_206_47#_c_344_n Y 9.02341e-19 $X=4.215 $Y=1.41 $X2=0 $Y2=0
cc_332 N_A_206_47#_c_342_n Y 0.0307725f $X=4.235 $Y=1.19 $X2=0 $Y2=0
cc_333 N_A_206_47#_c_350_n Y 0.00184817f $X=4.415 $Y=1.19 $X2=0 $Y2=0
cc_334 N_A_206_47#_c_384_n Y 0.0141847f $X=5.39 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_206_47#_M1002_g N_Y_c_830_n 0.00208161f $X=4.19 $Y=0.56 $X2=0 $Y2=0
cc_336 N_A_206_47#_M1002_g N_VGND_c_981_n 0.00357877f $X=4.19 $Y=0.56 $X2=0
+ $Y2=0
cc_337 N_A_206_47#_M1008_g N_VGND_c_981_n 0.00357877f $X=4.66 $Y=0.56 $X2=0
+ $Y2=0
cc_338 N_A_206_47#_M1025_g N_VGND_c_981_n 0.00357877f $X=5.13 $Y=0.56 $X2=0
+ $Y2=0
cc_339 N_A_206_47#_M1028_g N_VGND_c_981_n 0.00357877f $X=5.65 $Y=0.56 $X2=0
+ $Y2=0
cc_340 N_A_206_47#_c_340_n N_VGND_c_981_n 0.048343f $X=1.675 $Y=0.36 $X2=0 $Y2=0
cc_341 N_A_206_47#_M1013_d N_VGND_c_987_n 0.00421526f $X=1.03 $Y=0.235 $X2=0
+ $Y2=0
cc_342 N_A_206_47#_M1002_g N_VGND_c_987_n 0.00538422f $X=4.19 $Y=0.56 $X2=0
+ $Y2=0
cc_343 N_A_206_47#_M1008_g N_VGND_c_987_n 0.00548399f $X=4.66 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_206_47#_M1025_g N_VGND_c_987_n 0.00560377f $X=5.13 $Y=0.56 $X2=0
+ $Y2=0
cc_345 N_A_206_47#_M1028_g N_VGND_c_987_n 0.00680287f $X=5.65 $Y=0.56 $X2=0
+ $Y2=0
cc_346 N_A_206_47#_c_340_n N_VGND_c_987_n 0.0274952f $X=1.675 $Y=0.36 $X2=0
+ $Y2=0
cc_347 N_A_206_47#_c_340_n N_VGND_c_988_n 0.0142192f $X=1.675 $Y=0.36 $X2=0
+ $Y2=0
cc_348 N_A_206_47#_c_341_n N_A_395_47#_c_1077_n 0.031056f $X=1.76 $Y=1.075 $X2=0
+ $Y2=0
cc_349 N_A_206_47#_c_342_n N_A_395_47#_c_1077_n 0.00443762f $X=4.235 $Y=1.19
+ $X2=0 $Y2=0
cc_350 N_A_206_47#_c_378_n N_A_395_47#_c_1077_n 2.20995e-19 $X=2.025 $Y=1.19
+ $X2=0 $Y2=0
cc_351 N_A_206_47#_c_381_n N_A_395_47#_c_1077_n 6.33188e-19 $X=1.88 $Y=1.19
+ $X2=0 $Y2=0
cc_352 N_A_206_47#_c_340_n N_A_395_47#_c_1090_n 0.0193049f $X=1.675 $Y=0.36
+ $X2=0 $Y2=0
cc_353 N_A_206_47#_c_341_n N_A_395_47#_c_1090_n 0.00161596f $X=1.76 $Y=1.075
+ $X2=0 $Y2=0
cc_354 N_A_206_47#_M1002_g N_A_395_47#_c_1078_n 0.0124699f $X=4.19 $Y=0.56 $X2=0
+ $Y2=0
cc_355 N_A_206_47#_M1008_g N_A_395_47#_c_1078_n 0.00958923f $X=4.66 $Y=0.56
+ $X2=0 $Y2=0
cc_356 N_A_206_47#_M1025_g N_A_395_47#_c_1078_n 0.00994068f $X=5.13 $Y=0.56
+ $X2=0 $Y2=0
cc_357 N_A_206_47#_M1028_g N_A_395_47#_c_1078_n 0.00994068f $X=5.65 $Y=0.56
+ $X2=0 $Y2=0
cc_358 N_A_206_47#_c_384_n N_A_395_47#_c_1078_n 0.00125702f $X=5.39 $Y=1.16
+ $X2=0 $Y2=0
cc_359 N_A_206_47#_M1002_g N_A_853_47#_c_1120_n 0.0039189f $X=4.19 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_206_47#_M1008_g N_A_853_47#_c_1120_n 0.0111698f $X=4.66 $Y=0.56 $X2=0
+ $Y2=0
cc_361 N_A_206_47#_M1025_g N_A_853_47#_c_1120_n 0.0111976f $X=5.13 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_206_47#_M1028_g N_A_853_47#_c_1120_n 0.0156905f $X=5.65 $Y=0.56 $X2=0
+ $Y2=0
cc_363 N_A_206_47#_c_350_n N_A_853_47#_c_1120_n 0.00810938f $X=4.415 $Y=1.19
+ $X2=0 $Y2=0
cc_364 N_A_206_47#_c_384_n N_A_853_47#_c_1120_n 0.093932f $X=5.39 $Y=1.16 $X2=0
+ $Y2=0
cc_365 N_A_206_47#_c_343_n N_A_853_47#_c_1120_n 0.010834f $X=5.625 $Y=1.217
+ $X2=0 $Y2=0
cc_366 N_C_M1020_g N_D_M1016_g 0.0230736f $X=8.08 $Y=0.56 $X2=0 $Y2=0
cc_367 N_C_c_482_n N_D_c_555_n 0.0231619f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_368 N_C_c_477_n D 0.00910677f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_369 N_C_c_478_n D 0.00195998f $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_370 N_C_c_478_n N_D_c_553_n 0.0230736f $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_371 N_C_c_479_n N_VPWR_c_629_n 0.0199746f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_372 N_C_c_480_n N_VPWR_c_630_n 0.0052072f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_373 N_C_c_481_n N_VPWR_c_630_n 0.004751f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_374 N_C_c_482_n N_VPWR_c_631_n 0.0052072f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_375 N_C_c_479_n N_VPWR_c_637_n 0.00597712f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_376 N_C_c_480_n N_VPWR_c_637_n 0.00673617f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_377 N_C_c_481_n N_VPWR_c_639_n 0.00597712f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_378 N_C_c_482_n N_VPWR_c_639_n 0.00673617f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_379 N_C_c_479_n N_VPWR_c_622_n 0.0114792f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_380 N_C_c_480_n N_VPWR_c_622_n 0.0118438f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_381 N_C_c_481_n N_VPWR_c_622_n 0.00999457f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_382 N_C_c_482_n N_VPWR_c_622_n 0.011869f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_383 N_C_c_479_n N_Y_c_793_n 0.0139912f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_384 N_C_c_476_n N_Y_c_793_n 0.00729564f $X=6.545 $Y=1.16 $X2=0 $Y2=0
cc_385 N_C_c_477_n N_Y_c_793_n 0.0459683f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_386 N_C_c_478_n N_Y_c_793_n 2.73568e-19 $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_387 N_C_c_479_n N_Y_c_867_n 0.0183309f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_388 N_C_c_480_n N_Y_c_867_n 0.0106251f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_389 N_C_c_481_n N_Y_c_867_n 6.24674e-19 $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_390 N_C_c_480_n N_Y_c_794_n 0.0153933f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_391 N_C_c_481_n N_Y_c_794_n 0.0113962f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_392 N_C_c_477_n N_Y_c_794_n 0.040258f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_393 N_C_c_478_n N_Y_c_794_n 0.00725062f $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_394 N_C_c_480_n N_Y_c_874_n 6.48386e-19 $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_395 N_C_c_481_n N_Y_c_874_n 0.0130707f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_396 N_C_c_482_n N_Y_c_874_n 0.0106251f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_397 N_C_c_482_n N_Y_c_795_n 0.0199153f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_398 N_C_c_478_n N_Y_c_795_n 4.93319e-19 $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_399 N_C_c_482_n N_Y_c_879_n 6.48386e-19 $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_400 N_C_c_479_n N_Y_c_799_n 0.00292783f $X=6.645 $Y=1.41 $X2=0 $Y2=0
cc_401 N_C_c_480_n N_Y_c_799_n 0.00116723f $X=7.115 $Y=1.41 $X2=0 $Y2=0
cc_402 N_C_c_477_n N_Y_c_799_n 0.0305808f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_403 N_C_c_478_n N_Y_c_799_n 0.0074788f $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_404 N_C_c_481_n N_Y_c_800_n 0.00292783f $X=7.585 $Y=1.41 $X2=0 $Y2=0
cc_405 N_C_c_482_n N_Y_c_800_n 0.00116723f $X=8.055 $Y=1.41 $X2=0 $Y2=0
cc_406 N_C_c_477_n N_Y_c_800_n 0.0305808f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_407 N_C_c_478_n N_Y_c_800_n 0.0074788f $X=8.055 $Y=1.217 $X2=0 $Y2=0
cc_408 N_C_M1000_g N_VGND_c_981_n 0.00357877f $X=6.67 $Y=0.56 $X2=0 $Y2=0
cc_409 N_C_M1009_g N_VGND_c_981_n 0.00357877f $X=7.14 $Y=0.56 $X2=0 $Y2=0
cc_410 N_C_M1011_g N_VGND_c_981_n 0.00357877f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_411 N_C_M1020_g N_VGND_c_981_n 0.00357877f $X=8.08 $Y=0.56 $X2=0 $Y2=0
cc_412 N_C_M1000_g N_VGND_c_987_n 0.00668309f $X=6.67 $Y=0.56 $X2=0 $Y2=0
cc_413 N_C_M1009_g N_VGND_c_987_n 0.00548399f $X=7.14 $Y=0.56 $X2=0 $Y2=0
cc_414 N_C_M1011_g N_VGND_c_987_n 0.00548399f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_415 N_C_M1020_g N_VGND_c_987_n 0.00542415f $X=8.08 $Y=0.56 $X2=0 $Y2=0
cc_416 N_C_M1000_g N_A_853_47#_c_1120_n 0.013837f $X=6.67 $Y=0.56 $X2=0 $Y2=0
cc_417 N_C_M1009_g N_A_853_47#_c_1120_n 0.0111698f $X=7.14 $Y=0.56 $X2=0 $Y2=0
cc_418 N_C_M1011_g N_A_853_47#_c_1120_n 0.0111698f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_419 N_C_M1020_g N_A_853_47#_c_1120_n 0.00337098f $X=8.08 $Y=0.56 $X2=0 $Y2=0
cc_420 N_C_c_476_n N_A_853_47#_c_1120_n 0.00896085f $X=6.545 $Y=1.16 $X2=0 $Y2=0
cc_421 N_C_c_477_n N_A_853_47#_c_1120_n 0.143676f $X=7.82 $Y=1.16 $X2=0 $Y2=0
cc_422 N_C_c_478_n N_A_853_47#_c_1120_n 0.00968149f $X=8.055 $Y=1.217 $X2=0
+ $Y2=0
cc_423 N_C_M1000_g N_A_1251_47#_c_1156_n 0.00958923f $X=6.67 $Y=0.56 $X2=0 $Y2=0
cc_424 N_C_M1009_g N_A_1251_47#_c_1156_n 0.00958923f $X=7.14 $Y=0.56 $X2=0 $Y2=0
cc_425 N_C_M1011_g N_A_1251_47#_c_1156_n 0.00951434f $X=7.61 $Y=0.56 $X2=0 $Y2=0
cc_426 N_C_M1020_g N_A_1251_47#_c_1156_n 0.0149383f $X=8.08 $Y=0.56 $X2=0 $Y2=0
cc_427 N_D_c_555_n N_VPWR_c_631_n 0.004751f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_428 N_D_c_556_n N_VPWR_c_632_n 0.0052072f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_429 N_D_c_557_n N_VPWR_c_632_n 0.004751f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_430 N_D_c_558_n N_VPWR_c_634_n 0.00962132f $X=9.935 $Y=1.41 $X2=0 $Y2=0
cc_431 D N_VPWR_c_634_n 0.0207117f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_432 N_D_c_554_n N_VPWR_c_634_n 0.00593966f $X=10.17 $Y=1.16 $X2=0 $Y2=0
cc_433 N_D_c_555_n N_VPWR_c_641_n 0.00597712f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_434 N_D_c_556_n N_VPWR_c_641_n 0.00673617f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_435 N_D_c_557_n N_VPWR_c_647_n 0.00597712f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_436 N_D_c_558_n N_VPWR_c_647_n 0.00673617f $X=9.935 $Y=1.41 $X2=0 $Y2=0
cc_437 N_D_c_555_n N_VPWR_c_622_n 0.0100198f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_438 N_D_c_556_n N_VPWR_c_622_n 0.0118438f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_439 N_D_c_557_n N_VPWR_c_622_n 0.00999457f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_440 N_D_c_558_n N_VPWR_c_622_n 0.0128678f $X=9.935 $Y=1.41 $X2=0 $Y2=0
cc_441 N_D_c_555_n N_Y_c_874_n 6.24674e-19 $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_442 N_D_c_555_n N_Y_c_795_n 0.0113403f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_443 D N_Y_c_795_n 0.0107369f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_444 N_D_c_553_n N_Y_c_795_n 3.10838e-19 $X=10.035 $Y=1.165 $X2=0 $Y2=0
cc_445 N_D_c_555_n N_Y_c_879_n 0.0130707f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_446 N_D_c_556_n N_Y_c_879_n 0.0106251f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_447 N_D_c_557_n N_Y_c_879_n 6.24674e-19 $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_448 N_D_c_556_n N_Y_c_796_n 0.0153933f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_449 N_D_c_557_n N_Y_c_796_n 0.0113962f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_450 D N_Y_c_796_n 0.040258f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_451 N_D_c_553_n N_Y_c_796_n 0.00725062f $X=10.035 $Y=1.165 $X2=0 $Y2=0
cc_452 N_D_c_557_n N_Y_c_797_n 0.00292783f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_453 N_D_c_558_n N_Y_c_797_n 0.00349846f $X=9.935 $Y=1.41 $X2=0 $Y2=0
cc_454 D N_Y_c_797_n 0.0305808f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_455 N_D_c_553_n N_Y_c_797_n 0.0074788f $X=10.035 $Y=1.165 $X2=0 $Y2=0
cc_456 N_D_c_556_n N_Y_c_903_n 6.48386e-19 $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_457 N_D_c_557_n N_Y_c_903_n 0.0130707f $X=9.465 $Y=1.41 $X2=0 $Y2=0
cc_458 N_D_c_558_n N_Y_c_903_n 0.0100147f $X=9.935 $Y=1.41 $X2=0 $Y2=0
cc_459 N_D_c_555_n N_Y_c_801_n 0.00292783f $X=8.525 $Y=1.41 $X2=0 $Y2=0
cc_460 N_D_c_556_n N_Y_c_801_n 0.00116723f $X=8.995 $Y=1.41 $X2=0 $Y2=0
cc_461 D N_Y_c_801_n 0.0305808f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_462 N_D_c_553_n N_Y_c_801_n 0.0074788f $X=10.035 $Y=1.165 $X2=0 $Y2=0
cc_463 N_D_M1016_g N_VGND_c_979_n 0.00312892f $X=8.5 $Y=0.56 $X2=0 $Y2=0
cc_464 N_D_M1018_g N_VGND_c_979_n 0.00908276f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_465 N_D_M1026_g N_VGND_c_979_n 0.00121428f $X=9.44 $Y=0.56 $X2=0 $Y2=0
cc_466 N_D_M1026_g N_VGND_c_980_n 0.00167984f $X=9.44 $Y=0.56 $X2=0 $Y2=0
cc_467 N_D_M1030_g N_VGND_c_980_n 0.0160648f $X=9.91 $Y=0.56 $X2=0 $Y2=0
cc_468 N_D_M1016_g N_VGND_c_981_n 0.00428022f $X=8.5 $Y=0.56 $X2=0 $Y2=0
cc_469 N_D_M1018_g N_VGND_c_983_n 0.00341689f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_470 N_D_M1026_g N_VGND_c_983_n 0.00428022f $X=9.44 $Y=0.56 $X2=0 $Y2=0
cc_471 N_D_M1030_g N_VGND_c_986_n 0.00341689f $X=9.91 $Y=0.56 $X2=0 $Y2=0
cc_472 N_D_M1016_g N_VGND_c_987_n 0.00583939f $X=8.5 $Y=0.56 $X2=0 $Y2=0
cc_473 N_D_M1018_g N_VGND_c_987_n 0.00415805f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_474 N_D_M1026_g N_VGND_c_987_n 0.005943f $X=9.44 $Y=0.56 $X2=0 $Y2=0
cc_475 N_D_M1030_g N_VGND_c_987_n 0.00516698f $X=9.91 $Y=0.56 $X2=0 $Y2=0
cc_476 N_D_M1016_g N_A_853_47#_c_1120_n 4.63093e-19 $X=8.5 $Y=0.56 $X2=0 $Y2=0
cc_477 N_D_M1016_g N_A_1251_47#_c_1160_n 0.0114457f $X=8.5 $Y=0.56 $X2=0 $Y2=0
cc_478 N_D_M1018_g N_A_1251_47#_c_1160_n 0.0102148f $X=8.97 $Y=0.56 $X2=0 $Y2=0
cc_479 N_D_M1026_g N_A_1251_47#_c_1160_n 0.0105988f $X=9.44 $Y=0.56 $X2=0 $Y2=0
cc_480 N_D_M1030_g N_A_1251_47#_c_1160_n 0.01027f $X=9.91 $Y=0.56 $X2=0 $Y2=0
cc_481 D N_A_1251_47#_c_1160_n 0.0867497f $X=10.125 $Y=1.105 $X2=0 $Y2=0
cc_482 N_D_c_553_n N_A_1251_47#_c_1160_n 0.0156419f $X=10.035 $Y=1.165 $X2=0
+ $Y2=0
cc_483 N_VPWR_c_622_n N_Y_M1004_s 0.00439555f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_484 N_VPWR_c_622_n N_Y_M1022_s 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_485 N_VPWR_c_622_n N_Y_M1003_d 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_486 N_VPWR_c_622_n N_Y_M1019_d 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_487 N_VPWR_c_622_n N_Y_M1005_d 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_488 N_VPWR_c_622_n N_Y_M1027_d 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_489 N_VPWR_c_622_n N_Y_M1006_s 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_490 N_VPWR_c_622_n N_Y_M1017_s 0.00231261f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_491 N_VPWR_c_624_n N_Y_c_808_n 0.058597f $X=2.1 $Y=1.66 $X2=0 $Y2=0
cc_492 N_VPWR_c_625_n N_Y_c_808_n 0.048204f $X=3.04 $Y=2 $X2=0 $Y2=0
cc_493 N_VPWR_c_645_n N_Y_c_808_n 0.0187893f $X=2.825 $Y=2.72 $X2=0 $Y2=0
cc_494 N_VPWR_c_622_n N_Y_c_808_n 0.0110885f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_M1010_d N_Y_c_789_n 0.00184299f $X=2.895 $Y=1.485 $X2=0 $Y2=0
cc_496 N_VPWR_c_625_n N_Y_c_789_n 0.0189896f $X=3.04 $Y=2 $X2=0 $Y2=0
cc_497 N_VPWR_c_624_n N_Y_c_790_n 0.0133617f $X=2.1 $Y=1.66 $X2=0 $Y2=0
cc_498 N_VPWR_c_625_n N_Y_c_817_n 0.0490625f $X=3.04 $Y=2 $X2=0 $Y2=0
cc_499 N_VPWR_c_626_n N_Y_c_817_n 0.0223557f $X=3.895 $Y=2.72 $X2=0 $Y2=0
cc_500 N_VPWR_c_627_n N_Y_c_817_n 0.0385613f $X=3.98 $Y=2 $X2=0 $Y2=0
cc_501 N_VPWR_c_622_n N_Y_c_817_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_502 N_VPWR_c_627_n N_Y_c_820_n 0.0470327f $X=3.98 $Y=2 $X2=0 $Y2=0
cc_503 N_VPWR_c_628_n N_Y_c_820_n 0.0385613f $X=4.92 $Y=2 $X2=0 $Y2=0
cc_504 N_VPWR_c_635_n N_Y_c_820_n 0.0223557f $X=4.835 $Y=2.72 $X2=0 $Y2=0
cc_505 N_VPWR_c_622_n N_Y_c_820_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_506 N_VPWR_M1015_s N_Y_c_791_n 0.00180012f $X=4.775 $Y=1.485 $X2=0 $Y2=0
cc_507 N_VPWR_c_628_n N_Y_c_791_n 0.0139097f $X=4.92 $Y=2 $X2=0 $Y2=0
cc_508 N_VPWR_M1034_d N_Y_c_792_n 0.00180012f $X=3.835 $Y=1.485 $X2=0 $Y2=0
cc_509 N_VPWR_c_627_n N_Y_c_792_n 0.0135105f $X=3.98 $Y=2 $X2=0 $Y2=0
cc_510 N_VPWR_c_628_n N_Y_c_848_n 0.0470327f $X=4.92 $Y=2 $X2=0 $Y2=0
cc_511 N_VPWR_c_629_n N_Y_c_848_n 0.0365216f $X=6.255 $Y=2 $X2=0 $Y2=0
cc_512 N_VPWR_c_646_n N_Y_c_848_n 0.0223557f $X=5.825 $Y=2.72 $X2=0 $Y2=0
cc_513 N_VPWR_c_622_n N_Y_c_848_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_514 N_VPWR_M1031_s N_Y_c_793_n 0.015056f $X=5.715 $Y=1.485 $X2=0 $Y2=0
cc_515 N_VPWR_c_629_n N_Y_c_793_n 0.0528236f $X=6.255 $Y=2 $X2=0 $Y2=0
cc_516 N_VPWR_c_629_n N_Y_c_867_n 0.045928f $X=6.255 $Y=2 $X2=0 $Y2=0
cc_517 N_VPWR_c_630_n N_Y_c_867_n 0.0385613f $X=7.35 $Y=2 $X2=0 $Y2=0
cc_518 N_VPWR_c_637_n N_Y_c_867_n 0.0223557f $X=7.265 $Y=2.72 $X2=0 $Y2=0
cc_519 N_VPWR_c_622_n N_Y_c_867_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_520 N_VPWR_M1023_s N_Y_c_794_n 0.00180012f $X=7.205 $Y=1.485 $X2=0 $Y2=0
cc_521 N_VPWR_c_630_n N_Y_c_794_n 0.0139097f $X=7.35 $Y=2 $X2=0 $Y2=0
cc_522 N_VPWR_c_630_n N_Y_c_874_n 0.0470327f $X=7.35 $Y=2 $X2=0 $Y2=0
cc_523 N_VPWR_c_631_n N_Y_c_874_n 0.0385613f $X=8.29 $Y=2 $X2=0 $Y2=0
cc_524 N_VPWR_c_639_n N_Y_c_874_n 0.0223557f $X=8.205 $Y=2.72 $X2=0 $Y2=0
cc_525 N_VPWR_c_622_n N_Y_c_874_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_526 N_VPWR_M1029_s N_Y_c_795_n 0.00180012f $X=8.145 $Y=1.485 $X2=0 $Y2=0
cc_527 N_VPWR_c_631_n N_Y_c_795_n 0.0139097f $X=8.29 $Y=2 $X2=0 $Y2=0
cc_528 N_VPWR_c_631_n N_Y_c_879_n 0.0470327f $X=8.29 $Y=2 $X2=0 $Y2=0
cc_529 N_VPWR_c_632_n N_Y_c_879_n 0.0385613f $X=9.23 $Y=2 $X2=0 $Y2=0
cc_530 N_VPWR_c_641_n N_Y_c_879_n 0.0223557f $X=9.145 $Y=2.72 $X2=0 $Y2=0
cc_531 N_VPWR_c_622_n N_Y_c_879_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_532 N_VPWR_M1012_d N_Y_c_796_n 0.00180012f $X=9.085 $Y=1.485 $X2=0 $Y2=0
cc_533 N_VPWR_c_632_n N_Y_c_796_n 0.0139097f $X=9.23 $Y=2 $X2=0 $Y2=0
cc_534 N_VPWR_c_634_n N_Y_c_797_n 0.0147124f $X=10.17 $Y=1.66 $X2=0 $Y2=0
cc_535 N_VPWR_c_632_n N_Y_c_903_n 0.0470327f $X=9.23 $Y=2 $X2=0 $Y2=0
cc_536 N_VPWR_c_634_n N_Y_c_903_n 0.050728f $X=10.17 $Y=1.66 $X2=0 $Y2=0
cc_537 N_VPWR_c_647_n N_Y_c_903_n 0.0223557f $X=10.085 $Y=2.72 $X2=0 $Y2=0
cc_538 N_VPWR_c_622_n N_Y_c_903_n 0.0140101f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_539 N_VPWR_c_624_n N_A_395_47#_c_1077_n 0.00237022f $X=2.1 $Y=1.66 $X2=0
+ $Y2=0
cc_540 N_Y_M1007_d N_VGND_c_987_n 0.00256987f $X=2.435 $Y=0.235 $X2=0 $Y2=0
cc_541 N_Y_M1033_d N_VGND_c_987_n 0.00256987f $X=3.375 $Y=0.235 $X2=0 $Y2=0
cc_542 N_Y_c_787_n N_A_395_47#_M1032_s 0.00214463f $X=3.665 $Y=0.78 $X2=0 $Y2=0
cc_543 N_Y_c_830_n N_A_395_47#_M1035_s 0.00337005f $X=3.84 $Y=0.905 $X2=0 $Y2=0
cc_544 N_Y_c_787_n N_A_395_47#_c_1077_n 0.0195173f $X=3.665 $Y=0.78 $X2=0 $Y2=0
cc_545 N_Y_M1007_d N_A_395_47#_c_1078_n 0.00401739f $X=2.435 $Y=0.235 $X2=0
+ $Y2=0
cc_546 N_Y_M1033_d N_A_395_47#_c_1078_n 0.00401739f $X=3.375 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_Y_c_787_n N_A_395_47#_c_1078_n 0.0706773f $X=3.665 $Y=0.78 $X2=0 $Y2=0
cc_548 N_Y_c_830_n N_A_395_47#_c_1078_n 0.0199047f $X=3.84 $Y=0.905 $X2=0 $Y2=0
cc_549 N_Y_c_793_n N_A_853_47#_c_1120_n 0.0161561f $X=6.665 $Y=1.555 $X2=0 $Y2=0
cc_550 N_Y_c_795_n N_A_853_47#_c_1120_n 7.56209e-19 $X=8.545 $Y=1.555 $X2=0
+ $Y2=0
cc_551 N_Y_c_830_n N_A_853_47#_c_1120_n 0.0177762f $X=3.84 $Y=0.905 $X2=0 $Y2=0
cc_552 N_Y_c_795_n N_A_1251_47#_c_1166_n 0.00528716f $X=8.545 $Y=1.555 $X2=0
+ $Y2=0
cc_553 N_VGND_c_987_n N_A_395_47#_M1007_s 0.00389984f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_554 N_VGND_c_987_n N_A_395_47#_M1032_s 0.00255381f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_555 N_VGND_c_987_n N_A_395_47#_M1035_s 0.00215227f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_556 N_VGND_c_987_n N_A_395_47#_M1008_d 0.00255381f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_557 N_VGND_c_987_n N_A_395_47#_M1028_d 0.00209344f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_558 N_VGND_c_981_n N_A_395_47#_c_1090_n 0.0119155f $X=8.595 $Y=0 $X2=0 $Y2=0
cc_559 N_VGND_c_987_n N_A_395_47#_c_1090_n 0.00653933f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_560 N_VGND_c_981_n N_A_395_47#_c_1078_n 0.219099f $X=8.595 $Y=0 $X2=0 $Y2=0
cc_561 N_VGND_c_987_n N_A_395_47#_c_1078_n 0.137997f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_562 N_VGND_c_987_n N_A_853_47#_M1002_s 0.00256987f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_563 N_VGND_c_987_n N_A_853_47#_M1025_s 0.00297142f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_564 N_VGND_c_987_n N_A_853_47#_M1000_s 0.00256987f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_565 N_VGND_c_987_n N_A_853_47#_M1011_s 0.00256987f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_566 N_VGND_c_981_n N_A_853_47#_c_1120_n 0.00431692f $X=8.595 $Y=0 $X2=0 $Y2=0
cc_567 N_VGND_c_987_n N_A_853_47#_c_1120_n 0.0135976f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_568 N_VGND_c_987_n N_A_1251_47#_M1000_d 0.00278873f $X=10.35 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_569 N_VGND_c_987_n N_A_1251_47#_M1009_d 0.00255381f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_570 N_VGND_c_987_n N_A_1251_47#_M1020_d 0.00236502f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_571 N_VGND_c_987_n N_A_1251_47#_M1018_d 0.00382975f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_572 N_VGND_c_987_n N_A_1251_47#_M1030_d 0.00468341f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_573 N_VGND_c_981_n N_A_1251_47#_c_1156_n 0.122382f $X=8.595 $Y=0 $X2=0 $Y2=0
cc_574 N_VGND_c_987_n N_A_1251_47#_c_1156_n 0.0762982f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_575 N_VGND_M1016_s N_A_1251_47#_c_1160_n 0.00433058f $X=8.575 $Y=0.235 $X2=0
+ $Y2=0
cc_576 N_VGND_M1026_s N_A_1251_47#_c_1160_n 0.00433058f $X=9.515 $Y=0.235 $X2=0
+ $Y2=0
cc_577 N_VGND_c_979_n N_A_1251_47#_c_1160_n 0.0178569f $X=8.76 $Y=0.4 $X2=0
+ $Y2=0
cc_578 N_VGND_c_980_n N_A_1251_47#_c_1160_n 0.0178569f $X=9.7 $Y=0.4 $X2=0 $Y2=0
cc_579 N_VGND_c_981_n N_A_1251_47#_c_1160_n 0.0029785f $X=8.595 $Y=0 $X2=0 $Y2=0
cc_580 N_VGND_c_983_n N_A_1251_47#_c_1160_n 0.00888403f $X=9.535 $Y=0 $X2=0
+ $Y2=0
cc_581 N_VGND_c_986_n N_A_1251_47#_c_1160_n 0.00646047f $X=10.35 $Y=0 $X2=0
+ $Y2=0
cc_582 N_VGND_c_987_n N_A_1251_47#_c_1160_n 0.0348928f $X=10.35 $Y=0 $X2=0 $Y2=0
cc_583 N_A_395_47#_c_1078_n N_A_853_47#_M1002_s 0.00398854f $X=5.86 $Y=0.4
+ $X2=-0.19 $Y2=-0.24
cc_584 N_A_395_47#_c_1078_n N_A_853_47#_M1025_s 0.00510139f $X=5.86 $Y=0.4 $X2=0
+ $Y2=0
cc_585 N_A_395_47#_M1008_d N_A_853_47#_c_1120_n 0.00214463f $X=4.735 $Y=0.235
+ $X2=0 $Y2=0
cc_586 N_A_395_47#_M1028_d N_A_853_47#_c_1120_n 0.00312742f $X=5.725 $Y=0.235
+ $X2=0 $Y2=0
cc_587 N_A_395_47#_c_1078_n N_A_853_47#_c_1120_n 0.0984028f $X=5.86 $Y=0.4 $X2=0
+ $Y2=0
cc_588 N_A_395_47#_c_1078_n N_A_1251_47#_c_1156_n 0.0163246f $X=5.86 $Y=0.4
+ $X2=0 $Y2=0
cc_589 N_A_853_47#_c_1120_n N_A_1251_47#_M1000_d 0.00505104f $X=7.845 $Y=0.74
+ $X2=-0.19 $Y2=-0.24
cc_590 N_A_853_47#_c_1120_n N_A_1251_47#_M1009_d 0.00214463f $X=7.845 $Y=0.74
+ $X2=0 $Y2=0
cc_591 N_A_853_47#_M1000_s N_A_1251_47#_c_1156_n 0.00401739f $X=6.745 $Y=0.235
+ $X2=0 $Y2=0
cc_592 N_A_853_47#_M1011_s N_A_1251_47#_c_1156_n 0.00401739f $X=7.685 $Y=0.235
+ $X2=0 $Y2=0
cc_593 N_A_853_47#_c_1120_n N_A_1251_47#_c_1156_n 0.0955876f $X=7.845 $Y=0.74
+ $X2=0 $Y2=0
