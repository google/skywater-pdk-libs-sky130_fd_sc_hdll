# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a211oi_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a211oi_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 1.035000 3.305000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.100000 1.035000 1.535000 1.445000 ;
        RECT 0.100000 1.445000 3.975000 1.625000 ;
        RECT 3.595000 1.035000 3.975000 1.445000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.145000 1.035000 5.305000 1.275000 ;
        RECT 4.145000 1.275000 4.960000 1.615000 ;
        RECT 7.300000 0.995000 7.735000 1.325000 ;
        RECT 7.300000 1.325000 7.510000 1.655000 ;
      LAYER mcon ;
        RECT 4.285000 1.445000 4.455000 1.615000 ;
        RECT 7.340000 1.445000 7.510000 1.615000 ;
      LAYER met1 ;
        RECT 4.225000 1.415000 4.515000 1.460000 ;
        RECT 4.225000 1.460000 7.570000 1.600000 ;
        RECT 4.225000 1.600000 4.515000 1.645000 ;
        RECT 7.280000 1.415000 7.570000 1.460000 ;
        RECT 7.280000 1.600000 7.570000 1.645000 ;
    END
  END B1
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.550000 1.035000 7.050000 1.275000 ;
        RECT 6.830000 1.275000 7.050000 1.695000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  1.404000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 0.095000  0.085000 0.395000 0.585000 ;
        RECT 1.000000  0.085000 1.285000 0.525000 ;
        RECT 3.935000  0.085000 4.105000 0.525000 ;
        RECT 4.865000  0.085000 5.195000 0.445000 ;
        RECT 5.815000  0.085000 6.145000 0.445000 ;
        RECT 6.755000  0.085000 7.085000 0.445000 ;
        RECT 7.665000  0.085000 8.070000 0.445000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.160000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 0.515000 2.255000 0.895000 2.635000 ;
        RECT 1.455000 2.275000 1.835000 2.635000 ;
        RECT 2.395000 2.275000 2.775000 2.635000 ;
        RECT 3.335000 2.275000 3.715000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  1.985000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.925000 0.675000 3.680000 0.695000 ;
        RECT 1.925000 0.695000 8.160000 0.825000 ;
        RECT 1.925000 0.825000 7.055000 0.865000 ;
        RECT 4.275000 0.255000 4.645000 0.615000 ;
        RECT 4.275000 0.615000 5.595000 0.625000 ;
        RECT 4.275000 0.625000 8.160000 0.695000 ;
        RECT 5.425000 0.255000 5.595000 0.615000 ;
        RECT 5.720000 1.865000 8.160000 2.085000 ;
        RECT 6.365000 0.255000 6.535000 0.615000 ;
        RECT 6.365000 0.615000 8.160000 0.625000 ;
        RECT 7.680000 1.495000 8.160000 1.865000 ;
        RECT 7.905000 0.825000 8.160000 1.495000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.095000 1.795000 4.105000 2.085000 ;
      RECT 0.095000 2.085000 0.345000 2.465000 ;
      RECT 0.615000 0.530000 0.825000 0.695000 ;
      RECT 0.615000 0.695000 1.755000 0.865000 ;
      RECT 1.115000 2.085000 4.105000 2.105000 ;
      RECT 1.115000 2.105000 1.285000 2.465000 ;
      RECT 1.455000 0.255000 3.715000 0.505000 ;
      RECT 1.455000 0.505000 1.755000 0.695000 ;
      RECT 2.055000 2.105000 2.225000 2.465000 ;
      RECT 2.995000 2.105000 3.165000 2.465000 ;
      RECT 3.935000 2.105000 4.105000 2.255000 ;
      RECT 3.935000 2.255000 8.070000 2.465000 ;
      RECT 4.275000 1.785000 5.460000 2.085000 ;
      RECT 5.130000 1.445000 6.610000 1.695000 ;
      RECT 5.130000 1.695000 5.460000 1.785000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a211oi_4
