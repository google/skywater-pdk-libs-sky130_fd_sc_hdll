* File: sky130_fd_sc_hdll__isobufsrc_8.pex.spice
* Created: Thu Aug 27 19:10:13 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A 1 3 4 6 7 9 10 12 15 19 22
r45 22 23 35.6788 $w=3.58e-07 $l=2.65e-07 $layer=POLY_cond $X=1.015 $Y=1.202
+ $X2=1.28 $Y2=1.202
r46 21 22 27.6006 $w=3.58e-07 $l=2.05e-07 $layer=POLY_cond $X=0.81 $Y=1.202
+ $X2=1.015 $Y2=1.202
r47 20 21 42.4106 $w=3.58e-07 $l=3.15e-07 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.81 $Y2=1.202
r48 18 20 27.6006 $w=3.58e-07 $l=2.05e-07 $layer=POLY_cond $X=0.29 $Y=1.202
+ $X2=0.495 $Y2=1.202
r49 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.29
+ $Y=1.16 $X2=0.29 $Y2=1.16
r50 15 19 4.71454 $w=2.18e-07 $l=9e-08 $layer=LI1_cond $X=0.2 $Y=1.175 $X2=0.29
+ $Y2=1.175
r51 10 23 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.28 $Y=0.995
+ $X2=1.28 $Y2=1.202
r52 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.28 $Y=0.995
+ $X2=1.28 $Y2=0.56
r53 7 22 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.202
r54 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.015 $Y=1.41
+ $X2=1.015 $Y2=1.985
r55 4 21 23.1716 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.81 $Y=0.995
+ $X2=0.81 $Y2=1.202
r56 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.81 $Y=0.995 $X2=0.81
+ $Y2=0.56
r57 1 20 18.8375 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r58 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_117_297# 1 2 7 9 10 12 13 15 16 18
+ 19 21 22 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 57 63
+ 70 74 75 76 93
r174 93 94 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.395 $Y=1.202
+ $X2=5.42 $Y2=1.202
r175 90 91 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.9 $Y=1.202
+ $X2=4.925 $Y2=1.202
r176 89 90 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=4.455 $Y=1.202
+ $X2=4.9 $Y2=1.202
r177 88 89 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.43 $Y=1.202
+ $X2=4.455 $Y2=1.202
r178 87 88 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=3.985 $Y=1.202
+ $X2=4.43 $Y2=1.202
r179 86 87 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.96 $Y=1.202
+ $X2=3.985 $Y2=1.202
r180 85 86 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=3.515 $Y=1.202
+ $X2=3.96 $Y2=1.202
r181 84 85 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.49 $Y=1.202
+ $X2=3.515 $Y2=1.202
r182 83 84 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=3.045 $Y=1.202
+ $X2=3.49 $Y2=1.202
r183 82 83 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.02 $Y=1.202
+ $X2=3.045 $Y2=1.202
r184 81 82 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=2.575 $Y=1.202
+ $X2=3.02 $Y2=1.202
r185 80 81 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.55 $Y=1.202
+ $X2=2.575 $Y2=1.202
r186 77 78 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.08 $Y=1.202
+ $X2=2.105 $Y2=1.202
r187 74 75 7.16311 $w=4.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.62
+ $X2=0.73 $Y2=1.455
r188 71 93 17.6821 $w=3.68e-07 $l=1.35e-07 $layer=POLY_cond $X=5.26 $Y=1.202
+ $X2=5.395 $Y2=1.202
r189 71 91 43.8777 $w=3.68e-07 $l=3.35e-07 $layer=POLY_cond $X=5.26 $Y=1.202
+ $X2=4.925 $Y2=1.202
r190 70 71 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=5.26
+ $Y=1.16 $X2=5.26 $Y2=1.16
r191 68 80 47.1522 $w=3.68e-07 $l=3.6e-07 $layer=POLY_cond $X=2.19 $Y=1.202
+ $X2=2.55 $Y2=1.202
r192 68 78 11.1332 $w=3.68e-07 $l=8.5e-08 $layer=POLY_cond $X=2.19 $Y=1.202
+ $X2=2.105 $Y2=1.202
r193 67 70 162.139 $w=2.08e-07 $l=3.07e-06 $layer=LI1_cond $X=2.19 $Y=1.18
+ $X2=5.26 $Y2=1.18
r194 67 68 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=2.19
+ $Y=1.16 $X2=2.19 $Y2=1.16
r195 65 76 2.52678 $w=2.1e-07 $l=2.57488e-07 $layer=LI1_cond $X=1.235 $Y=1.18
+ $X2=0.98 $Y2=1.175
r196 65 67 50.4372 $w=2.08e-07 $l=9.55e-07 $layer=LI1_cond $X=1.235 $Y=1.18
+ $X2=2.19 $Y2=1.18
r197 61 76 3.91873 $w=2.9e-07 $l=1.42653e-07 $layer=LI1_cond $X=1.055 $Y=1.065
+ $X2=0.98 $Y2=1.175
r198 61 63 21.6083 $w=3.58e-07 $l=6.75e-07 $layer=LI1_cond $X=1.055 $Y=1.065
+ $X2=1.055 $Y2=0.39
r199 59 76 3.91873 $w=2.9e-07 $l=1.92289e-07 $layer=LI1_cond $X=0.835 $Y=1.285
+ $X2=0.98 $Y2=1.175
r200 59 75 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=0.835 $Y=1.285
+ $X2=0.835 $Y2=1.455
r201 55 74 1.34005 $w=4.28e-07 $l=5e-08 $layer=LI1_cond $X=0.73 $Y=1.67 $X2=0.73
+ $Y2=1.62
r202 55 57 16.8846 $w=4.28e-07 $l=6.3e-07 $layer=LI1_cond $X=0.73 $Y=1.67
+ $X2=0.73 $Y2=2.3
r203 52 94 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.42 $Y=0.995
+ $X2=5.42 $Y2=1.202
r204 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.42 $Y=0.995
+ $X2=5.42 $Y2=0.56
r205 49 93 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.395 $Y=1.41
+ $X2=5.395 $Y2=1.202
r206 49 51 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.395 $Y=1.41
+ $X2=5.395 $Y2=1.985
r207 46 91 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.925 $Y=1.41
+ $X2=4.925 $Y2=1.202
r208 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.925 $Y=1.41
+ $X2=4.925 $Y2=1.985
r209 43 90 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=1.202
r210 43 45 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.9 $Y=0.995
+ $X2=4.9 $Y2=0.56
r211 40 89 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.455 $Y2=1.202
r212 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.455 $Y=1.41
+ $X2=4.455 $Y2=1.985
r213 37 88 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=1.202
r214 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.43 $Y=0.995
+ $X2=4.43 $Y2=0.56
r215 34 87 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.985 $Y=1.41
+ $X2=3.985 $Y2=1.202
r216 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.985 $Y=1.41
+ $X2=3.985 $Y2=1.985
r217 31 86 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.96 $Y=0.995
+ $X2=3.96 $Y2=1.202
r218 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.96 $Y=0.995
+ $X2=3.96 $Y2=0.56
r219 28 85 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.515 $Y=1.41
+ $X2=3.515 $Y2=1.202
r220 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.515 $Y=1.41
+ $X2=3.515 $Y2=1.985
r221 25 84 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.49 $Y=0.995
+ $X2=3.49 $Y2=1.202
r222 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.49 $Y=0.995
+ $X2=3.49 $Y2=0.56
r223 22 83 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.045 $Y=1.41
+ $X2=3.045 $Y2=1.202
r224 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.045 $Y=1.41
+ $X2=3.045 $Y2=1.985
r225 19 82 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=1.202
r226 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.02 $Y=0.995
+ $X2=3.02 $Y2=0.56
r227 16 81 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.575 $Y=1.41
+ $X2=2.575 $Y2=1.202
r228 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.575 $Y=1.41
+ $X2=2.575 $Y2=1.985
r229 13 80 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=1.202
r230 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.55 $Y=0.995
+ $X2=2.55 $Y2=0.56
r231 10 78 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.202
r232 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.105 $Y=1.41
+ $X2=2.105 $Y2=1.985
r233 7 77 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=1.202
r234 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.08 $Y=0.995
+ $X2=2.08 $Y2=0.56
r235 2 74 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.62
r236 2 57 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.3
r237 1 63 91 $w=1.7e-07 $l=2.19203e-07 $layer=licon1_NDIFF $count=2 $X=0.885
+ $Y=0.235 $X2=1.04 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%SLEEP 1 3 4 6 7 9 10 12 13 15 16 18 19
+ 21 22 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 68 71 77
r139 71 72 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=9.155 $Y=1.202
+ $X2=9.18 $Y2=1.202
r140 70 71 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=8.685 $Y=1.202
+ $X2=9.155 $Y2=1.202
r141 69 70 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.66 $Y=1.202
+ $X2=8.685 $Y2=1.202
r142 68 77 95.6591 $w=1.98e-07 $l=1.725e-06 $layer=LI1_cond $X=8.645 $Y=1.175
+ $X2=6.92 $Y2=1.175
r143 67 69 1.96467 $w=3.68e-07 $l=1.5e-08 $layer=POLY_cond $X=8.645 $Y=1.202
+ $X2=8.66 $Y2=1.202
r144 67 68 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=8.645
+ $Y=1.16 $X2=8.645 $Y2=1.16
r145 65 67 56.3207 $w=3.68e-07 $l=4.3e-07 $layer=POLY_cond $X=8.215 $Y=1.202
+ $X2=8.645 $Y2=1.202
r146 64 65 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=8.19 $Y=1.202
+ $X2=8.215 $Y2=1.202
r147 63 64 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=7.745 $Y=1.202
+ $X2=8.19 $Y2=1.202
r148 62 63 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.72 $Y=1.202
+ $X2=7.745 $Y2=1.202
r149 61 62 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=7.275 $Y=1.202
+ $X2=7.72 $Y2=1.202
r150 60 61 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=7.25 $Y=1.202
+ $X2=7.275 $Y2=1.202
r151 59 60 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=6.805 $Y=1.202
+ $X2=7.25 $Y2=1.202
r152 58 59 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.78 $Y=1.202
+ $X2=6.805 $Y2=1.202
r153 57 58 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=6.335 $Y=1.202
+ $X2=6.78 $Y2=1.202
r154 56 57 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=6.31 $Y=1.202
+ $X2=6.335 $Y2=1.202
r155 54 56 45.1875 $w=3.68e-07 $l=3.45e-07 $layer=POLY_cond $X=5.965 $Y=1.202
+ $X2=6.31 $Y2=1.202
r156 54 55 36.32 $w=1.7e-07 $l=6.8e-07 $layer=licon1_POLY $count=4 $X=5.965
+ $Y=1.16 $X2=5.965 $Y2=1.16
r157 52 54 13.0978 $w=3.68e-07 $l=1e-07 $layer=POLY_cond $X=5.865 $Y=1.202
+ $X2=5.965 $Y2=1.202
r158 51 52 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.84 $Y=1.202
+ $X2=5.865 $Y2=1.202
r159 49 77 33.2727 $w=1.98e-07 $l=6e-07 $layer=LI1_cond $X=6.32 $Y=1.175
+ $X2=6.92 $Y2=1.175
r160 49 55 19.6864 $w=1.98e-07 $l=3.55e-07 $layer=LI1_cond $X=6.32 $Y=1.175
+ $X2=5.965 $Y2=1.175
r161 46 72 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.18 $Y=0.995
+ $X2=9.18 $Y2=1.202
r162 46 48 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.18 $Y=0.995
+ $X2=9.18 $Y2=0.56
r163 43 71 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=9.155 $Y=1.41
+ $X2=9.155 $Y2=1.202
r164 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.155 $Y=1.41
+ $X2=9.155 $Y2=1.985
r165 40 70 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.685 $Y=1.41
+ $X2=8.685 $Y2=1.202
r166 40 42 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.685 $Y=1.41
+ $X2=8.685 $Y2=1.985
r167 37 69 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.66 $Y2=1.202
r168 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.66 $Y=0.995
+ $X2=8.66 $Y2=0.56
r169 34 65 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=8.215 $Y=1.41
+ $X2=8.215 $Y2=1.202
r170 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.215 $Y=1.41
+ $X2=8.215 $Y2=1.985
r171 31 64 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=8.19 $Y=0.995
+ $X2=8.19 $Y2=1.202
r172 31 33 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=8.19 $Y=0.995
+ $X2=8.19 $Y2=0.56
r173 28 63 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.745 $Y=1.41
+ $X2=7.745 $Y2=1.202
r174 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.745 $Y=1.41
+ $X2=7.745 $Y2=1.985
r175 25 62 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.72 $Y=0.995
+ $X2=7.72 $Y2=1.202
r176 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.72 $Y=0.995
+ $X2=7.72 $Y2=0.56
r177 22 61 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=7.275 $Y=1.41
+ $X2=7.275 $Y2=1.202
r178 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.275 $Y=1.41
+ $X2=7.275 $Y2=1.985
r179 19 60 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=7.25 $Y=0.995
+ $X2=7.25 $Y2=1.202
r180 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=7.25 $Y=0.995
+ $X2=7.25 $Y2=0.56
r181 16 59 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.805 $Y=1.41
+ $X2=6.805 $Y2=1.202
r182 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.805 $Y=1.41
+ $X2=6.805 $Y2=1.985
r183 13 58 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.78 $Y2=1.202
r184 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.78 $Y=0.995
+ $X2=6.78 $Y2=0.56
r185 10 57 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.335 $Y=1.41
+ $X2=6.335 $Y2=1.202
r186 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.335 $Y=1.41
+ $X2=6.335 $Y2=1.985
r187 7 56 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.31 $Y=0.995
+ $X2=6.31 $Y2=1.202
r188 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.31 $Y=0.995
+ $X2=6.31 $Y2=0.56
r189 4 52 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.865 $Y=1.41
+ $X2=5.865 $Y2=1.202
r190 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.865 $Y=1.41
+ $X2=5.865 $Y2=1.985
r191 1 51 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.84 $Y=0.995
+ $X2=5.84 $Y2=1.202
r192 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.84 $Y=0.995
+ $X2=5.84 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VPWR 1 2 3 4 5 6 19 21 27 33 37 41 45
+ 48 49 51 52 54 55 57 58 60 61 62 84 85
r124 84 85 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r125 82 85 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=9.43 $Y2=2.72
r126 81 84 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=9.43 $Y2=2.72
r127 81 82 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r128 79 82 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r130 76 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r131 75 76 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r132 73 76 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r133 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r134 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r135 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r136 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r137 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r138 64 88 3.75277 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r139 64 66 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=1.15 $Y2=2.72
r140 62 67 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r141 62 88 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r142 60 78 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=4.83 $Y2=2.72
r143 60 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.035 $Y=2.72
+ $X2=5.16 $Y2=2.72
r144 59 81 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.29 $Y2=2.72
r145 59 61 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.285 $Y=2.72
+ $X2=5.16 $Y2=2.72
r146 57 75 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=3.91 $Y2=2.72
r147 57 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.095 $Y=2.72
+ $X2=4.22 $Y2=2.72
r148 56 78 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=4.83 $Y2=2.72
r149 56 58 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.345 $Y=2.72
+ $X2=4.22 $Y2=2.72
r150 54 72 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=2.99 $Y2=2.72
r151 54 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=3.28 $Y2=2.72
r152 53 75 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=3.405 $Y=2.72
+ $X2=3.91 $Y2=2.72
r153 53 55 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.405 $Y=2.72
+ $X2=3.28 $Y2=2.72
r154 51 69 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.07 $Y2=2.72
r155 51 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.215 $Y=2.72
+ $X2=2.34 $Y2=2.72
r156 50 72 34.2513 $w=1.68e-07 $l=5.25e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.99 $Y2=2.72
r157 50 52 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.465 $Y=2.72
+ $X2=2.34 $Y2=2.72
r158 48 66 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.15 $Y2=2.72
r159 48 49 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=1.312 $Y2=2.72
r160 47 69 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=2.07 $Y2=2.72
r161 47 49 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=1.46 $Y=2.72
+ $X2=1.312 $Y2=2.72
r162 43 61 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.16 $Y=2.635
+ $X2=5.16 $Y2=2.72
r163 43 45 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=5.16 $Y=2.635
+ $X2=5.16 $Y2=2
r164 39 58 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.22 $Y=2.635
+ $X2=4.22 $Y2=2.72
r165 39 41 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.22 $Y=2.635
+ $X2=4.22 $Y2=2
r166 35 55 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.28 $Y=2.635
+ $X2=3.28 $Y2=2.72
r167 35 37 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.28 $Y=2.635
+ $X2=3.28 $Y2=2
r168 31 52 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.34 $Y=2.635
+ $X2=2.34 $Y2=2.72
r169 31 33 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.34 $Y=2.635
+ $X2=2.34 $Y2=2
r170 27 30 27.3461 $w=2.93e-07 $l=7e-07 $layer=LI1_cond $X=1.312 $Y=1.64
+ $X2=1.312 $Y2=2.34
r171 25 49 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.312 $Y=2.635
+ $X2=1.312 $Y2=2.72
r172 25 30 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=1.312 $Y=2.635
+ $X2=1.312 $Y2=2.34
r173 21 24 36.6686 $w=2.18e-07 $l=7e-07 $layer=LI1_cond $X=0.235 $Y=1.64
+ $X2=0.235 $Y2=2.34
r174 19 88 3.21046 $w=2.2e-07 $l=1.12161e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.172 $Y2=2.72
r175 19 24 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.235 $Y=2.635
+ $X2=0.235 $Y2=2.34
r176 6 45 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.015
+ $Y=1.485 $X2=5.16 $Y2=2
r177 5 41 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.075
+ $Y=1.485 $X2=4.22 $Y2=2
r178 4 37 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.135
+ $Y=1.485 $X2=3.28 $Y2=2
r179 3 33 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.195
+ $Y=1.485 $X2=2.34 $Y2=2
r180 2 30 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=2.34
r181 2 27 400 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.105
+ $Y=1.485 $X2=1.25 $Y2=1.64
r182 1 24 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r183 1 21 400 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.64
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%A_345_297# 1 2 3 4 5 6 7 8 9 28 30 32
+ 36 38 42 44 48 50 52 53 54 58 60 64 66 70 72 76 81 83 85 90 91 92
r104 74 76 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=9.39 $Y=2.295
+ $X2=9.39 $Y2=1.96
r105 73 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.575 $Y=2.38
+ $X2=8.45 $Y2=2.38
r106 72 74 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=9.265 $Y=2.38
+ $X2=9.39 $Y2=2.295
r107 72 73 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=9.265 $Y=2.38
+ $X2=8.575 $Y2=2.38
r108 68 92 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=2.295
+ $X2=8.45 $Y2=2.38
r109 68 70 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=8.45 $Y=2.295
+ $X2=8.45 $Y2=1.96
r110 67 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.635 $Y=2.38
+ $X2=7.51 $Y2=2.38
r111 66 92 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.325 $Y=2.38
+ $X2=8.45 $Y2=2.38
r112 66 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.325 $Y=2.38
+ $X2=7.635 $Y2=2.38
r113 62 91 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=2.295
+ $X2=7.51 $Y2=2.38
r114 62 64 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=7.51 $Y=2.295
+ $X2=7.51 $Y2=1.96
r115 61 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.695 $Y=2.38
+ $X2=6.57 $Y2=2.38
r116 60 91 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.385 $Y=2.38
+ $X2=7.51 $Y2=2.38
r117 60 61 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.385 $Y=2.38
+ $X2=6.695 $Y2=2.38
r118 56 90 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=2.295
+ $X2=6.57 $Y2=2.38
r119 56 58 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.57 $Y=2.295
+ $X2=6.57 $Y2=1.96
r120 55 89 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.755 $Y=2.38
+ $X2=5.63 $Y2=2.38
r121 54 90 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.445 $Y=2.38
+ $X2=6.57 $Y2=2.38
r122 54 55 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.445 $Y=2.38
+ $X2=5.755 $Y2=2.38
r123 53 89 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=2.295
+ $X2=5.63 $Y2=2.38
r124 52 87 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=5.63 $Y=1.665
+ $X2=5.63 $Y2=1.56
r125 52 53 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=5.63 $Y=1.665
+ $X2=5.63 $Y2=2.295
r126 51 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.815 $Y=1.56
+ $X2=4.69 $Y2=1.56
r127 50 87 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=5.505 $Y=1.56
+ $X2=5.63 $Y2=1.56
r128 50 51 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=5.505 $Y=1.56
+ $X2=4.815 $Y2=1.56
r129 46 85 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.69 $Y=1.665
+ $X2=4.69 $Y2=1.56
r130 46 48 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=4.69 $Y=1.665
+ $X2=4.69 $Y2=2.3
r131 45 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.875 $Y=1.56
+ $X2=3.75 $Y2=1.56
r132 44 85 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.565 $Y=1.56
+ $X2=4.69 $Y2=1.56
r133 44 45 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=4.565 $Y=1.56
+ $X2=3.875 $Y2=1.56
r134 40 83 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=3.75 $Y=1.665
+ $X2=3.75 $Y2=1.56
r135 40 42 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=3.75 $Y=1.665
+ $X2=3.75 $Y2=2.3
r136 39 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.935 $Y=1.56
+ $X2=2.81 $Y2=1.56
r137 38 83 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.625 $Y=1.56
+ $X2=3.75 $Y2=1.56
r138 38 39 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=3.625 $Y=1.56
+ $X2=2.935 $Y2=1.56
r139 34 81 0.72291 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=2.81 $Y=1.665
+ $X2=2.81 $Y2=1.56
r140 34 36 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=2.81 $Y=1.665
+ $X2=2.81 $Y2=2.3
r141 33 79 4.35048 $w=2.1e-07 $l=1.6e-07 $layer=LI1_cond $X=1.995 $Y=1.56
+ $X2=1.835 $Y2=1.56
r142 32 81 5.95752 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.685 $Y=1.56
+ $X2=2.81 $Y2=1.56
r143 32 33 36.4416 $w=2.08e-07 $l=6.9e-07 $layer=LI1_cond $X=2.685 $Y=1.56
+ $X2=1.995 $Y2=1.56
r144 28 79 2.855 $w=3.2e-07 $l=1.05e-07 $layer=LI1_cond $X=1.835 $Y=1.665
+ $X2=1.835 $Y2=1.56
r145 28 30 22.8688 $w=3.18e-07 $l=6.35e-07 $layer=LI1_cond $X=1.835 $Y=1.665
+ $X2=1.835 $Y2=2.3
r146 9 76 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=9.245
+ $Y=1.485 $X2=9.39 $Y2=1.96
r147 8 70 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=8.305
+ $Y=1.485 $X2=8.45 $Y2=1.96
r148 7 64 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=7.365
+ $Y=1.485 $X2=7.51 $Y2=1.96
r149 6 58 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.425
+ $Y=1.485 $X2=6.57 $Y2=1.96
r150 5 89 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.485 $X2=5.63 $Y2=2.3
r151 5 87 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.485
+ $Y=1.485 $X2=5.63 $Y2=1.62
r152 4 85 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.485 $X2=4.69 $Y2=1.62
r153 4 48 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.545
+ $Y=1.485 $X2=4.69 $Y2=2.3
r154 3 83 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.485 $X2=3.75 $Y2=1.62
r155 3 42 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.605
+ $Y=1.485 $X2=3.75 $Y2=2.3
r156 2 81 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.81 $Y2=1.62
r157 2 36 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.665
+ $Y=1.485 $X2=2.81 $Y2=2.3
r158 1 79 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.485 $X2=1.87 $Y2=1.62
r159 1 30 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.725
+ $Y=1.485 $X2=1.87 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%X 1 2 3 4 5 6 7 8 9 10 11 12 39 41 42
+ 45 47 51 53 57 59 63 67 69 70 71 75 79 81 83 87 91 93 95 99 101 102 103 104
+ 105 106 107 108 110 113
r222 112 113 9.96117 $w=6.83e-07 $l=5.4e-07 $layer=LI1_cond $X=9.307 $Y=0.905
+ $X2=9.307 $Y2=1.445
r223 110 112 12.2 $w=3.87e-07 $l=5.76914e-07 $layer=LI1_cond $X=8.92 $Y=0.49
+ $X2=9.307 $Y2=0.905
r224 97 113 2.52089 $w=3.82e-07 $l=2.995e-07 $layer=LI1_cond $X=8.92 $Y=1.615
+ $X2=9.18 $Y2=1.53
r225 97 99 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.92 $Y=1.615
+ $X2=8.92 $Y2=1.62
r226 96 107 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=8.145 $Y=0.815
+ $X2=7.955 $Y2=0.815
r227 95 110 10.2957 $w=3.87e-07 $l=4.18927e-07 $layer=LI1_cond $X=8.705 $Y=0.815
+ $X2=8.92 $Y2=0.49
r228 95 96 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=8.705 $Y=0.815
+ $X2=8.145 $Y2=0.815
r229 94 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.105 $Y=1.53
+ $X2=7.98 $Y2=1.53
r230 93 113 4.37228 $w=1.7e-07 $l=3.85e-07 $layer=LI1_cond $X=8.795 $Y=1.53
+ $X2=9.18 $Y2=1.53
r231 93 94 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=8.795 $Y=1.53
+ $X2=8.105 $Y2=1.53
r232 89 108 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.98 $Y=1.615
+ $X2=7.98 $Y2=1.53
r233 89 91 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=7.98 $Y=1.615
+ $X2=7.98 $Y2=1.62
r234 85 107 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.955 $Y=0.725
+ $X2=7.955 $Y2=0.815
r235 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.955 $Y=0.725
+ $X2=7.955 $Y2=0.39
r236 84 105 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.205 $Y=0.815
+ $X2=7.015 $Y2=0.815
r237 83 107 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=7.765 $Y=0.815
+ $X2=7.955 $Y2=0.815
r238 83 84 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=7.765 $Y=0.815
+ $X2=7.205 $Y2=0.815
r239 82 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.165 $Y=1.53
+ $X2=7.04 $Y2=1.53
r240 81 108 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.855 $Y=1.53
+ $X2=7.98 $Y2=1.53
r241 81 82 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=7.855 $Y=1.53
+ $X2=7.165 $Y2=1.53
r242 77 106 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.04 $Y=1.615
+ $X2=7.04 $Y2=1.53
r243 77 79 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=7.04 $Y=1.615
+ $X2=7.04 $Y2=1.62
r244 73 105 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=7.015 $Y=0.725
+ $X2=7.015 $Y2=0.815
r245 73 75 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.015 $Y=0.725
+ $X2=7.015 $Y2=0.39
r246 72 104 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.265 $Y=0.815
+ $X2=6.075 $Y2=0.815
r247 71 105 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=6.825 $Y=0.815
+ $X2=7.015 $Y2=0.815
r248 71 72 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.825 $Y=0.815
+ $X2=6.265 $Y2=0.815
r249 69 106 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.915 $Y=1.53
+ $X2=7.04 $Y2=1.53
r250 69 70 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=6.915 $Y=1.53
+ $X2=6.225 $Y2=1.53
r251 65 70 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.1 $Y=1.615
+ $X2=6.225 $Y2=1.53
r252 65 67 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=6.1 $Y=1.615 $X2=6.1
+ $Y2=1.62
r253 61 104 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=6.075 $Y=0.725
+ $X2=6.075 $Y2=0.815
r254 61 63 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.075 $Y=0.725
+ $X2=6.075 $Y2=0.39
r255 60 103 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.325 $Y=0.815
+ $X2=5.135 $Y2=0.815
r256 59 104 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=5.885 $Y=0.815
+ $X2=6.075 $Y2=0.815
r257 59 60 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.885 $Y=0.815
+ $X2=5.325 $Y2=0.815
r258 55 103 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.135 $Y=0.725
+ $X2=5.135 $Y2=0.815
r259 55 57 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.135 $Y=0.725
+ $X2=5.135 $Y2=0.39
r260 54 102 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.385 $Y=0.815
+ $X2=4.195 $Y2=0.815
r261 53 103 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.945 $Y=0.815
+ $X2=5.135 $Y2=0.815
r262 53 54 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.945 $Y=0.815
+ $X2=4.385 $Y2=0.815
r263 49 102 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.195 $Y=0.725
+ $X2=4.195 $Y2=0.815
r264 49 51 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.195 $Y=0.725
+ $X2=4.195 $Y2=0.39
r265 48 101 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.445 $Y=0.815
+ $X2=3.255 $Y2=0.815
r266 47 102 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=4.005 $Y=0.815
+ $X2=4.195 $Y2=0.815
r267 47 48 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=4.005 $Y=0.815
+ $X2=3.445 $Y2=0.815
r268 43 101 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=3.255 $Y=0.725
+ $X2=3.255 $Y2=0.815
r269 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.255 $Y=0.725
+ $X2=3.255 $Y2=0.39
r270 41 101 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=3.065 $Y=0.815
+ $X2=3.255 $Y2=0.815
r271 41 42 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=3.065 $Y=0.815
+ $X2=2.505 $Y2=0.815
r272 37 42 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=2.315 $Y=0.725
+ $X2=2.505 $Y2=0.815
r273 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.315 $Y=0.725
+ $X2=2.315 $Y2=0.39
r274 12 99 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=8.775
+ $Y=1.485 $X2=8.92 $Y2=1.62
r275 11 91 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=7.835
+ $Y=1.485 $X2=7.98 $Y2=1.62
r276 10 79 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=6.895
+ $Y=1.485 $X2=7.04 $Y2=1.62
r277 9 67 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=5.955
+ $Y=1.485 $X2=6.1 $Y2=1.62
r278 8 110 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=8.735
+ $Y=0.235 $X2=8.92 $Y2=0.39
r279 7 87 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=7.795
+ $Y=0.235 $X2=7.98 $Y2=0.39
r280 6 75 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=6.855
+ $Y=0.235 $X2=7.04 $Y2=0.39
r281 5 63 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.915
+ $Y=0.235 $X2=6.1 $Y2=0.39
r282 4 57 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.975
+ $Y=0.235 $X2=5.16 $Y2=0.39
r283 3 51 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.035
+ $Y=0.235 $X2=4.22 $Y2=0.39
r284 2 45 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.095
+ $Y=0.235 $X2=3.28 $Y2=0.39
r285 1 39 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.155
+ $Y=0.235 $X2=2.34 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__ISOBUFSRC_8%VGND 1 2 3 4 5 6 7 8 9 10 33 37 41 45
+ 49 53 57 61 65 67 69 72 73 75 76 78 79 81 82 84 85 87 88 90 91 93 94 95 101
+ 127 132 136
r165 135 136 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r166 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r167 130 136 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=0
+ $X2=9.43 $Y2=0
r168 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=0
+ $X2=8.97 $Y2=0
r169 127 135 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=9.482 $Y2=0
r170 127 129 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=9.305 $Y=0
+ $X2=8.97 $Y2=0
r171 126 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=8.97 $Y2=0
r172 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r173 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r174 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r175 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=7.13 $Y2=0
r176 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r177 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=6.21 $Y2=0
r178 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r179 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.29 $Y2=0
r180 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r181 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=4.37 $Y2=0
r182 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r183 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.45 $Y2=0
r184 108 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=1.61 $Y2=0
r185 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0
+ $X2=2.53 $Y2=0
r186 105 132 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.955 $Y=0
+ $X2=1.7 $Y2=0
r187 105 107 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=1.955 $Y=0
+ $X2=2.53 $Y2=0
r188 104 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=1.61 $Y2=0
r189 103 104 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r190 101 132 11.4275 $w=1.7e-07 $l=2.55e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=1.7 $Y2=0
r191 101 103 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.445 $Y=0
+ $X2=1.15 $Y2=0
r192 95 104 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r193 95 98 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r194 93 125 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.365 $Y=0
+ $X2=8.05 $Y2=0
r195 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.365 $Y=0 $X2=8.45
+ $Y2=0
r196 92 129 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=8.535 $Y=0
+ $X2=8.97 $Y2=0
r197 92 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.535 $Y=0 $X2=8.45
+ $Y2=0
r198 90 122 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.425 $Y=0
+ $X2=7.13 $Y2=0
r199 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.425 $Y=0 $X2=7.51
+ $Y2=0
r200 89 125 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=7.595 $Y=0
+ $X2=8.05 $Y2=0
r201 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.595 $Y=0 $X2=7.51
+ $Y2=0
r202 87 119 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=6.485 $Y=0
+ $X2=6.21 $Y2=0
r203 87 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=0 $X2=6.57
+ $Y2=0
r204 86 122 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=6.655 $Y=0
+ $X2=7.13 $Y2=0
r205 86 88 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.655 $Y=0 $X2=6.57
+ $Y2=0
r206 84 116 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=0
+ $X2=5.29 $Y2=0
r207 84 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.545 $Y=0 $X2=5.63
+ $Y2=0
r208 83 119 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=5.715 $Y=0
+ $X2=6.21 $Y2=0
r209 83 85 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.715 $Y=0 $X2=5.63
+ $Y2=0
r210 81 113 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=4.605 $Y=0
+ $X2=4.37 $Y2=0
r211 81 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.605 $Y=0 $X2=4.69
+ $Y2=0
r212 80 116 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=4.775 $Y=0
+ $X2=5.29 $Y2=0
r213 80 82 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.775 $Y=0 $X2=4.69
+ $Y2=0
r214 78 110 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=3.665 $Y=0
+ $X2=3.45 $Y2=0
r215 78 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.665 $Y=0 $X2=3.75
+ $Y2=0
r216 77 113 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.835 $Y=0
+ $X2=4.37 $Y2=0
r217 77 79 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.835 $Y=0 $X2=3.75
+ $Y2=0
r218 75 107 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=2.725 $Y=0
+ $X2=2.53 $Y2=0
r219 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.725 $Y=0 $X2=2.81
+ $Y2=0
r220 74 110 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.895 $Y=0
+ $X2=3.45 $Y2=0
r221 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.895 $Y=0 $X2=2.81
+ $Y2=0
r222 72 98 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.485 $Y=0
+ $X2=0.23 $Y2=0
r223 72 73 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.485 $Y=0 $X2=0.595
+ $Y2=0
r224 71 103 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=1.15 $Y2=0
r225 71 73 6.36606 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=0.705 $Y=0 $X2=0.595
+ $Y2=0
r226 67 135 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.482 $Y2=0
r227 67 69 13.0183 $w=2.68e-07 $l=3.05e-07 $layer=LI1_cond $X=9.44 $Y=0.085
+ $X2=9.44 $Y2=0.39
r228 63 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0
r229 63 65 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.45 $Y=0.085
+ $X2=8.45 $Y2=0.39
r230 59 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0
r231 59 61 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=7.51 $Y=0.085
+ $X2=7.51 $Y2=0.39
r232 55 88 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0
r233 55 57 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.57 $Y=0.085
+ $X2=6.57 $Y2=0.39
r234 51 85 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0
r235 51 53 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.63 $Y=0.085
+ $X2=5.63 $Y2=0.39
r236 47 82 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.69 $Y=0.085
+ $X2=4.69 $Y2=0
r237 47 49 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.69 $Y=0.085
+ $X2=4.69 $Y2=0.39
r238 43 79 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0
r239 43 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.75 $Y=0.085
+ $X2=3.75 $Y2=0.39
r240 39 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0
r241 39 41 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.81 $Y=0.085
+ $X2=2.81 $Y2=0.39
r242 35 132 2.12513 $w=5.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0
r243 35 37 7.15302 $w=5.08e-07 $l=3.05e-07 $layer=LI1_cond $X=1.7 $Y=0.085
+ $X2=1.7 $Y2=0.39
r244 31 73 0.432806 $w=2.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.595 $Y=0.085
+ $X2=0.595 $Y2=0
r245 31 33 15.9771 $w=2.18e-07 $l=3.05e-07 $layer=LI1_cond $X=0.595 $Y=0.085
+ $X2=0.595 $Y2=0.39
r246 10 69 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=9.255
+ $Y=0.235 $X2=9.39 $Y2=0.39
r247 9 65 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=8.265
+ $Y=0.235 $X2=8.45 $Y2=0.39
r248 8 61 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=7.325
+ $Y=0.235 $X2=7.51 $Y2=0.39
r249 7 57 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=6.385
+ $Y=0.235 $X2=6.57 $Y2=0.39
r250 6 53 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.495
+ $Y=0.235 $X2=5.63 $Y2=0.39
r251 5 49 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=4.505
+ $Y=0.235 $X2=4.69 $Y2=0.39
r252 4 45 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.565
+ $Y=0.235 $X2=3.75 $Y2=0.39
r253 3 41 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.81 $Y2=0.39
r254 2 37 45.5 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_NDIFF $count=4 $X=1.355
+ $Y=0.235 $X2=1.87 $Y2=0.39
r255 1 33 91 $w=1.7e-07 $l=2.61247e-07 $layer=licon1_NDIFF $count=2 $X=0.375
+ $Y=0.235 $X2=0.57 $Y2=0.39
.ends

