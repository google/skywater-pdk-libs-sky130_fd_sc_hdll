* File: sky130_fd_sc_hdll__and4b_4.pex.spice
* Created: Wed Sep  2 08:23:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%A_N 2 3 5 8 10 11 12 17
c40 8 0 1.33735e-19 $X=0.52 $Y=0.445
c41 2 0 1.69423e-19 $X=0.495 $Y=1.89
r42 17 20 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.16
+ $X2=0.55 $Y2=1.325
r43 17 19 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.55 $Y=1.16
+ $X2=0.55 $Y2=0.995
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.525
+ $Y=1.16 $X2=0.525 $Y2=1.16
r45 11 12 9.79577 $w=3.98e-07 $l=3.4e-07 $layer=LI1_cond $X=0.64 $Y=1.19
+ $X2=0.64 $Y2=1.53
r46 11 18 0.864332 $w=3.98e-07 $l=3e-08 $layer=LI1_cond $X=0.64 $Y=1.19 $X2=0.64
+ $Y2=1.16
r47 10 18 8.93143 $w=3.98e-07 $l=3.1e-07 $layer=LI1_cond $X=0.64 $Y=0.85
+ $X2=0.64 $Y2=1.16
r48 8 19 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.445
+ $X2=0.52 $Y2=0.995
r49 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r50 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r51 2 20 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%A_184_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 43 44 45 51 52 54 64
c123 34 0 6.1784e-20 $X=2.53 $Y=1.16
r124 64 65 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=2.405 $Y=1.202
+ $X2=2.43 $Y2=1.202
r125 61 62 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=1.935 $Y=1.202
+ $X2=1.96 $Y2=1.202
r126 58 59 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=1.465 $Y=1.202
+ $X2=1.49 $Y2=1.202
r127 57 58 58.1274 $w=3.69e-07 $l=4.45e-07 $layer=POLY_cond $X=1.02 $Y=1.202
+ $X2=1.465 $Y2=1.202
r128 56 57 3.26558 $w=3.69e-07 $l=2.5e-08 $layer=POLY_cond $X=0.995 $Y=1.202
+ $X2=1.02 $Y2=1.202
r129 52 54 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.53 $Y=0.725
+ $X2=4.735 $Y2=0.725
r130 50 52 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.445 $Y=0.81
+ $X2=4.53 $Y2=0.725
r131 50 51 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=4.445 $Y=0.81
+ $X2=4.445 $Y2=1.545
r132 47 49 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=3.255 $Y=1.63
+ $X2=4.28 $Y2=1.63
r133 45 47 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=2.7 $Y=1.63
+ $X2=3.255 $Y2=1.63
r134 44 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.36 $Y=1.63
+ $X2=4.445 $Y2=1.545
r135 44 49 5.21925 $w=1.68e-07 $l=8e-08 $layer=LI1_cond $X=4.36 $Y=1.63 $X2=4.28
+ $Y2=1.63
r136 43 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.615 $Y=1.545
+ $X2=2.7 $Y2=1.63
r137 42 43 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.615 $Y=1.325
+ $X2=2.615 $Y2=1.545
r138 41 64 7.8374 $w=3.69e-07 $l=6e-08 $layer=POLY_cond $X=2.345 $Y=1.202
+ $X2=2.405 $Y2=1.202
r139 41 62 50.29 $w=3.69e-07 $l=3.85e-07 $layer=POLY_cond $X=2.345 $Y=1.202
+ $X2=1.96 $Y2=1.202
r140 40 41 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.345
+ $Y=1.16 $X2=2.345 $Y2=1.16
r141 37 61 41.7995 $w=3.69e-07 $l=3.2e-07 $layer=POLY_cond $X=1.615 $Y=1.202
+ $X2=1.935 $Y2=1.202
r142 37 59 16.3279 $w=3.69e-07 $l=1.25e-07 $layer=POLY_cond $X=1.615 $Y=1.202
+ $X2=1.49 $Y2=1.202
r143 36 40 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=1.615 $Y=1.16
+ $X2=2.345 $Y2=1.16
r144 36 37 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.615
+ $Y=1.16 $X2=1.615 $Y2=1.16
r145 34 42 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.615 $Y2=1.325
r146 34 40 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=2.53 $Y=1.16
+ $X2=2.345 $Y2=1.16
r147 31 65 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.202
r148 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.43 $Y=1.41
+ $X2=2.43 $Y2=1.985
r149 28 64 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.405 $Y=0.995
+ $X2=2.405 $Y2=1.202
r150 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.405 $Y=0.995
+ $X2=2.405 $Y2=0.56
r151 25 62 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.202
r152 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.96 $Y=1.41
+ $X2=1.96 $Y2=1.985
r153 22 61 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.935 $Y=0.995
+ $X2=1.935 $Y2=1.202
r154 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.935 $Y=0.995
+ $X2=1.935 $Y2=0.56
r155 19 59 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.202
r156 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.985
r157 16 58 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=1.202
r158 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=0.56
r159 13 57 19.55 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.202
r160 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.02 $Y=1.41
+ $X2=1.02 $Y2=1.985
r161 10 56 23.9013 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=1.202
r162 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.995 $Y=0.995
+ $X2=0.995 $Y2=0.56
r163 3 49 600 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_PDIFF $count=1 $X=4.11
+ $Y=1.485 $X2=4.28 $Y2=1.63
r164 2 47 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.11
+ $Y=1.485 $X2=3.255 $Y2=1.63
r165 1 54 182 $w=1.7e-07 $l=5.53399e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.235 $X2=4.735 $Y2=0.725
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%D 1 3 4 6 7 15
c28 15 0 1.24891e-19 $X=2.995 $Y=1.19
c29 1 0 1.02236e-19 $X=3.02 $Y=1.41
r30 7 15 1.3969 $w=3.28e-07 $l=4e-08 $layer=LI1_cond $X=2.955 $Y=1.16 $X2=2.995
+ $Y2=1.16
r31 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r32 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.045 $Y=0.995
+ $X2=2.96 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.045 $Y=0.995
+ $X2=3.045 $Y2=0.56
r34 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=3.02 $Y=1.41
+ $X2=2.96 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.02 $Y=1.41 $X2=3.02
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%C 1 3 4 6 7 8
c29 7 0 6.1784e-20 $X=3.455 $Y=0.85
r30 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.465
+ $Y=1.16 $X2=3.465 $Y2=1.16
r31 7 8 11.5244 $w=3.08e-07 $l=3.1e-07 $layer=LI1_cond $X=3.485 $Y=0.85
+ $X2=3.485 $Y2=1.16
r32 4 12 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.515 $Y=0.995
+ $X2=3.49 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.515 $Y=0.995
+ $X2=3.515 $Y2=0.56
r34 1 12 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=3.49 $Y=1.41
+ $X2=3.49 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=1.41 $X2=3.49
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%B 1 3 4 6 7 8
r35 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.055
+ $Y=1.16 $X2=4.055 $Y2=1.16
r36 8 13 0.909823 $w=3.78e-07 $l=3e-08 $layer=LI1_cond $X=4 $Y=1.19 $X2=4
+ $Y2=1.16
r37 7 13 9.40151 $w=3.78e-07 $l=3.1e-07 $layer=LI1_cond $X=4 $Y=0.85 $X2=4
+ $Y2=1.16
r38 4 12 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=4.02 $Y=1.41
+ $X2=4.08 $Y2=1.16
r39 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.02 $Y=1.41 $X2=4.02
+ $Y2=1.985
r40 1 12 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=4.08 $Y2=1.16
r41 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.995 $Y=0.995
+ $X2=3.995 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%A_27_47# 1 2 7 9 10 12 14 17 19 23 27 30
+ 32
r82 31 32 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.525 $Y=1.202
+ $X2=4.55 $Y2=1.202
r83 27 29 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.42
+ $X2=0.215 $Y2=0.585
r84 24 32 33.0137 $w=3.65e-07 $l=2.5e-07 $layer=POLY_cond $X=4.8 $Y=1.202
+ $X2=4.55 $Y2=1.202
r85 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.8
+ $Y=1.16 $X2=4.8 $Y2=1.16
r86 21 23 49.2567 $w=1.68e-07 $l=7.55e-07 $layer=LI1_cond $X=4.8 $Y=1.915
+ $X2=4.8 $Y2=1.16
r87 20 30 2.24312 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.345 $Y=2 $X2=0.215
+ $Y2=2
r88 19 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.715 $Y=2
+ $X2=4.8 $Y2=1.915
r89 19 20 285.102 $w=1.68e-07 $l=4.37e-06 $layer=LI1_cond $X=4.715 $Y=2
+ $X2=0.345 $Y2=2
r90 15 30 4.18896 $w=2.17e-07 $l=8.5e-08 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2
r91 15 17 9.52982 $w=2.58e-07 $l=2.15e-07 $layer=LI1_cond $X=0.215 $Y=2.085
+ $X2=0.215 $Y2=2.3
r92 14 30 4.18896 $w=2.17e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.215 $Y2=2
r93 14 29 84.2909 $w=1.73e-07 $l=1.33e-06 $layer=LI1_cond $X=0.172 $Y=1.915
+ $X2=0.172 $Y2=0.585
r94 10 32 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.55 $Y=1.41
+ $X2=4.55 $Y2=1.202
r95 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.55 $Y=1.41
+ $X2=4.55 $Y2=1.985
r96 7 31 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.525 $Y=0.995
+ $X2=4.525 $Y2=1.202
r97 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.525 $Y=0.995
+ $X2=4.525 $Y2=0.56
r98 2 17 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.3
r99 1 27 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%VPWR 1 2 3 4 5 16 19 22 25 27 32 41 46 53
+ 60 69 70
r75 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r76 67 69 11.1981 $w=4.14e-07 $l=3.8e-07 $layer=LI1_cond $X=4.815 $Y=2.34
+ $X2=4.815 $Y2=2.72
r77 63 64 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r78 60 63 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=2.64 $Y=2.34
+ $X2=2.64 $Y2=2.72
r79 57 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r81 53 56 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.7 $Y=2.34 $X2=1.7
+ $Y2=2.72
r82 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r83 46 49 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=2.34
+ $X2=0.705 $Y2=2.72
r84 44 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r85 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r86 41 69 5.98801 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=4.57 $Y=2.72
+ $X2=4.815 $Y2=2.72
r87 41 43 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.57 $Y=2.72 $X2=4.37
+ $Y2=2.72
r88 40 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r89 40 64 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r90 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r91 37 63 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.83 $Y=2.72 $X2=2.64
+ $Y2=2.72
r92 37 39 40.4492 $w=1.68e-07 $l=6.2e-07 $layer=LI1_cond $X=2.83 $Y=2.72
+ $X2=3.45 $Y2=2.72
r93 36 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r94 36 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r96 33 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r97 33 35 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 32 56 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=2.72 $X2=1.7
+ $Y2=2.72
r99 32 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r100 27 49 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r101 27 29 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r102 25 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r103 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r104 23 43 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.89 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 22 39 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.51 $Y=2.72 $X2=3.45
+ $Y2=2.72
r106 21 23 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.89
+ $Y2=2.72
r107 21 22 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.7 $Y=2.72 $X2=3.51
+ $Y2=2.72
r108 19 21 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.7 $Y=2.34 $X2=3.7
+ $Y2=2.72
r109 17 56 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=2.72 $X2=1.7
+ $Y2=2.72
r110 16 63 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=2.64 $Y2=2.72
r111 16 17 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=1.89 $Y2=2.72
r112 5 67 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.64
+ $Y=1.485 $X2=4.785 $Y2=2.34
r113 4 19 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=2.34
r114 3 60 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.52
+ $Y=1.485 $X2=2.665 $Y2=2.34
r115 2 53 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.485 $X2=1.725 $Y2=2.34
r116 1 46 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%X 1 2 3 4 15 17 21 25 27 28 29 36 38 46
c49 38 0 3.03158e-19 $X=1.155 $Y=0.85
c50 21 0 1.02236e-19 $X=2.195 $Y=1.63
r51 36 46 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=1.195 $Y=1.545
+ $X2=1.195 $Y2=1.53
r52 35 38 1.04768 $w=3.28e-07 $l=3e-08 $layer=LI1_cond $X=1.195 $Y=0.82
+ $X2=1.195 $Y2=0.85
r53 29 36 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=1.63
+ $X2=1.195 $Y2=1.545
r54 29 46 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=1.195 $Y=1.495
+ $X2=1.195 $Y2=1.53
r55 28 29 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.195 $Y=1.19
+ $X2=1.195 $Y2=1.495
r56 27 35 2.96976 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.195 $Y=0.735
+ $X2=1.195 $Y2=0.82
r57 27 28 10.9307 $w=3.28e-07 $l=3.13e-07 $layer=LI1_cond $X=1.195 $Y=0.877
+ $X2=1.195 $Y2=1.19
r58 27 38 0.942908 $w=3.28e-07 $l=2.7e-08 $layer=LI1_cond $X=1.195 $Y=0.877
+ $X2=1.195 $Y2=0.85
r59 23 25 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.195 $Y=0.65
+ $X2=2.195 $Y2=0.42
r60 19 29 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=1.63
+ $X2=1.195 $Y2=1.63
r61 19 21 54.4759 $w=1.68e-07 $l=8.35e-07 $layer=LI1_cond $X=1.36 $Y=1.63
+ $X2=2.195 $Y2=1.63
r62 18 27 3.69268 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.36 $Y=0.735
+ $X2=1.195 $Y2=0.735
r63 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=2.195 $Y2=0.65
r64 17 18 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.11 $Y=0.735
+ $X2=1.36 $Y2=0.735
r65 13 27 2.96976 $w=3.2e-07 $l=8.9861e-08 $layer=LI1_cond $X=1.185 $Y=0.65
+ $X2=1.195 $Y2=0.735
r66 13 15 8.55038 $w=3.08e-07 $l=2.3e-07 $layer=LI1_cond $X=1.185 $Y=0.65
+ $X2=1.185 $Y2=0.42
r67 4 21 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.485 $X2=2.195 $Y2=1.63
r68 3 29 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.11
+ $Y=1.485 $X2=1.255 $Y2=1.63
r69 2 25 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=2.01
+ $Y=0.235 $X2=2.195 $Y2=0.42
r70 1 15 182 $w=1.7e-07 $l=2.6163e-07 $layer=licon1_NDIFF $count=1 $X=1.07
+ $Y=0.235 $X2=1.255 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND4B_4%VGND 1 2 3 12 16 20 23 24 25 27 32 45 46
+ 49 52
r73 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r74 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r75 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r76 43 46 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r77 42 45 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=4.83
+ $Y2=0
r78 42 43 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r79 40 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r80 40 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r81 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r82 37 52 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=1.7
+ $Y2=0
r83 37 39 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=1.89 $Y=0 $X2=2.53
+ $Y2=0
r84 36 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r85 36 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r86 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r87 33 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.69
+ $Y2=0
r88 33 35 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r89 32 52 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.7
+ $Y2=0
r90 32 35 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=0 $X2=1.15
+ $Y2=0
r91 27 49 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.69
+ $Y2=0
r92 27 29 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.23
+ $Y2=0
r93 25 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r94 25 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r95 23 39 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.53
+ $Y2=0
r96 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.535 $Y=0 $X2=2.7
+ $Y2=0
r97 22 42 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.99
+ $Y2=0
r98 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.865 $Y=0 $X2=2.7
+ $Y2=0
r99 18 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.7 $Y=0.085 $X2=2.7
+ $Y2=0
r100 18 20 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.7 $Y=0.085
+ $X2=2.7 $Y2=0.36
r101 14 52 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0
r102 14 16 9.09823 $w=3.78e-07 $l=3e-07 $layer=LI1_cond $X=1.7 $Y=0.085 $X2=1.7
+ $Y2=0.385
r103 10 49 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0
r104 10 12 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.69 $Y=0.085
+ $X2=0.69 $Y2=0.38
r105 3 20 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=2.48
+ $Y=0.235 $X2=2.7 $Y2=0.36
r106 2 16 182 $w=1.7e-07 $l=2.48948e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.725 $Y2=0.385
r107 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

