* NGSPICE file created from sky130_fd_sc_hdll__o31ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
M1000 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=5.4e+11p ps=5.08e+06u
M1001 VGND A2 a_119_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=3.76e+06u as=5.33e+11p ps=4.24e+06u
M1002 Y B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=2.535e+11p pd=2.08e+06u as=0p ps=0u
M1003 Y A3 a_213_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.8e+11p pd=3.16e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_119_47# A3 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_119_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_213_297# A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

