# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__xor2_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__xor2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.075000 1.500000 1.275000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 0.995000 0.775000 1.445000 ;
        RECT 0.425000 1.445000 1.890000 1.615000 ;
        RECT 1.720000 1.075000 2.155000 1.245000 ;
        RECT 1.720000 1.245000 1.890000 1.445000 ;
    END
  END B
  PIN VGND
    ANTENNADIFFAREA  0.728000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.315000 3.085000 0.485000 ;
        RECT 2.915000 0.485000 3.085000 1.365000 ;
        RECT 2.915000 1.365000 3.545000 1.535000 ;
        RECT 3.225000 1.535000 3.545000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.085000  0.655000 2.745000 0.825000 ;
      RECT 0.085000  0.825000 0.255000 1.785000 ;
      RECT 0.085000  1.785000 0.465000 2.465000 ;
      RECT 0.135000  0.085000 0.465000 0.475000 ;
      RECT 0.685000  0.335000 0.855000 0.655000 ;
      RECT 1.035000  0.085000 1.415000 0.475000 ;
      RECT 1.165000  1.785000 1.335000 2.635000 ;
      RECT 1.505000  1.785000 2.855000 1.955000 ;
      RECT 1.505000  1.955000 1.885000 2.465000 ;
      RECT 2.115000  2.125000 2.285000 2.635000 ;
      RECT 2.455000  1.955000 2.855000 2.465000 ;
      RECT 2.515000  0.825000 2.745000 1.325000 ;
      RECT 3.255000  0.085000 3.545000 0.920000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__xor2_1
END LIBRARY
