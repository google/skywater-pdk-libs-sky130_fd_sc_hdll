* File: sky130_fd_sc_hdll__o21a_1.pex.spice
* Created: Wed Sep  2 08:43:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21A_1%A_83_21# 1 2 7 9 10 12 16 18 19 20 22 24 26
r61 24 33 2.8558 $w=3.3e-07 $l=1.08e-07 $layer=LI1_cond $X=1.645 $Y=1.69
+ $X2=1.645 $Y2=1.582
r62 24 26 22.6996 $w=3.28e-07 $l=6.5e-07 $layer=LI1_cond $X=1.645 $Y=1.69
+ $X2=1.645 $Y2=2.34
r63 20 22 10.0839 $w=3.58e-07 $l=3.15e-07 $layer=LI1_cond $X=1.205 $Y=0.715
+ $X2=1.205 $Y2=0.4
r64 18 33 4.36303 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=1.48 $Y=1.582
+ $X2=1.645 $Y2=1.582
r65 18 19 31.8932 $w=2.13e-07 $l=5.95e-07 $layer=LI1_cond $X=1.48 $Y=1.582
+ $X2=0.885 $Y2=1.582
r66 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.685
+ $Y=1.16 $X2=0.685 $Y2=1.16
r67 14 19 6.99171 $w=2.15e-07 $l=1.89077e-07 $layer=LI1_cond $X=0.742 $Y=1.475
+ $X2=0.885 $Y2=1.582
r68 14 16 12.7375 $w=2.83e-07 $l=3.15e-07 $layer=LI1_cond $X=0.742 $Y=1.475
+ $X2=0.742 $Y2=1.16
r69 13 20 27.0268 $w=1.88e-07 $l=4.63e-07 $layer=LI1_cond $X=0.742 $Y=0.81
+ $X2=1.205 $Y2=0.81
r70 13 16 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.742 $Y=0.905
+ $X2=0.742 $Y2=1.16
r71 10 17 45.4477 $w=3.63e-07 $l=2.96648e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.617 $Y2=1.16
r72 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r73 7 17 38.952 $w=3.63e-07 $l=2.19499e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.617 $Y2=1.16
r74 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
r75 2 33 400 $w=1.7e-07 $l=2.89569e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.485 $X2=1.645 $Y2=1.66
r76 2 26 400 $w=1.7e-07 $l=9.56478e-07 $layer=licon1_PDIFF $count=1 $X=1.43
+ $Y=1.485 $X2=1.645 $Y2=2.34
r77 1 22 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=1.095
+ $Y=0.235 $X2=1.22 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%B1 1 3 4 6 7 11 15 17
c29 4 0 1.57444e-19 $X=1.435 $Y=0.995
c30 1 0 1.21202e-19 $X=1.34 $Y=1.41
r31 15 17 0.0501062 $w=2.28e-07 $l=1e-09 $layer=LI1_cond $X=1.26 $Y=1.19
+ $X2=1.261 $Y2=1.19
r32 11 17 5.71211 $w=2.28e-07 $l=1.14e-07 $layer=LI1_cond $X=1.375 $Y=1.19
+ $X2=1.261 $Y2=1.19
r33 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.375
+ $Y=1.16 $X2=1.375 $Y2=1.16
r34 7 15 4.50956 $w=2.28e-07 $l=9e-08 $layer=LI1_cond $X=1.17 $Y=1.19 $X2=1.26
+ $Y2=1.19
r35 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.435 $Y=0.995
+ $X2=1.375 $Y2=1.16
r36 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.435 $Y=0.995
+ $X2=1.435 $Y2=0.56
r37 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.34 $Y=1.41
+ $X2=1.375 $Y2=1.16
r38 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.34 $Y=1.41 $X2=1.34
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%A2 1 3 4 6 7 16 21
c40 16 0 1.21202e-19 $X=2.07 $Y=1.275
c41 1 0 6.76182e-20 $X=1.855 $Y=0.995
r42 16 21 1.68994 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=2.07 $Y=1.275 $X2=2.07
+ $Y2=1.175
r43 7 21 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=1.905 $Y=1.175 $X2=2.07
+ $Y2=1.175
r44 7 16 0.908161 $w=1.113e-06 $l=8.3e-08 $layer=LI1_cond $X=1.987 $Y=1.832
+ $X2=2.07 $Y2=1.832
r45 7 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.915
+ $Y=1.16 $X2=1.915 $Y2=1.16
r46 4 11 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.88 $Y=1.41
+ $X2=1.915 $Y2=1.16
r47 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.88 $Y=1.41 $X2=1.88
+ $Y2=1.985
r48 1 11 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.915 $Y2=1.16
r49 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.855 $Y=0.995
+ $X2=1.855 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%A1 1 3 4 6 7 11
r25 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.49
+ $Y=1.16 $X2=2.49 $Y2=1.16
r26 7 11 12.183 $w=3.48e-07 $l=3.7e-07 $layer=LI1_cond $X=2.5 $Y=1.53 $X2=2.5
+ $Y2=1.16
r27 4 10 46.0897 $w=3.39e-07 $l=2.88097e-07 $layer=POLY_cond $X=2.36 $Y=1.41
+ $X2=2.442 $Y2=1.16
r28 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.36 $Y=1.41 $X2=2.36
+ $Y2=1.985
r29 1 10 38.6704 $w=3.39e-07 $l=2.11849e-07 $layer=POLY_cond $X=2.335 $Y=0.995
+ $X2=2.442 $Y2=1.16
r30 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.335 $Y=0.995
+ $X2=2.335 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%X 1 2 9 12 13 16
r20 13 20 17.6982 $w=2.78e-07 $l=4.3e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=2.3
r21 13 16 10.2897 $w=2.78e-07 $l=2.5e-07 $layer=LI1_cond $X=0.225 $Y=1.87
+ $X2=0.225 $Y2=1.62
r22 12 16 24.2836 $w=2.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.225 $Y=1.03
+ $X2=0.225 $Y2=1.62
r23 7 12 6.15521 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=1.03
r24 7 9 15.7614 $w=3.38e-07 $l=4.65e-07 $layer=LI1_cond $X=0.255 $Y=0.86
+ $X2=0.255 $Y2=0.395
r25 2 20 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r26 2 16 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r27 1 9 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%VPWR 1 2 9 11 13 18 24 29 30
r38 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r39 27 29 11.8383 $w=7.42e-07 $l=7.2e-07 $layer=LI1_cond $X=2.8 $Y=2 $X2=2.8
+ $Y2=2.72
r40 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r41 22 30 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r42 22 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r43 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r44 19 24 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=0.9 $Y2=2.72
r45 19 21 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=1.265 $Y=2.72
+ $X2=2.07 $Y2=2.72
r46 18 29 9.70684 $w=1.7e-07 $l=4.2e-07 $layer=LI1_cond $X=2.38 $Y=2.72 $X2=2.8
+ $Y2=2.72
r47 18 21 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=2.38 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 13 24 13.9655 $w=1.7e-07 $l=3.65e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.9 $Y2=2.72
r49 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.535 $Y=2.72
+ $X2=0.23 $Y2=2.72
r50 11 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 11 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r52 7 24 2.94957 $w=7.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.9 $Y=2.635 $X2=0.9
+ $Y2=2.72
r53 7 9 10.4042 $w=7.28e-07 $l=6.35e-07 $layer=LI1_cond $X=0.9 $Y=2.635 $X2=0.9
+ $Y2=2
r54 2 27 150 $w=1.7e-07 $l=7.17635e-07 $layer=licon1_PDIFF $count=4 $X=2.45
+ $Y=1.485 $X2=2.935 $Y2=2
r55 1 9 150 $w=1.7e-07 $l=7.21214e-07 $layer=licon1_PDIFF $count=4 $X=0.605
+ $Y=1.485 $X2=1.1 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%VGND 1 2 11 15 17 19 26 27 30 33
r42 33 34 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r43 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r44 27 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r45 26 27 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r46 24 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.065
+ $Y2=0
r47 24 26 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.15 $Y=0 $X2=2.99
+ $Y2=0
r48 23 34 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r49 23 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r50 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r51 20 30 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r52 20 22 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.61
+ $Y2=0
r53 19 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.98 $Y=0 $X2=2.065
+ $Y2=0
r54 19 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=0 $X2=1.61
+ $Y2=0
r55 17 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r56 13 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.065 $Y=0.085
+ $X2=2.065 $Y2=0
r57 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.065 $Y=0.085
+ $X2=2.065 $Y2=0.38
r58 9 30 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r59 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.38
r60 2 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.93
+ $Y=0.235 $X2=2.065 $Y2=0.38
r61 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_1%A_302_47# 1 2 7 11 14
c26 14 0 2.25062e-19 $X=1.645 $Y=0.72
r27 14 16 4.75325 $w=2.08e-07 $l=9e-08 $layer=LI1_cond $X=1.66 $Y=0.72 $X2=1.66
+ $Y2=0.81
r28 9 11 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=2.545 $Y=0.715
+ $X2=2.545 $Y2=0.4
r29 8 16 1.31963 $w=1.9e-07 $l=1.05e-07 $layer=LI1_cond $X=1.765 $Y=0.81
+ $X2=1.66 $Y2=0.81
r30 7 9 7.47963 $w=1.9e-07 $l=2.07123e-07 $layer=LI1_cond $X=2.38 $Y=0.81
+ $X2=2.545 $Y2=0.715
r31 7 8 35.8995 $w=1.88e-07 $l=6.15e-07 $layer=LI1_cond $X=2.38 $Y=0.81
+ $X2=1.765 $Y2=0.81
r32 2 11 91 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=2 $X=2.41
+ $Y=0.235 $X2=2.545 $Y2=0.4
r33 1 14 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.235 $X2=1.645 $Y2=0.72
.ends

