# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a221oi_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a221oi_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.680000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.985000 0.675000 2.350000 1.075000 ;
        RECT 1.985000 1.075000 2.425000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.670000 0.995000 3.075000 1.325000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.325000 1.075000 1.815000 1.285000 ;
        RECT 1.525000 0.675000 1.815000 1.075000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.605000 1.075000 1.155000 1.285000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.435000 1.285000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  0.432250 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.680000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.560000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 3.680000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  0.874500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.170000 0.255000 0.345000 0.735000 ;
        RECT 0.170000 0.735000 1.335000 0.905000 ;
        RECT 0.175000 1.455000 2.450000 1.495000 ;
        RECT 0.175000 1.495000 3.535000 1.625000 ;
        RECT 0.175000 1.625000 0.345000 2.465000 ;
        RECT 1.165000 0.255000 2.780000 0.505000 ;
        RECT 1.165000 0.505000 1.335000 0.735000 ;
        RECT 2.300000 1.625000 3.535000 1.665000 ;
        RECT 2.580000 0.505000 2.780000 0.655000 ;
        RECT 2.580000 0.655000 3.535000 0.825000 ;
        RECT 3.255000 0.825000 3.535000 1.495000 ;
    END
  END Y
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 3.870000 2.910000 ;
    END
  END VPB
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 3.680000 0.085000 ;
      RECT 0.000000  2.635000 3.680000 2.805000 ;
      RECT 0.515000  0.085000 0.895000 0.565000 ;
      RECT 0.515000  1.795000 0.815000 2.295000 ;
      RECT 0.515000  2.295000 1.835000 2.465000 ;
      RECT 1.115000  1.795000 2.175000 1.835000 ;
      RECT 1.115000  1.835000 2.825000 2.045000 ;
      RECT 1.115000  2.045000 1.340000 2.125000 ;
      RECT 1.455000  2.255000 1.835000 2.295000 ;
      RECT 2.025000  2.215000 2.355000 2.635000 ;
      RECT 2.575000  2.045000 2.825000 2.465000 ;
      RECT 3.030000  0.085000 3.360000 0.485000 ;
      RECT 3.045000  1.875000 3.375000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a221oi_1
END LIBRARY
