* File: sky130_fd_sc_hdll__bufinv_8.pxi.spice
* Created: Wed Sep  2 08:25:05 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%A N_A_c_119_n N_A_M1009_g N_A_c_120_n
+ N_A_M1015_g A PM_SKY130_FD_SC_HDLL__BUFINV_8%A
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%A_117_297# N_A_117_297#_M1015_d
+ N_A_117_297#_M1009_d N_A_117_297#_M1007_g N_A_117_297#_c_151_n
+ N_A_117_297#_M1010_g N_A_117_297#_M1016_g N_A_117_297#_c_152_n
+ N_A_117_297#_M1013_g N_A_117_297#_c_153_n N_A_117_297#_M1018_g
+ N_A_117_297#_M1023_g N_A_117_297#_c_144_n N_A_117_297#_c_154_n
+ N_A_117_297#_c_145_n N_A_117_297#_c_146_n N_A_117_297#_c_147_n
+ N_A_117_297#_c_155_n N_A_117_297#_c_148_n N_A_117_297#_c_149_n
+ N_A_117_297#_c_150_n PM_SKY130_FD_SC_HDLL__BUFINV_8%A_117_297#
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%A_225_47# N_A_225_47#_M1007_s
+ N_A_225_47#_M1016_s N_A_225_47#_M1010_s N_A_225_47#_M1013_s
+ N_A_225_47#_M1002_g N_A_225_47#_c_257_n N_A_225_47#_M1000_g
+ N_A_225_47#_M1005_g N_A_225_47#_c_258_n N_A_225_47#_M1001_g
+ N_A_225_47#_M1006_g N_A_225_47#_c_259_n N_A_225_47#_M1003_g
+ N_A_225_47#_M1008_g N_A_225_47#_c_260_n N_A_225_47#_M1004_g
+ N_A_225_47#_M1012_g N_A_225_47#_c_261_n N_A_225_47#_M1011_g
+ N_A_225_47#_M1014_g N_A_225_47#_c_262_n N_A_225_47#_M1017_g
+ N_A_225_47#_M1020_g N_A_225_47#_c_263_n N_A_225_47#_M1019_g
+ N_A_225_47#_c_264_n N_A_225_47#_M1022_g N_A_225_47#_M1021_g
+ N_A_225_47#_c_247_n N_A_225_47#_c_265_n N_A_225_47#_c_248_n
+ N_A_225_47#_c_249_n N_A_225_47#_c_266_n N_A_225_47#_c_267_n
+ N_A_225_47#_c_296_n N_A_225_47#_c_298_n N_A_225_47#_c_250_n
+ N_A_225_47#_c_268_n N_A_225_47#_c_251_n N_A_225_47#_c_252_n
+ N_A_225_47#_c_253_n N_A_225_47#_c_254_n N_A_225_47#_c_270_n
+ N_A_225_47#_c_255_n N_A_225_47#_c_256_n
+ PM_SKY130_FD_SC_HDLL__BUFINV_8%A_225_47#
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%VPWR N_VPWR_M1009_s N_VPWR_M1010_d
+ N_VPWR_M1018_d N_VPWR_M1001_s N_VPWR_M1004_s N_VPWR_M1017_s N_VPWR_M1022_s
+ N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n N_VPWR_c_492_n
+ N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n N_VPWR_c_497_n
+ N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_500_n N_VPWR_c_501_n N_VPWR_c_502_n
+ N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n
+ VPWR N_VPWR_c_508_n N_VPWR_c_487_n PM_SKY130_FD_SC_HDLL__BUFINV_8%VPWR
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%Y N_Y_M1002_s N_Y_M1006_s N_Y_M1012_s
+ N_Y_M1020_s N_Y_M1000_d N_Y_M1003_d N_Y_M1011_d N_Y_M1019_d N_Y_c_614_n
+ N_Y_c_615_n N_Y_c_595_n N_Y_c_596_n N_Y_c_604_n N_Y_c_605_n N_Y_c_641_n
+ N_Y_c_645_n N_Y_c_597_n N_Y_c_606_n N_Y_c_657_n N_Y_c_661_n N_Y_c_598_n
+ N_Y_c_607_n N_Y_c_673_n N_Y_c_675_n N_Y_c_599_n N_Y_c_608_n N_Y_c_600_n
+ N_Y_c_609_n N_Y_c_601_n N_Y_c_610_n N_Y_c_602_n N_Y_c_611_n Y Y
+ PM_SKY130_FD_SC_HDLL__BUFINV_8%Y
x_PM_SKY130_FD_SC_HDLL__BUFINV_8%VGND N_VGND_M1015_s N_VGND_M1007_d
+ N_VGND_M1023_d N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1014_d N_VGND_M1021_d
+ N_VGND_c_774_n N_VGND_c_775_n N_VGND_c_776_n N_VGND_c_777_n N_VGND_c_778_n
+ N_VGND_c_779_n N_VGND_c_780_n N_VGND_c_781_n N_VGND_c_782_n N_VGND_c_783_n
+ N_VGND_c_784_n N_VGND_c_785_n N_VGND_c_786_n N_VGND_c_787_n N_VGND_c_788_n
+ N_VGND_c_789_n N_VGND_c_790_n N_VGND_c_791_n N_VGND_c_792_n N_VGND_c_793_n
+ VGND N_VGND_c_794_n N_VGND_c_795_n PM_SKY130_FD_SC_HDLL__BUFINV_8%VGND
cc_1 VNB N_A_c_119_n 0.0482365f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_c_120_n 0.0247935f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB A 0.00900655f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_117_297#_M1007_g 0.0221524f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_5 VNB N_A_117_297#_M1016_g 0.0188756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_117_297#_M1023_g 0.0185511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_297#_c_144_n 0.00434074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_117_297#_c_145_n 0.00444855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_117_297#_c_146_n 0.0210275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_117_297#_c_147_n 0.00366951f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_c_148_n 8.20462e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_117_297#_c_149_n 0.00253509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_117_297#_c_150_n 0.0684039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_225_47#_M1002_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_225_47#_M1005_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_225_47#_M1006_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_225_47#_M1008_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_47#_M1012_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_225_47#_M1014_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_47#_M1020_g 0.0188782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_225_47#_M1021_g 0.0218826f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_225_47#_c_247_n 0.00451034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_225_47#_c_248_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_225_47#_c_249_n 0.004399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_225_47#_c_250_n 0.00102469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_225_47#_c_251_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_225_47#_c_252_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_225_47#_c_253_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_225_47#_c_254_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_225_47#_c_255_n 0.00153756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_225_47#_c_256_n 0.185466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VPWR_c_487_n 0.288713f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_595_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_596_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_597_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_598_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_599_n 0.0143792f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_600_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_601_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_602_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB Y 0.023733f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_774_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_775_n 0.00656836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_776_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_777_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_778_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_779_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_780_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_781_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_782_n 0.0334789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_783_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_784_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_785_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_786_n 0.0200002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_787_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_788_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_789_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_790_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_791_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_792_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_793_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_794_n 0.0136226f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_795_n 0.34616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VPB N_A_c_119_n 0.0443612f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB N_A_117_297#_c_151_n 0.0194367f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_66 VPB N_A_117_297#_c_152_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_117_297#_c_153_n 0.0159693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_117_297#_c_154_n 0.00682118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_117_297#_c_155_n 0.0017029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_117_297#_c_148_n 0.0051786f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_117_297#_c_150_n 0.0203235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_225_47#_c_257_n 0.0162292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A_225_47#_c_258_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A_225_47#_c_259_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_225_47#_c_260_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A_225_47#_c_261_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_A_225_47#_c_262_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_A_225_47#_c_263_n 0.0158863f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_A_225_47#_c_264_n 0.0191859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_A_225_47#_c_265_n 0.00788153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_225_47#_c_266_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_225_47#_c_267_n 0.00454699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_225_47#_c_268_n 0.00100785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_225_47#_c_252_n 0.00252324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_225_47#_c_270_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_225_47#_c_256_n 0.0514916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_488_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_489_n 0.00757198f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_490_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_491_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_492_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_493_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_494_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_495_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_496_n 0.03408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_497_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_498_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_499_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_500_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_501_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_502_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_503_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_504_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_505_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_506_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_507_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_508_n 0.014713f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_487_n 0.0648491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_Y_c_604_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_Y_c_605_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_Y_c_606_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_Y_c_607_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_Y_c_608_n 0.00178474f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_Y_c_609_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_Y_c_610_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_Y_c_611_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB Y 0.00852491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB Y 0.01924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 N_A_c_120_n N_A_117_297#_c_144_n 0.00719164f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_120 N_A_c_119_n N_A_117_297#_c_154_n 0.0111529f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_c_120_n N_A_117_297#_c_145_n 0.00646196f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_120_n N_A_117_297#_c_147_n 0.00526894f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_119_n N_A_117_297#_c_155_n 0.00463593f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_119_n N_A_117_297#_c_148_n 0.00762945f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_c_119_n N_A_117_297#_c_149_n 0.00550394f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_126 A N_A_117_297#_c_149_n 0.0140451f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_127 N_A_c_120_n N_A_225_47#_c_249_n 3.65437e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_119_n N_VPWR_c_489_n 0.012741f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 A N_VPWR_c_489_n 0.0136987f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_130 N_A_c_119_n N_VPWR_c_496_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_c_119_n N_VPWR_c_487_n 0.0121883f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_132 N_A_c_119_n N_VGND_c_775_n 0.00431355f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_120_n N_VGND_c_775_n 0.00643264f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_134 A N_VGND_c_775_n 0.0136981f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_135 N_A_c_120_n N_VGND_c_782_n 0.00466005f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_120_n N_VGND_c_795_n 0.0101005f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_117_297#_M1023_g N_A_225_47#_M1002_g 0.0207193f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_138 N_A_117_297#_c_153_n N_A_225_47#_c_257_n 0.0215651f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_139 N_A_117_297#_M1007_g N_A_225_47#_c_247_n 0.00693104f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_140 N_A_117_297#_M1016_g N_A_225_47#_c_247_n 5.47935e-19 $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_141 N_A_117_297#_c_144_n N_A_225_47#_c_247_n 0.0368926f $X=0.73 $Y=0.4 $X2=0
+ $Y2=0
cc_142 N_A_117_297#_c_151_n N_A_225_47#_c_265_n 0.0112091f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_143 N_A_117_297#_c_152_n N_A_225_47#_c_265_n 7.06303e-19 $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_144 N_A_117_297#_c_155_n N_A_225_47#_c_265_n 0.0660799f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_145 N_A_117_297#_M1007_g N_A_225_47#_c_248_n 0.00879805f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_146 N_A_117_297#_M1016_g N_A_225_47#_c_248_n 0.00879805f $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_147 N_A_117_297#_c_146_n N_A_225_47#_c_248_n 0.03957f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_148 N_A_117_297#_c_150_n N_A_225_47#_c_248_n 0.0031956f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_149 N_A_117_297#_M1007_g N_A_225_47#_c_249_n 0.00126794f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_150 N_A_117_297#_c_146_n N_A_225_47#_c_249_n 0.0278128f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_151 N_A_117_297#_c_147_n N_A_225_47#_c_249_n 0.0140416f $X=0.705 $Y=0.905
+ $X2=0 $Y2=0
cc_152 N_A_117_297#_c_151_n N_A_225_47#_c_266_n 0.0137916f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_153 N_A_117_297#_c_152_n N_A_225_47#_c_266_n 0.0101048f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_154 N_A_117_297#_c_146_n N_A_225_47#_c_266_n 0.0394547f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_117_297#_c_150_n N_A_225_47#_c_266_n 0.00720931f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_156 N_A_117_297#_c_151_n N_A_225_47#_c_267_n 0.00138874f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_157 N_A_117_297#_c_146_n N_A_225_47#_c_267_n 0.0279779f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_158 N_A_117_297#_c_148_n N_A_225_47#_c_267_n 0.0135536f $X=0.705 $Y=1.545
+ $X2=0 $Y2=0
cc_159 N_A_117_297#_c_150_n N_A_225_47#_c_267_n 3.20658e-19 $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_160 N_A_117_297#_M1007_g N_A_225_47#_c_296_n 5.25882e-19 $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_161 N_A_117_297#_M1016_g N_A_225_47#_c_296_n 0.00657592f $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_162 N_A_117_297#_c_151_n N_A_225_47#_c_298_n 7.33057e-19 $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_163 N_A_117_297#_c_152_n N_A_225_47#_c_298_n 0.0137692f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_164 N_A_117_297#_c_153_n N_A_225_47#_c_298_n 0.0112091f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_165 N_A_117_297#_M1023_g N_A_225_47#_c_250_n 0.0116573f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_166 N_A_117_297#_c_153_n N_A_225_47#_c_268_n 0.0151183f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_167 N_A_117_297#_c_150_n N_A_225_47#_c_268_n 3.58038e-19 $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_168 N_A_117_297#_M1023_g N_A_225_47#_c_251_n 0.00410511f $X=2.45 $Y=0.56
+ $X2=0 $Y2=0
cc_169 N_A_117_297#_c_153_n N_A_225_47#_c_252_n 8.16926e-19 $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_170 N_A_117_297#_c_150_n N_A_225_47#_c_252_n 0.00327205f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_171 N_A_117_297#_M1016_g N_A_225_47#_c_254_n 0.0011682f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_172 N_A_117_297#_c_146_n N_A_225_47#_c_254_n 0.0307156f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_173 N_A_117_297#_c_150_n N_A_225_47#_c_254_n 0.00450461f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_174 N_A_117_297#_c_152_n N_A_225_47#_c_270_n 0.00259297f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_175 N_A_117_297#_c_153_n N_A_225_47#_c_270_n 0.00107777f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_176 N_A_117_297#_c_146_n N_A_225_47#_c_270_n 0.0305808f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_177 N_A_117_297#_c_150_n N_A_225_47#_c_270_n 0.00723098f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_178 N_A_117_297#_c_146_n N_A_225_47#_c_255_n 0.014524f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_179 N_A_117_297#_c_150_n N_A_225_47#_c_255_n 0.00220849f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_180 N_A_117_297#_c_150_n N_A_225_47#_c_256_n 0.0207193f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_181 N_A_117_297#_c_155_n N_VPWR_c_489_n 0.0686444f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_182 N_A_117_297#_c_148_n N_VPWR_c_489_n 0.00410807f $X=0.705 $Y=1.545 $X2=0
+ $Y2=0
cc_183 N_A_117_297#_c_151_n N_VPWR_c_490_n 0.00547044f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_117_297#_c_152_n N_VPWR_c_490_n 0.00497803f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_117_297#_c_153_n N_VPWR_c_491_n 0.00547044f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_117_297#_c_151_n N_VPWR_c_496_n 0.00673617f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_117_297#_c_154_n N_VPWR_c_496_n 0.0244686f $X=0.73 $Y=2.31 $X2=0
+ $Y2=0
cc_188 N_A_117_297#_c_152_n N_VPWR_c_498_n 0.00597712f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_117_297#_c_153_n N_VPWR_c_498_n 0.00673617f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_117_297#_M1009_d N_VPWR_c_487_n 0.00217517f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_117_297#_c_151_n N_VPWR_c_487_n 0.0131262f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_117_297#_c_152_n N_VPWR_c_487_n 0.00999457f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_117_297#_c_153_n N_VPWR_c_487_n 0.011869f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_117_297#_c_154_n N_VPWR_c_487_n 0.0141694f $X=0.73 $Y=2.31 $X2=0
+ $Y2=0
cc_195 N_A_117_297#_M1023_g N_Y_c_614_n 5.33681e-19 $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_196 N_A_117_297#_c_153_n N_Y_c_615_n 7.33057e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_117_297#_c_144_n N_VGND_c_775_n 0.0481407f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_198 N_A_117_297#_M1007_g N_VGND_c_776_n 0.00390178f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_M1016_g N_VGND_c_776_n 0.00276126f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_200 N_A_117_297#_M1023_g N_VGND_c_777_n 0.00268723f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_M1007_g N_VGND_c_782_n 0.00424619f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_c_144_n N_VGND_c_782_n 0.023651f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_203 N_A_117_297#_M1016_g N_VGND_c_784_n 0.00424619f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_M1023_g N_VGND_c_784_n 0.00439206f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_M1015_d N_VGND_c_795_n 0.0020946f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_M1007_g N_VGND_c_795_n 0.00731205f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_207 N_A_117_297#_M1016_g N_VGND_c_795_n 0.00610552f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_208 N_A_117_297#_M1023_g N_VGND_c_795_n 0.00618081f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_209 N_A_117_297#_c_144_n N_VGND_c_795_n 0.0140774f $X=0.73 $Y=0.4 $X2=0 $Y2=0
cc_210 N_A_225_47#_c_266_n N_VPWR_M1010_d 0.00178587f $X=1.975 $Y=1.53 $X2=0
+ $Y2=0
cc_211 N_A_225_47#_c_268_n N_VPWR_M1018_d 0.00324655f $X=2.575 $Y=1.53 $X2=0
+ $Y2=0
cc_212 N_A_225_47#_c_265_n N_VPWR_c_490_n 0.0411685f $X=1.25 $Y=1.63 $X2=0 $Y2=0
cc_213 N_A_225_47#_c_266_n N_VPWR_c_490_n 0.0136682f $X=1.975 $Y=1.53 $X2=0
+ $Y2=0
cc_214 N_A_225_47#_c_298_n N_VPWR_c_490_n 0.0507655f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_215 N_A_225_47#_c_257_n N_VPWR_c_491_n 0.00497803f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_225_47#_c_298_n N_VPWR_c_491_n 0.0416217f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_217 N_A_225_47#_c_268_n N_VPWR_c_491_n 0.0151472f $X=2.575 $Y=1.53 $X2=0
+ $Y2=0
cc_218 N_A_225_47#_c_258_n N_VPWR_c_492_n 0.0052072f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_225_47#_c_259_n N_VPWR_c_492_n 0.004751f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A_225_47#_c_260_n N_VPWR_c_493_n 0.0052072f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_225_47#_c_261_n N_VPWR_c_493_n 0.004751f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_225_47#_c_262_n N_VPWR_c_494_n 0.0052072f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_225_47#_c_263_n N_VPWR_c_494_n 0.004751f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_225_47#_c_264_n N_VPWR_c_495_n 0.00688901f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_225_47#_c_265_n N_VPWR_c_496_n 0.0210596f $X=1.25 $Y=1.63 $X2=0 $Y2=0
cc_226 N_A_225_47#_c_298_n N_VPWR_c_498_n 0.0223557f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_227 N_A_225_47#_c_257_n N_VPWR_c_500_n 0.00597712f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_225_47#_c_258_n N_VPWR_c_500_n 0.00673617f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_225_47#_c_259_n N_VPWR_c_502_n 0.00597712f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_225_47#_c_260_n N_VPWR_c_502_n 0.00673617f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_225_47#_c_261_n N_VPWR_c_504_n 0.00597712f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_232 N_A_225_47#_c_262_n N_VPWR_c_504_n 0.00673617f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A_225_47#_c_263_n N_VPWR_c_506_n 0.00597712f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_225_47#_c_264_n N_VPWR_c_506_n 0.00673617f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_235 N_A_225_47#_M1010_s N_VPWR_c_487_n 0.00217517f $X=1.125 $Y=1.485 $X2=0
+ $Y2=0
cc_236 N_A_225_47#_M1013_s N_VPWR_c_487_n 0.00231261f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_237 N_A_225_47#_c_257_n N_VPWR_c_487_n 0.0100198f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_225_47#_c_258_n N_VPWR_c_487_n 0.0118438f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_225_47#_c_259_n N_VPWR_c_487_n 0.00999457f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_240 N_A_225_47#_c_260_n N_VPWR_c_487_n 0.0118438f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A_225_47#_c_261_n N_VPWR_c_487_n 0.00999457f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_225_47#_c_262_n N_VPWR_c_487_n 0.0118438f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_243 N_A_225_47#_c_263_n N_VPWR_c_487_n 0.00999457f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_244 N_A_225_47#_c_264_n N_VPWR_c_487_n 0.0129051f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_225_47#_c_265_n N_VPWR_c_487_n 0.0124725f $X=1.25 $Y=1.63 $X2=0 $Y2=0
cc_246 N_A_225_47#_c_298_n N_VPWR_c_487_n 0.0140101f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_247 N_A_225_47#_M1002_g N_Y_c_614_n 0.0065059f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_248 N_A_225_47#_M1005_g N_Y_c_614_n 0.00693104f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_249 N_A_225_47#_M1006_g N_Y_c_614_n 5.47131e-19 $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_250 N_A_225_47#_c_257_n N_Y_c_615_n 0.0137692f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_225_47#_c_258_n N_Y_c_615_n 0.0115459f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_225_47#_c_259_n N_Y_c_615_n 7.68612e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_225_47#_c_298_n N_Y_c_615_n 0.00486061f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_254 N_A_225_47#_M1005_g N_Y_c_595_n 0.00879805f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_225_47#_M1006_g N_Y_c_595_n 0.00879805f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_256 N_A_225_47#_c_253_n N_Y_c_595_n 0.03957f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_257 N_A_225_47#_c_256_n N_Y_c_595_n 0.0031956f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_258 N_A_225_47#_M1002_g N_Y_c_596_n 0.00243606f $X=2.87 $Y=0.56 $X2=0 $Y2=0
cc_259 N_A_225_47#_M1005_g N_Y_c_596_n 0.00113891f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_260 N_A_225_47#_c_250_n N_Y_c_596_n 0.00808484f $X=2.575 $Y=0.82 $X2=0 $Y2=0
cc_261 N_A_225_47#_c_253_n N_Y_c_596_n 0.030582f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_262 N_A_225_47#_c_256_n N_Y_c_596_n 0.00331919f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_263 N_A_225_47#_c_258_n N_Y_c_604_n 0.0137916f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_225_47#_c_259_n N_Y_c_604_n 0.0101048f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_225_47#_c_253_n N_Y_c_604_n 0.0394547f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_266 N_A_225_47#_c_256_n N_Y_c_604_n 0.00720931f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_267 N_A_225_47#_c_257_n N_Y_c_605_n 0.00386185f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_225_47#_c_258_n N_Y_c_605_n 0.00107777f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_225_47#_c_268_n N_Y_c_605_n 0.0149281f $X=2.575 $Y=1.53 $X2=0 $Y2=0
cc_270 N_A_225_47#_c_253_n N_Y_c_605_n 0.0305808f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_225_47#_c_256_n N_Y_c_605_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_272 N_A_225_47#_M1005_g N_Y_c_641_n 5.25882e-19 $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_273 N_A_225_47#_M1006_g N_Y_c_641_n 0.00657592f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_225_47#_M1008_g N_Y_c_641_n 0.00693104f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_275 N_A_225_47#_M1012_g N_Y_c_641_n 5.47131e-19 $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A_225_47#_c_258_n N_Y_c_645_n 8.07084e-19 $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_225_47#_c_259_n N_Y_c_645_n 0.0141618f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_225_47#_c_260_n N_Y_c_645_n 0.0115459f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_225_47#_c_261_n N_Y_c_645_n 7.68612e-19 $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_225_47#_M1008_g N_Y_c_597_n 0.00879805f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_225_47#_M1012_g N_Y_c_597_n 0.00879805f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_225_47#_c_253_n N_Y_c_597_n 0.03957f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_225_47#_c_256_n N_Y_c_597_n 0.0031956f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_284 N_A_225_47#_c_260_n N_Y_c_606_n 0.0137916f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_285 N_A_225_47#_c_261_n N_Y_c_606_n 0.0101048f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A_225_47#_c_253_n N_Y_c_606_n 0.0394547f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_287 N_A_225_47#_c_256_n N_Y_c_606_n 0.00720931f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_288 N_A_225_47#_M1008_g N_Y_c_657_n 5.25882e-19 $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_225_47#_M1012_g N_Y_c_657_n 0.00657592f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_225_47#_M1014_g N_Y_c_657_n 0.00693104f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_291 N_A_225_47#_M1020_g N_Y_c_657_n 5.47131e-19 $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_292 N_A_225_47#_c_260_n N_Y_c_661_n 8.07084e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_293 N_A_225_47#_c_261_n N_Y_c_661_n 0.0141618f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_294 N_A_225_47#_c_262_n N_Y_c_661_n 0.0115459f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_295 N_A_225_47#_c_263_n N_Y_c_661_n 7.68612e-19 $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_225_47#_M1014_g N_Y_c_598_n 0.00879805f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A_225_47#_M1020_g N_Y_c_598_n 0.00879805f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_225_47#_c_253_n N_Y_c_598_n 0.03957f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_225_47#_c_256_n N_Y_c_598_n 0.0031956f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_300 N_A_225_47#_c_262_n N_Y_c_607_n 0.0137916f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_225_47#_c_263_n N_Y_c_607_n 0.0101048f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_225_47#_c_253_n N_Y_c_607_n 0.0394547f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_225_47#_c_256_n N_Y_c_607_n 0.00720931f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_304 N_A_225_47#_M1014_g N_Y_c_673_n 5.25882e-19 $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A_225_47#_M1020_g N_Y_c_673_n 0.00657592f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_225_47#_c_262_n N_Y_c_675_n 8.07084e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_307 N_A_225_47#_c_263_n N_Y_c_675_n 0.0141618f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_308 N_A_225_47#_c_264_n N_Y_c_675_n 0.017566f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_309 N_A_225_47#_M1021_g N_Y_c_599_n 0.0127467f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A_225_47#_c_253_n N_Y_c_599_n 0.00896055f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_225_47#_c_264_n N_Y_c_608_n 0.0158923f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_312 N_A_225_47#_c_253_n N_Y_c_608_n 0.0088891f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_313 N_A_225_47#_c_256_n N_Y_c_608_n 3.58038e-19 $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_314 N_A_225_47#_M1006_g N_Y_c_600_n 0.00113891f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_315 N_A_225_47#_M1008_g N_Y_c_600_n 0.00113891f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_316 N_A_225_47#_c_253_n N_Y_c_600_n 0.030582f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_225_47#_c_256_n N_Y_c_600_n 0.00331919f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_318 N_A_225_47#_c_259_n N_Y_c_609_n 0.00260297f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_319 N_A_225_47#_c_260_n N_Y_c_609_n 0.00107777f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_320 N_A_225_47#_c_253_n N_Y_c_609_n 0.0305808f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_321 N_A_225_47#_c_256_n N_Y_c_609_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_322 N_A_225_47#_M1012_g N_Y_c_601_n 0.00113891f $X=4.75 $Y=0.56 $X2=0 $Y2=0
cc_323 N_A_225_47#_M1014_g N_Y_c_601_n 0.00113891f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_324 N_A_225_47#_c_253_n N_Y_c_601_n 0.030582f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_225_47#_c_256_n N_Y_c_601_n 0.00331919f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_326 N_A_225_47#_c_261_n N_Y_c_610_n 0.00260297f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_327 N_A_225_47#_c_262_n N_Y_c_610_n 0.00107777f $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A_225_47#_c_253_n N_Y_c_610_n 0.0305808f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_225_47#_c_256_n N_Y_c_610_n 0.0074788f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_330 N_A_225_47#_M1020_g N_Y_c_602_n 0.0011682f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_331 N_A_225_47#_c_253_n N_Y_c_602_n 0.0307156f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_332 N_A_225_47#_c_256_n N_Y_c_602_n 0.00450461f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_333 N_A_225_47#_c_263_n N_Y_c_611_n 0.00260297f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_334 N_A_225_47#_c_264_n N_Y_c_611_n 0.00107777f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_335 N_A_225_47#_c_253_n N_Y_c_611_n 0.0305808f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_336 N_A_225_47#_c_256_n N_Y_c_611_n 0.00723098f $X=6.185 $Y=1.217 $X2=0 $Y2=0
cc_337 N_A_225_47#_c_264_n Y 0.00135583f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_338 N_A_225_47#_M1021_g Y 0.0183546f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_339 N_A_225_47#_c_253_n Y 0.016826f $X=6.07 $Y=1.16 $X2=0 $Y2=0
cc_340 N_A_225_47#_c_248_n N_VGND_M1007_d 0.00251598f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_341 N_A_225_47#_c_250_n N_VGND_M1023_d 0.00193551f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_342 N_A_225_47#_c_247_n N_VGND_c_776_n 0.0184656f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_343 N_A_225_47#_c_248_n N_VGND_c_776_n 0.0127122f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_344 N_A_225_47#_M1002_g N_VGND_c_777_n 0.00268723f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_345 N_A_225_47#_c_250_n N_VGND_c_777_n 0.0135251f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_346 N_A_225_47#_M1005_g N_VGND_c_778_n 0.00390178f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_347 N_A_225_47#_M1006_g N_VGND_c_778_n 0.00276126f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_348 N_A_225_47#_M1008_g N_VGND_c_779_n 0.00390178f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_225_47#_M1012_g N_VGND_c_779_n 0.00276126f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_225_47#_M1014_g N_VGND_c_780_n 0.00390178f $X=5.22 $Y=0.56 $X2=0
+ $Y2=0
cc_351 N_A_225_47#_M1020_g N_VGND_c_780_n 0.00276126f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_352 N_A_225_47#_M1021_g N_VGND_c_781_n 0.00438629f $X=6.21 $Y=0.56 $X2=0
+ $Y2=0
cc_353 N_A_225_47#_c_247_n N_VGND_c_782_n 0.020318f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_354 N_A_225_47#_c_248_n N_VGND_c_782_n 0.00260082f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_355 N_A_225_47#_c_248_n N_VGND_c_784_n 0.00193763f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_356 N_A_225_47#_c_296_n N_VGND_c_784_n 0.022456f $X=2.19 $Y=0.4 $X2=0 $Y2=0
cc_357 N_A_225_47#_c_250_n N_VGND_c_784_n 0.00248202f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_358 N_A_225_47#_M1002_g N_VGND_c_786_n 0.00541562f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_359 N_A_225_47#_M1005_g N_VGND_c_786_n 0.00424619f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_360 N_A_225_47#_M1006_g N_VGND_c_788_n 0.00424619f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_361 N_A_225_47#_M1008_g N_VGND_c_788_n 0.00424619f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_225_47#_M1012_g N_VGND_c_790_n 0.00424619f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_363 N_A_225_47#_M1014_g N_VGND_c_790_n 0.00424619f $X=5.22 $Y=0.56 $X2=0
+ $Y2=0
cc_364 N_A_225_47#_M1020_g N_VGND_c_792_n 0.00424619f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_225_47#_M1021_g N_VGND_c_792_n 0.00439206f $X=6.21 $Y=0.56 $X2=0
+ $Y2=0
cc_366 N_A_225_47#_M1007_s N_VGND_c_795_n 0.0020946f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_367 N_A_225_47#_M1016_s N_VGND_c_795_n 0.00304616f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_368 N_A_225_47#_M1002_g N_VGND_c_795_n 0.00965588f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_369 N_A_225_47#_M1005_g N_VGND_c_795_n 0.00611295f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_370 N_A_225_47#_M1006_g N_VGND_c_795_n 0.00599018f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_371 N_A_225_47#_M1008_g N_VGND_c_795_n 0.00611295f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_372 N_A_225_47#_M1012_g N_VGND_c_795_n 0.00599018f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_373 N_A_225_47#_M1014_g N_VGND_c_795_n 0.00611295f $X=5.22 $Y=0.56 $X2=0
+ $Y2=0
cc_374 N_A_225_47#_M1020_g N_VGND_c_795_n 0.00610552f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_375 N_A_225_47#_M1021_g N_VGND_c_795_n 0.0072623f $X=6.21 $Y=0.56 $X2=0 $Y2=0
cc_376 N_A_225_47#_c_247_n N_VGND_c_795_n 0.0123792f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_377 N_A_225_47#_c_248_n N_VGND_c_795_n 0.00961016f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_378 N_A_225_47#_c_296_n N_VGND_c_795_n 0.0142976f $X=2.19 $Y=0.4 $X2=0 $Y2=0
cc_379 N_A_225_47#_c_250_n N_VGND_c_795_n 0.00561929f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_487_n N_Y_M1000_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_381 N_VPWR_c_487_n N_Y_M1003_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_382 N_VPWR_c_487_n N_Y_M1011_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_383 N_VPWR_c_487_n N_Y_M1019_d 0.00231261f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_384 N_VPWR_c_491_n N_Y_c_615_n 0.0507655f $X=2.66 $Y=2 $X2=0 $Y2=0
cc_385 N_VPWR_c_492_n N_Y_c_615_n 0.0385613f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_386 N_VPWR_c_500_n N_Y_c_615_n 0.0223557f $X=3.515 $Y=2.72 $X2=0 $Y2=0
cc_387 N_VPWR_c_487_n N_Y_c_615_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_388 N_VPWR_M1001_s N_Y_c_604_n 0.00199888f $X=3.455 $Y=1.485 $X2=0 $Y2=0
cc_389 N_VPWR_c_492_n N_Y_c_604_n 0.0112848f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_390 N_VPWR_c_492_n N_Y_c_645_n 0.0470327f $X=3.6 $Y=2 $X2=0 $Y2=0
cc_391 N_VPWR_c_493_n N_Y_c_645_n 0.0385613f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_392 N_VPWR_c_502_n N_Y_c_645_n 0.0223557f $X=4.455 $Y=2.72 $X2=0 $Y2=0
cc_393 N_VPWR_c_487_n N_Y_c_645_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_394 N_VPWR_M1004_s N_Y_c_606_n 0.00199888f $X=4.395 $Y=1.485 $X2=0 $Y2=0
cc_395 N_VPWR_c_493_n N_Y_c_606_n 0.0112848f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_396 N_VPWR_c_493_n N_Y_c_661_n 0.0470327f $X=4.54 $Y=2 $X2=0 $Y2=0
cc_397 N_VPWR_c_494_n N_Y_c_661_n 0.0385613f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_398 N_VPWR_c_504_n N_Y_c_661_n 0.0223557f $X=5.395 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_487_n N_Y_c_661_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_M1017_s N_Y_c_607_n 0.00199888f $X=5.335 $Y=1.485 $X2=0 $Y2=0
cc_401 N_VPWR_c_494_n N_Y_c_607_n 0.0112848f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_402 N_VPWR_c_494_n N_Y_c_675_n 0.0470327f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_403 N_VPWR_c_495_n N_Y_c_675_n 0.0385613f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_404 N_VPWR_c_506_n N_Y_c_675_n 0.0223557f $X=6.335 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_c_487_n N_Y_c_675_n 0.0140101f $X=6.67 $Y=2.72 $X2=0 $Y2=0
cc_406 N_VPWR_M1022_s N_Y_c_608_n 9.28053e-19 $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_407 N_VPWR_c_495_n N_Y_c_608_n 0.00527645f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_408 N_VPWR_M1022_s Y 0.0036007f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_409 N_VPWR_c_495_n Y 0.00661812f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_410 N_Y_c_595_n N_VGND_M1005_d 0.00251598f $X=3.855 $Y=0.82 $X2=0 $Y2=0
cc_411 N_Y_c_597_n N_VGND_M1008_d 0.00251598f $X=4.795 $Y=0.82 $X2=0 $Y2=0
cc_412 N_Y_c_598_n N_VGND_M1014_d 0.00251598f $X=5.735 $Y=0.82 $X2=0 $Y2=0
cc_413 N_Y_c_599_n N_VGND_M1021_d 0.0031882f $X=6.415 $Y=0.82 $X2=0 $Y2=0
cc_414 N_Y_c_614_n N_VGND_c_778_n 0.0186688f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_415 N_Y_c_595_n N_VGND_c_778_n 0.0127122f $X=3.855 $Y=0.82 $X2=0 $Y2=0
cc_416 N_Y_c_641_n N_VGND_c_779_n 0.0186688f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_417 N_Y_c_597_n N_VGND_c_779_n 0.0127122f $X=4.795 $Y=0.82 $X2=0 $Y2=0
cc_418 N_Y_c_657_n N_VGND_c_780_n 0.0186688f $X=5.01 $Y=0.4 $X2=0 $Y2=0
cc_419 N_Y_c_598_n N_VGND_c_780_n 0.0127122f $X=5.735 $Y=0.82 $X2=0 $Y2=0
cc_420 N_Y_c_599_n N_VGND_c_781_n 0.0134107f $X=6.415 $Y=0.82 $X2=0 $Y2=0
cc_421 N_Y_c_614_n N_VGND_c_786_n 0.0216617f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_422 N_Y_c_595_n N_VGND_c_786_n 0.00260082f $X=3.855 $Y=0.82 $X2=0 $Y2=0
cc_423 N_Y_c_595_n N_VGND_c_788_n 0.00193763f $X=3.855 $Y=0.82 $X2=0 $Y2=0
cc_424 N_Y_c_641_n N_VGND_c_788_n 0.0216617f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_425 N_Y_c_597_n N_VGND_c_788_n 0.00260082f $X=4.795 $Y=0.82 $X2=0 $Y2=0
cc_426 N_Y_c_597_n N_VGND_c_790_n 0.00193763f $X=4.795 $Y=0.82 $X2=0 $Y2=0
cc_427 N_Y_c_657_n N_VGND_c_790_n 0.0216617f $X=5.01 $Y=0.4 $X2=0 $Y2=0
cc_428 N_Y_c_598_n N_VGND_c_790_n 0.00260082f $X=5.735 $Y=0.82 $X2=0 $Y2=0
cc_429 N_Y_c_598_n N_VGND_c_792_n 0.00193763f $X=5.735 $Y=0.82 $X2=0 $Y2=0
cc_430 N_Y_c_673_n N_VGND_c_792_n 0.022456f $X=5.95 $Y=0.4 $X2=0 $Y2=0
cc_431 N_Y_c_599_n N_VGND_c_792_n 0.00248202f $X=6.415 $Y=0.82 $X2=0 $Y2=0
cc_432 N_Y_c_599_n N_VGND_c_794_n 0.00496764f $X=6.415 $Y=0.82 $X2=0 $Y2=0
cc_433 N_Y_M1002_s N_VGND_c_795_n 0.00255524f $X=2.945 $Y=0.235 $X2=0 $Y2=0
cc_434 N_Y_M1006_s N_VGND_c_795_n 0.00255524f $X=3.885 $Y=0.235 $X2=0 $Y2=0
cc_435 N_Y_M1012_s N_VGND_c_795_n 0.00255524f $X=4.825 $Y=0.235 $X2=0 $Y2=0
cc_436 N_Y_M1020_s N_VGND_c_795_n 0.00304616f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_437 N_Y_c_614_n N_VGND_c_795_n 0.0140924f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_438 N_Y_c_595_n N_VGND_c_795_n 0.00961016f $X=3.855 $Y=0.82 $X2=0 $Y2=0
cc_439 N_Y_c_641_n N_VGND_c_795_n 0.0140924f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_440 N_Y_c_597_n N_VGND_c_795_n 0.00961016f $X=4.795 $Y=0.82 $X2=0 $Y2=0
cc_441 N_Y_c_657_n N_VGND_c_795_n 0.0140924f $X=5.01 $Y=0.4 $X2=0 $Y2=0
cc_442 N_Y_c_598_n N_VGND_c_795_n 0.00961016f $X=5.735 $Y=0.82 $X2=0 $Y2=0
cc_443 N_Y_c_673_n N_VGND_c_795_n 0.0142976f $X=5.95 $Y=0.4 $X2=0 $Y2=0
cc_444 N_Y_c_599_n N_VGND_c_795_n 0.014027f $X=6.415 $Y=0.82 $X2=0 $Y2=0
