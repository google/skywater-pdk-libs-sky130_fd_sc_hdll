* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfrtn_1 CLK_N D RESET_B SCD SCE VGND VNB VPB VPWR Q
M1000 a_1428_47# a_1380_303# a_1322_47# VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=1.518e+11p ps=1.6e+06u
M1001 a_213_47# a_27_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=1.3533e+12p ps=1.268e+07u
M1002 VPWR a_1972_21# a_1951_413# VPB phighvt w=420000u l=180000u
+  ad=1.6398e+12p pd=1.569e+07u as=1.386e+11p ps=1.5e+06u
M1003 a_1972_21# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=1.344e+11p pd=1.48e+06u as=0p ps=0u
M1004 Q a_1972_21# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3.15e+11p pd=2.63e+06u as=0p ps=0u
M1005 a_2157_47# RESET_B VGND VNB nshort w=420000u l=150000u
+  ad=1.386e+11p pd=1.5e+06u as=0p ps=0u
M1006 VPWR SCD a_870_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=1.971e+11p ps=1.81e+06u
M1007 a_700_389# D a_631_119# VNB nshort w=420000u l=150000u
+  ad=3.3215e+11p pd=3.47e+06u as=1.302e+11p ps=1.46e+06u
M1008 a_1380_303# a_1202_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=2.541e+11p pd=2.37e+06u as=0p ps=0u
M1009 a_1202_413# a_213_47# a_700_389# VNB nshort w=360000u l=150000u
+  ad=1.44e+11p pd=1.52e+06u as=0p ps=0u
M1010 VPWR a_1757_47# a_1972_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_1972_21# a_1757_47# a_2157_47# VNB nshort w=420000u l=150000u
+  ad=1.365e+11p pd=1.49e+06u as=0p ps=0u
M1012 Q a_1972_21# VGND VNB nshort w=650000u l=150000u
+  ad=1.9825e+11p pd=1.91e+06u as=0p ps=0u
M1013 VPWR a_1380_303# a_1324_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=2.352e+11p ps=2.8e+06u
M1014 VPWR CLK_N a_27_47# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1015 a_618_389# SCE VPWR VPB phighvt w=540000u l=180000u
+  ad=1.242e+11p pd=1.54e+06u as=0p ps=0u
M1016 a_1951_413# a_27_47# a_1757_47# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.26e+11p ps=1.44e+06u
M1017 a_700_389# D a_618_389# VPB phighvt w=540000u l=180000u
+  ad=5.193e+11p pd=4.01e+06u as=0p ps=0u
M1018 a_631_119# a_331_66# VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VGND RESET_B a_1428_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1020 a_1324_413# RESET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1202_413# a_27_47# a_700_389# VPB phighvt w=420000u l=180000u
+  ad=1.806e+11p pd=1.7e+06u as=0p ps=0u
M1022 a_1324_413# a_213_47# a_1202_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_1866_47# a_213_47# a_1757_47# VNB nshort w=360000u l=150000u
+  ad=2.121e+11p pd=1.9e+06u as=1.422e+11p ps=1.51e+06u
M1024 a_1757_47# a_27_47# a_1380_303# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=1.87e+11p ps=1.93e+06u
M1025 VPWR SCE a_331_66# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=2.214e+11p ps=1.9e+06u
M1026 VGND CLK_N a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.015e+11p ps=1.92e+06u
M1027 VGND a_1972_21# a_1866_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_213_47# a_27_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.75e+11p pd=2.55e+06u as=0p ps=0u
M1029 a_899_66# SCE a_700_389# VNB nshort w=420000u l=500000u
+  ad=1.554e+11p pd=1.58e+06u as=0p ps=0u
M1030 a_1757_47# a_213_47# a_1380_303# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_1322_47# a_27_47# a_1202_413# VNB nshort w=360000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1032 VGND SCD a_899_66# VNB nshort w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1033 a_870_389# a_331_66# a_700_389# VPB phighvt w=540000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1034 VGND SCE a_331_66# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1035 a_1380_303# a_1202_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
