* File: sky130_fd_sc_hdll__nand3b_4.pxi.spice
* Created: Wed Sep  2 08:38:09 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%A_N N_A_N_M1023_g N_A_N_c_100_n N_A_N_M1007_g
+ A_N A_N PM_SKY130_FD_SC_HDLL__NAND3B_4%A_N
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%A_27_47# N_A_27_47#_M1023_s N_A_27_47#_M1007_s
+ N_A_27_47#_c_136_n N_A_27_47#_M1002_g N_A_27_47#_M1005_g N_A_27_47#_c_137_n
+ N_A_27_47#_M1009_g N_A_27_47#_M1006_g N_A_27_47#_c_138_n N_A_27_47#_M1014_g
+ N_A_27_47#_M1008_g N_A_27_47#_c_139_n N_A_27_47#_M1020_g N_A_27_47#_M1018_g
+ N_A_27_47#_c_129_n N_A_27_47#_c_140_n N_A_27_47#_c_141_n N_A_27_47#_c_130_n
+ N_A_27_47#_c_131_n N_A_27_47#_c_186_p N_A_27_47#_c_132_n N_A_27_47#_c_133_n
+ N_A_27_47#_c_134_n N_A_27_47#_c_135_n PM_SKY130_FD_SC_HDLL__NAND3B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%B N_B_M1003_g N_B_c_240_n N_B_M1001_g
+ N_B_M1004_g N_B_c_241_n N_B_M1013_g N_B_M1016_g N_B_c_242_n N_B_M1017_g
+ N_B_c_243_n N_B_M1025_g N_B_M1024_g B B B N_B_c_239_n B B B
+ PM_SKY130_FD_SC_HDLL__NAND3B_4%B
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%C N_C_c_314_n N_C_M1000_g N_C_M1011_g
+ N_C_c_315_n N_C_M1010_g N_C_M1012_g N_C_c_316_n N_C_M1015_g N_C_M1019_g
+ N_C_c_317_n N_C_M1021_g N_C_M1022_g C C C C N_C_c_311_n N_C_c_312_n
+ N_C_c_313_n C C C C PM_SKY130_FD_SC_HDLL__NAND3B_4%C
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%VPWR N_VPWR_M1007_d N_VPWR_M1002_d
+ N_VPWR_M1009_d N_VPWR_M1020_d N_VPWR_M1013_s N_VPWR_M1025_s N_VPWR_M1000_s
+ N_VPWR_M1010_s N_VPWR_M1021_s N_VPWR_c_385_n N_VPWR_c_386_n N_VPWR_c_387_n
+ N_VPWR_c_388_n N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n
+ N_VPWR_c_393_n N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n VPWR N_VPWR_c_401_n
+ N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n N_VPWR_c_384_n VPWR
+ PM_SKY130_FD_SC_HDLL__NAND3B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%Y N_Y_M1005_s N_Y_M1008_s N_Y_M1002_s
+ N_Y_M1014_s N_Y_M1001_d N_Y_M1017_d N_Y_M1000_d N_Y_M1015_d N_Y_c_502_n
+ N_Y_c_505_n N_Y_c_525_n N_Y_c_506_n N_Y_c_532_n N_Y_c_503_n N_Y_c_535_n
+ N_Y_c_507_n N_Y_c_504_n N_Y_c_555_n N_Y_c_509_n N_Y_c_569_n N_Y_c_510_n
+ N_Y_c_511_n N_Y_c_580_n N_Y_c_512_n N_Y_c_513_n Y Y
+ PM_SKY130_FD_SC_HDLL__NAND3B_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%VGND N_VGND_M1023_d N_VGND_M1011_d
+ N_VGND_M1012_d N_VGND_M1022_d N_VGND_c_646_n N_VGND_c_647_n N_VGND_c_648_n
+ N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n N_VGND_c_653_n
+ N_VGND_c_654_n VGND N_VGND_c_655_n N_VGND_c_656_n N_VGND_c_657_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND3B_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%A_225_47# N_A_225_47#_M1005_d
+ N_A_225_47#_M1006_d N_A_225_47#_M1018_d N_A_225_47#_M1004_d
+ N_A_225_47#_M1024_d N_A_225_47#_c_733_n
+ PM_SKY130_FD_SC_HDLL__NAND3B_4%A_225_47#
x_PM_SKY130_FD_SC_HDLL__NAND3B_4%A_683_47# N_A_683_47#_M1003_s
+ N_A_683_47#_M1016_s N_A_683_47#_M1011_s N_A_683_47#_M1019_s
+ N_A_683_47#_c_767_n N_A_683_47#_c_768_n N_A_683_47#_c_781_n
+ N_A_683_47#_c_769_n N_A_683_47#_c_787_n N_A_683_47#_c_770_n
+ N_A_683_47#_c_771_n PM_SKY130_FD_SC_HDLL__NAND3B_4%A_683_47#
cc_1 VNB N_A_N_M1023_g 0.0257996f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_N_c_100_n 0.0302727f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB A_N 0.00171958f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_4 VNB N_A_27_47#_M1005_g 0.0213354f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_5 VNB N_A_27_47#_M1006_g 0.0183665f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1008_g 0.0183647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1018_g 0.0180545f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_129_n 0.0183576f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_130_n 0.0100294f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_131_n 0.00415457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_132_n 0.00993195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_133_n 0.0188173f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_134_n 0.03161f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_135_n 0.0850182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B_M1003_g 0.0182033f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_16 VNB N_B_M1004_g 0.0183647f $X=-0.19 $Y=-0.24 $X2=0.602 $Y2=1.16
cc_17 VNB N_B_M1016_g 0.0188863f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_18 VNB N_B_M1024_g 0.0249344f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB B 0.00259229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_c_239_n 0.0890901f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_C_M1011_g 0.0244336f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_22 VNB N_C_M1012_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_23 VNB N_C_M1019_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_C_M1022_g 0.0244024f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_C_c_311_n 0.0304355f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_C_c_312_n 0.00425884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_C_c_313_n 0.0947773f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_384_n 0.326667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_Y_c_502_n 0.00833823f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_Y_c_503_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_504_n 0.00278804f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_646_n 0.00900466f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_33 VNB N_VGND_c_647_n 0.00878036f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_648_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_649_n 0.0138117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_650_n 0.0363821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_651_n 0.101225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_652_n 0.00477752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_653_n 0.0192454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_654_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_655_n 0.0200877f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_656_n 0.023298f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_657_n 0.379044f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_225_47#_c_733_n 0.00510926f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_683_47#_c_767_n 0.0107074f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.175
cc_46 VNB N_A_683_47#_c_768_n 0.00834731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_683_47#_c_769_n 0.00512293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_683_47#_c_770_n 0.00367221f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_683_47#_c_771_n 0.00233388f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VPB N_A_N_c_100_n 0.0413178f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_A_27_47#_c_136_n 0.0198486f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_52 VPB N_A_27_47#_c_137_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A_27_47#_c_138_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A_27_47#_c_139_n 0.015983f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A_27_47#_c_140_n 0.00865987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB N_A_27_47#_c_141_n 0.0336524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_27_47#_c_133_n 0.00666133f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_27_47#_c_135_n 0.0289602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_B_c_240_n 0.0156532f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_60 VPB N_B_c_241_n 0.0158787f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.16
cc_61 VPB N_B_c_242_n 0.0158686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_B_c_243_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_B_c_239_n 0.0277069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_C_c_314_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.015
cc_65 VPB N_C_c_315_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_66 VPB N_C_c_316_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.175
cc_67 VPB N_C_c_317_n 0.0198539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_C_c_313_n 0.0321197f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_385_n 0.0252173f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_386_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_387_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_388_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_389_n 0.0164978f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_390_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_391_n 0.0137858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_392_n 0.0508068f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_393_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_394_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_395_n 0.0199956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_396_n 0.00323937f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_397_n 0.0201854f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_398_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_399_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_400_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_401_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_402_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_403_n 0.0326056f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_404_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_384_n 0.0468182f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_Y_c_505_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_Y_c_506_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_507_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_Y_c_504_n 0.00720502f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_509_n 0.012664f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_510_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_511_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_Y_c_512_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_513_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 N_A_N_M1023_g N_A_27_47#_c_129_n 0.0112137f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_100 N_A_N_c_100_n N_A_27_47#_c_140_n 0.00376263f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_N_c_100_n N_A_27_47#_c_141_n 0.0106318f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_N_M1023_g N_A_27_47#_c_130_n 0.0112031f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_N_c_100_n N_A_27_47#_c_130_n 0.00643687f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 A_N N_A_27_47#_c_130_n 0.0288482f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_105 N_A_N_M1023_g N_A_27_47#_c_131_n 0.00277479f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_106 N_A_N_c_100_n N_A_27_47#_c_131_n 8.46056e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_107 A_N N_A_27_47#_c_131_n 0.0137035f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_108 N_A_N_M1023_g N_A_27_47#_c_132_n 0.00161631f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_109 N_A_N_M1023_g N_A_27_47#_c_133_n 0.0139959f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_110 A_N N_A_27_47#_c_133_n 0.0152087f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_111 N_A_N_c_100_n N_A_27_47#_c_134_n 0.0153114f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_112 A_N N_A_27_47#_c_134_n 7.44645e-19 $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_113 N_A_N_c_100_n N_A_27_47#_c_135_n 2.90262e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_N_c_100_n N_VPWR_c_385_n 0.0147779f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_115 A_N N_VPWR_c_385_n 0.0150811f $X=0.695 $Y=1.19 $X2=0 $Y2=0
cc_116 N_A_N_c_100_n N_VPWR_c_403_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_N_c_100_n N_VPWR_c_384_n 0.0140376f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_N_M1023_g N_VGND_c_646_n 0.00548508f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_119 N_A_N_M1023_g N_VGND_c_656_n 0.00422241f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_120 N_A_N_M1023_g N_VGND_c_657_n 0.0080996f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_121 N_A_27_47#_M1018_g N_B_M1003_g 0.0216625f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_122 N_A_27_47#_c_139_n N_B_c_240_n 0.0374064f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_27_47#_c_135_n N_B_c_239_n 0.0216625f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_124 N_A_27_47#_c_136_n N_VPWR_c_385_n 0.00989303f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_125 N_A_27_47#_c_140_n N_VPWR_c_385_n 0.0690564f $X=0.255 $Y=1.615 $X2=0
+ $Y2=0
cc_126 N_A_27_47#_c_130_n N_VPWR_c_385_n 0.00855453f $X=1.055 $Y=0.81 $X2=0
+ $Y2=0
cc_127 N_A_27_47#_c_131_n N_VPWR_c_385_n 0.0244885f $X=1.195 $Y=1.075 $X2=0
+ $Y2=0
cc_128 N_A_27_47#_c_134_n N_VPWR_c_385_n 0.00639477f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_129 N_A_27_47#_c_137_n N_VPWR_c_386_n 0.0052072f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_27_47#_c_138_n N_VPWR_c_386_n 0.00474848f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_131 N_A_27_47#_c_139_n N_VPWR_c_387_n 0.00402622f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_132 N_A_27_47#_c_136_n N_VPWR_c_393_n 0.00597712f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A_27_47#_c_137_n N_VPWR_c_393_n 0.00673617f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_27_47#_c_138_n N_VPWR_c_395_n 0.00597712f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_135 N_A_27_47#_c_139_n N_VPWR_c_395_n 0.00563331f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_136 N_A_27_47#_c_141_n N_VPWR_c_403_n 0.0217765f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_137 N_A_27_47#_M1007_s N_VPWR_c_384_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_138 N_A_27_47#_c_136_n N_VPWR_c_384_n 0.0112769f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_27_47#_c_137_n N_VPWR_c_384_n 0.0118438f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_27_47#_c_138_n N_VPWR_c_384_n 0.00999457f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_27_47#_c_139_n N_VPWR_c_384_n 0.00839257f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_27_47#_c_141_n N_VPWR_c_384_n 0.0128576f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_143 N_A_27_47#_M1005_g N_Y_c_502_n 0.00922668f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_144 N_A_27_47#_M1006_g N_Y_c_502_n 0.0117281f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_145 N_A_27_47#_M1008_g N_Y_c_502_n 0.0117222f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_146 N_A_27_47#_M1018_g N_Y_c_502_n 0.0121451f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_147 N_A_27_47#_c_130_n N_Y_c_502_n 0.0165524f $X=1.055 $Y=0.81 $X2=0 $Y2=0
cc_148 N_A_27_47#_c_186_p N_Y_c_502_n 0.0976508f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_27_47#_c_135_n N_Y_c_502_n 0.00970138f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_150 N_A_27_47#_c_136_n N_Y_c_505_n 0.0046976f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_27_47#_c_137_n N_Y_c_505_n 0.00116723f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_27_47#_c_186_p N_Y_c_505_n 0.0305808f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_135_n N_Y_c_505_n 0.0074788f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_136_n N_Y_c_525_n 0.0121679f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_137_n N_Y_c_525_n 0.0106224f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A_27_47#_c_138_n N_Y_c_525_n 6.24491e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_137_n N_Y_c_506_n 0.0153933f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_138_n N_Y_c_506_n 0.0113962f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_186_p N_Y_c_506_n 0.040258f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_135_n N_Y_c_506_n 0.00725062f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_138_n N_Y_c_532_n 0.00699422f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_139_n N_Y_c_532_n 0.00665381f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_27_47#_M1018_g N_Y_c_503_n 0.00410511f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_139_n N_Y_c_535_n 5.5123e-19 $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_137_n N_Y_c_504_n 5.15343e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_138_n N_Y_c_504_n 0.00902851f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_139_n N_Y_c_504_n 0.0247886f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_186_p N_Y_c_504_n 0.044778f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_135_n N_Y_c_504_n 0.0140587f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_130_n N_VGND_M1023_d 0.00420907f $X=1.055 $Y=0.81 $X2=-0.19
+ $Y2=-0.24
cc_171 N_A_27_47#_M1005_g N_VGND_c_646_n 0.0021243f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_129_n N_VGND_c_646_n 0.0181155f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_130_n N_VGND_c_646_n 0.0196192f $X=1.055 $Y=0.81 $X2=0 $Y2=0
cc_174 N_A_27_47#_M1005_g N_VGND_c_651_n 0.00357877f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_175 N_A_27_47#_M1006_g N_VGND_c_651_n 0.00357877f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_176 N_A_27_47#_M1008_g N_VGND_c_651_n 0.00357877f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1018_g N_VGND_c_651_n 0.00357877f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_130_n N_VGND_c_651_n 0.00300337f $X=1.055 $Y=0.81 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_129_n N_VGND_c_656_n 0.0217307f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_130_n N_VGND_c_656_n 0.00273345f $X=1.055 $Y=0.81 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_M1023_s N_VGND_c_657_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_M1005_g N_VGND_c_657_n 0.00668309f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1006_g N_VGND_c_657_n 0.00548399f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1008_g N_VGND_c_657_n 0.00548399f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1018_g N_VGND_c_657_n 0.00538422f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_129_n N_VGND_c_657_n 0.0128045f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_130_n N_VGND_c_657_n 0.0121755f $X=1.055 $Y=0.81 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_130_n N_A_225_47#_M1005_d 0.00555397f $X=1.055 $Y=0.81
+ $X2=-0.19 $Y2=-0.24
cc_189 N_A_27_47#_M1005_g N_A_225_47#_c_733_n 0.00999874f $X=1.51 $Y=0.56 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1006_g N_A_225_47#_c_733_n 0.00903374f $X=1.98 $Y=0.56 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_M1008_g N_A_225_47#_c_733_n 0.00903374f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_192 N_A_27_47#_M1018_g N_A_225_47#_c_733_n 0.00903374f $X=2.92 $Y=0.56 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_130_n N_A_225_47#_c_733_n 0.0139638f $X=1.055 $Y=0.81 $X2=0
+ $Y2=0
cc_194 N_A_27_47#_c_186_p N_A_225_47#_c_733_n 0.00348368f $X=2.66 $Y=1.16 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_134_n N_A_225_47#_c_733_n 0.00249878f $X=1.385 $Y=1.16 $X2=0
+ $Y2=0
cc_196 B N_C_c_311_n 6.97286e-19 $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_197 N_B_c_239_n N_C_c_311_n 0.00741568f $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_198 B N_C_c_312_n 0.0139438f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_199 N_B_c_239_n N_C_c_312_n 8.43693e-19 $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_200 N_B_c_240_n N_VPWR_c_387_n 0.00381622f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_241_n N_VPWR_c_388_n 0.00520479f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_242_n N_VPWR_c_388_n 0.004751f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_243_n N_VPWR_c_389_n 0.00825342f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_240_n N_VPWR_c_397_n 0.00537104f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_c_241_n N_VPWR_c_397_n 0.00673617f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_242_n N_VPWR_c_401_n 0.00597712f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_243_n N_VPWR_c_401_n 0.00673617f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_240_n N_VPWR_c_384_n 0.00812353f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_241_n N_VPWR_c_384_n 0.0118438f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_242_n N_VPWR_c_384_n 0.00999457f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_243_n N_VPWR_c_384_n 0.0131262f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_M1003_g N_Y_c_502_n 0.00121164f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_213 N_B_c_240_n N_Y_c_532_n 5.16456e-19 $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B_M1003_g N_Y_c_503_n 0.00410511f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_215 N_B_c_240_n N_Y_c_535_n 0.00832135f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B_c_241_n N_Y_c_535_n 0.00551548f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B_c_241_n N_Y_c_507_n 0.0153933f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_242_n N_Y_c_507_n 0.0113962f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_219 B N_Y_c_507_n 0.040258f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_220 N_B_c_239_n N_Y_c_507_n 0.00725062f $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_221 N_B_c_240_n N_Y_c_504_n 0.0193107f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_222 N_B_c_241_n N_Y_c_504_n 0.00718431f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_242_n N_Y_c_504_n 4.76697e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_224 B N_Y_c_504_n 0.0195734f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_225 N_B_c_239_n N_Y_c_504_n 0.0326746f $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_226 N_B_c_241_n N_Y_c_555_n 6.4818e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_227 N_B_c_242_n N_Y_c_555_n 0.0130681f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_228 N_B_c_243_n N_Y_c_555_n 0.0153658f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_243_n N_Y_c_509_n 0.0179883f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_230 B N_Y_c_509_n 0.016181f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_231 N_B_c_239_n N_Y_c_509_n 3.10838e-19 $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_232 N_B_c_242_n N_Y_c_512_n 0.00292783f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B_c_243_n N_Y_c_512_n 0.00116723f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_234 B N_Y_c_512_n 0.0305808f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_235 N_B_c_239_n N_Y_c_512_n 0.00723098f $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_236 N_B_M1024_g N_VGND_c_647_n 0.00231165f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_237 N_B_M1003_g N_VGND_c_651_n 0.00357877f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_238 N_B_M1004_g N_VGND_c_651_n 0.00357877f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_239 N_B_M1016_g N_VGND_c_651_n 0.00357877f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_240 N_B_M1024_g N_VGND_c_651_n 0.00357877f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_241 N_B_M1003_g N_VGND_c_657_n 0.00538422f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_242 N_B_M1004_g N_VGND_c_657_n 0.00548399f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_243 N_B_M1016_g N_VGND_c_657_n 0.00560377f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_244 N_B_M1024_g N_VGND_c_657_n 0.00680287f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_245 N_B_M1003_g N_A_225_47#_c_733_n 0.0106952f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_246 N_B_M1004_g N_A_225_47#_c_733_n 0.00903374f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_247 N_B_M1016_g N_A_225_47#_c_733_n 0.00935436f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_248 N_B_M1024_g N_A_225_47#_c_733_n 0.00935436f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_249 N_B_M1003_g N_A_683_47#_c_767_n 0.00386108f $X=3.34 $Y=0.56 $X2=0 $Y2=0
cc_250 N_B_M1004_g N_A_683_47#_c_767_n 0.0117281f $X=3.81 $Y=0.56 $X2=0 $Y2=0
cc_251 N_B_M1016_g N_A_683_47#_c_767_n 0.0117558f $X=4.28 $Y=0.56 $X2=0 $Y2=0
cc_252 N_B_M1024_g N_A_683_47#_c_767_n 0.014325f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_253 B N_A_683_47#_c_767_n 0.0889433f $X=4.745 $Y=1.105 $X2=0 $Y2=0
cc_254 N_B_c_239_n N_A_683_47#_c_767_n 0.0112736f $X=4.775 $Y=1.217 $X2=0 $Y2=0
cc_255 N_C_c_314_n N_VPWR_c_389_n 0.00762417f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_256 N_C_c_315_n N_VPWR_c_390_n 0.0052072f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_257 N_C_c_316_n N_VPWR_c_390_n 0.004751f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_258 N_C_c_317_n N_VPWR_c_392_n 0.0297018f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_259 N_C_c_314_n N_VPWR_c_399_n 0.00597712f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_260 N_C_c_315_n N_VPWR_c_399_n 0.00673617f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_261 N_C_c_316_n N_VPWR_c_402_n 0.00597712f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_262 N_C_c_317_n N_VPWR_c_402_n 0.00673617f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_263 N_C_c_314_n N_VPWR_c_384_n 0.0112769f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_264 N_C_c_315_n N_VPWR_c_384_n 0.0118438f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_265 N_C_c_316_n N_VPWR_c_384_n 0.00999457f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_266 N_C_c_317_n N_VPWR_c_384_n 0.0129848f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_267 N_C_c_314_n N_Y_c_509_n 0.0139912f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_268 N_C_c_311_n N_Y_c_509_n 0.00729564f $X=5.665 $Y=1.16 $X2=0 $Y2=0
cc_269 N_C_c_312_n N_Y_c_509_n 0.0444134f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_270 N_C_c_313_n N_Y_c_509_n 2.73568e-19 $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_271 N_C_c_314_n N_Y_c_569_n 0.0178402f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_272 N_C_c_315_n N_Y_c_569_n 0.0106251f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_273 N_C_c_316_n N_Y_c_569_n 6.24674e-19 $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_274 N_C_c_315_n N_Y_c_510_n 0.0153933f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_275 N_C_c_316_n N_Y_c_510_n 0.0113962f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_276 N_C_c_312_n N_Y_c_510_n 0.040258f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_277 N_C_c_313_n N_Y_c_510_n 0.00725062f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_278 N_C_c_316_n N_Y_c_511_n 0.00292783f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_279 N_C_c_317_n N_Y_c_511_n 0.00356328f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_280 N_C_c_312_n N_Y_c_511_n 0.0301956f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_281 N_C_c_313_n N_Y_c_511_n 0.0074788f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_282 N_C_c_315_n N_Y_c_580_n 6.48386e-19 $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_283 N_C_c_316_n N_Y_c_580_n 0.0130707f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_284 N_C_c_317_n N_Y_c_580_n 0.0100147f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_285 N_C_c_314_n N_Y_c_513_n 0.00292783f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_286 N_C_c_315_n N_Y_c_513_n 0.00116723f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_287 N_C_c_312_n N_Y_c_513_n 0.0305808f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_288 N_C_c_313_n N_Y_c_513_n 0.0074788f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_289 N_C_M1011_g N_VGND_c_647_n 0.0052731f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_290 N_C_M1012_g N_VGND_c_648_n 0.00276126f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_291 N_C_M1019_g N_VGND_c_648_n 0.0035663f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_292 N_C_M1022_g N_VGND_c_650_n 0.0175467f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_293 N_C_M1011_g N_VGND_c_653_n 0.00395968f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_294 N_C_M1012_g N_VGND_c_653_n 0.00436487f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_295 N_C_M1019_g N_VGND_c_655_n 0.00395968f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_296 N_C_M1022_g N_VGND_c_655_n 0.00585385f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_297 N_C_M1011_g N_VGND_c_657_n 0.0070025f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_298 N_C_M1012_g N_VGND_c_657_n 0.0061161f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_299 N_C_M1019_g N_VGND_c_657_n 0.0058034f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_300 N_C_M1022_g N_VGND_c_657_n 0.0118511f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_301 N_C_M1011_g N_A_683_47#_c_768_n 0.0084307f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_302 N_C_c_311_n N_A_683_47#_c_768_n 0.00889913f $X=5.665 $Y=1.16 $X2=0 $Y2=0
cc_303 N_C_c_312_n N_A_683_47#_c_768_n 0.0440565f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_304 N_C_M1011_g N_A_683_47#_c_781_n 0.0111702f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_305 N_C_M1012_g N_A_683_47#_c_769_n 0.0111881f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_306 N_C_M1019_g N_A_683_47#_c_769_n 0.0091819f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_307 N_C_M1022_g N_A_683_47#_c_769_n 2.01812e-19 $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_308 N_C_c_312_n N_A_683_47#_c_769_n 0.0700927f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_309 N_C_c_313_n N_A_683_47#_c_769_n 0.00652443f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_310 N_C_M1012_g N_A_683_47#_c_787_n 5.79378e-19 $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_311 N_C_M1019_g N_A_683_47#_c_787_n 0.00837042f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_312 N_C_M1011_g N_A_683_47#_c_770_n 0.00129432f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_313 N_C_M1011_g N_A_683_47#_c_771_n 0.00281161f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_314 N_C_c_312_n N_A_683_47#_c_771_n 0.030512f $X=6.935 $Y=1.16 $X2=0 $Y2=0
cc_315 N_C_c_313_n N_A_683_47#_c_771_n 0.00332f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_316 N_VPWR_c_384_n N_Y_M1002_s 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_317 N_VPWR_c_384_n N_Y_M1014_s 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_384_n N_Y_M1001_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_319 N_VPWR_c_384_n N_Y_M1017_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_384_n N_Y_M1000_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_321 N_VPWR_c_384_n N_Y_M1015_d 0.00231261f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_c_385_n N_Y_c_505_n 0.0192276f $X=0.73 $Y=1.66 $X2=0 $Y2=0
cc_323 N_VPWR_c_385_n N_Y_c_525_n 0.066442f $X=0.73 $Y=1.66 $X2=0 $Y2=0
cc_324 N_VPWR_c_386_n N_Y_c_525_n 0.0385613f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_c_393_n N_Y_c_525_n 0.0223557f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_326 N_VPWR_c_384_n N_Y_c_525_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_M1009_d N_Y_c_506_n 0.00180012f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_328 N_VPWR_c_386_n N_Y_c_506_n 0.0139097f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_329 N_VPWR_c_386_n N_Y_c_532_n 0.034303f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_330 N_VPWR_c_387_n N_Y_c_532_n 0.0177504f $X=3.13 $Y=2.34 $X2=0 $Y2=0
cc_331 N_VPWR_c_395_n N_Y_c_532_n 0.0223557f $X=3.045 $Y=2.72 $X2=0 $Y2=0
cc_332 N_VPWR_c_384_n N_Y_c_532_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_333 N_VPWR_c_387_n N_Y_c_535_n 0.02165f $X=3.13 $Y=2.34 $X2=0 $Y2=0
cc_334 N_VPWR_c_388_n N_Y_c_535_n 0.0281247f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_335 N_VPWR_c_397_n N_Y_c_535_n 0.0223557f $X=3.985 $Y=2.72 $X2=0 $Y2=0
cc_336 N_VPWR_c_384_n N_Y_c_535_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_337 N_VPWR_M1013_s N_Y_c_507_n 0.00180012f $X=3.925 $Y=1.485 $X2=0 $Y2=0
cc_338 N_VPWR_c_388_n N_Y_c_507_n 0.0139097f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_339 N_VPWR_M1020_d N_Y_c_504_n 0.00181151f $X=2.985 $Y=1.485 $X2=0 $Y2=0
cc_340 N_VPWR_c_386_n N_Y_c_504_n 0.0133617f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_341 N_VPWR_c_387_n N_Y_c_504_n 0.0144908f $X=3.13 $Y=2.34 $X2=0 $Y2=0
cc_342 N_VPWR_c_388_n N_Y_c_504_n 0.0109394f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_343 N_VPWR_c_395_n N_Y_c_504_n 0.00214482f $X=3.045 $Y=2.72 $X2=0 $Y2=0
cc_344 N_VPWR_c_397_n N_Y_c_504_n 0.001415f $X=3.985 $Y=2.72 $X2=0 $Y2=0
cc_345 N_VPWR_c_384_n N_Y_c_504_n 0.00810304f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_346 N_VPWR_c_388_n N_Y_c_555_n 0.0470327f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_347 N_VPWR_c_389_n N_Y_c_555_n 0.0429581f $X=5.01 $Y=2 $X2=0 $Y2=0
cc_348 N_VPWR_c_401_n N_Y_c_555_n 0.0223557f $X=4.925 $Y=2.72 $X2=0 $Y2=0
cc_349 N_VPWR_c_384_n N_Y_c_555_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_350 N_VPWR_M1025_s N_Y_c_509_n 0.00313113f $X=4.865 $Y=1.485 $X2=0 $Y2=0
cc_351 N_VPWR_M1000_s N_Y_c_509_n 0.00313113f $X=5.405 $Y=1.485 $X2=0 $Y2=0
cc_352 N_VPWR_c_389_n N_Y_c_509_n 0.0578207f $X=5.01 $Y=2 $X2=0 $Y2=0
cc_353 N_VPWR_c_389_n N_Y_c_569_n 0.0523533f $X=5.01 $Y=2 $X2=0 $Y2=0
cc_354 N_VPWR_c_390_n N_Y_c_569_n 0.0385613f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_355 N_VPWR_c_399_n N_Y_c_569_n 0.0223557f $X=6.385 $Y=2.72 $X2=0 $Y2=0
cc_356 N_VPWR_c_384_n N_Y_c_569_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_357 N_VPWR_M1010_s N_Y_c_510_n 0.00180012f $X=6.325 $Y=1.485 $X2=0 $Y2=0
cc_358 N_VPWR_c_390_n N_Y_c_510_n 0.0139097f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_359 N_VPWR_c_392_n N_Y_c_511_n 0.0149111f $X=7.49 $Y=1.66 $X2=0 $Y2=0
cc_360 N_VPWR_c_390_n N_Y_c_580_n 0.0470327f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_361 N_VPWR_c_392_n N_Y_c_580_n 0.05144f $X=7.49 $Y=1.66 $X2=0 $Y2=0
cc_362 N_VPWR_c_402_n N_Y_c_580_n 0.0223557f $X=7.325 $Y=2.72 $X2=0 $Y2=0
cc_363 N_VPWR_c_384_n N_Y_c_580_n 0.0140101f $X=7.59 $Y=2.72 $X2=0 $Y2=0
cc_364 N_VPWR_c_392_n N_VGND_c_650_n 0.0137178f $X=7.49 $Y=1.66 $X2=0 $Y2=0
cc_365 N_Y_M1005_s N_VGND_c_657_n 0.00256987f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_366 N_Y_M1008_s N_VGND_c_657_n 0.00256987f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_367 N_Y_c_502_n N_A_225_47#_M1006_d 0.00214196f $X=3.045 $Y=0.77 $X2=0 $Y2=0
cc_368 N_Y_c_502_n N_A_225_47#_M1018_d 0.00206479f $X=3.045 $Y=0.77 $X2=0 $Y2=0
cc_369 N_Y_M1005_s N_A_225_47#_c_733_n 0.00401386f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_370 N_Y_M1008_s N_A_225_47#_c_733_n 0.00401386f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_371 N_Y_c_502_n N_A_225_47#_c_733_n 0.0925712f $X=3.045 $Y=0.77 $X2=0 $Y2=0
cc_372 N_Y_c_504_n N_A_225_47#_c_733_n 0.00415296f $X=3.765 $Y=1.555 $X2=0 $Y2=0
cc_373 N_Y_c_502_n N_A_683_47#_c_767_n 0.0121859f $X=3.045 $Y=0.77 $X2=0 $Y2=0
cc_374 N_Y_c_504_n N_A_683_47#_c_767_n 0.0205179f $X=3.765 $Y=1.555 $X2=0 $Y2=0
cc_375 N_Y_c_509_n N_A_683_47#_c_767_n 0.00906097f $X=5.785 $Y=1.555 $X2=0 $Y2=0
cc_376 N_VGND_c_657_n N_A_225_47#_M1005_d 0.00250339f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_377 N_VGND_c_657_n N_A_225_47#_M1006_d 0.00255381f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_378 N_VGND_c_657_n N_A_225_47#_M1018_d 0.00215227f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_379 N_VGND_c_657_n N_A_225_47#_M1004_d 0.00255381f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_380 N_VGND_c_657_n N_A_225_47#_M1024_d 0.00209344f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_381 N_VGND_c_646_n N_A_225_47#_c_733_n 0.0166763f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_382 N_VGND_c_647_n N_A_225_47#_c_733_n 0.0166762f $X=5.53 $Y=0.38 $X2=0 $Y2=0
cc_383 N_VGND_c_651_n N_A_225_47#_c_733_n 0.234075f $X=5.365 $Y=0 $X2=0 $Y2=0
cc_384 N_VGND_c_657_n N_A_225_47#_c_733_n 0.147f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_385 N_VGND_c_657_n N_A_683_47#_M1003_s 0.00256987f $X=7.59 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_386 N_VGND_c_657_n N_A_683_47#_M1016_s 0.00297142f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_387 N_VGND_c_657_n N_A_683_47#_M1011_s 0.0026371f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_388 N_VGND_c_657_n N_A_683_47#_M1019_s 0.00324782f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_389 N_VGND_M1011_d N_A_683_47#_c_768_n 0.00420907f $X=5.405 $Y=0.235 $X2=0
+ $Y2=0
cc_390 N_VGND_c_647_n N_A_683_47#_c_768_n 0.0196192f $X=5.53 $Y=0.38 $X2=0 $Y2=0
cc_391 N_VGND_c_651_n N_A_683_47#_c_768_n 0.00296114f $X=5.365 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_653_n N_A_683_47#_c_768_n 0.0020445f $X=6.385 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_657_n N_A_683_47#_c_768_n 0.0102777f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_647_n N_A_683_47#_c_781_n 0.0222763f $X=5.53 $Y=0.38 $X2=0 $Y2=0
cc_395 N_VGND_c_653_n N_A_683_47#_c_781_n 0.023074f $X=6.385 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_657_n N_A_683_47#_c_781_n 0.0141066f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_M1012_d N_A_683_47#_c_769_n 0.0025045f $X=6.335 $Y=0.235 $X2=0
+ $Y2=0
cc_398 N_VGND_c_648_n N_A_683_47#_c_769_n 0.0127393f $X=6.47 $Y=0.38 $X2=0 $Y2=0
cc_399 N_VGND_c_650_n N_A_683_47#_c_769_n 0.00140016f $X=7.49 $Y=0.38 $X2=0
+ $Y2=0
cc_400 N_VGND_c_653_n N_A_683_47#_c_769_n 0.00260993f $X=6.385 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_655_n N_A_683_47#_c_769_n 0.0020445f $X=7.325 $Y=0 $X2=0 $Y2=0
cc_402 N_VGND_c_657_n N_A_683_47#_c_769_n 0.00988931f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_403 N_VGND_c_648_n N_A_683_47#_c_787_n 0.0216501f $X=6.47 $Y=0.38 $X2=0 $Y2=0
cc_404 N_VGND_c_655_n N_A_683_47#_c_787_n 0.023074f $X=7.325 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_657_n N_A_683_47#_c_787_n 0.0141066f $X=7.59 $Y=0 $X2=0 $Y2=0
cc_406 N_A_225_47#_c_733_n N_A_683_47#_M1003_s 0.00401386f $X=5.01 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_407 N_A_225_47#_c_733_n N_A_683_47#_M1016_s 0.00508685f $X=5.01 $Y=0.38 $X2=0
+ $Y2=0
cc_408 N_A_225_47#_M1004_d N_A_683_47#_c_767_n 0.00214196f $X=3.885 $Y=0.235
+ $X2=0 $Y2=0
cc_409 N_A_225_47#_M1024_d N_A_683_47#_c_767_n 0.00111257f $X=4.875 $Y=0.235
+ $X2=0 $Y2=0
cc_410 N_A_225_47#_c_733_n N_A_683_47#_c_767_n 0.0983164f $X=5.01 $Y=0.38 $X2=0
+ $Y2=0
cc_411 N_A_225_47#_M1024_d N_A_683_47#_c_770_n 0.00209037f $X=4.875 $Y=0.235
+ $X2=0 $Y2=0
