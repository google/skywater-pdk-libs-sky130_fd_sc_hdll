* File: sky130_fd_sc_hdll__o21a_1.pxi.spice
* Created: Wed Sep  2 08:43:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21A_1%A_83_21# N_A_83_21#_M1003_s N_A_83_21#_M1005_d
+ N_A_83_21#_c_46_n N_A_83_21#_M1002_g N_A_83_21#_c_47_n N_A_83_21#_M1000_g
+ N_A_83_21#_c_48_n N_A_83_21#_c_53_n N_A_83_21#_c_82_p N_A_83_21#_c_49_n
+ N_A_83_21#_c_50_n N_A_83_21#_c_54_n N_A_83_21#_c_70_p
+ PM_SKY130_FD_SC_HDLL__O21A_1%A_83_21#
x_PM_SKY130_FD_SC_HDLL__O21A_1%B1 N_B1_c_107_n N_B1_M1005_g N_B1_c_108_n
+ N_B1_M1003_g B1 N_B1_c_109_n B1 N_B1_X9_noxref_CONDUCTOR
+ PM_SKY130_FD_SC_HDLL__O21A_1%B1
x_PM_SKY130_FD_SC_HDLL__O21A_1%A2 N_A2_c_136_n N_A2_M1004_g N_A2_c_137_n
+ N_A2_M1001_g A2 N_A2_c_138_n N_A2_c_139_n PM_SKY130_FD_SC_HDLL__O21A_1%A2
x_PM_SKY130_FD_SC_HDLL__O21A_1%A1 N_A1_c_176_n N_A1_M1007_g N_A1_c_177_n
+ N_A1_M1006_g A1 N_A1_c_178_n PM_SKY130_FD_SC_HDLL__O21A_1%A1
x_PM_SKY130_FD_SC_HDLL__O21A_1%X N_X_M1002_s N_X_M1000_s N_X_c_201_n N_X_c_202_n
+ X N_X_c_203_n PM_SKY130_FD_SC_HDLL__O21A_1%X
x_PM_SKY130_FD_SC_HDLL__O21A_1%VPWR N_VPWR_M1000_d N_VPWR_M1006_d N_VPWR_c_222_n
+ VPWR N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_226_n
+ N_VPWR_c_221_n PM_SKY130_FD_SC_HDLL__O21A_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O21A_1%VGND N_VGND_M1002_d N_VGND_M1004_d N_VGND_c_261_n
+ N_VGND_c_262_n VGND N_VGND_c_263_n N_VGND_c_264_n N_VGND_c_265_n
+ N_VGND_c_266_n N_VGND_c_267_n PM_SKY130_FD_SC_HDLL__O21A_1%VGND
x_PM_SKY130_FD_SC_HDLL__O21A_1%A_302_47# N_A_302_47#_M1003_d N_A_302_47#_M1007_d
+ N_A_302_47#_c_303_n N_A_302_47#_c_304_n N_A_302_47#_c_305_n
+ PM_SKY130_FD_SC_HDLL__O21A_1%A_302_47#
cc_1 VNB N_A_83_21#_c_46_n 0.0230738f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_83_21#_c_47_n 0.0345033f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_3 VNB N_A_83_21#_c_48_n 0.00503065f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_4 VNB N_A_83_21#_c_49_n 0.00979926f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.715
cc_5 VNB N_A_83_21#_c_50_n 0.00613503f $X=-0.19 $Y=-0.24 $X2=1.22 $Y2=0.4
cc_6 VNB N_B1_c_107_n 0.0224608f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.235
cc_7 VNB N_B1_c_108_n 0.0200494f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B1_c_109_n 0.00840093f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_9 VNB N_A2_c_136_n 0.0167728f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.235
cc_10 VNB N_A2_c_137_n 0.0200686f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A2_c_138_n 4.71823e-19 $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_12 VNB N_A2_c_139_n 0.00470838f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.4
cc_13 VNB N_A1_c_176_n 0.0222311f $X=-0.19 $Y=-0.24 $X2=1.095 $Y2=0.235
cc_14 VNB N_A1_c_177_n 0.0329435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_178_n 0.00909117f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_16 VNB N_X_c_201_n 0.0240441f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.56
cc_17 VNB N_X_c_202_n 0.00923964f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_18 VNB N_X_c_203_n 0.0137431f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.16
cc_19 VNB N_VPWR_c_221_n 0.136896f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.81
cc_20 VNB N_VGND_c_261_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_21 VNB N_VGND_c_262_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0.742 $Y2=1.16
cc_22 VNB N_VGND_c_263_n 0.0316376f $X=-0.19 $Y=-0.24 $X2=0.885 $Y2=1.582
cc_23 VNB N_VGND_c_264_n 0.0320977f $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=2.34
cc_24 VNB N_VGND_c_265_n 0.201121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_266_n 0.0216012f $X=-0.19 $Y=-0.24 $X2=1.205 $Y2=0.81
cc_26 VNB N_VGND_c_267_n 0.0032427f $X=-0.19 $Y=-0.24 $X2=1.645 $Y2=1.66
cc_27 VNB N_A_302_47#_c_303_n 0.0166886f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_28 VNB N_A_302_47#_c_304_n 0.0180521f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.985
cc_29 VNB N_A_302_47#_c_305_n 0.0031677f $X=-0.19 $Y=-0.24 $X2=0.742 $Y2=1.475
cc_30 VPB N_A_83_21#_c_47_n 0.0342049f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_31 VPB N_A_83_21#_c_48_n 0.00202704f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_32 VPB N_A_83_21#_c_53_n 0.00439336f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.582
cc_33 VPB N_A_83_21#_c_54_n 0.00389781f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.69
cc_34 VPB N_B1_c_107_n 0.0285447f $X=-0.19 $Y=1.305 $X2=1.095 $Y2=0.235
cc_35 VPB N_A2_c_137_n 0.0264118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A2_c_138_n 0.00245533f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_37 VPB N_A1_c_177_n 0.0321953f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_A1_c_178_n 0.00675685f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.985
cc_39 VPB N_X_c_203_n 0.0475183f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=1.16
cc_40 VPB N_VPWR_c_222_n 0.00206262f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=0.56
cc_41 VPB N_VPWR_c_223_n 0.0155059f $X=-0.19 $Y=1.305 $X2=0.742 $Y2=0.905
cc_42 VPB N_VPWR_c_224_n 0.0287285f $X=-0.19 $Y=1.305 $X2=1.48 $Y2=1.582
cc_43 VPB N_VPWR_c_225_n 0.011382f $X=-0.19 $Y=1.305 $X2=1.645 $Y2=1.69
cc_44 VPB N_VPWR_c_226_n 0.0489168f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB N_VPWR_c_221_n 0.0442805f $X=-0.19 $Y=1.305 $X2=1.205 $Y2=0.81
cc_46 N_A_83_21#_c_47_n N_B1_c_107_n 0.0170768f $X=0.515 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_47 N_A_83_21#_c_48_n N_B1_c_107_n 0.00571992f $X=0.685 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_48 N_A_83_21#_c_53_n N_B1_c_107_n 0.0227877f $X=1.48 $Y=1.582 $X2=-0.19
+ $Y2=-0.24
cc_49 N_A_83_21#_c_49_n N_B1_c_107_n 0.00345035f $X=1.205 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_50 N_A_83_21#_c_54_n N_B1_c_107_n 8.36819e-19 $X=1.645 $Y=1.69 $X2=-0.19
+ $Y2=-0.24
cc_51 N_A_83_21#_c_48_n N_B1_c_108_n 0.00236697f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_52 N_A_83_21#_c_49_n N_B1_c_108_n 0.00281855f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_53 N_A_83_21#_c_50_n N_B1_c_108_n 0.00740708f $X=1.22 $Y=0.4 $X2=0 $Y2=0
cc_54 N_A_83_21#_c_47_n N_B1_c_109_n 8.05495e-19 $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_83_21#_c_48_n N_B1_c_109_n 0.019476f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_56 N_A_83_21#_c_53_n N_B1_c_109_n 0.0316569f $X=1.48 $Y=1.582 $X2=0 $Y2=0
cc_57 N_A_83_21#_c_49_n N_B1_c_109_n 0.0249787f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_58 N_A_83_21#_c_54_n N_B1_c_109_n 0.00634969f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_59 N_A_83_21#_c_50_n N_A2_c_136_n 9.04416e-19 $X=1.22 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_60 N_A_83_21#_c_54_n N_A2_c_137_n 0.00305536f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_61 N_A_83_21#_c_70_p N_A2_c_137_n 0.00898749f $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_62 N_A_83_21#_c_54_n N_A2_c_138_n 0.00922326f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_63 N_A_83_21#_c_54_n N_A2_c_139_n 0.00626176f $X=1.645 $Y=1.69 $X2=0 $Y2=0
cc_64 N_A_83_21#_c_70_p N_A1_c_177_n 3.95309e-19 $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_65 N_A_83_21#_c_46_n N_X_c_201_n 0.00778053f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_66 N_A_83_21#_c_49_n N_X_c_201_n 0.0077405f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_67 N_A_83_21#_c_50_n N_X_c_201_n 0.00523487f $X=1.22 $Y=0.4 $X2=0 $Y2=0
cc_68 N_A_83_21#_c_46_n N_X_c_202_n 0.0035265f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A_83_21#_c_47_n N_X_c_202_n 0.00168031f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A_83_21#_c_48_n N_X_c_202_n 0.00940917f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_71 N_A_83_21#_c_47_n N_X_c_203_n 0.0186919f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_83_21#_c_48_n N_X_c_203_n 0.0269108f $X=0.685 $Y=1.16 $X2=0 $Y2=0
cc_73 N_A_83_21#_c_82_p N_X_c_203_n 0.0136425f $X=0.885 $Y=1.582 $X2=0 $Y2=0
cc_74 N_A_83_21#_c_53_n N_VPWR_M1000_d 0.00523862f $X=1.48 $Y=1.582 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_83_21#_c_82_p N_VPWR_M1000_d 0.0034447f $X=0.885 $Y=1.582 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_83_21#_c_47_n N_VPWR_c_222_n 0.0208306f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_83_21#_c_53_n N_VPWR_c_222_n 0.026465f $X=1.48 $Y=1.582 $X2=0 $Y2=0
cc_78 N_A_83_21#_c_82_p N_VPWR_c_222_n 0.0204447f $X=0.885 $Y=1.582 $X2=0 $Y2=0
cc_79 N_A_83_21#_c_47_n N_VPWR_c_223_n 0.00427505f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_83_21#_c_70_p N_VPWR_c_224_n 0.0207969f $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_81 N_A_83_21#_c_70_p N_VPWR_c_226_n 0.00224253f $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_82 N_A_83_21#_M1005_d N_VPWR_c_221_n 0.00465323f $X=1.43 $Y=1.485 $X2=0 $Y2=0
cc_83 N_A_83_21#_c_47_n N_VPWR_c_221_n 0.00825932f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_83_21#_c_70_p N_VPWR_c_221_n 0.0124725f $X=1.645 $Y=2.34 $X2=0 $Y2=0
cc_85 N_A_83_21#_c_49_n N_VGND_M1002_d 0.00355962f $X=1.205 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_83_21#_c_46_n N_VGND_c_261_n 0.00438629f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_83_21#_c_49_n N_VGND_c_261_n 0.0127393f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_88 N_A_83_21#_c_50_n N_VGND_c_261_n 0.0177842f $X=1.22 $Y=0.4 $X2=0 $Y2=0
cc_89 N_A_83_21#_c_49_n N_VGND_c_263_n 0.0037506f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_90 N_A_83_21#_c_50_n N_VGND_c_263_n 0.0226055f $X=1.22 $Y=0.4 $X2=0 $Y2=0
cc_91 N_A_83_21#_M1003_s N_VGND_c_265_n 0.00213418f $X=1.095 $Y=0.235 $X2=0
+ $Y2=0
cc_92 N_A_83_21#_c_46_n N_VGND_c_265_n 0.0125402f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_83_21#_c_49_n N_VGND_c_265_n 0.00756473f $X=1.205 $Y=0.715 $X2=0 $Y2=0
cc_94 N_A_83_21#_c_50_n N_VGND_c_265_n 0.0134689f $X=1.22 $Y=0.4 $X2=0 $Y2=0
cc_95 N_A_83_21#_c_46_n N_VGND_c_266_n 0.00571722f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_83_21#_c_49_n N_A_302_47#_c_305_n 0.00862159f $X=1.205 $Y=0.715 $X2=0
+ $Y2=0
cc_97 N_A_83_21#_c_54_n N_A_302_47#_c_305_n 0.00647563f $X=1.645 $Y=1.69 $X2=0
+ $Y2=0
cc_98 N_B1_c_108_n N_A2_c_136_n 0.02069f $X=1.435 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_99 N_B1_c_107_n N_A2_c_137_n 0.0450221f $X=1.34 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B1_c_109_n N_A2_c_137_n 9.48492e-19 $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_101 N_B1_c_109_n N_A2_c_138_n 0.00110461f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B1_c_107_n N_A2_c_139_n 6.43496e-19 $X=1.34 $Y=1.41 $X2=0 $Y2=0
cc_103 N_B1_c_109_n N_A2_c_139_n 0.0175102f $X=1.375 $Y=1.16 $X2=0 $Y2=0
cc_104 N_B1_c_107_n N_VPWR_c_222_n 0.0130774f $X=1.34 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B1_c_107_n N_VPWR_c_224_n 0.00642146f $X=1.34 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B1_c_107_n N_VPWR_c_221_n 0.0109755f $X=1.34 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B1_c_108_n N_VGND_c_261_n 0.00192994f $X=1.435 $Y=0.995 $X2=0 $Y2=0
cc_108 N_B1_c_108_n N_VGND_c_263_n 0.00547957f $X=1.435 $Y=0.995 $X2=0 $Y2=0
cc_109 N_B1_c_108_n N_VGND_c_265_n 0.0111934f $X=1.435 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A2_c_136_n N_A1_c_176_n 0.0209659f $X=1.855 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A2_c_137_n N_A1_c_177_n 0.066552f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A2_c_138_n N_A1_c_177_n 0.0124531f $X=2.07 $Y=1.275 $X2=0 $Y2=0
cc_113 N_A2_c_139_n N_A1_c_177_n 0.00132453f $X=2.07 $Y=1.175 $X2=0 $Y2=0
cc_114 N_A2_c_137_n N_A1_c_178_n 2.26415e-19 $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A2_c_138_n N_A1_c_178_n 0.0255193f $X=2.07 $Y=1.275 $X2=0 $Y2=0
cc_116 N_A2_c_139_n N_A1_c_178_n 0.0161492f $X=2.07 $Y=1.175 $X2=0 $Y2=0
cc_117 N_A2_c_137_n N_VPWR_c_222_n 9.47269e-19 $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A2_c_137_n N_VPWR_c_224_n 0.00673617f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A2_c_138_n N_VPWR_c_224_n 0.00706536f $X=2.07 $Y=1.275 $X2=0 $Y2=0
cc_120 N_A2_c_137_n N_VPWR_c_226_n 0.00159846f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A2_c_138_n N_VPWR_c_226_n 0.0302455f $X=2.07 $Y=1.275 $X2=0 $Y2=0
cc_122 N_A2_c_137_n N_VPWR_c_221_n 0.0122525f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A2_c_138_n N_VPWR_c_221_n 0.00629072f $X=2.07 $Y=1.275 $X2=0 $Y2=0
cc_124 N_A2_c_138_n A_394_297# 0.0163643f $X=2.07 $Y=1.275 $X2=-0.19 $Y2=-0.24
cc_125 N_A2_c_136_n N_VGND_c_262_n 0.00277568f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A2_c_136_n N_VGND_c_263_n 0.00436487f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A2_c_136_n N_VGND_c_265_n 0.00610249f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A2_c_136_n N_A_302_47#_c_303_n 0.0110016f $X=1.855 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A2_c_137_n N_A_302_47#_c_303_n 0.00314948f $X=1.88 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A2_c_139_n N_A_302_47#_c_303_n 0.0283717f $X=2.07 $Y=1.175 $X2=0 $Y2=0
cc_131 N_A2_c_136_n N_A_302_47#_c_304_n 5.71745e-19 $X=1.855 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_A2_c_139_n N_A_302_47#_c_305_n 0.00315792f $X=2.07 $Y=1.175 $X2=0 $Y2=0
cc_133 N_A1_c_178_n N_VPWR_M1006_d 0.00798567f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A1_c_177_n N_VPWR_c_224_n 0.00427505f $X=2.36 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A1_c_177_n N_VPWR_c_226_n 0.019039f $X=2.36 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A1_c_178_n N_VPWR_c_226_n 0.0133678f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A1_c_177_n N_VPWR_c_221_n 0.00740991f $X=2.36 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A1_c_176_n N_VGND_c_262_n 0.00373921f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A1_c_176_n N_VGND_c_264_n 0.00422241f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A1_c_176_n N_VGND_c_265_n 0.0073132f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A1_c_176_n N_A_302_47#_c_303_n 0.0125771f $X=2.335 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A1_c_177_n N_A_302_47#_c_303_n 0.00573167f $X=2.36 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A1_c_178_n N_A_302_47#_c_303_n 0.0298014f $X=2.49 $Y=1.16 $X2=0 $Y2=0
cc_144 N_A1_c_176_n N_A_302_47#_c_304_n 0.00697687f $X=2.335 $Y=0.995 $X2=0
+ $Y2=0
cc_145 N_X_c_203_n N_VPWR_c_222_n 0.0490385f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_146 N_X_c_203_n N_VPWR_c_223_n 0.0196165f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_147 N_X_M1000_s N_VPWR_c_221_n 0.00442207f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_148 N_X_c_203_n N_VPWR_c_221_n 0.0107063f $X=0.28 $Y=1.62 $X2=0 $Y2=0
cc_149 N_X_M1002_s N_VGND_c_265_n 0.00225715f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_150 N_X_c_201_n N_VGND_c_265_n 0.0129034f $X=0.26 $Y=0.395 $X2=0 $Y2=0
cc_151 N_X_c_201_n N_VGND_c_266_n 0.0217979f $X=0.26 $Y=0.395 $X2=0 $Y2=0
cc_152 N_VPWR_c_221_n A_394_297# 0.00696385f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_153 N_VGND_c_265_n N_A_302_47#_M1003_d 0.00435306f $X=2.99 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_154 N_VGND_c_265_n N_A_302_47#_M1007_d 0.00209319f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_155 N_VGND_M1004_d N_A_302_47#_c_303_n 0.00269535f $X=1.93 $Y=0.235 $X2=0
+ $Y2=0
cc_156 N_VGND_c_262_n N_A_302_47#_c_303_n 0.0127393f $X=2.065 $Y=0.38 $X2=0
+ $Y2=0
cc_157 N_VGND_c_263_n N_A_302_47#_c_303_n 0.00257016f $X=1.98 $Y=0 $X2=0 $Y2=0
cc_158 N_VGND_c_264_n N_A_302_47#_c_303_n 0.00288236f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_159 N_VGND_c_265_n N_A_302_47#_c_303_n 0.0111492f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_160 N_VGND_c_262_n N_A_302_47#_c_304_n 0.0169696f $X=2.065 $Y=0.38 $X2=0
+ $Y2=0
cc_161 N_VGND_c_264_n N_A_302_47#_c_304_n 0.0209752f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_162 N_VGND_c_265_n N_A_302_47#_c_304_n 0.0124119f $X=2.99 $Y=0 $X2=0 $Y2=0
cc_163 N_VGND_c_263_n N_A_302_47#_c_305_n 0.00408973f $X=1.98 $Y=0 $X2=0 $Y2=0
cc_164 N_VGND_c_265_n N_A_302_47#_c_305_n 0.00644927f $X=2.99 $Y=0 $X2=0 $Y2=0
