* File: sky130_fd_sc_hdll__xor3_4.pxi.spice
* Created: Wed Sep  2 08:55:00 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_80_207# N_A_80_207#_M1005_d N_A_80_207#_M1007_d
+ N_A_80_207#_c_177_n N_A_80_207#_M1002_g N_A_80_207#_c_188_n
+ N_A_80_207#_M1000_g N_A_80_207#_c_178_n N_A_80_207#_M1016_g
+ N_A_80_207#_c_189_n N_A_80_207#_M1011_g N_A_80_207#_c_179_n
+ N_A_80_207#_M1017_g N_A_80_207#_c_190_n N_A_80_207#_M1012_g
+ N_A_80_207#_c_180_n N_A_80_207#_M1025_g N_A_80_207#_c_191_n
+ N_A_80_207#_M1019_g N_A_80_207#_c_181_n N_A_80_207#_c_192_n
+ N_A_80_207#_c_203_p N_A_80_207#_c_230_p N_A_80_207#_c_182_n
+ N_A_80_207#_c_183_n N_A_80_207#_c_193_n N_A_80_207#_c_194_n
+ N_A_80_207#_c_195_n N_A_80_207#_c_184_n N_A_80_207#_c_185_n
+ N_A_80_207#_c_212_p N_A_80_207#_c_186_n N_A_80_207#_c_187_n
+ PM_SKY130_FD_SC_HDLL__XOR3_4%A_80_207#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%C N_C_c_324_n N_C_M1020_g N_C_c_325_n N_C_M1023_g
+ N_C_c_326_n N_C_c_327_n N_C_M1007_g N_C_c_328_n N_C_M1005_g C N_C_c_329_n C
+ PM_SKY130_FD_SC_HDLL__XOR3_4%C
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_528_297# N_A_528_297#_M1023_d
+ N_A_528_297#_M1020_d N_A_528_297#_c_387_n N_A_528_297#_M1001_g
+ N_A_528_297#_c_388_n N_A_528_297#_M1013_g N_A_528_297#_c_400_n
+ N_A_528_297#_c_389_n N_A_528_297#_c_393_n N_A_528_297#_c_394_n
+ N_A_528_297#_c_390_n PM_SKY130_FD_SC_HDLL__XOR3_4%A_528_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_1109_297# N_A_1109_297#_M1004_d
+ N_A_1109_297#_M1022_d N_A_1109_297#_c_472_n N_A_1109_297#_M1014_g
+ N_A_1109_297#_M1021_g N_A_1109_297#_c_459_n N_A_1109_297#_c_460_n
+ N_A_1109_297#_c_474_n N_A_1109_297#_M1006_g N_A_1109_297#_c_461_n
+ N_A_1109_297#_M1027_g N_A_1109_297#_c_462_n N_A_1109_297#_c_463_n
+ N_A_1109_297#_c_477_n N_A_1109_297#_c_464_n N_A_1109_297#_c_465_n
+ N_A_1109_297#_c_481_p N_A_1109_297#_c_466_n N_A_1109_297#_c_467_n
+ N_A_1109_297#_c_468_n N_A_1109_297#_c_469_n N_A_1109_297#_c_470_n
+ N_A_1109_297#_c_471_n PM_SKY130_FD_SC_HDLL__XOR3_4%A_1109_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%B N_B_c_644_n N_B_M1022_g N_B_M1004_g N_B_c_637_n
+ N_B_c_638_n N_B_M1018_g N_B_M1003_g N_B_c_647_n N_B_c_648_n N_B_M1026_g
+ N_B_c_649_n N_B_c_650_n N_B_M1008_g N_B_c_640_n B N_B_c_641_n N_B_c_642_n
+ N_B_c_643_n B PM_SKY130_FD_SC_HDLL__XOR3_4%B
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A N_A_c_765_n N_A_M1009_g N_A_c_766_n N_A_M1015_g
+ A PM_SKY130_FD_SC_HDLL__XOR3_4%A
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_1225_365# N_A_1225_365#_M1003_s
+ N_A_1225_365#_M1027_d N_A_1225_365#_M1018_s N_A_1225_365#_M1006_d
+ N_A_1225_365#_c_802_n N_A_1225_365#_M1010_g N_A_1225_365#_c_803_n
+ N_A_1225_365#_M1024_g N_A_1225_365#_c_804_n N_A_1225_365#_c_812_n
+ N_A_1225_365#_c_805_n N_A_1225_365#_c_806_n N_A_1225_365#_c_807_n
+ N_A_1225_365#_c_813_n N_A_1225_365#_c_823_n N_A_1225_365#_c_808_n
+ N_A_1225_365#_c_809_n N_A_1225_365#_c_836_n N_A_1225_365#_c_837_n
+ PM_SKY130_FD_SC_HDLL__XOR3_4%A_1225_365#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%VPWR N_VPWR_M1000_d N_VPWR_M1011_d N_VPWR_M1019_d
+ N_VPWR_M1022_s N_VPWR_M1009_d N_VPWR_c_932_n N_VPWR_c_933_n N_VPWR_c_934_n
+ N_VPWR_c_935_n N_VPWR_c_936_n N_VPWR_c_937_n N_VPWR_c_938_n N_VPWR_c_939_n
+ N_VPWR_c_940_n N_VPWR_c_941_n N_VPWR_c_942_n N_VPWR_c_943_n VPWR
+ N_VPWR_c_944_n N_VPWR_c_945_n N_VPWR_c_931_n N_VPWR_c_947_n N_VPWR_c_948_n
+ N_VPWR_X31_noxref_CONDUCTOR VPWR PM_SKY130_FD_SC_HDLL__XOR3_4%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR3_4%X N_X_M1002_s N_X_M1017_s N_X_M1000_s N_X_M1012_s
+ N_X_c_1061_n N_X_c_1091_n N_X_c_1055_n N_X_c_1056_n N_X_c_1057_n N_X_c_1075_n
+ N_X_c_1095_n N_X_c_1058_n X X N_X_c_1060_n PM_SKY130_FD_SC_HDLL__XOR3_4%X
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_652_325# N_A_652_325#_M1013_d
+ N_A_652_325#_M1026_d N_A_652_325#_M1007_s N_A_652_325#_M1018_d
+ N_A_652_325#_c_1121_n N_A_652_325#_c_1141_n N_A_652_325#_c_1119_n
+ N_A_652_325#_c_1123_n N_A_652_325#_c_1159_n N_A_652_325#_c_1124_n
+ N_A_652_325#_c_1120_n N_A_652_325#_c_1252_p N_A_652_325#_c_1172_n
+ N_A_652_325#_c_1173_n N_A_652_325#_c_1193_n N_A_652_325#_c_1126_n
+ N_A_652_325#_c_1127_n N_A_652_325#_c_1128_n N_A_652_325#_c_1129_n
+ PM_SKY130_FD_SC_HDLL__XOR3_4%A_652_325#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_658_49# N_A_658_49#_M1005_s N_A_658_49#_M1003_d
+ N_A_658_49#_M1001_d N_A_658_49#_M1008_d N_A_658_49#_c_1266_n
+ N_A_658_49#_c_1290_n N_A_658_49#_c_1267_n N_A_658_49#_c_1291_n
+ N_A_658_49#_c_1273_n N_A_658_49#_c_1274_n N_A_658_49#_c_1275_n
+ N_A_658_49#_c_1268_n N_A_658_49#_c_1269_n N_A_658_49#_c_1277_n
+ N_A_658_49#_c_1278_n N_A_658_49#_c_1279_n N_A_658_49#_c_1280_n
+ N_A_658_49#_c_1270_n N_A_658_49#_c_1282_n N_A_658_49#_c_1327_n
+ N_A_658_49#_c_1283_n N_A_658_49#_c_1271_n N_A_658_49#_c_1284_n
+ N_A_658_49#_c_1272_n N_A_658_49#_c_1285_n
+ PM_SKY130_FD_SC_HDLL__XOR3_4%A_658_49#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%A_1510_297# N_A_1510_297#_M1021_d
+ N_A_1510_297#_M1024_d N_A_1510_297#_M1014_d N_A_1510_297#_M1010_d
+ N_A_1510_297#_c_1451_n N_A_1510_297#_c_1463_n N_A_1510_297#_c_1455_n
+ N_A_1510_297#_c_1452_n N_A_1510_297#_c_1464_n N_A_1510_297#_c_1457_n
+ N_A_1510_297#_c_1453_n PM_SKY130_FD_SC_HDLL__XOR3_4%A_1510_297#
x_PM_SKY130_FD_SC_HDLL__XOR3_4%VGND N_VGND_M1002_d N_VGND_M1016_d N_VGND_M1025_d
+ N_VGND_M1004_s N_VGND_M1015_d N_VGND_c_1515_n N_VGND_c_1516_n N_VGND_c_1517_n
+ N_VGND_c_1518_n N_VGND_c_1519_n N_VGND_c_1520_n N_VGND_c_1521_n
+ N_VGND_c_1522_n N_VGND_c_1523_n N_VGND_c_1524_n VGND N_VGND_c_1525_n
+ N_VGND_c_1526_n N_VGND_c_1527_n N_VGND_c_1528_n N_VGND_c_1529_n VGND
+ PM_SKY130_FD_SC_HDLL__XOR3_4%VGND
cc_1 VNB N_A_80_207#_c_177_n 0.0224465f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_80_207#_c_178_n 0.0160466f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A_80_207#_c_179_n 0.015981f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_4 VNB N_A_80_207#_c_180_n 0.0202761f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_A_80_207#_c_181_n 0.00125562f $X=-0.19 $Y=-0.24 $X2=2.105 $Y2=1.16
cc_6 VNB N_A_80_207#_c_182_n 3.43171e-19 $X=-0.19 $Y=-0.24 $X2=2.48 $Y2=0.695
cc_7 VNB N_A_80_207#_c_183_n 7.26786e-19 $X=-0.19 $Y=-0.24 $X2=2.565 $Y2=0.34
cc_8 VNB N_A_80_207#_c_184_n 0.00433686f $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=0.865
cc_9 VNB N_A_80_207#_c_185_n 8.6207e-19 $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=1.325
cc_10 VNB N_A_80_207#_c_186_n 0.0148792f $X=-0.19 $Y=-0.24 $X2=3.66 $Y2=0.355
cc_11 VNB N_A_80_207#_c_187_n 0.100463f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.202
cc_12 VNB N_C_c_324_n 0.0186017f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.245
cc_13 VNB N_C_c_325_n 0.0209904f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_C_c_326_n 0.0450449f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_15 VNB N_C_c_327_n 0.012954f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.41
cc_16 VNB N_C_c_328_n 0.0220325f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_17 VNB N_C_c_329_n 0.00241009f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.41
cc_18 VNB N_A_528_297#_c_387_n 0.0277403f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_19 VNB N_A_528_297#_c_388_n 0.021936f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.41
cc_20 VNB N_A_528_297#_c_389_n 0.00256019f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_21 VNB N_A_528_297#_c_390_n 0.00598209f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_22 VNB N_A_1109_297#_M1021_g 0.0360507f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.985
cc_23 VNB N_A_1109_297#_c_459_n 0.029369f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_24 VNB N_A_1109_297#_c_460_n 0.001407f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_25 VNB N_A_1109_297#_c_461_n 0.0195477f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_26 VNB N_A_1109_297#_c_462_n 0.0291443f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.41
cc_27 VNB N_A_1109_297#_c_463_n 0.0176862f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.985
cc_28 VNB N_A_1109_297#_c_464_n 0.00230039f $X=-0.19 $Y=-0.24 $X2=2.105 $Y2=1.16
cc_29 VNB N_A_1109_297#_c_465_n 0.00817223f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.875
cc_30 VNB N_A_1109_297#_c_466_n 0.0128206f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=1.96
cc_31 VNB N_A_1109_297#_c_467_n 0.00133954f $X=-0.19 $Y=-0.24 $X2=2.48 $Y2=0.425
cc_32 VNB N_A_1109_297#_c_468_n 0.00303586f $X=-0.19 $Y=-0.24 $X2=3.9 $Y2=2.32
cc_33 VNB N_A_1109_297#_c_469_n 0.00230082f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_1109_297#_c_470_n 0.00779728f $X=-0.19 $Y=-0.24 $X2=2.132
+ $Y2=0.865
cc_35 VNB N_A_1109_297#_c_471_n 0.00253923f $X=-0.19 $Y=-0.24 $X2=0.595
+ $Y2=1.202
cc_36 VNB N_B_M1004_g 0.0302599f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_B_c_637_n 0.056013f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_38 VNB N_B_c_638_n 0.0314614f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_39 VNB N_B_M1003_g 0.0287687f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.41
cc_40 VNB N_B_c_640_n 0.0103656f $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=1.077
cc_41 VNB N_B_c_641_n 0.0298429f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.875
cc_42 VNB N_B_c_642_n 0.00130221f $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=1.96
cc_43 VNB N_B_c_643_n 0.021241f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=1.96
cc_44 VNB N_A_c_765_n 0.0230531f $X=-0.19 $Y=-0.24 $X2=3.76 $Y2=0.245
cc_45 VNB N_A_c_766_n 0.0185643f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB A 0.00406657f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_47 VNB N_A_1225_365#_c_802_n 0.0262706f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_48 VNB N_A_1225_365#_c_803_n 0.0201779f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.41
cc_49 VNB N_A_1225_365#_c_804_n 0.0064095f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_50 VNB N_A_1225_365#_c_805_n 0.00275527f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_51 VNB N_A_1225_365#_c_806_n 0.0020163f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.41
cc_52 VNB N_A_1225_365#_c_807_n 0.00310506f $X=-0.19 $Y=-0.24 $X2=2.005
+ $Y2=1.985
cc_53 VNB N_A_1225_365#_c_808_n 0.0020298f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.875
cc_54 VNB N_A_1225_365#_c_809_n 0.00505355f $X=-0.19 $Y=-0.24 $X2=2.48 $Y2=0.425
cc_55 VNB N_VPWR_c_931_n 0.440529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_X_c_1055_n 0.00274486f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_57 VNB N_X_c_1056_n 0.00326222f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.41
cc_58 VNB N_X_c_1057_n 0.00136406f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.985
cc_59 VNB N_X_c_1058_n 0.00198529f $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=1.16
cc_60 VNB N_A_652_325#_c_1119_n 0.00944527f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_61 VNB N_A_652_325#_c_1120_n 0.0097913f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.985
cc_62 VNB N_A_658_49#_c_1266_n 0.00251794f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_63 VNB N_A_658_49#_c_1267_n 0.00850511f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.995
cc_64 VNB N_A_658_49#_c_1268_n 0.013524f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_65 VNB N_A_658_49#_c_1269_n 0.0025441f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.41
cc_66 VNB N_A_658_49#_c_1270_n 0.0023252f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.325
cc_67 VNB N_A_658_49#_c_1271_n 0.0108826f $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=0.865
cc_68 VNB N_A_658_49#_c_1272_n 3.39774e-19 $X=-0.19 $Y=-0.24 $X2=3.895 $Y2=0.355
cc_69 VNB N_A_1510_297#_c_1451_n 0.00788636f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_70 VNB N_A_1510_297#_c_1452_n 0.0308726f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_71 VNB N_A_1510_297#_c_1453_n 0.0129899f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.325
cc_72 VNB N_VGND_c_1515_n 0.0110259f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.41
cc_73 VNB N_VGND_c_1516_n 0.00418552f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.985
cc_74 VNB N_VGND_c_1517_n 0.0196683f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_75 VNB N_VGND_c_1518_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.985
cc_76 VNB N_VGND_c_1519_n 0.00647657f $X=-0.19 $Y=-0.24 $X2=2.005 $Y2=1.41
cc_77 VNB N_VGND_c_1520_n 0.00474148f $X=-0.19 $Y=-0.24 $X2=2.132 $Y2=1.213
cc_78 VNB N_VGND_c_1521_n 0.071988f $X=-0.19 $Y=-0.24 $X2=2.105 $Y2=1.16
cc_79 VNB N_VGND_c_1522_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=2.16 $Y2=1.325
cc_80 VNB N_VGND_c_1523_n 0.110135f $X=-0.19 $Y=-0.24 $X2=2.575 $Y2=1.96
cc_81 VNB N_VGND_c_1524_n 0.00324324f $X=-0.19 $Y=-0.24 $X2=2.245 $Y2=1.96
cc_82 VNB N_VGND_c_1525_n 0.0172377f $X=-0.19 $Y=-0.24 $X2=3.66 $Y2=0.34
cc_83 VNB N_VGND_c_1526_n 0.0220539f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.202
cc_84 VNB N_VGND_c_1527_n 0.5261f $X=-0.19 $Y=-0.24 $X2=1.535 $Y2=1.202
cc_85 VNB N_VGND_c_1528_n 0.00850314f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1529_n 0.00324214f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VPB N_A_80_207#_c_188_n 0.0210716f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.41
cc_88 VPB N_A_80_207#_c_189_n 0.0156597f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.41
cc_89 VPB N_A_80_207#_c_190_n 0.0155948f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.41
cc_90 VPB N_A_80_207#_c_191_n 0.0178805f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.41
cc_91 VPB N_A_80_207#_c_192_n 0.00148444f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=1.875
cc_92 VPB N_A_80_207#_c_193_n 0.0038652f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=2.235
cc_93 VPB N_A_80_207#_c_194_n 0.00116793f $X=-0.19 $Y=1.305 $X2=2.795 $Y2=2.32
cc_94 VPB N_A_80_207#_c_195_n 0.012572f $X=-0.19 $Y=1.305 $X2=3.9 $Y2=2.32
cc_95 VPB N_A_80_207#_c_187_n 0.061607f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.202
cc_96 VPB N_C_c_324_n 0.00946979f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=0.245
cc_97 VPB N_C_M1020_g 0.0311106f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_C_c_326_n 0.0216091f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_99 VPB N_C_c_327_n 0.0395735f $X=-0.19 $Y=1.305 $X2=0.595 $Y2=1.41
cc_100 VPB N_C_c_329_n 6.20239e-19 $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.41
cc_101 VPB N_A_528_297#_c_387_n 0.0399788f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_102 VPB N_A_528_297#_c_389_n 0.00361092f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_103 VPB N_A_528_297#_c_393_n 0.016535f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.985
cc_104 VPB N_A_528_297#_c_394_n 0.00230347f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_105 VPB N_A_528_297#_c_390_n 9.95022e-19 $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_106 VPB N_A_1109_297#_c_472_n 0.0204718f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_107 VPB N_A_1109_297#_c_460_n 0.0105904f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_108 VPB N_A_1109_297#_c_474_n 0.0249586f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.41
cc_109 VPB N_A_1109_297#_c_462_n 0.0105826f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.41
cc_110 VPB N_A_1109_297#_c_463_n 0.00766821f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_111 VPB N_A_1109_297#_c_477_n 0.00590189f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_112 VPB N_A_1109_297#_c_471_n 0.0032041f $X=-0.19 $Y=1.305 $X2=0.595
+ $Y2=1.202
cc_113 VPB N_B_c_644_n 0.0216572f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=0.245
cc_114 VPB N_B_c_638_n 0.00747973f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_115 VPB N_B_M1018_g 0.0155307f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_116 VPB N_B_c_647_n 0.12486f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.985
cc_117 VPB N_B_c_648_n 0.0170126f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.995
cc_118 VPB N_B_c_649_n 0.0101708f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.985
cc_119 VPB N_B_c_650_n 0.00720353f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_120 VPB N_B_M1008_g 0.0131171f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.41
cc_121 VPB N_B_c_640_n 0.0087608f $X=-0.19 $Y=1.305 $X2=2.132 $Y2=1.077
cc_122 VPB B 0.00763142f $X=-0.19 $Y=1.305 $X2=2.132 $Y2=1.16
cc_123 VPB N_B_c_641_n 0.0052573f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=1.875
cc_124 VPB N_B_c_642_n 0.00107001f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.96
cc_125 VPB N_A_c_765_n 0.0278895f $X=-0.19 $Y=1.305 $X2=3.76 $Y2=0.245
cc_126 VPB A 0.00142645f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_127 VPB N_A_1225_365#_c_802_n 0.0294091f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_128 VPB N_A_1225_365#_c_804_n 0.00277419f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_129 VPB N_A_1225_365#_c_812_n 0.00214671f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_130 VPB N_A_1225_365#_c_813_n 0.00156472f $X=-0.19 $Y=1.305 $X2=2.005
+ $Y2=1.985
cc_131 VPB N_VPWR_c_932_n 0.00474148f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.985
cc_132 VPB N_VPWR_c_933_n 0.0185674f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_133 VPB N_VPWR_c_934_n 4.12476e-19 $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.985
cc_134 VPB N_VPWR_c_935_n 0.00711287f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.41
cc_135 VPB N_VPWR_c_936_n 0.00804433f $X=-0.19 $Y=1.305 $X2=2.132 $Y2=1.213
cc_136 VPB N_VPWR_c_937_n 0.00285927f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=1.325
cc_137 VPB N_VPWR_c_938_n 0.0108943f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.96
cc_138 VPB N_VPWR_c_939_n 0.00324376f $X=-0.19 $Y=1.305 $X2=2.245 $Y2=1.96
cc_139 VPB N_VPWR_c_940_n 0.0149748f $X=-0.19 $Y=1.305 $X2=2.48 $Y2=0.695
cc_140 VPB N_VPWR_c_941_n 0.00513322f $X=-0.19 $Y=1.305 $X2=3.66 $Y2=0.34
cc_141 VPB N_VPWR_c_942_n 0.0995635f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=2.045
cc_142 VPB N_VPWR_c_943_n 0.00512961f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=2.235
cc_143 VPB N_VPWR_c_944_n 0.0646337f $X=-0.19 $Y=1.305 $X2=3.66 $Y2=0.355
cc_144 VPB N_VPWR_c_945_n 0.0178464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_931_n 0.0795543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_947_n 0.0043639f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_948_n 0.00513206f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_X_c_1057_n 0.00113396f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.985
cc_149 VPB N_X_c_1060_n 0.00503395f $X=-0.19 $Y=1.305 $X2=2.685 $Y2=2.045
cc_150 VPB N_A_652_325#_c_1121_n 0.004249f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_151 VPB N_A_652_325#_c_1119_n 0.00162471f $X=-0.19 $Y=1.305 $X2=1.46 $Y2=0.56
cc_152 VPB N_A_652_325#_c_1123_n 0.00269586f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_153 VPB N_A_652_325#_c_1124_n 8.54813e-19 $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_154 VPB N_A_652_325#_c_1120_n 0.0021572f $X=-0.19 $Y=1.305 $X2=2.005
+ $Y2=1.985
cc_155 VPB N_A_652_325#_c_1126_n 0.0149543f $X=-0.19 $Y=1.305 $X2=2.575 $Y2=1.96
cc_156 VPB N_A_652_325#_c_1127_n 0.00318498f $X=-0.19 $Y=1.305 $X2=2.245
+ $Y2=1.96
cc_157 VPB N_A_652_325#_c_1128_n 0.00154035f $X=-0.19 $Y=1.305 $X2=2.685
+ $Y2=2.235
cc_158 VPB N_A_652_325#_c_1129_n 0.0207022f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_658_49#_c_1273_n 0.0026444f $X=-0.19 $Y=1.305 $X2=1.535 $Y2=1.41
cc_160 VPB N_A_658_49#_c_1274_n 0.00579762f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_161 VPB N_A_658_49#_c_1275_n 8.62166e-19 $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_162 VPB N_A_658_49#_c_1269_n 0.00847729f $X=-0.19 $Y=1.305 $X2=2.005 $Y2=1.41
cc_163 VPB N_A_658_49#_c_1277_n 0.00306425f $X=-0.19 $Y=1.305 $X2=2.005
+ $Y2=1.985
cc_164 VPB N_A_658_49#_c_1278_n 0.00301837f $X=-0.19 $Y=1.305 $X2=2.132
+ $Y2=1.213
cc_165 VPB N_A_658_49#_c_1279_n 0.0104899f $X=-0.19 $Y=1.305 $X2=2.132 $Y2=1.16
cc_166 VPB N_A_658_49#_c_1280_n 0.00185607f $X=-0.19 $Y=1.305 $X2=2.105 $Y2=1.16
cc_167 VPB N_A_658_49#_c_1270_n 0.00156022f $X=-0.19 $Y=1.305 $X2=2.16 $Y2=1.325
cc_168 VPB N_A_658_49#_c_1282_n 0.024688f $X=-0.19 $Y=1.305 $X2=2.245 $Y2=1.96
cc_169 VPB N_A_658_49#_c_1283_n 0.00221665f $X=-0.19 $Y=1.305 $X2=3.9 $Y2=2.32
cc_170 VPB N_A_658_49#_c_1284_n 2.86933e-19 $X=-0.19 $Y=1.305 $X2=2.132
+ $Y2=1.325
cc_171 VPB N_A_658_49#_c_1285_n 2.28173e-19 $X=-0.19 $Y=1.305 $X2=3.66 $Y2=0.355
cc_172 VPB N_A_1510_297#_c_1451_n 0.00468519f $X=-0.19 $Y=1.305 $X2=0.99
+ $Y2=0.56
cc_173 VPB N_A_1510_297#_c_1455_n 0.0141756f $X=-0.19 $Y=1.305 $X2=1.535
+ $Y2=1.985
cc_174 VPB N_A_1510_297#_c_1452_n 0.0227839f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_175 VPB N_A_1510_297#_c_1457_n 0.00990626f $X=-0.19 $Y=1.305 $X2=2.132
+ $Y2=1.077
cc_176 N_A_80_207#_c_181_n N_C_c_324_n 0.00316117f $X=2.105 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_177 N_A_80_207#_c_184_n N_C_c_324_n 0.00567528f $X=2.132 $Y=0.865 $X2=-0.19
+ $Y2=-0.24
cc_178 N_A_80_207#_c_186_n N_C_c_324_n 6.72752e-19 $X=3.66 $Y=0.355 $X2=-0.19
+ $Y2=-0.24
cc_179 N_A_80_207#_c_187_n N_C_c_324_n 0.024764f $X=2.005 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_180 N_A_80_207#_c_191_n N_C_M1020_g 0.022858f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_80_207#_c_192_n N_C_M1020_g 0.00597276f $X=2.16 $Y=1.875 $X2=0 $Y2=0
cc_182 N_A_80_207#_c_203_p N_C_M1020_g 0.016545f $X=2.575 $Y=1.96 $X2=0 $Y2=0
cc_183 N_A_80_207#_c_193_n N_C_M1020_g 0.0073266f $X=2.685 $Y=2.235 $X2=0 $Y2=0
cc_184 N_A_80_207#_c_194_n N_C_M1020_g 0.00730512f $X=2.795 $Y=2.32 $X2=0 $Y2=0
cc_185 N_A_80_207#_c_180_n N_C_c_325_n 0.00651061f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_186 N_A_80_207#_c_182_n N_C_c_325_n 0.00299032f $X=2.48 $Y=0.695 $X2=0 $Y2=0
cc_187 N_A_80_207#_c_184_n N_C_c_325_n 0.00117465f $X=2.132 $Y=0.865 $X2=0 $Y2=0
cc_188 N_A_80_207#_c_186_n N_C_c_325_n 0.01362f $X=3.66 $Y=0.355 $X2=0 $Y2=0
cc_189 N_A_80_207#_c_186_n N_C_c_326_n 0.00684077f $X=3.66 $Y=0.355 $X2=0 $Y2=0
cc_190 N_A_80_207#_c_195_n N_C_c_327_n 0.0112964f $X=3.9 $Y=2.32 $X2=0 $Y2=0
cc_191 N_A_80_207#_c_212_p N_C_c_328_n 0.00537539f $X=3.895 $Y=0.37 $X2=0 $Y2=0
cc_192 N_A_80_207#_c_186_n N_C_c_328_n 0.00603149f $X=3.66 $Y=0.355 $X2=0 $Y2=0
cc_193 N_A_80_207#_c_186_n N_C_c_329_n 0.00331115f $X=3.66 $Y=0.355 $X2=0 $Y2=0
cc_194 N_A_80_207#_c_203_p N_A_528_297#_M1020_d 0.0041981f $X=2.575 $Y=1.96
+ $X2=0 $Y2=0
cc_195 N_A_80_207#_c_193_n N_A_528_297#_M1020_d 0.00267049f $X=2.685 $Y=2.235
+ $X2=0 $Y2=0
cc_196 N_A_80_207#_c_195_n N_A_528_297#_c_387_n 0.00841967f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_197 N_A_80_207#_c_212_p N_A_528_297#_c_388_n 0.00165143f $X=3.895 $Y=0.37
+ $X2=0 $Y2=0
cc_198 N_A_80_207#_c_192_n N_A_528_297#_c_400_n 0.00809417f $X=2.16 $Y=1.875
+ $X2=0 $Y2=0
cc_199 N_A_80_207#_c_203_p N_A_528_297#_c_400_n 0.0130455f $X=2.575 $Y=1.96
+ $X2=0 $Y2=0
cc_200 N_A_80_207#_c_195_n N_A_528_297#_c_400_n 0.00596778f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_201 N_A_80_207#_c_181_n N_A_528_297#_c_389_n 0.0143175f $X=2.105 $Y=1.16
+ $X2=0 $Y2=0
cc_202 N_A_80_207#_c_184_n N_A_528_297#_c_389_n 0.00648081f $X=2.132 $Y=0.865
+ $X2=0 $Y2=0
cc_203 N_A_80_207#_c_186_n N_A_528_297#_c_389_n 0.0127861f $X=3.66 $Y=0.355
+ $X2=0 $Y2=0
cc_204 N_A_80_207#_c_187_n N_A_528_297#_c_389_n 2.69065e-19 $X=2.005 $Y=1.202
+ $X2=0 $Y2=0
cc_205 N_A_80_207#_M1007_d N_A_528_297#_c_393_n 0.00327687f $X=3.71 $Y=1.625
+ $X2=0 $Y2=0
cc_206 N_A_80_207#_c_195_n N_A_528_297#_c_393_n 0.00613544f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_207 N_A_80_207#_c_192_n N_VPWR_M1019_d 0.00460371f $X=2.16 $Y=1.875 $X2=0
+ $Y2=0
cc_208 N_A_80_207#_c_203_p N_VPWR_M1019_d 0.0076537f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_209 N_A_80_207#_c_230_p N_VPWR_M1019_d 9.86211e-19 $X=2.245 $Y=1.96 $X2=0
+ $Y2=0
cc_210 N_A_80_207#_c_188_n N_VPWR_c_932_n 0.00620807f $X=0.595 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_80_207#_c_188_n N_VPWR_c_933_n 0.00702461f $X=0.595 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_80_207#_c_189_n N_VPWR_c_933_n 0.00458723f $X=1.065 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_80_207#_c_188_n N_VPWR_c_934_n 0.0010752f $X=0.595 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_80_207#_c_189_n N_VPWR_c_934_n 0.00831343f $X=1.065 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_80_207#_c_190_n N_VPWR_c_934_n 0.00736445f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_80_207#_c_191_n N_VPWR_c_934_n 5.15829e-19 $X=2.005 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_80_207#_c_190_n N_VPWR_c_935_n 5.15829e-19 $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_80_207#_c_191_n N_VPWR_c_935_n 0.00839108f $X=2.005 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_80_207#_c_203_p N_VPWR_c_935_n 0.0122785f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_220 N_A_80_207#_c_230_p N_VPWR_c_935_n 0.00937215f $X=2.245 $Y=1.96 $X2=0
+ $Y2=0
cc_221 N_A_80_207#_c_193_n N_VPWR_c_935_n 0.00150207f $X=2.685 $Y=2.235 $X2=0
+ $Y2=0
cc_222 N_A_80_207#_c_194_n N_VPWR_c_935_n 0.0142215f $X=2.795 $Y=2.32 $X2=0
+ $Y2=0
cc_223 N_A_80_207#_c_190_n N_VPWR_c_940_n 0.00458723f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_80_207#_c_191_n N_VPWR_c_940_n 0.00622633f $X=2.005 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_80_207#_c_203_p N_VPWR_c_944_n 0.00218776f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_226 N_A_80_207#_c_194_n N_VPWR_c_944_n 0.0109858f $X=2.795 $Y=2.32 $X2=0
+ $Y2=0
cc_227 N_A_80_207#_c_195_n N_VPWR_c_944_n 0.0617415f $X=3.9 $Y=2.32 $X2=0 $Y2=0
cc_228 N_A_80_207#_c_188_n N_VPWR_c_931_n 0.0135015f $X=0.595 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_80_207#_c_189_n N_VPWR_c_931_n 0.00523894f $X=1.065 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_80_207#_c_190_n N_VPWR_c_931_n 0.00523894f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_80_207#_c_191_n N_VPWR_c_931_n 0.0104011f $X=2.005 $Y=1.41 $X2=0
+ $Y2=0
cc_232 N_A_80_207#_c_203_p N_VPWR_c_931_n 0.00523504f $X=2.575 $Y=1.96 $X2=0
+ $Y2=0
cc_233 N_A_80_207#_c_230_p N_VPWR_c_931_n 7.83888e-19 $X=2.245 $Y=1.96 $X2=0
+ $Y2=0
cc_234 N_A_80_207#_c_194_n N_VPWR_c_931_n 0.00809722f $X=2.795 $Y=2.32 $X2=0
+ $Y2=0
cc_235 N_A_80_207#_c_195_n N_VPWR_c_931_n 0.0495864f $X=3.9 $Y=2.32 $X2=0 $Y2=0
cc_236 N_A_80_207#_c_178_n N_X_c_1061_n 0.00398532f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A_80_207#_c_178_n N_X_c_1055_n 0.0152628f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_80_207#_c_187_n N_X_c_1055_n 0.00181533f $X=2.005 $Y=1.202 $X2=0
+ $Y2=0
cc_239 N_A_80_207#_c_177_n N_X_c_1056_n 0.00188945f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_80_207#_c_187_n N_X_c_1056_n 0.00513503f $X=2.005 $Y=1.202 $X2=0
+ $Y2=0
cc_241 N_A_80_207#_c_178_n N_X_c_1057_n 0.0017485f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_80_207#_c_189_n N_X_c_1057_n 8.15909e-19 $X=1.065 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_80_207#_c_179_n N_X_c_1057_n 0.0019079f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A_80_207#_c_190_n N_X_c_1057_n 9.5783e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_245 N_A_80_207#_c_180_n N_X_c_1057_n 5.72848e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_80_207#_c_181_n N_X_c_1057_n 0.00825007f $X=2.105 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A_80_207#_c_192_n N_X_c_1057_n 0.00334517f $X=2.16 $Y=1.875 $X2=0 $Y2=0
cc_248 N_A_80_207#_c_184_n N_X_c_1057_n 0.00546783f $X=2.132 $Y=0.865 $X2=0
+ $Y2=0
cc_249 N_A_80_207#_c_187_n N_X_c_1057_n 0.0486346f $X=2.005 $Y=1.202 $X2=0 $Y2=0
cc_250 N_A_80_207#_c_180_n N_X_c_1075_n 0.00185065f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_251 N_A_80_207#_c_182_n N_X_c_1075_n 0.0035889f $X=2.48 $Y=0.695 $X2=0 $Y2=0
cc_252 N_A_80_207#_c_179_n N_X_c_1058_n 0.0124594f $X=1.46 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A_80_207#_c_180_n N_X_c_1058_n 0.00254012f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A_80_207#_c_182_n N_X_c_1058_n 0.00102903f $X=2.48 $Y=0.695 $X2=0 $Y2=0
cc_255 N_A_80_207#_c_184_n N_X_c_1058_n 0.0125513f $X=2.132 $Y=0.865 $X2=0 $Y2=0
cc_256 N_A_80_207#_c_187_n N_X_c_1058_n 0.0041816f $X=2.005 $Y=1.202 $X2=0 $Y2=0
cc_257 N_A_80_207#_c_188_n N_X_c_1060_n 0.0167037f $X=0.595 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_80_207#_c_189_n N_X_c_1060_n 0.0263799f $X=1.065 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_80_207#_c_190_n N_X_c_1060_n 0.0233053f $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_80_207#_c_191_n N_X_c_1060_n 0.00303371f $X=2.005 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_80_207#_c_192_n N_X_c_1060_n 0.02768f $X=2.16 $Y=1.875 $X2=0 $Y2=0
cc_262 N_A_80_207#_c_230_p N_X_c_1060_n 0.0122124f $X=2.245 $Y=1.96 $X2=0 $Y2=0
cc_263 N_A_80_207#_c_187_n N_X_c_1060_n 0.0181857f $X=2.005 $Y=1.202 $X2=0 $Y2=0
cc_264 N_A_80_207#_c_195_n N_A_652_325#_M1007_s 0.00537509f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_265 N_A_80_207#_M1007_d N_A_652_325#_c_1121_n 0.00649326f $X=3.71 $Y=1.625
+ $X2=0 $Y2=0
cc_266 N_A_80_207#_c_203_p N_A_652_325#_c_1121_n 0.0082675f $X=2.575 $Y=1.96
+ $X2=0 $Y2=0
cc_267 N_A_80_207#_c_193_n N_A_652_325#_c_1121_n 9.46755e-19 $X=2.685 $Y=2.235
+ $X2=0 $Y2=0
cc_268 N_A_80_207#_c_195_n N_A_652_325#_c_1121_n 0.0614522f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_269 N_A_80_207#_c_186_n N_A_658_49#_M1005_s 0.00669207f $X=3.66 $Y=0.355
+ $X2=-0.19 $Y2=-0.24
cc_270 N_A_80_207#_M1005_d N_A_658_49#_c_1266_n 0.0130594f $X=3.76 $Y=0.245
+ $X2=0 $Y2=0
cc_271 N_A_80_207#_c_212_p N_A_658_49#_c_1266_n 0.0203761f $X=3.895 $Y=0.37
+ $X2=0 $Y2=0
cc_272 N_A_80_207#_c_186_n N_A_658_49#_c_1266_n 0.0191047f $X=3.66 $Y=0.355
+ $X2=0 $Y2=0
cc_273 N_A_80_207#_c_212_p N_A_658_49#_c_1290_n 0.002195f $X=3.895 $Y=0.37 $X2=0
+ $Y2=0
cc_274 N_A_80_207#_c_212_p N_A_658_49#_c_1291_n 0.0147713f $X=3.895 $Y=0.37
+ $X2=0 $Y2=0
cc_275 N_A_80_207#_c_195_n N_A_658_49#_c_1283_n 0.0100105f $X=3.9 $Y=2.32 $X2=0
+ $Y2=0
cc_276 N_A_80_207#_c_182_n N_VGND_M1025_d 0.00445136f $X=2.48 $Y=0.695 $X2=0
+ $Y2=0
cc_277 N_A_80_207#_c_183_n N_VGND_M1025_d 0.00243608f $X=2.565 $Y=0.34 $X2=0
+ $Y2=0
cc_278 N_A_80_207#_c_184_n N_VGND_M1025_d 0.0197712f $X=2.132 $Y=0.865 $X2=0
+ $Y2=0
cc_279 N_A_80_207#_c_177_n N_VGND_c_1516_n 0.00453301f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_80_207#_c_179_n N_VGND_c_1517_n 0.00428601f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_80_207#_c_180_n N_VGND_c_1517_n 0.00585385f $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_80_207#_c_180_n N_VGND_c_1518_n 0.00438629f $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_80_207#_c_182_n N_VGND_c_1518_n 0.00722699f $X=2.48 $Y=0.695 $X2=0
+ $Y2=0
cc_284 N_A_80_207#_c_183_n N_VGND_c_1518_n 0.0138309f $X=2.565 $Y=0.34 $X2=0
+ $Y2=0
cc_285 N_A_80_207#_c_184_n N_VGND_c_1518_n 0.0134844f $X=2.132 $Y=0.865 $X2=0
+ $Y2=0
cc_286 N_A_80_207#_c_187_n N_VGND_c_1518_n 7.03336e-19 $X=2.005 $Y=1.202 $X2=0
+ $Y2=0
cc_287 N_A_80_207#_c_183_n N_VGND_c_1521_n 0.0119943f $X=2.565 $Y=0.34 $X2=0
+ $Y2=0
cc_288 N_A_80_207#_c_184_n N_VGND_c_1521_n 0.00264854f $X=2.132 $Y=0.865 $X2=0
+ $Y2=0
cc_289 N_A_80_207#_c_186_n N_VGND_c_1521_n 0.0921862f $X=3.66 $Y=0.355 $X2=0
+ $Y2=0
cc_290 N_A_80_207#_c_177_n N_VGND_c_1525_n 0.00585385f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_80_207#_c_178_n N_VGND_c_1525_n 0.00200081f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_292 N_A_80_207#_c_177_n N_VGND_c_1527_n 0.0118665f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_80_207#_c_178_n N_VGND_c_1527_n 0.00279397f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_80_207#_c_179_n N_VGND_c_1527_n 0.00595274f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_80_207#_c_180_n N_VGND_c_1527_n 0.0120709f $X=1.93 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_80_207#_c_183_n N_VGND_c_1527_n 0.00652842f $X=2.565 $Y=0.34 $X2=0
+ $Y2=0
cc_297 N_A_80_207#_c_184_n N_VGND_c_1527_n 0.00535855f $X=2.132 $Y=0.865 $X2=0
+ $Y2=0
cc_298 N_A_80_207#_c_186_n N_VGND_c_1527_n 0.0550361f $X=3.66 $Y=0.355 $X2=0
+ $Y2=0
cc_299 N_A_80_207#_c_177_n N_VGND_c_1528_n 9.42918e-19 $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_300 N_A_80_207#_c_178_n N_VGND_c_1528_n 0.0107476f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_301 N_A_80_207#_c_179_n N_VGND_c_1528_n 0.00317372f $X=1.46 $Y=0.995 $X2=0
+ $Y2=0
cc_302 N_A_80_207#_c_187_n N_VGND_c_1528_n 4.41839e-19 $X=2.005 $Y=1.202 $X2=0
+ $Y2=0
cc_303 N_C_c_327_n N_A_528_297#_c_387_n 0.0495097f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_304 N_C_c_329_n N_A_528_297#_c_387_n 0.001133f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_305 N_C_c_327_n N_A_528_297#_c_388_n 3.1776e-19 $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_306 N_C_c_328_n N_A_528_297#_c_388_n 0.0194799f $X=3.685 $Y=0.985 $X2=0 $Y2=0
cc_307 N_C_c_324_n N_A_528_297#_c_400_n 0.00477143f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_308 N_C_M1020_g N_A_528_297#_c_400_n 0.00696208f $X=2.55 $Y=1.805 $X2=0 $Y2=0
cc_309 N_C_c_324_n N_A_528_297#_c_389_n 0.00212943f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_310 N_C_M1020_g N_A_528_297#_c_389_n 0.00211239f $X=2.55 $Y=1.805 $X2=0 $Y2=0
cc_311 N_C_c_325_n N_A_528_297#_c_389_n 0.00292931f $X=2.665 $Y=0.995 $X2=0
+ $Y2=0
cc_312 N_C_c_326_n N_A_528_297#_c_389_n 0.0226128f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_313 N_C_c_327_n N_A_528_297#_c_389_n 0.00495404f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_314 N_C_c_328_n N_A_528_297#_c_389_n 0.00292894f $X=3.685 $Y=0.985 $X2=0
+ $Y2=0
cc_315 N_C_c_329_n N_A_528_297#_c_389_n 0.0250009f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_316 N_C_c_326_n N_A_528_297#_c_393_n 0.0145971f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_317 N_C_c_327_n N_A_528_297#_c_393_n 0.0166507f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_318 N_C_c_329_n N_A_528_297#_c_393_n 0.0433481f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_319 N_C_c_327_n N_A_528_297#_c_394_n 0.00411747f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_320 N_C_c_327_n N_A_528_297#_c_390_n 0.0010471f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_321 N_C_c_329_n N_A_528_297#_c_390_n 0.0296672f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_322 N_C_M1020_g N_VPWR_c_935_n 0.00197057f $X=2.55 $Y=1.805 $X2=0 $Y2=0
cc_323 N_C_M1020_g N_VPWR_c_944_n 0.00515602f $X=2.55 $Y=1.805 $X2=0 $Y2=0
cc_324 N_C_c_327_n N_VPWR_c_944_n 0.00427564f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_325 N_C_M1020_g N_VPWR_c_931_n 0.00682402f $X=2.55 $Y=1.805 $X2=0 $Y2=0
cc_326 N_C_c_327_n N_VPWR_c_931_n 0.00728509f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_327 N_C_M1020_g N_A_652_325#_c_1121_n 9.33413e-19 $X=2.55 $Y=1.805 $X2=0
+ $Y2=0
cc_328 N_C_c_327_n N_A_652_325#_c_1121_n 0.0104309f $X=3.62 $Y=1.55 $X2=0 $Y2=0
cc_329 N_C_c_326_n N_A_658_49#_c_1266_n 0.00625753f $X=3.52 $Y=1.16 $X2=0 $Y2=0
cc_330 N_C_c_328_n N_A_658_49#_c_1266_n 0.0094194f $X=3.685 $Y=0.985 $X2=0 $Y2=0
cc_331 N_C_c_329_n N_A_658_49#_c_1266_n 0.0382257f $X=3.58 $Y=1.16 $X2=0 $Y2=0
cc_332 N_C_c_328_n N_A_658_49#_c_1290_n 7.51336e-19 $X=3.685 $Y=0.985 $X2=0
+ $Y2=0
cc_333 N_C_c_325_n N_VGND_c_1518_n 3.76925e-19 $X=2.665 $Y=0.995 $X2=0 $Y2=0
cc_334 N_C_c_325_n N_VGND_c_1521_n 7.74126e-19 $X=2.665 $Y=0.995 $X2=0 $Y2=0
cc_335 N_C_c_328_n N_VGND_c_1521_n 0.00357877f $X=3.685 $Y=0.985 $X2=0 $Y2=0
cc_336 N_C_c_328_n N_VGND_c_1527_n 0.00706369f $X=3.685 $Y=0.985 $X2=0 $Y2=0
cc_337 N_A_528_297#_c_387_n N_VPWR_c_944_n 0.00455111f $X=4.2 $Y=1.55 $X2=0
+ $Y2=0
cc_338 N_A_528_297#_c_387_n N_VPWR_c_931_n 0.00760152f $X=4.2 $Y=1.55 $X2=0
+ $Y2=0
cc_339 N_A_528_297#_c_393_n N_A_652_325#_M1007_s 0.00272894f $X=3.985 $Y=1.62
+ $X2=0 $Y2=0
cc_340 N_A_528_297#_c_387_n N_A_652_325#_c_1121_n 0.017225f $X=4.2 $Y=1.55 $X2=0
+ $Y2=0
cc_341 N_A_528_297#_c_393_n N_A_652_325#_c_1121_n 0.0561298f $X=3.985 $Y=1.62
+ $X2=0 $Y2=0
cc_342 N_A_528_297#_c_390_n N_A_652_325#_c_1121_n 0.00522966f $X=4.175 $Y=1.16
+ $X2=0 $Y2=0
cc_343 N_A_528_297#_c_387_n N_A_652_325#_c_1141_n 0.00748858f $X=4.2 $Y=1.55
+ $X2=0 $Y2=0
cc_344 N_A_528_297#_c_393_n N_A_652_325#_c_1141_n 6.13389e-19 $X=3.985 $Y=1.62
+ $X2=0 $Y2=0
cc_345 N_A_528_297#_c_387_n N_A_652_325#_c_1119_n 0.00294142f $X=4.2 $Y=1.55
+ $X2=0 $Y2=0
cc_346 N_A_528_297#_c_388_n N_A_652_325#_c_1119_n 0.006614f $X=4.285 $Y=0.995
+ $X2=0 $Y2=0
cc_347 N_A_528_297#_c_394_n N_A_652_325#_c_1119_n 0.00166649f $X=4.07 $Y=1.535
+ $X2=0 $Y2=0
cc_348 N_A_528_297#_c_390_n N_A_652_325#_c_1119_n 0.0225705f $X=4.175 $Y=1.16
+ $X2=0 $Y2=0
cc_349 N_A_528_297#_c_393_n N_A_652_325#_c_1127_n 4.56942e-19 $X=3.985 $Y=1.62
+ $X2=0 $Y2=0
cc_350 N_A_528_297#_c_394_n N_A_652_325#_c_1127_n 6.00479e-19 $X=4.07 $Y=1.535
+ $X2=0 $Y2=0
cc_351 N_A_528_297#_c_387_n N_A_652_325#_c_1129_n 0.00700676f $X=4.2 $Y=1.55
+ $X2=0 $Y2=0
cc_352 N_A_528_297#_c_393_n N_A_652_325#_c_1129_n 0.0109044f $X=3.985 $Y=1.62
+ $X2=0 $Y2=0
cc_353 N_A_528_297#_c_394_n N_A_652_325#_c_1129_n 0.00528578f $X=4.07 $Y=1.535
+ $X2=0 $Y2=0
cc_354 N_A_528_297#_c_390_n N_A_652_325#_c_1129_n 0.00232363f $X=4.175 $Y=1.16
+ $X2=0 $Y2=0
cc_355 N_A_528_297#_c_387_n N_A_658_49#_c_1266_n 0.0041059f $X=4.2 $Y=1.55 $X2=0
+ $Y2=0
cc_356 N_A_528_297#_c_388_n N_A_658_49#_c_1266_n 0.0104524f $X=4.285 $Y=0.995
+ $X2=0 $Y2=0
cc_357 N_A_528_297#_c_389_n N_A_658_49#_c_1266_n 0.00976986f $X=2.875 $Y=0.76
+ $X2=0 $Y2=0
cc_358 N_A_528_297#_c_390_n N_A_658_49#_c_1266_n 0.0282776f $X=4.175 $Y=1.16
+ $X2=0 $Y2=0
cc_359 N_A_528_297#_c_388_n N_A_658_49#_c_1290_n 0.00969442f $X=4.285 $Y=0.995
+ $X2=0 $Y2=0
cc_360 N_A_528_297#_c_388_n N_A_658_49#_c_1291_n 0.00814783f $X=4.285 $Y=0.995
+ $X2=0 $Y2=0
cc_361 N_A_528_297#_c_387_n N_A_658_49#_c_1273_n 0.00452598f $X=4.2 $Y=1.55
+ $X2=0 $Y2=0
cc_362 N_A_528_297#_c_387_n N_A_658_49#_c_1275_n 7.6183e-19 $X=4.2 $Y=1.55 $X2=0
+ $Y2=0
cc_363 N_A_528_297#_c_388_n N_A_658_49#_c_1268_n 0.00103799f $X=4.285 $Y=0.995
+ $X2=0 $Y2=0
cc_364 N_A_528_297#_c_387_n N_A_658_49#_c_1283_n 0.00354471f $X=4.2 $Y=1.55
+ $X2=0 $Y2=0
cc_365 N_A_528_297#_c_388_n N_VGND_c_1521_n 0.00367048f $X=4.285 $Y=0.995 $X2=0
+ $Y2=0
cc_366 N_A_528_297#_c_388_n N_VGND_c_1527_n 0.00715174f $X=4.285 $Y=0.995 $X2=0
+ $Y2=0
cc_367 N_A_1109_297#_c_477_n N_B_c_644_n 0.00851867f $X=5.845 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_368 N_A_1109_297#_c_471_n N_B_c_644_n 8.21886e-19 $X=5.905 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_369 N_A_1109_297#_c_481_p N_B_M1004_g 0.00363512f $X=5.985 $Y=0.85 $X2=0
+ $Y2=0
cc_370 N_A_1109_297#_c_471_n N_B_M1004_g 0.0173433f $X=5.905 $Y=0.72 $X2=0 $Y2=0
cc_371 N_A_1109_297#_c_465_n N_B_c_637_n 0.0050801f $X=7.125 $Y=0.85 $X2=0 $Y2=0
cc_372 N_A_1109_297#_c_471_n N_B_c_637_n 0.0122189f $X=5.905 $Y=0.72 $X2=0 $Y2=0
cc_373 N_A_1109_297#_c_477_n N_B_c_638_n 0.00731407f $X=5.845 $Y=1.58 $X2=0
+ $Y2=0
cc_374 N_A_1109_297#_c_471_n N_B_c_638_n 0.00956129f $X=5.905 $Y=0.72 $X2=0
+ $Y2=0
cc_375 N_A_1109_297#_c_472_n N_B_M1018_g 0.0117785f $X=7.46 $Y=1.41 $X2=0 $Y2=0
cc_376 N_A_1109_297#_M1021_g N_B_M1003_g 0.0101671f $X=7.485 $Y=0.455 $X2=0
+ $Y2=0
cc_377 N_A_1109_297#_c_462_n N_B_M1003_g 0.021215f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_378 N_A_1109_297#_c_464_n N_B_M1003_g 0.00182991f $X=7.247 $Y=0.995 $X2=0
+ $Y2=0
cc_379 N_A_1109_297#_c_465_n N_B_M1003_g 0.00123925f $X=7.125 $Y=0.85 $X2=0
+ $Y2=0
cc_380 N_A_1109_297#_c_467_n N_B_M1003_g 6.73467e-19 $X=7.415 $Y=0.85 $X2=0
+ $Y2=0
cc_381 N_A_1109_297#_c_468_n N_B_M1003_g 0.00122412f $X=7.27 $Y=0.85 $X2=0 $Y2=0
cc_382 N_A_1109_297#_c_472_n N_B_c_647_n 0.0105804f $X=7.46 $Y=1.41 $X2=0 $Y2=0
cc_383 N_A_1109_297#_c_474_n N_B_c_647_n 0.00616735f $X=8.95 $Y=1.57 $X2=0 $Y2=0
cc_384 N_A_1109_297#_c_460_n N_B_c_649_n 0.00390956f $X=8.95 $Y=1.47 $X2=0 $Y2=0
cc_385 N_A_1109_297#_c_474_n N_B_c_650_n 0.00390956f $X=8.95 $Y=1.57 $X2=0 $Y2=0
cc_386 N_A_1109_297#_c_474_n N_B_M1008_g 0.0248649f $X=8.95 $Y=1.57 $X2=0 $Y2=0
cc_387 N_A_1109_297#_c_463_n N_B_c_640_n 0.0017886f $X=7.46 $Y=1.202 $X2=0 $Y2=0
cc_388 N_A_1109_297#_c_460_n B 0.00195994f $X=8.95 $Y=1.47 $X2=0 $Y2=0
cc_389 N_A_1109_297#_c_474_n B 4.37948e-19 $X=8.95 $Y=1.57 $X2=0 $Y2=0
cc_390 N_A_1109_297#_c_466_n B 0.00421862f $X=8.605 $Y=0.85 $X2=0 $Y2=0
cc_391 N_A_1109_297#_c_469_n B 0.00123911f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_392 N_A_1109_297#_c_459_n N_B_c_641_n 0.0192205f $X=8.95 $Y=1.28 $X2=0 $Y2=0
cc_393 N_A_1109_297#_c_463_n N_B_c_641_n 0.00774829f $X=7.46 $Y=1.202 $X2=0
+ $Y2=0
cc_394 N_A_1109_297#_c_466_n N_B_c_641_n 0.00133312f $X=8.605 $Y=0.85 $X2=0
+ $Y2=0
cc_395 N_A_1109_297#_c_470_n N_B_c_641_n 0.00172718f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_396 N_A_1109_297#_c_459_n N_B_c_642_n 0.00126991f $X=8.95 $Y=1.28 $X2=0 $Y2=0
cc_397 N_A_1109_297#_c_466_n N_B_c_642_n 0.00715618f $X=8.605 $Y=0.85 $X2=0
+ $Y2=0
cc_398 N_A_1109_297#_c_470_n N_B_c_642_n 0.021521f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_399 N_A_1109_297#_M1021_g N_B_c_643_n 0.00774829f $X=7.485 $Y=0.455 $X2=0
+ $Y2=0
cc_400 N_A_1109_297#_c_459_n N_B_c_643_n 0.00135777f $X=8.95 $Y=1.28 $X2=0 $Y2=0
cc_401 N_A_1109_297#_c_461_n N_B_c_643_n 0.0134808f $X=8.98 $Y=0.945 $X2=0 $Y2=0
cc_402 N_A_1109_297#_c_466_n N_B_c_643_n 0.00736426f $X=8.605 $Y=0.85 $X2=0
+ $Y2=0
cc_403 N_A_1109_297#_c_469_n N_B_c_643_n 0.0014125f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_404 N_A_1109_297#_c_470_n N_B_c_643_n 0.00207369f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_405 N_A_1109_297#_c_459_n N_A_c_765_n 0.0181958f $X=8.95 $Y=1.28 $X2=-0.19
+ $Y2=-0.24
cc_406 N_A_1109_297#_c_460_n N_A_c_765_n 0.0104505f $X=8.95 $Y=1.47 $X2=-0.19
+ $Y2=-0.24
cc_407 N_A_1109_297#_c_474_n N_A_c_765_n 0.031579f $X=8.95 $Y=1.57 $X2=-0.19
+ $Y2=-0.24
cc_408 N_A_1109_297#_c_470_n N_A_c_765_n 6.45074e-19 $X=8.75 $Y=0.85 $X2=-0.19
+ $Y2=-0.24
cc_409 N_A_1109_297#_c_461_n N_A_c_766_n 0.0188728f $X=8.98 $Y=0.945 $X2=0 $Y2=0
cc_410 N_A_1109_297#_c_470_n N_A_c_766_n 2.38541e-19 $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_411 N_A_1109_297#_c_459_n A 0.0015686f $X=8.95 $Y=1.28 $X2=0 $Y2=0
cc_412 N_A_1109_297#_c_460_n A 0.00114147f $X=8.95 $Y=1.47 $X2=0 $Y2=0
cc_413 N_A_1109_297#_c_470_n A 0.0133858f $X=8.75 $Y=0.85 $X2=0 $Y2=0
cc_414 N_A_1109_297#_c_465_n N_A_1225_365#_M1003_s 9.57955e-19 $X=7.125 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_415 N_A_1109_297#_c_477_n N_A_1225_365#_c_804_n 0.0199218f $X=5.845 $Y=1.58
+ $X2=0 $Y2=0
cc_416 N_A_1109_297#_c_465_n N_A_1225_365#_c_804_n 0.0125056f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_417 N_A_1109_297#_c_481_p N_A_1225_365#_c_804_n 6.65751e-19 $X=5.985 $Y=0.85
+ $X2=0 $Y2=0
cc_418 N_A_1109_297#_c_471_n N_A_1225_365#_c_804_n 0.0617069f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_419 N_A_1109_297#_c_474_n N_A_1225_365#_c_812_n 0.00468351f $X=8.95 $Y=1.57
+ $X2=0 $Y2=0
cc_420 N_A_1109_297#_c_461_n N_A_1225_365#_c_806_n 0.00187335f $X=8.98 $Y=0.945
+ $X2=0 $Y2=0
cc_421 N_A_1109_297#_c_469_n N_A_1225_365#_c_806_n 0.00537182f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_422 N_A_1109_297#_c_470_n N_A_1225_365#_c_806_n 0.00520032f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_423 N_A_1109_297#_M1021_g N_A_1225_365#_c_823_n 0.00614563f $X=7.485 $Y=0.455
+ $X2=0 $Y2=0
cc_424 N_A_1109_297#_c_461_n N_A_1225_365#_c_823_n 0.0087978f $X=8.98 $Y=0.945
+ $X2=0 $Y2=0
cc_425 N_A_1109_297#_c_464_n N_A_1225_365#_c_823_n 3.7129e-19 $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_426 N_A_1109_297#_c_465_n N_A_1225_365#_c_823_n 0.0530453f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_427 N_A_1109_297#_c_466_n N_A_1225_365#_c_823_n 0.0955498f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_428 N_A_1109_297#_c_467_n N_A_1225_365#_c_823_n 0.0266362f $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_429 N_A_1109_297#_c_468_n N_A_1225_365#_c_823_n 0.00318096f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_430 N_A_1109_297#_c_469_n N_A_1225_365#_c_823_n 0.0266136f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_431 N_A_1109_297#_c_470_n N_A_1225_365#_c_823_n 0.00475288f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_432 N_A_1109_297#_c_465_n N_A_1225_365#_c_808_n 0.0261136f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_433 N_A_1109_297#_c_471_n N_A_1225_365#_c_808_n 0.00677952f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_434 N_A_1109_297#_c_465_n N_A_1225_365#_c_809_n 0.00119953f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_435 N_A_1109_297#_c_471_n N_A_1225_365#_c_809_n 0.0118823f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_436 N_A_1109_297#_c_461_n N_A_1225_365#_c_836_n 0.00156626f $X=8.98 $Y=0.945
+ $X2=0 $Y2=0
cc_437 N_A_1109_297#_c_461_n N_A_1225_365#_c_837_n 0.00809859f $X=8.98 $Y=0.945
+ $X2=0 $Y2=0
cc_438 N_A_1109_297#_c_474_n N_VPWR_c_942_n 0.00434439f $X=8.95 $Y=1.57 $X2=0
+ $Y2=0
cc_439 N_A_1109_297#_M1022_d N_VPWR_c_931_n 0.00359518f $X=5.545 $Y=1.485 $X2=0
+ $Y2=0
cc_440 N_A_1109_297#_c_474_n N_VPWR_c_931_n 0.00650675f $X=8.95 $Y=1.57 $X2=0
+ $Y2=0
cc_441 N_A_1109_297#_c_466_n N_A_652_325#_M1026_d 0.00140408f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_442 N_A_1109_297#_c_469_n N_A_652_325#_M1026_d 0.00214439f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_443 N_A_1109_297#_c_470_n N_A_652_325#_M1026_d 0.00513165f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_444 N_A_1109_297#_c_462_n N_A_652_325#_c_1123_n 0.00894291f $X=7.36 $Y=1.16
+ $X2=0 $Y2=0
cc_445 N_A_1109_297#_c_464_n N_A_652_325#_c_1123_n 0.0270839f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_446 N_A_1109_297#_c_465_n N_A_652_325#_c_1123_n 5.63647e-19 $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_447 N_A_1109_297#_c_472_n N_A_652_325#_c_1159_n 0.00385601f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_448 N_A_1109_297#_c_472_n N_A_652_325#_c_1124_n 0.0175866f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_449 N_A_1109_297#_c_462_n N_A_652_325#_c_1124_n 7.42472e-19 $X=7.36 $Y=1.16
+ $X2=0 $Y2=0
cc_450 N_A_1109_297#_c_463_n N_A_652_325#_c_1124_n 9.0109e-19 $X=7.46 $Y=1.202
+ $X2=0 $Y2=0
cc_451 N_A_1109_297#_c_464_n N_A_652_325#_c_1124_n 0.00152864f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_452 N_A_1109_297#_c_466_n N_A_652_325#_c_1124_n 0.00419686f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_453 N_A_1109_297#_c_467_n N_A_652_325#_c_1124_n 6.55203e-19 $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_454 N_A_1109_297#_c_472_n N_A_652_325#_c_1120_n 0.00139259f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_455 N_A_1109_297#_M1021_g N_A_652_325#_c_1120_n 0.0164123f $X=7.485 $Y=0.455
+ $X2=0 $Y2=0
cc_456 N_A_1109_297#_c_464_n N_A_652_325#_c_1120_n 0.0173003f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_457 N_A_1109_297#_c_466_n N_A_652_325#_c_1120_n 0.0173494f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_458 N_A_1109_297#_c_467_n N_A_652_325#_c_1120_n 0.00232583f $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_459 N_A_1109_297#_c_468_n N_A_652_325#_c_1120_n 0.0185429f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_460 N_A_1109_297#_c_466_n N_A_652_325#_c_1172_n 0.00166303f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_461 N_A_1109_297#_c_461_n N_A_652_325#_c_1173_n 0.00333256f $X=8.98 $Y=0.945
+ $X2=0 $Y2=0
cc_462 N_A_1109_297#_c_469_n N_A_652_325#_c_1173_n 3.55136e-19 $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_463 N_A_1109_297#_c_470_n N_A_652_325#_c_1173_n 0.00528249f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_464 N_A_1109_297#_c_477_n N_A_652_325#_c_1126_n 0.0270997f $X=5.845 $Y=1.58
+ $X2=0 $Y2=0
cc_465 N_A_1109_297#_c_464_n N_A_652_325#_c_1126_n 8.37577e-19 $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_466 N_A_1109_297#_c_465_n N_A_652_325#_c_1126_n 0.0507283f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_467 N_A_1109_297#_c_481_p N_A_652_325#_c_1126_n 0.0145572f $X=5.985 $Y=0.85
+ $X2=0 $Y2=0
cc_468 N_A_1109_297#_c_471_n N_A_652_325#_c_1126_n 0.00231601f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_469 N_A_1109_297#_c_472_n N_A_652_325#_c_1128_n 0.00348597f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_470 N_A_1109_297#_c_462_n N_A_652_325#_c_1128_n 0.00431105f $X=7.36 $Y=1.16
+ $X2=0 $Y2=0
cc_471 N_A_1109_297#_c_463_n N_A_652_325#_c_1128_n 2.0806e-19 $X=7.46 $Y=1.202
+ $X2=0 $Y2=0
cc_472 N_A_1109_297#_c_464_n N_A_652_325#_c_1128_n 0.00243787f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_473 N_A_1109_297#_c_467_n N_A_652_325#_c_1128_n 0.0154521f $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_474 N_A_1109_297#_c_465_n N_A_658_49#_M1003_d 0.00139415f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_475 N_A_1109_297#_c_467_n N_A_658_49#_M1003_d 5.07779e-19 $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_476 N_A_1109_297#_c_468_n N_A_658_49#_M1003_d 0.00662486f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_477 N_A_1109_297#_c_481_p N_A_658_49#_c_1268_n 0.00193559f $X=5.985 $Y=0.85
+ $X2=0 $Y2=0
cc_478 N_A_1109_297#_c_471_n N_A_658_49#_c_1268_n 0.00327327f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_479 N_A_1109_297#_c_477_n N_A_658_49#_c_1269_n 0.0144112f $X=5.845 $Y=1.58
+ $X2=0 $Y2=0
cc_480 N_A_1109_297#_c_471_n N_A_658_49#_c_1269_n 0.00933598f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_481 N_A_1109_297#_M1022_d N_A_658_49#_c_1277_n 0.0074794f $X=5.545 $Y=1.485
+ $X2=0 $Y2=0
cc_482 N_A_1109_297#_c_477_n N_A_658_49#_c_1277_n 0.0314935f $X=5.845 $Y=1.58
+ $X2=0 $Y2=0
cc_483 N_A_1109_297#_M1022_d N_A_658_49#_c_1278_n 0.00302314f $X=5.545 $Y=1.485
+ $X2=0 $Y2=0
cc_484 N_A_1109_297#_M1022_d N_A_658_49#_c_1280_n 0.00298868f $X=5.545 $Y=1.485
+ $X2=0 $Y2=0
cc_485 N_A_1109_297#_c_472_n N_A_658_49#_c_1270_n 0.00133682f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_486 N_A_1109_297#_c_462_n N_A_658_49#_c_1270_n 6.73654e-19 $X=7.36 $Y=1.16
+ $X2=0 $Y2=0
cc_487 N_A_1109_297#_c_463_n N_A_658_49#_c_1270_n 4.04864e-19 $X=7.46 $Y=1.202
+ $X2=0 $Y2=0
cc_488 N_A_1109_297#_c_464_n N_A_658_49#_c_1270_n 0.0165874f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_489 N_A_1109_297#_c_465_n N_A_658_49#_c_1270_n 0.00618113f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_490 N_A_1109_297#_c_467_n N_A_658_49#_c_1270_n 0.00105795f $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_491 N_A_1109_297#_c_468_n N_A_658_49#_c_1270_n 0.00274672f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_492 N_A_1109_297#_c_472_n N_A_658_49#_c_1282_n 0.00258134f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_493 N_A_1109_297#_c_474_n N_A_658_49#_c_1282_n 0.00822576f $X=8.95 $Y=1.57
+ $X2=0 $Y2=0
cc_494 N_A_1109_297#_M1021_g N_A_658_49#_c_1327_n 0.0022242f $X=7.485 $Y=0.455
+ $X2=0 $Y2=0
cc_495 N_A_1109_297#_c_468_n N_A_658_49#_c_1327_n 0.00181204f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_496 N_A_1109_297#_c_471_n N_A_658_49#_c_1271_n 0.00628163f $X=5.905 $Y=0.72
+ $X2=0 $Y2=0
cc_497 N_A_1109_297#_c_462_n N_A_658_49#_c_1272_n 2.22283e-19 $X=7.36 $Y=1.16
+ $X2=0 $Y2=0
cc_498 N_A_1109_297#_c_464_n N_A_658_49#_c_1272_n 0.00265833f $X=7.247 $Y=0.995
+ $X2=0 $Y2=0
cc_499 N_A_1109_297#_c_465_n N_A_658_49#_c_1272_n 0.0168776f $X=7.125 $Y=0.85
+ $X2=0 $Y2=0
cc_500 N_A_1109_297#_c_467_n N_A_658_49#_c_1272_n 0.00133834f $X=7.415 $Y=0.85
+ $X2=0 $Y2=0
cc_501 N_A_1109_297#_c_468_n N_A_658_49#_c_1272_n 0.0141874f $X=7.27 $Y=0.85
+ $X2=0 $Y2=0
cc_502 N_A_1109_297#_c_466_n N_A_1510_297#_M1021_d 0.00166227f $X=8.605 $Y=0.85
+ $X2=-0.19 $Y2=-0.24
cc_503 N_A_1109_297#_c_472_n N_A_1510_297#_c_1451_n 0.00686704f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_504 N_A_1109_297#_c_466_n N_A_1510_297#_c_1451_n 0.0181022f $X=8.605 $Y=0.85
+ $X2=0 $Y2=0
cc_505 N_A_1109_297#_c_469_n N_A_1510_297#_c_1451_n 0.0020738f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_506 N_A_1109_297#_c_470_n N_A_1510_297#_c_1451_n 0.00517339f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_507 N_A_1109_297#_c_472_n N_A_1510_297#_c_1463_n 0.00431165f $X=7.46 $Y=1.41
+ $X2=0 $Y2=0
cc_508 N_A_1109_297#_c_459_n N_A_1510_297#_c_1464_n 4.12581e-19 $X=8.95 $Y=1.28
+ $X2=0 $Y2=0
cc_509 N_A_1109_297#_c_474_n N_A_1510_297#_c_1464_n 0.0167368f $X=8.95 $Y=1.57
+ $X2=0 $Y2=0
cc_510 N_A_1109_297#_c_470_n N_A_1510_297#_c_1464_n 0.00745833f $X=8.75 $Y=0.85
+ $X2=0 $Y2=0
cc_511 N_A_1109_297#_c_481_p N_VGND_c_1519_n 0.00432343f $X=5.985 $Y=0.85 $X2=0
+ $Y2=0
cc_512 N_A_1109_297#_c_471_n N_VGND_c_1519_n 0.0251293f $X=5.905 $Y=0.72 $X2=0
+ $Y2=0
cc_513 N_A_1109_297#_M1021_g N_VGND_c_1523_n 0.00575161f $X=7.485 $Y=0.455 $X2=0
+ $Y2=0
cc_514 N_A_1109_297#_c_461_n N_VGND_c_1523_n 0.00585385f $X=8.98 $Y=0.945 $X2=0
+ $Y2=0
cc_515 N_A_1109_297#_c_468_n N_VGND_c_1523_n 0.00348958f $X=7.27 $Y=0.85 $X2=0
+ $Y2=0
cc_516 N_A_1109_297#_c_470_n N_VGND_c_1523_n 0.00104987f $X=8.75 $Y=0.85 $X2=0
+ $Y2=0
cc_517 N_A_1109_297#_c_471_n N_VGND_c_1523_n 0.0088551f $X=5.905 $Y=0.72 $X2=0
+ $Y2=0
cc_518 N_A_1109_297#_M1004_d N_VGND_c_1527_n 0.00194539f $X=5.77 $Y=0.235 $X2=0
+ $Y2=0
cc_519 N_A_1109_297#_M1021_g N_VGND_c_1527_n 0.00669445f $X=7.485 $Y=0.455 $X2=0
+ $Y2=0
cc_520 N_A_1109_297#_c_461_n N_VGND_c_1527_n 0.00635456f $X=8.98 $Y=0.945 $X2=0
+ $Y2=0
cc_521 N_A_1109_297#_c_465_n N_VGND_c_1527_n 0.00899211f $X=7.125 $Y=0.85 $X2=0
+ $Y2=0
cc_522 N_A_1109_297#_c_481_p N_VGND_c_1527_n 0.0173285f $X=5.985 $Y=0.85 $X2=0
+ $Y2=0
cc_523 N_A_1109_297#_c_471_n N_VGND_c_1527_n 0.0044502f $X=5.905 $Y=0.72 $X2=0
+ $Y2=0
cc_524 N_B_c_644_n N_A_1225_365#_c_804_n 0.00363086f $X=5.455 $Y=1.41 $X2=0
+ $Y2=0
cc_525 N_B_M1004_g N_A_1225_365#_c_804_n 0.00120086f $X=5.695 $Y=0.56 $X2=0
+ $Y2=0
cc_526 N_B_c_637_n N_A_1225_365#_c_804_n 0.0146583f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_527 N_B_M1018_g N_A_1225_365#_c_804_n 0.00433609f $X=6.65 $Y=1.905 $X2=0
+ $Y2=0
cc_528 N_B_M1003_g N_A_1225_365#_c_804_n 0.00358418f $X=6.675 $Y=0.565 $X2=0
+ $Y2=0
cc_529 N_B_c_640_n N_A_1225_365#_c_804_n 0.00113811f $X=6.65 $Y=1.16 $X2=0 $Y2=0
cc_530 B N_A_1225_365#_c_812_n 0.00522506f $X=8.42 $Y=1.445 $X2=0 $Y2=0
cc_531 N_B_M1003_g N_A_1225_365#_c_823_n 0.00201366f $X=6.675 $Y=0.565 $X2=0
+ $Y2=0
cc_532 N_B_c_643_n N_A_1225_365#_c_823_n 0.00325658f $X=8.365 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_B_M1004_g N_A_1225_365#_c_808_n 4.1997e-19 $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_534 N_B_M1003_g N_A_1225_365#_c_808_n 9.1979e-19 $X=6.675 $Y=0.565 $X2=0
+ $Y2=0
cc_535 N_B_M1004_g N_A_1225_365#_c_809_n 0.00489085f $X=5.695 $Y=0.56 $X2=0
+ $Y2=0
cc_536 N_B_c_637_n N_A_1225_365#_c_809_n 0.00321312f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_537 N_B_c_644_n N_VPWR_c_936_n 0.0113699f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_538 N_B_c_644_n N_VPWR_c_942_n 0.00455828f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_539 N_B_c_648_n N_VPWR_c_942_n 0.0408107f $X=6.75 $Y=2.54 $X2=0 $Y2=0
cc_540 N_B_c_644_n N_VPWR_c_931_n 0.00656627f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_541 N_B_c_647_n N_VPWR_c_931_n 0.0413158f $X=8.285 $Y=2.54 $X2=0 $Y2=0
cc_542 N_B_c_648_n N_VPWR_c_931_n 0.00712076f $X=6.75 $Y=2.54 $X2=0 $Y2=0
cc_543 N_B_M1018_g N_A_652_325#_c_1123_n 0.00142554f $X=6.65 $Y=1.905 $X2=0
+ $Y2=0
cc_544 N_B_M1018_g N_A_652_325#_c_1159_n 0.00438122f $X=6.65 $Y=1.905 $X2=0
+ $Y2=0
cc_545 N_B_c_643_n N_A_652_325#_c_1120_n 0.0026019f $X=8.365 $Y=0.995 $X2=0
+ $Y2=0
cc_546 N_B_c_641_n N_A_652_325#_c_1172_n 4.30216e-19 $X=8.34 $Y=1.16 $X2=0 $Y2=0
cc_547 N_B_c_642_n N_A_652_325#_c_1172_n 0.00286315f $X=8.34 $Y=1.16 $X2=0 $Y2=0
cc_548 N_B_c_643_n N_A_652_325#_c_1172_n 0.00498906f $X=8.365 $Y=0.995 $X2=0
+ $Y2=0
cc_549 N_B_c_641_n N_A_652_325#_c_1173_n 0.00110831f $X=8.34 $Y=1.16 $X2=0 $Y2=0
cc_550 N_B_c_643_n N_A_652_325#_c_1193_n 0.00521263f $X=8.365 $Y=0.995 $X2=0
+ $Y2=0
cc_551 N_B_c_644_n N_A_652_325#_c_1126_n 0.00482215f $X=5.455 $Y=1.41 $X2=0
+ $Y2=0
cc_552 N_B_c_637_n N_A_652_325#_c_1126_n 0.0051668f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_553 N_B_c_638_n N_A_652_325#_c_1126_n 2.58451e-19 $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_554 N_B_M1018_g N_A_652_325#_c_1126_n 0.00401754f $X=6.65 $Y=1.905 $X2=0
+ $Y2=0
cc_555 N_B_c_640_n N_A_652_325#_c_1126_n 2.29578e-19 $X=6.65 $Y=1.16 $X2=0 $Y2=0
cc_556 N_B_M1018_g N_A_652_325#_c_1128_n 4.47596e-19 $X=6.65 $Y=1.905 $X2=0
+ $Y2=0
cc_557 N_B_c_644_n N_A_658_49#_c_1273_n 0.00287893f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_558 N_B_M1004_g N_A_658_49#_c_1268_n 0.00290426f $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_559 N_B_c_644_n N_A_658_49#_c_1269_n 0.0127864f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_560 N_B_c_638_n N_A_658_49#_c_1269_n 0.00534214f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_561 N_B_c_644_n N_A_658_49#_c_1277_n 0.0174362f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_562 N_B_c_644_n N_A_658_49#_c_1278_n 0.00608631f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_563 N_B_M1018_g N_A_658_49#_c_1278_n 9.07378e-19 $X=6.65 $Y=1.905 $X2=0 $Y2=0
cc_564 N_B_c_644_n N_A_658_49#_c_1280_n 0.00366198f $X=5.455 $Y=1.41 $X2=0 $Y2=0
cc_565 N_B_c_637_n N_A_658_49#_c_1270_n 0.00307814f $X=6.55 $Y=1.16 $X2=0 $Y2=0
cc_566 N_B_M1018_g N_A_658_49#_c_1270_n 0.0320054f $X=6.65 $Y=1.905 $X2=0 $Y2=0
cc_567 N_B_M1003_g N_A_658_49#_c_1270_n 0.00658469f $X=6.675 $Y=0.565 $X2=0
+ $Y2=0
cc_568 N_B_c_640_n N_A_658_49#_c_1270_n 0.0107758f $X=6.65 $Y=1.16 $X2=0 $Y2=0
cc_569 N_B_M1018_g N_A_658_49#_c_1282_n 0.00712819f $X=6.65 $Y=1.905 $X2=0 $Y2=0
cc_570 N_B_c_647_n N_A_658_49#_c_1282_n 0.0365765f $X=8.285 $Y=2.54 $X2=0 $Y2=0
cc_571 N_B_c_648_n N_A_658_49#_c_1282_n 2.38151e-19 $X=6.75 $Y=2.54 $X2=0 $Y2=0
cc_572 N_B_M1008_g N_A_658_49#_c_1282_n 0.0102069f $X=8.385 $Y=1.965 $X2=0 $Y2=0
cc_573 N_B_M1003_g N_A_658_49#_c_1327_n 5.72667e-19 $X=6.675 $Y=0.565 $X2=0
+ $Y2=0
cc_574 N_B_M1004_g N_A_658_49#_c_1271_n 8.66132e-19 $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_575 N_B_c_638_n N_A_658_49#_c_1271_n 0.00389387f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_576 N_B_M1003_g N_A_658_49#_c_1272_n 0.0132636f $X=6.675 $Y=0.565 $X2=0 $Y2=0
cc_577 N_B_M1018_g N_A_658_49#_c_1285_n 0.00754618f $X=6.65 $Y=1.905 $X2=0 $Y2=0
cc_578 N_B_c_648_n N_A_658_49#_c_1285_n 2.51585e-19 $X=6.75 $Y=2.54 $X2=0 $Y2=0
cc_579 N_B_c_649_n N_A_1510_297#_c_1451_n 0.00158574f $X=8.385 $Y=1.47 $X2=0
+ $Y2=0
cc_580 N_B_M1008_g N_A_1510_297#_c_1451_n 0.00915065f $X=8.385 $Y=1.965 $X2=0
+ $Y2=0
cc_581 B N_A_1510_297#_c_1451_n 0.0135447f $X=8.42 $Y=1.445 $X2=0 $Y2=0
cc_582 N_B_c_642_n N_A_1510_297#_c_1451_n 0.0332687f $X=8.34 $Y=1.16 $X2=0 $Y2=0
cc_583 N_B_c_643_n N_A_1510_297#_c_1451_n 0.0105486f $X=8.365 $Y=0.995 $X2=0
+ $Y2=0
cc_584 N_B_M1008_g N_A_1510_297#_c_1464_n 0.0111978f $X=8.385 $Y=1.965 $X2=0
+ $Y2=0
cc_585 B N_A_1510_297#_c_1464_n 0.0147778f $X=8.42 $Y=1.445 $X2=0 $Y2=0
cc_586 N_B_c_641_n N_A_1510_297#_c_1464_n 0.00114355f $X=8.34 $Y=1.16 $X2=0
+ $Y2=0
cc_587 N_B_M1004_g N_VGND_c_1519_n 0.0194419f $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_588 N_B_c_638_n N_VGND_c_1519_n 0.00530155f $X=5.77 $Y=1.16 $X2=0 $Y2=0
cc_589 N_B_M1004_g N_VGND_c_1523_n 0.00494995f $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_590 N_B_M1003_g N_VGND_c_1523_n 0.00427876f $X=6.675 $Y=0.565 $X2=0 $Y2=0
cc_591 N_B_c_643_n N_VGND_c_1523_n 0.00357877f $X=8.365 $Y=0.995 $X2=0 $Y2=0
cc_592 N_B_M1004_g N_VGND_c_1527_n 0.00933567f $X=5.695 $Y=0.56 $X2=0 $Y2=0
cc_593 N_B_M1003_g N_VGND_c_1527_n 0.00718941f $X=6.675 $Y=0.565 $X2=0 $Y2=0
cc_594 N_B_c_643_n N_VGND_c_1527_n 0.00613199f $X=8.365 $Y=0.995 $X2=0 $Y2=0
cc_595 N_A_c_765_n N_A_1225_365#_c_802_n 0.0575966f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_596 A N_A_1225_365#_c_802_n 8.4217e-19 $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_597 N_A_c_766_n N_A_1225_365#_c_803_n 0.0174128f $X=9.53 $Y=0.995 $X2=0 $Y2=0
cc_598 N_A_c_765_n N_A_1225_365#_c_812_n 0.0147059f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_599 A N_A_1225_365#_c_812_n 0.0301432f $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_600 N_A_c_765_n N_A_1225_365#_c_805_n 5.76324e-19 $X=9.505 $Y=1.41 $X2=0
+ $Y2=0
cc_601 N_A_c_766_n N_A_1225_365#_c_805_n 0.0116619f $X=9.53 $Y=0.995 $X2=0 $Y2=0
cc_602 A N_A_1225_365#_c_805_n 0.0142387f $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_603 N_A_c_765_n N_A_1225_365#_c_806_n 0.00444032f $X=9.505 $Y=1.41 $X2=0
+ $Y2=0
cc_604 A N_A_1225_365#_c_806_n 0.0205785f $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_605 N_A_c_765_n N_A_1225_365#_c_807_n 7.08841e-19 $X=9.505 $Y=1.41 $X2=0
+ $Y2=0
cc_606 N_A_c_766_n N_A_1225_365#_c_807_n 0.00356706f $X=9.53 $Y=0.995 $X2=0
+ $Y2=0
cc_607 A N_A_1225_365#_c_807_n 0.0208188f $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_608 N_A_c_765_n N_A_1225_365#_c_813_n 0.00343171f $X=9.505 $Y=1.41 $X2=0
+ $Y2=0
cc_609 A N_A_1225_365#_c_836_n 9.51454e-19 $X=9.35 $Y=1.105 $X2=0 $Y2=0
cc_610 N_A_c_765_n N_VPWR_c_937_n 0.00315802f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_611 N_A_c_765_n N_VPWR_c_942_n 0.00506535f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_612 N_A_c_765_n N_VPWR_c_931_n 0.00688028f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_613 N_A_c_765_n N_A_658_49#_c_1282_n 0.00163845f $X=9.505 $Y=1.41 $X2=0 $Y2=0
cc_614 N_A_c_765_n N_A_1510_297#_c_1464_n 0.0144611f $X=9.505 $Y=1.41 $X2=0
+ $Y2=0
cc_615 N_A_c_766_n N_VGND_c_1520_n 0.00471691f $X=9.53 $Y=0.995 $X2=0 $Y2=0
cc_616 N_A_c_766_n N_VGND_c_1523_n 0.00439206f $X=9.53 $Y=0.995 $X2=0 $Y2=0
cc_617 N_A_c_766_n N_VGND_c_1527_n 0.00661448f $X=9.53 $Y=0.995 $X2=0 $Y2=0
cc_618 N_A_1225_365#_c_812_n N_VPWR_M1009_d 0.00546234f $X=9.805 $Y=1.6 $X2=0
+ $Y2=0
cc_619 N_A_1225_365#_c_802_n N_VPWR_c_937_n 0.00802533f $X=10.015 $Y=1.41 $X2=0
+ $Y2=0
cc_620 N_A_1225_365#_c_802_n N_VPWR_c_945_n 0.00449565f $X=10.015 $Y=1.41 $X2=0
+ $Y2=0
cc_621 N_A_1225_365#_M1006_d N_VPWR_c_931_n 0.00402227f $X=9.04 $Y=1.645 $X2=0
+ $Y2=0
cc_622 N_A_1225_365#_c_802_n N_VPWR_c_931_n 0.00605666f $X=10.015 $Y=1.41 $X2=0
+ $Y2=0
cc_623 N_A_1225_365#_c_823_n N_A_652_325#_M1026_d 0.00427772f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_624 N_A_1225_365#_c_823_n N_A_652_325#_c_1120_n 0.014738f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_625 N_A_1225_365#_c_823_n N_A_652_325#_c_1172_n 0.00610486f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_626 N_A_1225_365#_c_823_n N_A_652_325#_c_1173_n 0.00980954f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_627 N_A_1225_365#_c_836_n N_A_652_325#_c_1173_n 0.0012274f $X=9.26 $Y=0.51
+ $X2=0 $Y2=0
cc_628 N_A_1225_365#_c_837_n N_A_652_325#_c_1173_n 0.00676874f $X=9.26 $Y=0.51
+ $X2=0 $Y2=0
cc_629 N_A_1225_365#_c_823_n N_A_652_325#_c_1193_n 0.0119237f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_630 N_A_1225_365#_M1018_s N_A_652_325#_c_1126_n 0.00840572f $X=6.125 $Y=1.825
+ $X2=0 $Y2=0
cc_631 N_A_1225_365#_c_804_n N_A_652_325#_c_1126_n 0.0184168f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_632 N_A_1225_365#_c_823_n N_A_658_49#_M1003_d 0.00606718f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_633 N_A_1225_365#_c_804_n N_A_658_49#_c_1277_n 0.0138372f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_634 N_A_1225_365#_c_804_n N_A_658_49#_c_1278_n 0.0028603f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_635 N_A_1225_365#_M1018_s N_A_658_49#_c_1279_n 0.0104901f $X=6.125 $Y=1.825
+ $X2=0 $Y2=0
cc_636 N_A_1225_365#_c_804_n N_A_658_49#_c_1279_n 0.0128549f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_637 N_A_1225_365#_c_804_n N_A_658_49#_c_1270_n 0.0619836f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_638 N_A_1225_365#_M1006_d N_A_658_49#_c_1282_n 0.00281879f $X=9.04 $Y=1.645
+ $X2=0 $Y2=0
cc_639 N_A_1225_365#_c_823_n N_A_658_49#_c_1327_n 0.0125744f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_640 N_A_1225_365#_c_808_n N_A_658_49#_c_1327_n 0.00143452f $X=6.445 $Y=0.51
+ $X2=0 $Y2=0
cc_641 N_A_1225_365#_c_809_n N_A_658_49#_c_1327_n 0.00335094f $X=6.3 $Y=0.51
+ $X2=0 $Y2=0
cc_642 N_A_1225_365#_M1003_s N_A_658_49#_c_1272_n 0.00143708f $X=6.29 $Y=0.245
+ $X2=0 $Y2=0
cc_643 N_A_1225_365#_c_804_n N_A_658_49#_c_1272_n 0.0110368f $X=6.25 $Y=1.94
+ $X2=0 $Y2=0
cc_644 N_A_1225_365#_c_823_n N_A_658_49#_c_1272_n 0.00357405f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_645 N_A_1225_365#_c_809_n N_A_658_49#_c_1272_n 0.00104769f $X=6.3 $Y=0.51
+ $X2=0 $Y2=0
cc_646 N_A_1225_365#_c_823_n N_A_1510_297#_M1021_d 0.00653094f $X=9.115 $Y=0.51
+ $X2=-0.19 $Y2=-0.24
cc_647 N_A_1225_365#_c_823_n N_A_1510_297#_c_1451_n 0.00162336f $X=9.115 $Y=0.51
+ $X2=0 $Y2=0
cc_648 N_A_1225_365#_c_802_n N_A_1510_297#_c_1452_n 0.020342f $X=10.015 $Y=1.41
+ $X2=0 $Y2=0
cc_649 N_A_1225_365#_c_803_n N_A_1510_297#_c_1452_n 0.0102506f $X=10.04 $Y=0.995
+ $X2=0 $Y2=0
cc_650 N_A_1225_365#_c_812_n N_A_1510_297#_c_1452_n 0.0112209f $X=9.805 $Y=1.6
+ $X2=0 $Y2=0
cc_651 N_A_1225_365#_c_807_n N_A_1510_297#_c_1452_n 0.0335352f $X=9.89 $Y=1.325
+ $X2=0 $Y2=0
cc_652 N_A_1225_365#_c_813_n N_A_1510_297#_c_1452_n 0.00830245f $X=9.89 $Y=1.495
+ $X2=0 $Y2=0
cc_653 N_A_1225_365#_M1006_d N_A_1510_297#_c_1464_n 0.00774465f $X=9.04 $Y=1.645
+ $X2=0 $Y2=0
cc_654 N_A_1225_365#_c_802_n N_A_1510_297#_c_1464_n 2.11775e-19 $X=10.015
+ $Y=1.41 $X2=0 $Y2=0
cc_655 N_A_1225_365#_c_812_n N_A_1510_297#_c_1464_n 0.0377124f $X=9.805 $Y=1.6
+ $X2=0 $Y2=0
cc_656 N_A_1225_365#_c_802_n N_A_1510_297#_c_1457_n 0.0156096f $X=10.015 $Y=1.41
+ $X2=0 $Y2=0
cc_657 N_A_1225_365#_c_812_n N_A_1510_297#_c_1457_n 0.00381196f $X=9.805 $Y=1.6
+ $X2=0 $Y2=0
cc_658 N_A_1225_365#_c_807_n N_A_1510_297#_c_1457_n 0.0016745f $X=9.89 $Y=1.325
+ $X2=0 $Y2=0
cc_659 N_A_1225_365#_c_805_n N_VGND_M1015_d 0.00176133f $X=9.805 $Y=0.82 $X2=0
+ $Y2=0
cc_660 N_A_1225_365#_c_807_n N_VGND_M1015_d 0.00151302f $X=9.89 $Y=1.325 $X2=0
+ $Y2=0
cc_661 N_A_1225_365#_c_802_n N_VGND_c_1520_n 2.16114e-19 $X=10.015 $Y=1.41 $X2=0
+ $Y2=0
cc_662 N_A_1225_365#_c_803_n N_VGND_c_1520_n 0.00419914f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_663 N_A_1225_365#_c_805_n N_VGND_c_1520_n 0.00851939f $X=9.805 $Y=0.82 $X2=0
+ $Y2=0
cc_664 N_A_1225_365#_c_807_n N_VGND_c_1520_n 0.00511527f $X=9.89 $Y=1.325 $X2=0
+ $Y2=0
cc_665 N_A_1225_365#_c_836_n N_VGND_c_1520_n 0.00111658f $X=9.26 $Y=0.51 $X2=0
+ $Y2=0
cc_666 N_A_1225_365#_c_805_n N_VGND_c_1523_n 0.00300328f $X=9.805 $Y=0.82 $X2=0
+ $Y2=0
cc_667 N_A_1225_365#_c_823_n N_VGND_c_1523_n 0.00575847f $X=9.115 $Y=0.51 $X2=0
+ $Y2=0
cc_668 N_A_1225_365#_c_808_n N_VGND_c_1523_n 2.49898e-19 $X=6.445 $Y=0.51 $X2=0
+ $Y2=0
cc_669 N_A_1225_365#_c_809_n N_VGND_c_1523_n 0.0254286f $X=6.3 $Y=0.51 $X2=0
+ $Y2=0
cc_670 N_A_1225_365#_c_836_n N_VGND_c_1523_n 3.63685e-19 $X=9.26 $Y=0.51 $X2=0
+ $Y2=0
cc_671 N_A_1225_365#_c_837_n N_VGND_c_1523_n 0.0149689f $X=9.26 $Y=0.51 $X2=0
+ $Y2=0
cc_672 N_A_1225_365#_c_803_n N_VGND_c_1526_n 0.0057563f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_673 N_A_1225_365#_c_807_n N_VGND_c_1526_n 0.00124625f $X=9.89 $Y=1.325 $X2=0
+ $Y2=0
cc_674 N_A_1225_365#_M1027_d N_VGND_c_1527_n 0.00240207f $X=9.055 $Y=0.235 $X2=0
+ $Y2=0
cc_675 N_A_1225_365#_c_803_n N_VGND_c_1527_n 0.0116259f $X=10.04 $Y=0.995 $X2=0
+ $Y2=0
cc_676 N_A_1225_365#_c_805_n N_VGND_c_1527_n 0.00646188f $X=9.805 $Y=0.82 $X2=0
+ $Y2=0
cc_677 N_A_1225_365#_c_807_n N_VGND_c_1527_n 0.00327885f $X=9.89 $Y=1.325 $X2=0
+ $Y2=0
cc_678 N_A_1225_365#_c_823_n N_VGND_c_1527_n 0.232956f $X=9.115 $Y=0.51 $X2=0
+ $Y2=0
cc_679 N_A_1225_365#_c_808_n N_VGND_c_1527_n 0.0285546f $X=6.445 $Y=0.51 $X2=0
+ $Y2=0
cc_680 N_A_1225_365#_c_809_n N_VGND_c_1527_n 0.00396297f $X=6.3 $Y=0.51 $X2=0
+ $Y2=0
cc_681 N_A_1225_365#_c_836_n N_VGND_c_1527_n 0.0285254f $X=9.26 $Y=0.51 $X2=0
+ $Y2=0
cc_682 N_A_1225_365#_c_837_n N_VGND_c_1527_n 0.0036194f $X=9.26 $Y=0.51 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_931_n N_X_M1000_s 0.0061735f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_684 N_VPWR_c_931_n N_X_M1012_s 0.0061735f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_685 N_VPWR_c_932_n N_X_c_1091_n 0.0157757f $X=0.36 $Y=2.3 $X2=0 $Y2=0
cc_686 N_VPWR_c_933_n N_X_c_1091_n 0.0118139f $X=1.135 $Y=2.72 $X2=0 $Y2=0
cc_687 N_VPWR_c_934_n N_X_c_1091_n 0.0151355f $X=1.3 $Y=2.3 $X2=0 $Y2=0
cc_688 N_VPWR_c_931_n N_X_c_1091_n 0.00646998f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_689 N_VPWR_c_934_n N_X_c_1095_n 0.0151355f $X=1.3 $Y=2.3 $X2=0 $Y2=0
cc_690 N_VPWR_c_935_n N_X_c_1095_n 0.0151355f $X=2.24 $Y=2.3 $X2=0 $Y2=0
cc_691 N_VPWR_c_940_n N_X_c_1095_n 0.0118139f $X=2.075 $Y=2.72 $X2=0 $Y2=0
cc_692 N_VPWR_c_931_n N_X_c_1095_n 0.00646998f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_693 N_VPWR_M1011_d N_X_c_1060_n 0.00188666f $X=1.155 $Y=1.485 $X2=0 $Y2=0
cc_694 N_VPWR_c_933_n N_X_c_1060_n 0.00268748f $X=1.135 $Y=2.72 $X2=0 $Y2=0
cc_695 N_VPWR_c_934_n N_X_c_1060_n 0.0179606f $X=1.3 $Y=2.3 $X2=0 $Y2=0
cc_696 N_VPWR_c_940_n N_X_c_1060_n 0.00269999f $X=2.075 $Y=2.72 $X2=0 $Y2=0
cc_697 N_VPWR_c_931_n N_X_c_1060_n 0.00979924f $X=10.35 $Y=2.72 $X2=0 $Y2=0
cc_698 N_VPWR_c_944_n N_A_652_325#_c_1121_n 0.00407465f $X=5.055 $Y=2.72 $X2=0
+ $Y2=0
cc_699 N_VPWR_c_931_n N_A_652_325#_c_1121_n 0.0092333f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_700 N_VPWR_M1022_s N_A_652_325#_c_1126_n 0.00109947f $X=5.095 $Y=1.485 $X2=0
+ $Y2=0
cc_701 N_VPWR_c_931_n N_A_658_49#_M1008_d 0.00241089f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_702 N_VPWR_c_936_n N_A_658_49#_c_1274_n 0.00147971f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_703 N_VPWR_c_944_n N_A_658_49#_c_1274_n 0.00296166f $X=5.055 $Y=2.72 $X2=0
+ $Y2=0
cc_704 N_VPWR_c_931_n N_A_658_49#_c_1274_n 0.00485654f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_705 N_VPWR_M1022_s N_A_658_49#_c_1269_n 0.00659923f $X=5.095 $Y=1.485 $X2=0
+ $Y2=0
cc_706 N_VPWR_M1022_s N_A_658_49#_c_1277_n 0.00155527f $X=5.095 $Y=1.485 $X2=0
+ $Y2=0
cc_707 N_VPWR_c_936_n N_A_658_49#_c_1277_n 0.00612755f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_708 N_VPWR_c_942_n N_A_658_49#_c_1277_n 0.00666556f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_709 N_VPWR_c_931_n N_A_658_49#_c_1277_n 0.0119497f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_710 N_VPWR_c_936_n N_A_658_49#_c_1278_n 0.00140976f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_711 N_VPWR_c_942_n N_A_658_49#_c_1279_n 0.0305955f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_712 N_VPWR_c_931_n N_A_658_49#_c_1279_n 0.0196786f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_713 N_VPWR_c_936_n N_A_658_49#_c_1280_n 0.00679194f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_714 N_VPWR_c_942_n N_A_658_49#_c_1280_n 0.0105745f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_715 N_VPWR_c_931_n N_A_658_49#_c_1280_n 0.00644066f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_716 N_VPWR_c_942_n N_A_658_49#_c_1282_n 0.134152f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_717 N_VPWR_c_931_n N_A_658_49#_c_1282_n 0.0807991f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_718 N_VPWR_c_936_n N_A_658_49#_c_1283_n 0.0142739f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_719 N_VPWR_c_944_n N_A_658_49#_c_1283_n 0.0186431f $X=5.055 $Y=2.72 $X2=0
+ $Y2=0
cc_720 N_VPWR_c_931_n N_A_658_49#_c_1283_n 0.0145279f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_721 N_VPWR_M1022_s N_A_658_49#_c_1284_n 0.00243878f $X=5.095 $Y=1.485 $X2=0
+ $Y2=0
cc_722 N_VPWR_c_936_n N_A_658_49#_c_1284_n 0.0143988f $X=5.22 $Y=2.32 $X2=0
+ $Y2=0
cc_723 N_VPWR_c_931_n N_A_658_49#_c_1284_n 8.22076e-19 $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_724 N_VPWR_c_942_n N_A_658_49#_c_1285_n 0.0102998f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_725 N_VPWR_c_931_n N_A_658_49#_c_1285_n 0.0058084f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_726 N_VPWR_c_931_n N_A_1510_297#_M1010_d 0.00237688f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_727 N_VPWR_c_937_n N_A_1510_297#_c_1455_n 0.0118776f $X=9.78 $Y=2.36 $X2=0
+ $Y2=0
cc_728 N_VPWR_c_945_n N_A_1510_297#_c_1455_n 0.0173928f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_729 N_VPWR_c_931_n N_A_1510_297#_c_1455_n 0.00977915f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_730 N_VPWR_M1009_d N_A_1510_297#_c_1464_n 0.00475729f $X=9.595 $Y=1.485 $X2=0
+ $Y2=0
cc_731 N_VPWR_c_937_n N_A_1510_297#_c_1464_n 0.0177094f $X=9.78 $Y=2.36 $X2=0
+ $Y2=0
cc_732 N_VPWR_c_942_n N_A_1510_297#_c_1464_n 0.00831891f $X=9.615 $Y=2.72 $X2=0
+ $Y2=0
cc_733 N_VPWR_c_931_n N_A_1510_297#_c_1464_n 0.0168826f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_734 N_VPWR_c_945_n N_A_1510_297#_c_1457_n 0.00344451f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_735 N_VPWR_c_931_n N_A_1510_297#_c_1457_n 0.00563469f $X=10.35 $Y=2.72 $X2=0
+ $Y2=0
cc_736 N_X_c_1055_n N_VGND_M1016_d 9.03344e-19 $X=1.205 $Y=0.792 $X2=0 $Y2=0
cc_737 N_X_c_1058_n N_VGND_M1016_d 0.00139194f $X=1.48 $Y=0.792 $X2=0 $Y2=0
cc_738 N_X_c_1075_n N_VGND_c_1517_n 0.00709805f $X=1.67 $Y=0.56 $X2=0 $Y2=0
cc_739 N_X_c_1058_n N_VGND_c_1517_n 0.00318227f $X=1.48 $Y=0.792 $X2=0 $Y2=0
cc_740 N_X_c_1061_n N_VGND_c_1525_n 0.00709805f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_741 N_X_c_1055_n N_VGND_c_1525_n 0.00235507f $X=1.205 $Y=0.792 $X2=0 $Y2=0
cc_742 N_X_M1002_s N_VGND_c_1527_n 0.00481217f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_743 N_X_M1017_s N_VGND_c_1527_n 0.00632802f $X=1.535 $Y=0.235 $X2=0 $Y2=0
cc_744 N_X_c_1061_n N_VGND_c_1527_n 0.00611294f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_745 N_X_c_1055_n N_VGND_c_1527_n 0.00546587f $X=1.205 $Y=0.792 $X2=0 $Y2=0
cc_746 N_X_c_1075_n N_VGND_c_1527_n 0.00611294f $X=1.67 $Y=0.56 $X2=0 $Y2=0
cc_747 N_X_c_1058_n N_VGND_c_1527_n 0.00647762f $X=1.48 $Y=0.792 $X2=0 $Y2=0
cc_748 N_X_c_1061_n N_VGND_c_1528_n 0.00858539f $X=0.73 $Y=0.56 $X2=0 $Y2=0
cc_749 N_X_c_1055_n N_VGND_c_1528_n 0.0108868f $X=1.205 $Y=0.792 $X2=0 $Y2=0
cc_750 N_X_c_1058_n N_VGND_c_1528_n 0.00922799f $X=1.48 $Y=0.792 $X2=0 $Y2=0
cc_751 N_A_652_325#_c_1121_n N_A_658_49#_M1001_d 0.00619557f $X=4.375 $Y=1.98
+ $X2=0 $Y2=0
cc_752 N_A_652_325#_c_1141_n N_A_658_49#_M1001_d 0.00677252f $X=4.46 $Y=1.895
+ $X2=0 $Y2=0
cc_753 N_A_652_325#_c_1129_n N_A_658_49#_M1001_d 0.00697789f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_754 N_A_652_325#_M1013_d N_A_658_49#_c_1266_n 0.00334341f $X=4.36 $Y=0.245
+ $X2=0 $Y2=0
cc_755 N_A_652_325#_c_1119_n N_A_658_49#_c_1266_n 0.0138308f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_756 N_A_652_325#_M1013_d N_A_658_49#_c_1290_n 0.00348437f $X=4.36 $Y=0.245
+ $X2=0 $Y2=0
cc_757 N_A_652_325#_c_1119_n N_A_658_49#_c_1290_n 0.00440606f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_758 N_A_652_325#_M1013_d N_A_658_49#_c_1267_n 0.0175141f $X=4.36 $Y=0.245
+ $X2=0 $Y2=0
cc_759 N_A_652_325#_c_1119_n N_A_658_49#_c_1267_n 0.0128008f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_760 N_A_652_325#_M1013_d N_A_658_49#_c_1291_n 3.2099e-19 $X=4.36 $Y=0.245
+ $X2=0 $Y2=0
cc_761 N_A_652_325#_c_1126_n N_A_658_49#_c_1274_n 0.00437461f $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_762 N_A_652_325#_c_1127_n N_A_658_49#_c_1274_n 0.00277011f $X=4.965 $Y=1.53
+ $X2=0 $Y2=0
cc_763 N_A_652_325#_c_1129_n N_A_658_49#_c_1274_n 0.00125154f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_764 N_A_652_325#_c_1121_n N_A_658_49#_c_1275_n 0.0153275f $X=4.375 $Y=1.98
+ $X2=0 $Y2=0
cc_765 N_A_652_325#_c_1127_n N_A_658_49#_c_1275_n 0.00119193f $X=4.965 $Y=1.53
+ $X2=0 $Y2=0
cc_766 N_A_652_325#_c_1129_n N_A_658_49#_c_1275_n 0.0114314f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_767 N_A_652_325#_c_1119_n N_A_658_49#_c_1268_n 0.0327079f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_768 N_A_652_325#_c_1141_n N_A_658_49#_c_1269_n 0.00649967f $X=4.46 $Y=1.895
+ $X2=0 $Y2=0
cc_769 N_A_652_325#_c_1119_n N_A_658_49#_c_1269_n 0.00889026f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_770 N_A_652_325#_c_1126_n N_A_658_49#_c_1269_n 0.0221806f $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_771 N_A_652_325#_c_1127_n N_A_658_49#_c_1269_n 0.00275249f $X=4.965 $Y=1.53
+ $X2=0 $Y2=0
cc_772 N_A_652_325#_c_1129_n N_A_658_49#_c_1269_n 0.0233325f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_773 N_A_652_325#_c_1126_n N_A_658_49#_c_1277_n 0.011487f $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_774 N_A_652_325#_c_1123_n N_A_658_49#_c_1270_n 0.00911487f $X=7.122 $Y=1.615
+ $X2=0 $Y2=0
cc_775 N_A_652_325#_c_1159_n N_A_658_49#_c_1270_n 0.0264421f $X=7.09 $Y=1.62
+ $X2=0 $Y2=0
cc_776 N_A_652_325#_c_1126_n N_A_658_49#_c_1270_n 0.0195229f $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_777 N_A_652_325#_c_1128_n N_A_658_49#_c_1270_n 0.00128822f $X=7.27 $Y=1.53
+ $X2=0 $Y2=0
cc_778 N_A_652_325#_M1018_d N_A_658_49#_c_1282_n 0.0094538f $X=6.74 $Y=1.485
+ $X2=0 $Y2=0
cc_779 N_A_652_325#_c_1159_n N_A_658_49#_c_1282_n 0.0238103f $X=7.09 $Y=1.62
+ $X2=0 $Y2=0
cc_780 N_A_652_325#_c_1124_n N_A_658_49#_c_1282_n 0.0100462f $X=7.575 $Y=1.53
+ $X2=0 $Y2=0
cc_781 N_A_652_325#_c_1120_n N_A_658_49#_c_1327_n 0.00250545f $X=7.66 $Y=1.445
+ $X2=0 $Y2=0
cc_782 N_A_652_325#_c_1121_n N_A_658_49#_c_1283_n 0.0049241f $X=4.375 $Y=1.98
+ $X2=0 $Y2=0
cc_783 N_A_652_325#_c_1127_n N_A_658_49#_c_1283_n 2.48159e-19 $X=4.965 $Y=1.53
+ $X2=0 $Y2=0
cc_784 N_A_652_325#_c_1129_n N_A_658_49#_c_1283_n 0.00535873f $X=4.705 $Y=1.535
+ $X2=0 $Y2=0
cc_785 N_A_652_325#_c_1119_n N_A_658_49#_c_1271_n 0.0133806f $X=4.705 $Y=0.76
+ $X2=0 $Y2=0
cc_786 N_A_652_325#_c_1126_n N_A_658_49#_c_1271_n 0.0053051f $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_787 N_A_652_325#_c_1127_n N_A_658_49#_c_1271_n 2.6396e-19 $X=4.965 $Y=1.53
+ $X2=0 $Y2=0
cc_788 N_A_652_325#_c_1123_n N_A_658_49#_c_1272_n 2.53366e-19 $X=7.122 $Y=1.615
+ $X2=0 $Y2=0
cc_789 N_A_652_325#_c_1126_n N_A_658_49#_c_1272_n 7.5408e-19 $X=7.125 $Y=1.53
+ $X2=0 $Y2=0
cc_790 N_A_652_325#_c_1120_n N_A_1510_297#_M1021_d 0.00729398f $X=7.66 $Y=1.445
+ $X2=-0.19 $Y2=-0.24
cc_791 N_A_652_325#_c_1252_p N_A_1510_297#_M1021_d 0.0024562f $X=7.745 $Y=0.34
+ $X2=-0.19 $Y2=-0.24
cc_792 N_A_652_325#_c_1193_n N_A_1510_297#_M1021_d 0.0107136f $X=8.255 $Y=0.36
+ $X2=-0.19 $Y2=-0.24
cc_793 N_A_652_325#_c_1124_n N_A_1510_297#_M1014_d 0.00443096f $X=7.575 $Y=1.53
+ $X2=0 $Y2=0
cc_794 N_A_652_325#_c_1159_n N_A_1510_297#_c_1451_n 0.00453141f $X=7.09 $Y=1.62
+ $X2=0 $Y2=0
cc_795 N_A_652_325#_c_1124_n N_A_1510_297#_c_1451_n 0.013519f $X=7.575 $Y=1.53
+ $X2=0 $Y2=0
cc_796 N_A_652_325#_c_1120_n N_A_1510_297#_c_1451_n 0.062318f $X=7.66 $Y=1.445
+ $X2=0 $Y2=0
cc_797 N_A_652_325#_c_1193_n N_A_1510_297#_c_1451_n 0.0106102f $X=8.255 $Y=0.36
+ $X2=0 $Y2=0
cc_798 N_A_652_325#_c_1128_n N_A_1510_297#_c_1451_n 0.00130235f $X=7.27 $Y=1.53
+ $X2=0 $Y2=0
cc_799 N_A_652_325#_c_1126_n N_VGND_c_1519_n 0.00568966f $X=7.125 $Y=1.53 $X2=0
+ $Y2=0
cc_800 N_A_652_325#_c_1252_p N_VGND_c_1523_n 0.0104913f $X=7.745 $Y=0.34 $X2=0
+ $Y2=0
cc_801 N_A_652_325#_c_1193_n N_VGND_c_1523_n 0.0617902f $X=8.255 $Y=0.36 $X2=0
+ $Y2=0
cc_802 N_A_652_325#_M1026_d N_VGND_c_1527_n 0.00231474f $X=8.355 $Y=0.245 $X2=0
+ $Y2=0
cc_803 N_A_652_325#_c_1252_p N_VGND_c_1527_n 0.00184693f $X=7.745 $Y=0.34 $X2=0
+ $Y2=0
cc_804 N_A_652_325#_c_1193_n N_VGND_c_1527_n 0.00974346f $X=8.255 $Y=0.36 $X2=0
+ $Y2=0
cc_805 N_A_658_49#_c_1282_n N_A_1510_297#_M1014_d 0.00563686f $X=8.705 $Y=2.36
+ $X2=0 $Y2=0
cc_806 N_A_658_49#_c_1282_n N_A_1510_297#_c_1463_n 0.0129278f $X=8.705 $Y=2.36
+ $X2=0 $Y2=0
cc_807 N_A_658_49#_M1008_d N_A_1510_297#_c_1464_n 0.00785854f $X=8.475 $Y=1.645
+ $X2=0 $Y2=0
cc_808 N_A_658_49#_c_1282_n N_A_1510_297#_c_1464_n 0.0533312f $X=8.705 $Y=2.36
+ $X2=0 $Y2=0
cc_809 N_A_658_49#_c_1267_n N_VGND_c_1519_n 0.0141318f $X=4.96 $Y=0.34 $X2=0
+ $Y2=0
cc_810 N_A_658_49#_c_1268_n N_VGND_c_1519_n 0.0336084f $X=5.045 $Y=1.035 $X2=0
+ $Y2=0
cc_811 N_A_658_49#_c_1266_n N_VGND_c_1521_n 0.00239374f $X=4.23 $Y=0.74 $X2=0
+ $Y2=0
cc_812 N_A_658_49#_c_1267_n N_VGND_c_1521_n 0.0445697f $X=4.96 $Y=0.34 $X2=0
+ $Y2=0
cc_813 N_A_658_49#_c_1291_n N_VGND_c_1521_n 0.0130641f $X=4.45 $Y=0.34 $X2=0
+ $Y2=0
cc_814 N_A_658_49#_c_1327_n N_VGND_c_1523_n 0.00800682f $X=6.885 $Y=0.545 $X2=0
+ $Y2=0
cc_815 N_A_658_49#_c_1272_n N_VGND_c_1523_n 0.00285234f $X=6.61 $Y=0.772 $X2=0
+ $Y2=0
cc_816 N_A_658_49#_c_1266_n N_VGND_c_1527_n 0.00649067f $X=4.23 $Y=0.74 $X2=0
+ $Y2=0
cc_817 N_A_658_49#_c_1267_n N_VGND_c_1527_n 0.0255342f $X=4.96 $Y=0.34 $X2=0
+ $Y2=0
cc_818 N_A_658_49#_c_1291_n N_VGND_c_1527_n 0.00783952f $X=4.45 $Y=0.34 $X2=0
+ $Y2=0
cc_819 N_A_658_49#_c_1327_n N_VGND_c_1527_n 0.0018012f $X=6.885 $Y=0.545 $X2=0
+ $Y2=0
cc_820 N_A_1510_297#_c_1453_n N_VGND_c_1526_n 0.0170867f $X=10.34 $Y=0.42 $X2=0
+ $Y2=0
cc_821 N_A_1510_297#_M1024_d N_VGND_c_1527_n 0.00379446f $X=10.115 $Y=0.235
+ $X2=0 $Y2=0
cc_822 N_A_1510_297#_c_1453_n N_VGND_c_1527_n 0.00982816f $X=10.34 $Y=0.42 $X2=0
+ $Y2=0
