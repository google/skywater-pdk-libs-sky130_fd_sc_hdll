* File: sky130_fd_sc_hdll__nor3b_2.pxi.spice
* Created: Wed Sep  2 08:40:42 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%A N_A_c_65_n N_A_M1006_g N_A_c_69_n N_A_M1001_g
+ N_A_c_70_n N_A_M1010_g N_A_c_66_n N_A_M1012_g A A N_A_c_68_n A
+ PM_SKY130_FD_SC_HDLL__NOR3B_2%A
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%B N_B_c_102_n N_B_M1007_g N_B_c_106_n
+ N_B_M1003_g N_B_c_107_n N_B_M1004_g N_B_c_103_n N_B_M1011_g B N_B_c_105_n B
+ PM_SKY130_FD_SC_HDLL__NOR3B_2%B
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%A_571_21# N_A_571_21#_M1002_s
+ N_A_571_21#_M1009_s N_A_571_21#_c_144_n N_A_571_21#_M1005_g
+ N_A_571_21#_c_152_n N_A_571_21#_M1000_g N_A_571_21#_c_145_n
+ N_A_571_21#_M1008_g N_A_571_21#_c_153_n N_A_571_21#_M1013_g
+ N_A_571_21#_c_146_n N_A_571_21#_c_147_n N_A_571_21#_c_148_n
+ N_A_571_21#_c_149_n N_A_571_21#_c_154_n N_A_571_21#_c_150_n
+ N_A_571_21#_c_151_n PM_SKY130_FD_SC_HDLL__NOR3B_2%A_571_21#
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%C_N N_C_N_c_206_n N_C_N_M1002_g N_C_N_c_207_n
+ N_C_N_M1009_g C_N C_N PM_SKY130_FD_SC_HDLL__NOR3B_2%C_N
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%A_27_297# N_A_27_297#_M1001_s
+ N_A_27_297#_M1010_s N_A_27_297#_M1004_d N_A_27_297#_c_231_n
+ N_A_27_297#_c_232_n N_A_27_297#_c_233_n N_A_27_297#_c_254_p
+ N_A_27_297#_c_234_n N_A_27_297#_c_235_n N_A_27_297#_c_236_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_2%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%VPWR N_VPWR_M1001_d N_VPWR_M1009_d
+ N_VPWR_c_272_n N_VPWR_c_273_n N_VPWR_c_274_n VPWR N_VPWR_c_275_n
+ N_VPWR_c_276_n N_VPWR_c_271_n PM_SKY130_FD_SC_HDLL__NOR3B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%A_309_297# N_A_309_297#_M1003_s
+ N_A_309_297#_M1000_s N_A_309_297#_M1013_s N_A_309_297#_c_327_n
+ N_A_309_297#_c_316_n N_A_309_297#_c_336_n N_A_309_297#_c_338_n
+ N_A_309_297#_c_317_n PM_SKY130_FD_SC_HDLL__NOR3B_2%A_309_297#
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%Y N_Y_M1006_d N_Y_M1007_s N_Y_M1005_s
+ N_Y_M1000_d N_Y_c_347_n N_Y_c_343_n N_Y_c_344_n N_Y_c_353_n N_Y_c_345_n
+ N_Y_c_359_n N_Y_c_346_n N_Y_c_372_n Y N_Y_c_375_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_2%Y
x_PM_SKY130_FD_SC_HDLL__NOR3B_2%VGND N_VGND_M1006_s N_VGND_M1012_s
+ N_VGND_M1011_d N_VGND_M1005_d N_VGND_M1008_d N_VGND_M1002_d N_VGND_c_411_n
+ N_VGND_c_412_n N_VGND_c_413_n N_VGND_c_414_n N_VGND_c_415_n N_VGND_c_416_n
+ N_VGND_c_417_n N_VGND_c_418_n N_VGND_c_419_n VGND N_VGND_c_420_n
+ N_VGND_c_421_n N_VGND_c_422_n N_VGND_c_423_n N_VGND_c_424_n
+ PM_SKY130_FD_SC_HDLL__NOR3B_2%VGND
cc_1 VNB N_A_c_65_n 0.0222857f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_66_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_3 VNB A 0.0163753f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_4 VNB N_A_c_68_n 0.0440201f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.202
cc_5 VNB N_B_c_102_n 0.0169338f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_6 VNB N_B_c_103_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=0.995
cc_7 VNB B 0.0096168f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_B_c_105_n 0.0426802f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_9 VNB N_A_571_21#_c_144_n 0.0215821f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_10 VNB N_A_571_21#_c_145_n 0.0198817f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_11 VNB N_A_571_21#_c_146_n 0.0108596f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.202
cc_12 VNB N_A_571_21#_c_147_n 0.00435791f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_571_21#_c_148_n 0.0133777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_571_21#_c_149_n 0.00241416f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_571_21#_c_150_n 4.69823e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_571_21#_c_151_n 0.0694535f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_C_N_c_206_n 0.021411f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_18 VNB N_C_N_c_207_n 0.0348547f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.41
cc_19 VNB C_N 0.0202773f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_20 VNB N_VPWR_c_271_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_Y_c_343_n 0.00355899f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_22 VNB N_Y_c_344_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_23 VNB N_Y_c_345_n 0.0262373f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_24 VNB N_Y_c_346_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_411_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.202
cc_26 VNB N_VGND_c_412_n 0.0335786f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.16
cc_27 VNB N_VGND_c_413_n 0.0199314f $X=-0.19 $Y=-0.24 $X2=1.01 $Y2=1.202
cc_28 VNB N_VGND_c_414_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_29 VNB N_VGND_c_415_n 0.00639354f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_416_n 0.0143182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_417_n 0.0348602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_418_n 0.0208833f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_419_n 0.00394313f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_420_n 0.0223166f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_421_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_422_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_423_n 0.0266115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_424_n 0.276615f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VPB N_A_c_69_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_40 VPB N_A_c_70_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_41 VPB N_A_c_68_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_42 VPB N_B_c_106_n 0.0161064f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_43 VPB N_B_c_107_n 0.0203249f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_44 VPB N_B_c_105_n 0.022695f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_45 VPB N_A_571_21#_c_152_n 0.0201936f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_46 VPB N_A_571_21#_c_153_n 0.0191031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_A_571_21#_c_154_n 0.00983079f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_A_571_21#_c_150_n 0.00394254f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A_571_21#_c_151_n 0.0345861f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_C_N_c_207_n 0.0368738f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_51 VPB N_A_27_297#_c_231_n 0.0103928f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.995
cc_52 VPB N_A_27_297#_c_232_n 0.0327764f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_53 VPB N_A_27_297#_c_233_n 0.0020765f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_54 VPB N_A_27_297#_c_234_n 0.00185169f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_55 VPB N_A_27_297#_c_235_n 0.00322557f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_56 VPB N_A_27_297#_c_236_n 0.0110427f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_VPWR_c_272_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.01 $Y2=0.56
cc_58 VPB N_VPWR_c_273_n 0.0147989f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_59 VPB N_VPWR_c_274_n 0.0486042f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_VPWR_c_275_n 0.0937623f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.202
cc_61 VPB N_VPWR_c_276_n 0.0238702f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.18
cc_62 VPB N_VPWR_c_271_n 0.0703905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_309_297#_c_316_n 0.0127436f $X=-0.19 $Y=1.305 $X2=0.66 $Y2=1.105
cc_64 VPB N_A_309_297#_c_317_n 0.00206719f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_65 N_A_c_66_n N_B_c_102_n 0.024264f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_66 N_A_c_70_n N_B_c_106_n 0.00985632f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_67 A B 0.0152605f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_68 N_A_c_68_n B 0.0018186f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_69 N_A_c_68_n N_B_c_105_n 0.024264f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_70 A N_A_27_297#_c_231_n 0.0252798f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_71 N_A_c_69_n N_A_27_297#_c_233_n 0.0158609f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_c_70_n N_A_27_297#_c_233_n 0.016363f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_73 A N_A_27_297#_c_233_n 0.0431894f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A_c_68_n N_A_27_297#_c_233_n 0.00794509f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_75 N_A_c_69_n N_VPWR_c_272_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_c_70_n N_VPWR_c_272_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_c_70_n N_VPWR_c_275_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_c_69_n N_VPWR_c_276_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_c_69_n N_VPWR_c_271_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_70_n N_VPWR_c_271_n 0.0124344f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_65_n N_Y_c_347_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_c_66_n N_Y_c_343_n 0.0114598f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_83 A N_Y_c_343_n 0.00695775f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A_c_65_n N_Y_c_344_n 0.00269085f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_85 A N_Y_c_344_n 0.030835f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_86 N_A_c_68_n N_Y_c_344_n 0.00486271f $X=0.985 $Y=1.202 $X2=0 $Y2=0
cc_87 N_A_c_66_n N_Y_c_353_n 5.32212e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_c_65_n N_VGND_c_412_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_89 A N_VGND_c_412_n 0.0217663f $X=0.66 $Y=1.105 $X2=0 $Y2=0
cc_90 N_A_c_65_n N_VGND_c_413_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_c_66_n N_VGND_c_413_n 0.00437852f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A_c_66_n N_VGND_c_414_n 0.00268723f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_65_n N_VGND_c_424_n 0.0107167f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_94 N_A_c_66_n N_VGND_c_424_n 0.00615622f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_95 B N_A_571_21#_c_151_n 0.00396852f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_96 N_B_c_106_n N_A_27_297#_c_234_n 0.0156202f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_107_n N_A_27_297#_c_234_n 0.0112811f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_98 B N_A_27_297#_c_234_n 0.0459115f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_99 N_B_c_105_n N_A_27_297#_c_234_n 0.00759056f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_100 B N_A_27_297#_c_235_n 0.00942636f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_101 N_B_c_106_n N_A_27_297#_c_236_n 5.04304e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_102 N_B_c_107_n N_A_27_297#_c_236_n 0.00739719f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_103 B N_A_27_297#_c_236_n 0.0171373f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_104 N_B_c_105_n N_A_27_297#_c_236_n 3.14831e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_105 N_B_c_106_n N_VPWR_c_275_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_c_107_n N_VPWR_c_275_n 0.00429453f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B_c_106_n N_VPWR_c_271_n 0.0126324f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B_c_107_n N_VPWR_c_271_n 0.00739666f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_109 N_B_c_107_n N_A_309_297#_c_316_n 0.0141207f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_110 N_B_c_102_n N_Y_c_343_n 0.00865686f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_111 B N_Y_c_343_n 0.0174927f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_112 N_B_c_102_n N_Y_c_353_n 0.00644736f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_113 N_B_c_103_n N_Y_c_345_n 0.01289f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_114 B N_Y_c_345_n 0.0252519f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_115 B N_Y_c_359_n 0.00634213f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_116 N_B_c_102_n N_Y_c_346_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 B N_Y_c_346_n 0.030835f $X=1.68 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B_c_105_n N_Y_c_346_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_119 N_B_c_102_n N_VGND_c_414_n 0.00268723f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_120 N_B_c_102_n N_VGND_c_422_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B_c_103_n N_VGND_c_422_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B_c_103_n N_VGND_c_423_n 0.00481673f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B_c_102_n N_VGND_c_424_n 0.00598581f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B_c_103_n N_VGND_c_424_n 0.00745263f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_125 N_A_571_21#_c_147_n N_C_N_c_206_n 0.00481607f $X=4.075 $Y=1.075 $X2=-0.19
+ $Y2=-0.24
cc_126 N_A_571_21#_c_148_n N_C_N_c_206_n 0.00356691f $X=4.22 $Y=0.66 $X2=-0.19
+ $Y2=-0.24
cc_127 N_A_571_21#_c_149_n N_C_N_c_207_n 8.89289e-19 $X=4.075 $Y=1.18 $X2=0
+ $Y2=0
cc_128 N_A_571_21#_c_154_n N_C_N_c_207_n 0.00184336f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_129 N_A_571_21#_c_150_n N_C_N_c_207_n 0.0053252f $X=4.167 $Y=1.455 $X2=0
+ $Y2=0
cc_130 N_A_571_21#_c_151_n N_C_N_c_207_n 0.00586563f $X=3.425 $Y=1.202 $X2=0
+ $Y2=0
cc_131 N_A_571_21#_c_148_n C_N 0.0011748f $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_132 N_A_571_21#_c_149_n C_N 0.0191447f $X=4.075 $Y=1.18 $X2=0 $Y2=0
cc_133 N_A_571_21#_c_154_n C_N 0.00115298f $X=4.22 $Y=1.705 $X2=0 $Y2=0
cc_134 N_A_571_21#_c_151_n C_N 4.54955e-19 $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_135 N_A_571_21#_c_152_n N_A_27_297#_c_236_n 0.00922102f $X=2.955 $Y=1.41
+ $X2=0 $Y2=0
cc_136 N_A_571_21#_c_152_n N_VPWR_c_275_n 0.00429453f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_137 N_A_571_21#_c_153_n N_VPWR_c_275_n 0.00429453f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_571_21#_c_152_n N_VPWR_c_271_n 0.00734734f $X=2.955 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_571_21#_c_153_n N_VPWR_c_271_n 0.00734734f $X=3.425 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_571_21#_c_154_n N_VPWR_c_271_n 0.0133729f $X=4.22 $Y=1.705 $X2=0
+ $Y2=0
cc_141 N_A_571_21#_c_152_n N_A_309_297#_c_316_n 0.0100504f $X=2.955 $Y=1.41
+ $X2=0 $Y2=0
cc_142 N_A_571_21#_c_153_n N_A_309_297#_c_316_n 0.0144985f $X=3.425 $Y=1.41
+ $X2=0 $Y2=0
cc_143 N_A_571_21#_c_153_n N_A_309_297#_c_317_n 7.2217e-19 $X=3.425 $Y=1.41
+ $X2=0 $Y2=0
cc_144 N_A_571_21#_c_146_n N_A_309_297#_c_317_n 0.0198783f $X=3.99 $Y=1.18 $X2=0
+ $Y2=0
cc_145 N_A_571_21#_c_154_n N_A_309_297#_c_317_n 0.0287258f $X=4.22 $Y=1.705
+ $X2=0 $Y2=0
cc_146 N_A_571_21#_c_151_n N_A_309_297#_c_317_n 0.0059411f $X=3.425 $Y=1.202
+ $X2=0 $Y2=0
cc_147 N_A_571_21#_c_144_n N_Y_c_345_n 0.00529831f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_148 N_A_571_21#_c_144_n N_Y_c_359_n 0.00593473f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_571_21#_c_152_n N_Y_c_359_n 0.0246629f $X=2.955 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_571_21#_c_145_n N_Y_c_359_n 0.003119f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_571_21#_c_153_n N_Y_c_359_n 0.0088412f $X=3.425 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_571_21#_c_146_n N_Y_c_359_n 0.0162029f $X=3.99 $Y=1.18 $X2=0 $Y2=0
cc_153 N_A_571_21#_c_147_n N_Y_c_359_n 0.00473951f $X=4.075 $Y=1.075 $X2=0 $Y2=0
cc_154 N_A_571_21#_c_150_n N_Y_c_359_n 0.00475909f $X=4.167 $Y=1.455 $X2=0 $Y2=0
cc_155 N_A_571_21#_c_151_n N_Y_c_359_n 0.0492924f $X=3.425 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_571_21#_c_144_n N_Y_c_372_n 0.00417236f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_157 N_A_571_21#_c_145_n N_Y_c_372_n 0.00257353f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_571_21#_c_148_n N_Y_c_372_n 3.08264e-19 $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_159 N_A_571_21#_c_144_n N_Y_c_375_n 0.0128481f $X=2.93 $Y=0.995 $X2=0 $Y2=0
cc_160 N_A_571_21#_c_145_n N_Y_c_375_n 0.00600712f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_161 N_A_571_21#_c_145_n N_VGND_c_415_n 0.00672154f $X=3.4 $Y=0.995 $X2=0
+ $Y2=0
cc_162 N_A_571_21#_c_146_n N_VGND_c_415_n 0.0159069f $X=3.99 $Y=1.18 $X2=0 $Y2=0
cc_163 N_A_571_21#_c_148_n N_VGND_c_415_n 0.0351615f $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_164 N_A_571_21#_c_151_n N_VGND_c_415_n 0.00518707f $X=3.425 $Y=1.202 $X2=0
+ $Y2=0
cc_165 N_A_571_21#_c_148_n N_VGND_c_417_n 0.0175451f $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_166 N_A_571_21#_c_144_n N_VGND_c_418_n 0.00401892f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_167 N_A_571_21#_c_145_n N_VGND_c_418_n 0.00541359f $X=3.4 $Y=0.995 $X2=0
+ $Y2=0
cc_168 N_A_571_21#_c_148_n N_VGND_c_420_n 0.0139405f $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_169 N_A_571_21#_c_144_n N_VGND_c_423_n 0.00599911f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_170 N_A_571_21#_c_144_n N_VGND_c_424_n 0.00704363f $X=2.93 $Y=0.995 $X2=0
+ $Y2=0
cc_171 N_A_571_21#_c_145_n N_VGND_c_424_n 0.0110773f $X=3.4 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_571_21#_c_148_n N_VGND_c_424_n 0.0126218f $X=4.22 $Y=0.66 $X2=0 $Y2=0
cc_173 N_C_N_c_207_n N_VPWR_c_274_n 0.0081971f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_174 C_N N_VPWR_c_274_n 0.0138817f $X=4.635 $Y=1.105 $X2=0 $Y2=0
cc_175 N_C_N_c_207_n N_VPWR_c_275_n 0.00393512f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_176 N_C_N_c_207_n N_VPWR_c_271_n 0.00500987f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_177 N_C_N_c_207_n N_A_309_297#_c_317_n 0.00413513f $X=4.455 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_C_N_c_206_n N_VGND_c_415_n 0.00172213f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_179 N_C_N_c_206_n N_VGND_c_417_n 0.00521921f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_180 N_C_N_c_207_n N_VGND_c_417_n 0.00280284f $X=4.455 $Y=1.41 $X2=0 $Y2=0
cc_181 C_N N_VGND_c_417_n 0.017914f $X=4.635 $Y=1.105 $X2=0 $Y2=0
cc_182 N_C_N_c_206_n N_VGND_c_420_n 0.00510437f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_183 N_C_N_c_206_n N_VGND_c_424_n 0.00512902f $X=4.43 $Y=0.995 $X2=0 $Y2=0
cc_184 N_A_27_297#_c_233_n N_VPWR_M1001_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_185 N_A_27_297#_c_233_n N_VPWR_c_272_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_186 N_A_27_297#_c_254_p N_VPWR_c_275_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_187 N_A_27_297#_c_232_n N_VPWR_c_276_n 0.0208166f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_188 N_A_27_297#_M1001_s N_VPWR_c_271_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_189 N_A_27_297#_M1010_s N_VPWR_c_271_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_27_297#_M1004_d N_VPWR_c_271_n 0.00234744f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_27_297#_c_232_n N_VPWR_c_271_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_192 N_A_27_297#_c_254_p N_VPWR_c_271_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_193 N_A_27_297#_c_234_n N_A_309_297#_M1003_s 0.00187091f $X=1.995 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_194 N_A_27_297#_c_234_n N_A_309_297#_c_327_n 0.0143018f $X=1.995 $Y=1.54
+ $X2=0 $Y2=0
cc_195 N_A_27_297#_M1004_d N_A_309_297#_c_316_n 0.00623749f $X=2.015 $Y=1.485
+ $X2=0 $Y2=0
cc_196 N_A_27_297#_c_234_n N_A_309_297#_c_316_n 0.00355499f $X=1.995 $Y=1.54
+ $X2=0 $Y2=0
cc_197 N_A_27_297#_c_236_n N_A_309_297#_c_316_n 0.0153216f $X=2.16 $Y=1.61 $X2=0
+ $Y2=0
cc_198 N_A_27_297#_c_233_n N_Y_c_343_n 0.00217122f $X=1.095 $Y=1.54 $X2=0 $Y2=0
cc_199 N_A_27_297#_c_235_n N_Y_c_343_n 0.00524452f $X=1.22 $Y=1.62 $X2=0 $Y2=0
cc_200 N_A_27_297#_c_236_n N_Y_c_345_n 0.00462221f $X=2.16 $Y=1.61 $X2=0 $Y2=0
cc_201 N_A_27_297#_c_236_n N_Y_c_359_n 0.0199903f $X=2.16 $Y=1.61 $X2=0 $Y2=0
cc_202 N_A_27_297#_c_231_n N_VGND_c_412_n 7.84254e-19 $X=0.247 $Y=1.625 $X2=0
+ $Y2=0
cc_203 N_VPWR_c_271_n N_A_309_297#_M1003_s 0.00297222f $X=4.83 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_204 N_VPWR_c_271_n N_A_309_297#_M1000_s 0.00233941f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_205 N_VPWR_c_271_n N_A_309_297#_M1013_s 0.00320704f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_206 N_VPWR_c_275_n N_A_309_297#_c_316_n 0.101366f $X=4.565 $Y=2.72 $X2=0
+ $Y2=0
cc_207 N_VPWR_c_271_n N_A_309_297#_c_316_n 0.0615382f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_208 N_VPWR_c_275_n N_A_309_297#_c_336_n 0.0149886f $X=4.565 $Y=2.72 $X2=0
+ $Y2=0
cc_209 N_VPWR_c_271_n N_A_309_297#_c_336_n 0.00962421f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_210 N_VPWR_c_275_n N_A_309_297#_c_338_n 0.0159047f $X=4.565 $Y=2.72 $X2=0
+ $Y2=0
cc_211 N_VPWR_c_271_n N_A_309_297#_c_338_n 0.00942493f $X=4.83 $Y=2.72 $X2=0
+ $Y2=0
cc_212 N_VPWR_c_271_n N_Y_M1000_d 0.00232895f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_213 N_A_309_297#_c_316_n N_Y_M1000_d 0.00380371f $X=3.535 $Y=2.37 $X2=0 $Y2=0
cc_214 N_A_309_297#_c_316_n N_Y_c_359_n 0.0209917f $X=3.535 $Y=2.37 $X2=0 $Y2=0
cc_215 N_A_309_297#_c_317_n N_Y_c_359_n 0.0235368f $X=3.66 $Y=1.62 $X2=0 $Y2=0
cc_216 N_Y_c_343_n N_VGND_M1012_s 0.00162089f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_217 N_Y_c_345_n N_VGND_M1011_d 0.00281828f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_218 N_Y_c_345_n N_VGND_M1005_d 0.00387807f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_219 N_Y_c_344_n N_VGND_c_412_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_220 N_Y_c_347_n N_VGND_c_413_n 0.0231806f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_221 N_Y_c_343_n N_VGND_c_413_n 0.00254521f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_222 N_Y_c_343_n N_VGND_c_414_n 0.0122559f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_223 N_Y_c_372_n N_VGND_c_415_n 0.0110997f $X=3.112 $Y=0.815 $X2=0 $Y2=0
cc_224 N_Y_c_375_n N_VGND_c_415_n 0.0293643f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_225 N_Y_c_345_n N_VGND_c_418_n 0.00110992f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_226 N_Y_c_372_n N_VGND_c_418_n 9.59101e-19 $X=3.112 $Y=0.815 $X2=0 $Y2=0
cc_227 N_Y_c_375_n N_VGND_c_418_n 0.0251471f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_228 N_Y_c_343_n N_VGND_c_422_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_229 N_Y_c_353_n N_VGND_c_422_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_230 N_Y_c_345_n N_VGND_c_422_n 0.00254521f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_231 N_Y_c_345_n N_VGND_c_423_n 0.0541915f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_232 N_Y_c_375_n N_VGND_c_423_n 0.025144f $X=3.19 $Y=0.39 $X2=0 $Y2=0
cc_233 N_Y_M1006_d N_VGND_c_424_n 0.00304143f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_234 N_Y_M1007_s N_VGND_c_424_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_235 N_Y_M1005_s N_VGND_c_424_n 0.0025535f $X=3.005 $Y=0.235 $X2=0 $Y2=0
cc_236 N_Y_c_347_n N_VGND_c_424_n 0.0143352f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_237 N_Y_c_343_n N_VGND_c_424_n 0.0094839f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_238 N_Y_c_353_n N_VGND_c_424_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_239 N_Y_c_345_n N_VGND_c_424_n 0.0102742f $X=2.87 $Y=0.815 $X2=0 $Y2=0
cc_240 N_Y_c_372_n N_VGND_c_424_n 0.00149581f $X=3.112 $Y=0.815 $X2=0 $Y2=0
cc_241 N_Y_c_375_n N_VGND_c_424_n 0.0155048f $X=3.19 $Y=0.39 $X2=0 $Y2=0
