* File: sky130_fd_sc_hdll__dlygate4sd1_1.pex.spice
* Created: Thu Aug 27 19:06:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A 3 7 9 10 18
c33 18 0 1.31538e-19 $X=0.52 $Y=1.16
r34 17 18 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=0.505 $Y=1.16
+ $X2=0.52 $Y2=1.16
r35 14 17 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=0.31 $Y=1.16
+ $X2=0.505 $Y2=1.16
r36 9 10 8.51056 $w=5.18e-07 $l=3.7e-07 $layer=LI1_cond $X=0.345 $Y=1.16
+ $X2=0.345 $Y2=1.53
r37 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.31
+ $Y=1.16 $X2=0.31 $Y2=1.16
r38 5 18 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r39 5 7 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r40 1 17 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=1.16
r41 1 3 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=0.505 $Y=1.325
+ $X2=0.505 $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_27_47# 1 2 9 13 17 21 23 24 25 26
+ 27 28 32
c71 32 0 3.81592e-20 $X=0.94 $Y=1.16
c72 27 0 1.89841e-19 $X=0.86 $Y=1.325
c73 25 0 1.31538e-19 $X=0.775 $Y=1.895
r74 32 35 40.7092 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=1.325
r75 32 34 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.16
+ $X2=0.965 $Y2=0.995
r76 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r77 29 31 18.0741 $w=2.43e-07 $l=3.6e-07 $layer=LI1_cond $X=0.927 $Y=0.8
+ $X2=0.927 $Y2=1.16
r78 27 31 9.39863 $w=2.43e-07 $l=1.95653e-07 $layer=LI1_cond $X=0.86 $Y=1.325
+ $X2=0.927 $Y2=1.16
r79 27 28 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.86 $Y=1.325
+ $X2=0.86 $Y2=1.785
r80 25 28 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.775 $Y=1.895
+ $X2=0.86 $Y2=1.785
r81 25 26 20.6916 $w=2.18e-07 $l=3.95e-07 $layer=LI1_cond $X=0.775 $Y=1.895
+ $X2=0.38 $Y2=1.895
r82 23 29 2.8297 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=0.775 $Y=0.8
+ $X2=0.927 $Y2=0.8
r83 23 24 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=0.775 $Y=0.8
+ $X2=0.38 $Y2=0.8
r84 19 24 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.38 $Y2=0.8
r85 19 21 8.2895 $w=2.83e-07 $l=2.05e-07 $layer=LI1_cond $X=0.237 $Y=0.715
+ $X2=0.237 $Y2=0.51
r86 15 26 7.00622 $w=2.2e-07 $l=1.95407e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.38 $Y2=1.895
r87 15 17 8.0085 $w=2.93e-07 $l=2.05e-07 $layer=LI1_cond $X=0.232 $Y=2.005
+ $X2=0.232 $Y2=2.21
r88 13 34 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.99 $Y=0.445
+ $X2=0.99 $Y2=0.995
r89 9 35 369.274 $w=1.8e-07 $l=9.5e-07 $layer=POLY_cond $X=0.975 $Y=2.275
+ $X2=0.975 $Y2=1.325
r90 2 17 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.21
r91 1 21 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_213_47# 1 2 7 9 10 12 14 16 19 25
+ 30 32 36
c63 36 0 1.89841e-19 $X=1.99 $Y=1.16
c64 19 0 1.94217e-19 $X=1.73 $Y=1.16
r65 35 36 2.62292 $w=3.3e-07 $l=1.5e-08 $layer=POLY_cond $X=1.975 $Y=1.16
+ $X2=1.99 $Y2=1.16
r66 28 30 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=2.32
+ $X2=1.335 $Y2=2.32
r67 23 25 5.36482 $w=2.88e-07 $l=1.35e-07 $layer=LI1_cond $X=1.2 $Y=0.4
+ $X2=1.335 $Y2=0.4
r68 20 35 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=1.73 $Y=1.16
+ $X2=1.975 $Y2=1.16
r69 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r70 17 32 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.42 $Y=1.175
+ $X2=1.335 $Y2=1.175
r71 17 19 17.1909 $w=1.98e-07 $l=3.1e-07 $layer=LI1_cond $X=1.42 $Y=1.175
+ $X2=1.73 $Y2=1.175
r72 16 30 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.335 $Y=2.175
+ $X2=1.335 $Y2=2.32
r73 15 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.335 $Y=1.275
+ $X2=1.335 $Y2=1.175
r74 15 16 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=1.335 $Y=1.275
+ $X2=1.335 $Y2=2.175
r75 14 32 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.335 $Y=1.075
+ $X2=1.335 $Y2=1.175
r76 13 25 3.86198 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=1.335 $Y=0.545
+ $X2=1.335 $Y2=0.4
r77 13 14 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=1.335 $Y=0.545
+ $X2=1.335 $Y2=1.075
r78 10 36 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=1.16
r79 10 12 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.99 $Y2=0.675
r80 7 35 16.9318 $w=1.8e-07 $l=1.65e-07 $layer=POLY_cond $X=1.975 $Y=1.325
+ $X2=1.975 $Y2=1.16
r81 7 9 157.989 $w=1.8e-07 $l=5.9e-07 $layer=POLY_cond $X=1.975 $Y=1.325
+ $X2=1.975 $Y2=1.915
r82 2 28 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=2.065 $X2=1.2 $Y2=2.34
r83 1 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%A_319_93# 1 2 9 13 16 19 21 22 23 24
+ 26 30 32
c65 30 0 3.88279e-19 $X=2.645 $Y=1.16
r66 30 33 40.7727 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.16
+ $X2=2.685 $Y2=1.325
r67 30 32 46.4315 $w=3.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.685 $Y=1.16
+ $X2=2.685 $Y2=0.995
r68 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.645
+ $Y=1.16 $X2=2.645 $Y2=1.16
r69 27 29 14.9747 $w=2.77e-07 $l=3.4e-07 $layer=LI1_cond $X=2.565 $Y=0.82
+ $X2=2.565 $Y2=1.16
r70 23 29 8.01 $w=2.77e-07 $l=1.92678e-07 $layer=LI1_cond $X=2.505 $Y=1.325
+ $X2=2.565 $Y2=1.16
r71 23 24 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=2.505 $Y=1.325
+ $X2=2.505 $Y2=1.575
r72 21 24 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.4 $Y=1.66
+ $X2=2.505 $Y2=1.575
r73 21 22 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.4 $Y=1.66 $X2=1.84
+ $Y2=1.66
r74 20 26 3.98913 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=1.84 $Y=0.82
+ $X2=1.727 $Y2=0.82
r75 19 27 3.59349 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.4 $Y=0.82
+ $X2=2.565 $Y2=0.82
r76 19 20 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.4 $Y=0.82 $X2=1.84
+ $Y2=0.82
r77 16 22 6.9898 $w=1.7e-07 $l=1.49579e-07 $layer=LI1_cond $X=1.727 $Y=1.745
+ $X2=1.84 $Y2=1.66
r78 16 18 5.69333 $w=2.25e-07 $l=1.05e-07 $layer=LI1_cond $X=1.727 $Y=1.745
+ $X2=1.727 $Y2=1.85
r79 13 32 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.735 $Y=0.56
+ $X2=2.735 $Y2=0.995
r80 9 33 256.548 $w=1.8e-07 $l=6.6e-07 $layer=POLY_cond $X=2.7 $Y=1.985 $X2=2.7
+ $Y2=1.325
r81 2 18 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.605
+ $Y=1.705 $X2=1.73 $Y2=1.85
r82 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.465 $X2=1.72 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
+ 42
r42 38 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 25 37 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=0.707 $Y2=2.72
r52 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 22 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r54 20 37 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.6 $Y=2.72
+ $X2=0.707 $Y2=2.72
r55 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=2.72 $X2=0.23
+ $Y2=2.72
r56 18 42 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 16 30 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 16 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.145 $Y=2.72
+ $X2=2.33 $Y2=2.72
r59 15 33 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 15 17 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.515 $Y=2.72
+ $X2=2.33 $Y2=2.72
r61 11 17 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.33 $Y=2.635
+ $X2=2.33 $Y2=2.72
r62 11 13 19.7784 $w=3.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.33 $Y=2.635
+ $X2=2.33 $Y2=2
r63 7 37 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=2.635
+ $X2=0.707 $Y2=2.72
r64 7 9 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.707 $Y=2.635
+ $X2=0.707 $Y2=2.34
r65 2 13 600 $w=1.7e-07 $l=4.06448e-07 $layer=licon1_PDIFF $count=1 $X=2.065
+ $Y=1.705 $X2=2.33 $Y2=2
r66 1 9 600 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_PDIFF $count=1 $X=0.595
+ $Y=2.065 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%X 1 2 10 11 12 13 14 15
r20 14 15 15.0704 $w=2.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.99 $Y=1.87
+ $X2=2.99 $Y2=2.21
r21 11 14 10.8596 $w=2.58e-07 $l=2.45e-07 $layer=LI1_cond $X=2.99 $Y=1.625
+ $X2=2.99 $Y2=1.87
r22 11 12 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.99 $Y=1.625
+ $X2=2.99 $Y2=1.495
r23 10 12 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.035 $Y=0.825
+ $X2=3.035 $Y2=1.495
r24 9 13 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.975 $Y=0.68
+ $X2=2.975 $Y2=0.51
r25 9 10 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=2.975 $Y=0.68
+ $X2=2.975 $Y2=0.825
r26 2 14 300 $w=1.7e-07 $l=4.55961e-07 $layer=licon1_PDIFF $count=2 $X=2.79
+ $Y=1.485 $X2=2.945 $Y2=1.87
r27 1 13 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=2.81
+ $Y=0.235 $X2=2.945 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLYGATE4SD1_1%VGND 1 2 9 13 16 17 18 20 33 34 37
+ 42
c47 13 0 1.94061e-19 $X=2.35 $Y=0.38
c48 9 0 3.81592e-20 $X=0.73 $Y=0.38
r49 38 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r50 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r52 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r53 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r54 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r55 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r56 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r57 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 25 37 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.707
+ $Y2=0
r59 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r60 22 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r61 20 37 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.707
+ $Y2=0
r62 20 22 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=0.6 $Y=0 $X2=0.23
+ $Y2=0
r63 18 42 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.225 $Y=0 $X2=0.23
+ $Y2=0
r64 16 30 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.07
+ $Y2=0
r65 16 17 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.145 $Y=0 $X2=2.35
+ $Y2=0
r66 15 33 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.99
+ $Y2=0
r67 15 17 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.555 $Y=0 $X2=2.35
+ $Y2=0
r68 11 17 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0
r69 11 13 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=2.35 $Y=0.085
+ $X2=2.35 $Y2=0.38
r70 7 37 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0
r71 7 9 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.707 $Y=0.085
+ $X2=0.707 $Y2=0.38
r72 2 13 182 $w=1.7e-07 $l=3.24731e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.465 $X2=2.35 $Y2=0.38
r73 1 9 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

