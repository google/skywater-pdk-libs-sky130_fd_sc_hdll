* File: sky130_fd_sc_hdll__sdfrtp_2.spice
* Created: Wed Sep  2 08:51:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfrtp_2.pex.spice"
.subckt sky130_fd_sc_hdll__sdfrtp_2  VNB VPB CLK D SCE SCD RESET_B VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* RESET_B	RESET_B
* SCD	SCD
* SCE	SCE
* D	D
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1027 N_VGND_M1027_d N_CLK_M1027_g N_A_27_47#_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1001 N_A_213_47#_M1001_d N_A_27_47#_M1001_g N_VGND_M1027_d VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1036 N_VGND_M1036_d N_SCE_M1036_g N_A_331_66#_M1036_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1092 AS=0.1302 PD=1.36 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1018 A_631_119# N_A_331_66#_M1018_g N_VGND_M1018_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0651 AS=0.1302 PD=0.73 PS=1.46 NRD=28.56 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1007 N_A_700_389#_M1007_d N_D_M1007_g A_631_119# VNB NSHORT L=0.15 W=0.42
+ AD=0.110275 AS=0.0651 PD=1.065 PS=0.73 NRD=0 NRS=28.56 M=1 R=2.8 SA=75000.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1031 A_899_66# N_SCE_M1031_g N_A_700_389#_M1007_d VNB NSHORT L=0.5 W=0.42
+ AD=0.0777 AS=0.110275 PD=0.79 PS=1.065 NRD=37.14 NRS=59.292 M=1 R=0.84
+ SA=250000 SB=250001 A=0.21 P=1.84 MULT=1
MM1034 N_VGND_M1034_d N_SCD_M1034_g A_899_66# VNB NSHORT L=0.18 W=0.42 AD=0.1197
+ AS=0.0777 PD=1.41 PS=0.79 NRD=0 NRS=37.14 M=1 R=2.33333 SA=90001.5 SB=90000.2
+ A=0.0756 P=1.2 MULT=1
MM1009 N_A_1202_413#_M1009_d N_A_27_47#_M1009_g N_A_700_389#_M1009_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.072 AS=0.1116 PD=0.76 PS=1.34 NRD=24.996 NRS=14.988 M=1
+ R=2.4 SA=75000.2 SB=75005.5 A=0.054 P=1.02 MULT=1
MM1033 A_1322_47# N_A_213_47#_M1033_g N_A_1202_413#_M1009_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0700615 AS=0.072 PD=0.738462 PS=0.76 NRD=46.536 NRS=14.988 M=1
+ R=2.4 SA=75000.8 SB=75004.9 A=0.054 P=1.02 MULT=1
MM1000 A_1428_47# N_A_1380_303#_M1000_g A_1322_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0546 AS=0.0817385 PD=0.68 PS=0.861538 NRD=21.42 NRS=39.888 M=1 R=2.8
+ SA=75001.2 SB=75003.9 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_RESET_B_M1020_g A_1428_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.127664 AS=0.0546 PD=0.990566 PS=0.68 NRD=47.136 NRS=21.42 M=1 R=2.8
+ SA=75001.6 SB=75003.5 A=0.063 P=1.14 MULT=1
MM1037 N_A_1380_303#_M1037_d N_A_1202_413#_M1037_g N_VGND_M1020_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.11968 AS=0.194536 PD=1.2352 PS=1.50943 NRD=0 NRS=30.936 M=1
+ R=4.26667 SA=75001.6 SB=75001.9 A=0.096 P=1.58 MULT=1
MM1025 N_A_1757_47#_M1025_d N_A_213_47#_M1025_g N_A_1380_303#_M1037_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0711 AS=0.06732 PD=0.755 PS=0.6948 NRD=6.66 NRS=16.656 M=1
+ R=2.4 SA=75003 SB=75002.7 A=0.054 P=1.02 MULT=1
MM1024 A_1866_47# N_A_27_47#_M1024_g N_A_1757_47#_M1025_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0978923 AS=0.0711 PD=0.876923 PS=0.755 NRD=72.3 NRS=31.656 M=1
+ R=2.4 SA=75003.5 SB=75002.2 A=0.054 P=1.02 MULT=1
MM1028 N_VGND_M1028_d N_A_1972_21#_M1028_g A_1866_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.13125 AS=0.114208 PD=1.045 PS=1.02308 NRD=12.852 NRS=61.968 M=1 R=2.8
+ SA=75003.6 SB=75001.5 A=0.063 P=1.14 MULT=1
MM1005 A_2157_47# N_RESET_B_M1005_g N_VGND_M1028_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.13125 PD=0.75 PS=1.045 NRD=31.428 NRS=85.704 M=1 R=2.8
+ SA=75004.4 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1011 N_A_1972_21#_M1011_d N_A_1757_47#_M1011_g A_2157_47# VNB NSHORT L=0.15
+ W=0.42 AD=0.1365 AS=0.0693 PD=1.49 PS=0.75 NRD=11.424 NRS=31.428 M=1 R=2.8
+ SA=75004.9 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1016 N_VGND_M1016_d N_A_1972_21#_M1016_g N_Q_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.299 AS=0.104 PD=2.22 PS=0.97 NRD=16.608 NRS=0 M=1 R=4.33333 SA=75000.4
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_A_1972_21#_M1019_g N_Q_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1013 N_VPWR_M1013_d N_CLK_M1013_g N_A_27_47#_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1525 AS=0.27 PD=1.305 PS=2.54 NRD=3.9203 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1029 N_A_213_47#_M1029_d N_A_27_47#_M1029_g N_VPWR_M1013_d VPB PHIGHVT L=0.18
+ W=1 AD=0.275 AS=0.1525 PD=2.55 PS=1.305 NRD=1.9503 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1026 N_VPWR_M1026_d N_SCE_M1026_g N_A_331_66#_M1026_s VPB PHIGHVT L=0.18
+ W=0.54 AD=0.0783 AS=0.2214 PD=0.83 PS=1.9 NRD=1.8124 NRS=1.8124 M=1 R=3
+ SA=90000.3 SB=90002.5 A=0.0972 P=1.44 MULT=1
MM1014 A_618_389# N_SCE_M1014_g N_VPWR_M1026_d VPB PHIGHVT L=0.18 W=0.54
+ AD=0.0621 AS=0.0783 PD=0.77 PS=0.83 NRD=21.8867 NRS=1.8124 M=1 R=3 SA=90000.8
+ SB=90002 A=0.0972 P=1.44 MULT=1
MM1017 N_A_700_389#_M1017_d N_D_M1017_g A_618_389# VPB PHIGHVT L=0.18 W=0.54
+ AD=0.1809 AS=0.0621 PD=1.21 PS=0.77 NRD=114.91 NRS=21.8867 M=1 R=3 SA=90001.2
+ SB=90001.6 A=0.0972 P=1.44 MULT=1
MM1035 A_870_389# N_A_331_66#_M1035_g N_A_700_389#_M1017_d VPB PHIGHVT L=0.18
+ W=0.54 AD=0.09855 AS=0.1809 PD=0.905 PS=1.21 NRD=46.5117 NRS=27.3436 M=1 R=3
+ SA=90002 SB=90000.7 A=0.0972 P=1.44 MULT=1
MM1006 N_VPWR_M1006_d N_SCD_M1006_g A_870_389# VPB PHIGHVT L=0.18 W=0.54
+ AD=0.1566 AS=0.09855 PD=1.66 PS=0.905 NRD=1.8124 NRS=46.5117 M=1 R=3
+ SA=90002.6 SB=90000.2 A=0.0972 P=1.44 MULT=1
MM1022 N_A_1202_413#_M1022_d N_A_213_47#_M1022_g N_A_700_389#_M1022_s VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0903 AS=0.1575 PD=0.85 PS=1.59 NRD=68.0044
+ NRS=2.3443 M=1 R=2.33333 SA=90000.3 SB=90001.9 A=0.0756 P=1.2 MULT=1
MM1023 N_A_1324_413#_M1023_d N_A_27_47#_M1023_g N_A_1202_413#_M1022_d VPB
+ PHIGHVT L=0.18 W=0.42 AD=0.0609 AS=0.0903 PD=0.71 PS=0.85 NRD=2.3443
+ NRS=2.3443 M=1 R=2.33333 SA=90000.9 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1012 N_VPWR_M1012_d N_A_1380_303#_M1012_g N_A_1324_413#_M1023_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1049 AS=0.0609 PD=0.96 PS=0.71 NRD=35.1645 NRS=2.3443 M=1
+ R=2.33333 SA=90001.4 SB=90000.8 A=0.0756 P=1.2 MULT=1
MM1021 N_A_1324_413#_M1021_d N_RESET_B_M1021_g N_VPWR_M1012_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.1049 PD=1.38 PS=0.96 NRD=2.3443 NRS=44.5417 M=1
+ R=2.33333 SA=90002 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1008 N_A_1380_303#_M1008_d N_A_1202_413#_M1008_g N_VPWR_M1008_s VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.1694 AS=0.2688 PD=1.58 PS=2.32 NRD=2.3443 NRS=1.1623 M=1
+ R=4.66667 SA=90000.2 SB=90001.5 A=0.1512 P=2.04 MULT=1
MM1032 N_A_1757_47#_M1032_d N_A_27_47#_M1032_g N_A_1380_303#_M1008_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.063 AS=0.0847 PD=0.72 PS=0.79 NRD=7.0329 NRS=25.7873 M=1
+ R=2.33333 SA=90000.8 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1015 A_1951_413# N_A_213_47#_M1015_g N_A_1757_47#_M1032_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0693 AS=0.063 PD=0.75 PS=0.72 NRD=51.5943 NRS=2.3443 M=1 R=2.33333
+ SA=90001.2 SB=90001.7 A=0.0756 P=1.2 MULT=1
MM1003 N_VPWR_M1003_d N_A_1972_21#_M1003_g A_1951_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0798 AS=0.0693 PD=0.8 PS=0.75 NRD=44.5417 NRS=51.5943 M=1 R=2.33333
+ SA=90001.7 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1004 N_A_1972_21#_M1004_d N_RESET_B_M1004_g N_VPWR_M1003_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0672 AS=0.0798 PD=0.74 PS=0.8 NRD=14.0658 NRS=2.3443 M=1 R=2.33333
+ SA=90002.3 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1757_47#_M1010_g N_A_1972_21#_M1004_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.1134 AS=0.0672 PD=1.38 PS=0.74 NRD=2.3443 NRS=4.6886 M=1
+ R=2.33333 SA=90002.8 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1002 N_Q_M1002_d N_A_1972_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.42 PD=1.29 PS=2.84 NRD=0.9653 NRS=9.8303 M=1 R=5.55556
+ SA=90000.3 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1030 N_Q_M1002_d N_A_1972_21#_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.8 SB=90000.2 A=0.18 P=2.36 MULT=1
DX38_noxref VNB VPB NWDIODE A=21.7404 P=30.89
c_246 VPB 0 2.92951e-19 $X=0.17 $Y=2.64
*
.include "sky130_fd_sc_hdll__sdfrtp_2.pxi.spice"
*
.ends
*
*
