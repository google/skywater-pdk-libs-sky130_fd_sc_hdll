* File: sky130_fd_sc_hdll__muxb16to1_4.spice
* Created: Wed Sep  2 08:35:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb16to1_4.pex.spice"
.subckt sky130_fd_sc_hdll__muxb16to1_4  VNB VPB D[0] D[8] S[0] S[8] S[1] S[9]
+ D[1] D[9] D[2] D[10] S[2] S[10] S[3] S[11] D[3] D[11] D[4] D[12] S[4] S[12]
+ S[5] S[13] D[5] D[13] D[6] D[14] S[6] S[14] S[7] S[15] D[7] D[15] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[15]	D[15]
* D[7]	D[7]
* S[15]	S[15]
* S[7]	S[7]
* S[14]	S[14]
* S[6]	S[6]
* D[14]	D[14]
* D[6]	D[6]
* D[13]	D[13]
* D[5]	D[5]
* S[13]	S[13]
* S[5]	S[5]
* S[12]	S[12]
* S[4]	S[4]
* D[12]	D[12]
* D[4]	D[4]
* D[11]	D[11]
* D[3]	D[3]
* S[11]	S[11]
* S[3]	S[3]
* S[10]	S[10]
* S[2]	S[2]
* D[10]	D[10]
* D[2]	D[2]
* D[9]	D[9]
* D[1]	D[1]
* S[9]	S[9]
* S[1]	S[1]
* S[8]	S[8]
* S[0]	S[0]
* D[8]	D[8]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1084 N_VGND_M1084_d N_D[0]_M1084_g N_A_119_47#_M1084_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1085 N_VGND_M1085_d N_D[8]_M1085_g N_A_119_911#_M1085_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1219 N_VGND_M1219_d N_D[0]_M1219_g N_A_119_47#_M1084_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1090 N_VGND_M1090_d N_D[8]_M1090_g N_A_119_911#_M1085_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1300 N_VGND_M1219_d N_D[0]_M1300_g N_A_119_47#_M1300_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1235 N_VGND_M1090_d N_D[8]_M1235_g N_A_119_911#_M1235_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1317 N_VGND_M1317_d N_D[0]_M1317_g N_A_119_47#_M1300_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1240 N_VGND_M1240_d N_D[8]_M1240_g N_A_119_911#_M1235_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1053 N_A_119_47#_M1053_d N_S[0]_M1053_g N_Z_M1053_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1070 N_Z_M1070_d N_S[8]_M1070_g N_A_119_911#_M1070_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1074 N_A_119_47#_M1074_d N_S[0]_M1074_g N_Z_M1053_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1159 N_Z_M1070_d N_S[8]_M1159_g N_A_119_911#_M1159_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1105 N_A_119_47#_M1074_d N_S[0]_M1105_g N_Z_M1105_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1236 N_Z_M1236_d N_S[8]_M1236_g N_A_119_911#_M1159_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1125 N_A_119_47#_M1125_d N_S[0]_M1125_g N_Z_M1105_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1302 N_Z_M1236_d N_S[8]_M1302_g N_A_119_911#_M1302_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1139 N_A_559_265#_M1139_d N_S[0]_M1139_g N_VGND_M1139_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1017 N_A_559_793#_M1017_d N_S[8]_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1192 N_A_559_265#_M1139_d N_S[0]_M1192_g N_VGND_M1192_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1078 N_A_559_793#_M1017_d N_S[8]_M1078_g N_VGND_M1078_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1241 N_VGND_M1241_d N_S[1]_M1241_g N_A_1430_325#_M1241_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1008 N_A_1430_599#_M1008_d N_S[9]_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1288 N_VGND_M1288_d N_S[1]_M1288_g N_A_1430_325#_M1241_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1107 N_A_1430_599#_M1008_d N_S[9]_M1107_g N_VGND_M1107_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1039 N_Z_M1039_d N_S[1]_M1039_g N_A_1693_66#_M1039_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1027 N_Z_M1027_d N_S[9]_M1027_g N_A_1693_918#_M1027_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1045 N_Z_M1039_d N_S[1]_M1045_g N_A_1693_66#_M1045_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1032 N_Z_M1027_d N_S[9]_M1032_g N_A_1693_918#_M1032_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1093 N_Z_M1093_d N_S[1]_M1093_g N_A_1693_66#_M1045_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1096 N_Z_M1096_d N_S[9]_M1096_g N_A_1693_918#_M1032_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1113 N_Z_M1093_d N_S[1]_M1113_g N_A_1693_66#_M1113_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1259 N_Z_M1096_d N_S[9]_M1259_g N_A_1693_918#_M1259_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1049 N_VGND_M1049_d N_D[1]_M1049_g N_A_1693_66#_M1049_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1019_d N_D[9]_M1019_g N_A_1693_918#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1098 N_VGND_M1098_d N_D[1]_M1098_g N_A_1693_66#_M1049_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1111 N_VGND_M1111_d N_D[9]_M1111_g N_A_1693_918#_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1167 N_VGND_M1098_d N_D[1]_M1167_g N_A_1693_66#_M1167_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1178 N_VGND_M1111_d N_D[9]_M1178_g N_A_1693_918#_M1178_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1315 N_VGND_M1315_d N_D[1]_M1315_g N_A_1693_66#_M1167_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1276 N_VGND_M1276_d N_D[9]_M1276_g N_A_1693_918#_M1178_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_2695_47#_M1001_d N_D[2]_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1033 N_VGND_M1033_d N_D[10]_M1033_g N_A_2695_911#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1062 N_A_2695_47#_M1001_d N_D[2]_M1062_g N_VGND_M1062_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1143 N_VGND_M1143_d N_D[10]_M1143_g N_A_2695_911#_M1033_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1110 N_A_2695_47#_M1110_d N_D[2]_M1110_g N_VGND_M1062_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1195 N_VGND_M1143_d N_D[10]_M1195_g N_A_2695_911#_M1195_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1182 N_A_2695_47#_M1110_d N_D[2]_M1182_g N_VGND_M1182_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1307 N_VGND_M1307_d N_D[10]_M1307_g N_A_2695_911#_M1195_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1035 N_Z_M1035_d N_S[2]_M1035_g N_A_2695_47#_M1035_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1010 N_A_2695_911#_M1010_d N_S[10]_M1010_g N_Z_M1010_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1036 N_Z_M1035_d N_S[2]_M1036_g N_A_2695_47#_M1036_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1214 N_A_2695_911#_M1214_d N_S[10]_M1214_g N_Z_M1010_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1108 N_Z_M1108_d N_S[2]_M1108_g N_A_2695_47#_M1036_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1263 N_A_2695_911#_M1214_d N_S[10]_M1263_g N_Z_M1263_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1306 N_Z_M1108_d N_S[2]_M1306_g N_A_2695_47#_M1306_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1268 N_A_2695_911#_M1268_d N_S[10]_M1268_g N_Z_M1263_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1222 N_VGND_M1222_d N_S[2]_M1222_g N_A_3135_265#_M1222_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1043 N_A_3135_793#_M1043_d N_S[10]_M1043_g N_VGND_M1043_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1239 N_VGND_M1239_d N_S[2]_M1239_g N_A_3135_265#_M1222_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1215 N_A_3135_793#_M1043_d N_S[10]_M1215_g N_VGND_M1215_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1234 N_VGND_M1234_d N_S[3]_M1234_g N_A_4006_325#_M1234_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1054 N_VGND_M1054_d N_S[11]_M1054_g N_A_4006_599#_M1054_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1291 N_VGND_M1291_d N_S[3]_M1291_g N_A_4006_325#_M1234_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1072 N_VGND_M1072_d N_S[11]_M1072_g N_A_4006_599#_M1054_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1030 N_A_4269_66#_M1030_d N_S[3]_M1030_g N_Z_M1030_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1047 N_A_4269_918#_M1047_d N_S[11]_M1047_g N_Z_M1047_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1031 N_A_4269_66#_M1031_d N_S[3]_M1031_g N_Z_M1030_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1160 N_A_4269_918#_M1160_d N_S[11]_M1160_g N_Z_M1047_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1059 N_A_4269_66#_M1031_d N_S[3]_M1059_g N_Z_M1059_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1316 N_A_4269_918#_M1160_d N_S[11]_M1316_g N_Z_M1316_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1106 N_A_4269_66#_M1106_d N_S[3]_M1106_g N_Z_M1059_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1318 N_A_4269_918#_M1318_d N_S[11]_M1318_g N_Z_M1316_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1041 N_VGND_M1041_d N_D[3]_M1041_g N_A_4269_66#_M1041_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1245 N_A_4269_918#_M1245_d N_D[11]_M1245_g N_VGND_M1245_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1100 N_VGND_M1100_d N_D[3]_M1100_g N_A_4269_66#_M1041_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1296 N_A_4269_918#_M1245_d N_D[11]_M1296_g N_VGND_M1296_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1135 N_VGND_M1100_d N_D[3]_M1135_g N_A_4269_66#_M1135_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1310 N_A_4269_918#_M1310_d N_D[11]_M1310_g N_VGND_M1296_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1193 N_VGND_M1193_d N_D[3]_M1193_g N_A_4269_66#_M1135_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1311 N_A_4269_918#_M1310_d N_D[11]_M1311_g N_VGND_M1311_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1021 N_VGND_M1021_d N_D[4]_M1021_g N_A_5363_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_D[12]_M1012_g N_A_5363_911#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1177 N_VGND_M1177_d N_D[4]_M1177_g N_A_5363_47#_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1128 N_VGND_M1128_d N_D[12]_M1128_g N_A_5363_911#_M1012_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1232 N_VGND_M1177_d N_D[4]_M1232_g N_A_5363_47#_M1232_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1187 N_VGND_M1128_d N_D[12]_M1187_g N_A_5363_911#_M1187_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1275 N_VGND_M1275_d N_D[4]_M1275_g N_A_5363_47#_M1232_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1267 N_VGND_M1267_d N_D[12]_M1267_g N_A_5363_911#_M1187_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1154 N_Z_M1154_d N_S[4]_M1154_g N_A_5363_47#_M1154_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1044 N_A_5363_911#_M1044_d N_S[12]_M1044_g N_Z_M1044_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1191 N_Z_M1154_d N_S[4]_M1191_g N_A_5363_47#_M1191_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1091 N_A_5363_911#_M1091_d N_S[12]_M1091_g N_Z_M1044_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1205 N_Z_M1205_d N_S[4]_M1205_g N_A_5363_47#_M1191_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1218 N_A_5363_911#_M1091_d N_S[12]_M1218_g N_Z_M1218_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1213 N_Z_M1205_d N_S[4]_M1213_g N_A_5363_47#_M1213_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1312 N_A_5363_911#_M1312_d N_S[12]_M1312_g N_Z_M1218_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1037 N_VGND_M1037_d N_S[4]_M1037_g N_A_5803_265#_M1037_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1188 N_A_5803_793#_M1188_d N_S[12]_M1188_g N_VGND_M1188_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1086 N_VGND_M1086_d N_S[4]_M1086_g N_A_5803_265#_M1037_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1283 N_A_5803_793#_M1188_d N_S[12]_M1283_g N_VGND_M1283_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1126 N_VGND_M1126_d N_S[5]_M1126_g N_A_6674_325#_M1126_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1060 N_VGND_M1060_d N_S[13]_M1060_g N_A_6674_599#_M1060_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1152 N_VGND_M1152_d N_S[5]_M1152_g N_A_6674_325#_M1126_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1211 N_VGND_M1211_d N_S[13]_M1211_g N_A_6674_599#_M1060_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1175 N_A_6937_66#_M1175_d N_S[5]_M1175_g N_Z_M1175_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1149 N_A_6937_918#_M1149_d N_S[13]_M1149_g N_Z_M1149_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1210 N_A_6937_66#_M1210_d N_S[5]_M1210_g N_Z_M1175_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1226 N_A_6937_918#_M1226_d N_S[13]_M1226_g N_Z_M1149_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1220 N_A_6937_66#_M1210_d N_S[5]_M1220_g N_Z_M1220_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1242 N_A_6937_918#_M1226_d N_S[13]_M1242_g N_Z_M1242_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1228 N_A_6937_66#_M1228_d N_S[5]_M1228_g N_Z_M1220_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1290 N_A_6937_918#_M1290_d N_S[13]_M1290_g N_Z_M1242_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1029 N_VGND_M1029_d N_D[5]_M1029_g N_A_6937_66#_M1029_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1132 N_VGND_M1132_d N_D[13]_M1132_g N_A_6937_918#_M1132_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1057 N_VGND_M1057_d N_D[5]_M1057_g N_A_6937_66#_M1029_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1136 N_VGND_M1136_d N_D[13]_M1136_g N_A_6937_918#_M1132_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1247 N_VGND_M1057_d N_D[5]_M1247_g N_A_6937_66#_M1247_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1274 N_VGND_M1136_d N_D[13]_M1274_g N_A_6937_918#_M1274_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1262 N_VGND_M1262_d N_D[5]_M1262_g N_A_6937_66#_M1247_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1298 N_VGND_M1298_d N_D[13]_M1298_g N_A_6937_918#_M1274_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1069 N_A_7939_47#_M1069_d N_D[6]_M1069_g N_VGND_M1069_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1004 N_A_7939_911#_M1004_d N_D[14]_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1122 N_A_7939_47#_M1069_d N_D[6]_M1122_g N_VGND_M1122_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1179 N_A_7939_911#_M1004_d N_D[14]_M1179_g N_VGND_M1179_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1147 N_A_7939_47#_M1147_d N_D[6]_M1147_g N_VGND_M1122_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1189 N_A_7939_911#_M1189_d N_D[14]_M1189_g N_VGND_M1179_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1258 N_A_7939_47#_M1147_d N_D[6]_M1258_g N_VGND_M1258_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1305 N_A_7939_911#_M1189_d N_D[14]_M1305_g N_VGND_M1305_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1202 N_A_7939_47#_M1202_d N_S[6]_M1202_g N_Z_M1202_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1005 N_A_7939_911#_M1005_d N_S[14]_M1005_g N_Z_M1005_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1212 N_A_7939_47#_M1212_d N_S[6]_M1212_g N_Z_M1202_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1064 N_A_7939_911#_M1064_d N_S[14]_M1064_g N_Z_M1005_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1244 N_A_7939_47#_M1212_d N_S[6]_M1244_g N_Z_M1244_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1162 N_A_7939_911#_M1064_d N_S[14]_M1162_g N_Z_M1162_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1254 N_A_7939_47#_M1254_d N_S[6]_M1254_g N_Z_M1244_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1230 N_A_7939_911#_M1230_d N_S[14]_M1230_g N_Z_M1162_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1009 N_A_8379_265#_M1009_d N_S[6]_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1028 N_A_8379_793#_M1028_d N_S[14]_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1075 N_A_8379_265#_M1009_d N_S[6]_M1075_g N_VGND_M1075_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1097 N_A_8379_793#_M1028_d N_S[14]_M1097_g N_VGND_M1097_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1141 N_A_9250_325#_M1141_d N_S[7]_M1141_g N_VGND_M1141_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1174 N_A_9250_599#_M1174_d N_S[15]_M1174_g N_VGND_M1174_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1198 N_A_9250_325#_M1141_d N_S[7]_M1198_g N_VGND_M1198_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1223 N_A_9250_599#_M1174_d N_S[15]_M1223_g N_VGND_M1223_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_A_9513_66#_M1003_d N_S[7]_M1003_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1104 N_Z_M1104_d N_S[15]_M1104_g N_A_9513_918#_M1104_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.4 A=0.078 P=1.34 MULT=1
MM1209 N_A_9513_66#_M1209_d N_S[7]_M1209_g N_Z_M1003_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1169 N_Z_M1104_d N_S[15]_M1169_g N_A_9513_918#_M1169_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001 A=0.078 P=1.34 MULT=1
MM1253 N_A_9513_66#_M1209_d N_S[7]_M1253_g N_Z_M1253_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1197 N_Z_M1197_d N_S[15]_M1197_g N_A_9513_918#_M1169_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1272 N_A_9513_66#_M1272_d N_S[7]_M1272_g N_Z_M1253_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1252 N_Z_M1197_d N_S[15]_M1252_g N_A_9513_918#_M1252_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.4 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1068 N_VGND_M1068_d N_D[7]_M1068_g N_A_9513_66#_M1068_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1073 N_A_9513_918#_M1073_d N_D[15]_M1073_g N_VGND_M1073_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1115 N_VGND_M1115_d N_D[7]_M1115_g N_A_9513_66#_M1068_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1144 N_A_9513_918#_M1073_d N_D[15]_M1144_g N_VGND_M1144_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1216 N_VGND_M1115_d N_D[7]_M1216_g N_A_9513_66#_M1216_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1190 N_A_9513_918#_M1190_d N_D[15]_M1190_g N_VGND_M1144_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1281 N_VGND_M1281_d N_D[7]_M1281_g N_A_9513_66#_M1216_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1278 N_A_9513_918#_M1190_d N_D[15]_M1278_g N_VGND_M1278_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1014 N_VPWR_M1014_d N_D[0]_M1014_g N_A_117_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1023_d N_D[8]_M1023_g N_A_117_591#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1146 N_VPWR_M1146_d N_D[0]_M1146_g N_A_117_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1155 N_VPWR_M1155_d N_D[8]_M1155_g N_A_117_591#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1208 N_VPWR_M1146_d N_D[0]_M1208_g N_A_117_297#_M1208_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1221 N_VPWR_M1155_d N_D[8]_M1221_g N_A_117_591#_M1221_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1294 N_VPWR_M1294_d N_D[0]_M1294_g N_A_117_297#_M1208_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1304 N_VPWR_M1304_d N_D[8]_M1304_g N_A_117_591#_M1221_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1137 N_A_117_297#_M1137_d N_A_559_265#_M1137_g N_Z_M1137_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1026 N_Z_M1026_d N_A_559_793#_M1026_g N_A_117_591#_M1026_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1207 N_A_117_297#_M1207_d N_A_559_265#_M1207_g N_Z_M1137_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1079 N_Z_M1026_d N_A_559_793#_M1079_g N_A_117_591#_M1079_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1249 N_A_117_297#_M1207_d N_A_559_265#_M1249_g N_Z_M1249_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1127 N_Z_M1127_d N_A_559_793#_M1127_g N_A_117_591#_M1079_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1299 N_A_117_297#_M1299_d N_A_559_265#_M1299_g N_Z_M1249_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1269 N_Z_M1127_d N_A_559_793#_M1269_g N_A_117_591#_M1269_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1018 N_VPWR_M1018_d N_S[0]_M1018_g N_A_559_265#_M1018_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1123 N_VPWR_M1123_d N_S[8]_M1123_g N_A_559_793#_M1123_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1061 N_VPWR_M1061_d N_S[0]_M1061_g N_A_559_265#_M1018_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1172 N_VPWR_M1172_d N_S[8]_M1172_g N_A_559_793#_M1123_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1133 N_VPWR_M1133_d N_S[1]_M1133_g N_A_1430_325#_M1133_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1225 N_VPWR_M1225_d N_S[9]_M1225_g N_A_1430_599#_M1225_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1180 N_VPWR_M1180_d N_S[1]_M1180_g N_A_1430_325#_M1133_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1266 N_VPWR_M1266_d N_S[9]_M1266_g N_A_1430_599#_M1225_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1007 N_Z_M1007_d N_A_1430_325#_M1007_g N_A_1643_311#_M1007_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1112 N_A_1643_613#_M1112_d N_A_1430_599#_M1112_g N_Z_M1112_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1048 N_Z_M1007_d N_A_1430_325#_M1048_g N_A_1643_311#_M1048_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1161 N_A_1643_613#_M1161_d N_A_1430_599#_M1161_g N_Z_M1112_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1140 N_Z_M1140_d N_A_1430_325#_M1140_g N_A_1643_311#_M1048_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1199 N_A_1643_613#_M1161_d N_A_1430_599#_M1199_g N_Z_M1199_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1284 N_Z_M1140_d N_A_1430_325#_M1284_g N_A_1643_311#_M1284_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1273 N_A_1643_613#_M1273_d N_A_1430_599#_M1273_g N_Z_M1199_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1002 N_A_1643_311#_M1002_d N_D[1]_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_A_1643_613#_M1011_d N_D[9]_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1038 N_A_1643_311#_M1002_d N_D[1]_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1051 N_A_1643_613#_M1011_d N_D[9]_M1051_g N_VPWR_M1051_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1134 N_A_1643_311#_M1134_d N_D[1]_M1134_g N_VPWR_M1038_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1148 N_A_1643_613#_M1148_d N_D[9]_M1148_g N_VPWR_M1051_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1271 N_A_1643_311#_M1134_d N_D[1]_M1271_g N_VPWR_M1271_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1285 N_A_1643_613#_M1148_d N_D[9]_M1285_g N_VPWR_M1285_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1020 N_A_2693_297#_M1020_d N_D[2]_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1024 N_A_2693_591#_M1024_d N_D[10]_M1024_g N_VPWR_M1024_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1067 N_A_2693_297#_M1020_d N_D[2]_M1067_g N_VPWR_M1067_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1076 N_A_2693_591#_M1024_d N_D[10]_M1076_g N_VPWR_M1076_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1157 N_A_2693_297#_M1157_d N_D[2]_M1157_g N_VPWR_M1067_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1164 N_A_2693_591#_M1164_d N_D[10]_M1164_g N_VPWR_M1076_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1301 N_A_2693_297#_M1157_d N_D[2]_M1301_g N_VPWR_M1301_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1309 N_A_2693_591#_M1164_d N_D[10]_M1309_g N_VPWR_M1309_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1082 N_A_2693_297#_M1082_d N_A_3135_265#_M1082_g N_Z_M1082_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1000 N_A_2693_591#_M1000_d N_A_3135_793#_M1000_g N_Z_M1000_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1138 N_A_2693_297#_M1138_d N_A_3135_265#_M1138_g N_Z_M1082_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1080 N_A_2693_591#_M1080_d N_A_3135_793#_M1080_g N_Z_M1000_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1181 N_A_2693_297#_M1138_d N_A_3135_265#_M1181_g N_Z_M1181_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1229 N_A_2693_591#_M1080_d N_A_3135_793#_M1229_g N_Z_M1229_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1250 N_A_2693_297#_M1250_d N_A_3135_265#_M1250_g N_Z_M1181_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1270 N_A_2693_591#_M1270_d N_A_3135_793#_M1270_g N_Z_M1229_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1065 N_A_3135_265#_M1065_d N_S[2]_M1065_g N_VPWR_M1065_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1083 N_VPWR_M1083_d N_S[10]_M1083_g N_A_3135_793#_M1083_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1308 N_A_3135_265#_M1065_d N_S[2]_M1308_g N_VPWR_M1308_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1173 N_VPWR_M1173_d N_S[10]_M1173_g N_A_3135_793#_M1083_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1150 N_A_4006_325#_M1150_d N_S[3]_M1150_g N_VPWR_M1150_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1066 N_VPWR_M1066_d N_S[11]_M1066_g N_A_4006_599#_M1066_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1280 N_A_4006_325#_M1150_d N_S[3]_M1280_g N_VPWR_M1280_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1237 N_VPWR_M1237_d N_S[11]_M1237_g N_A_4006_599#_M1066_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1121 N_A_4219_311#_M1121_d N_A_4006_325#_M1121_g N_Z_M1121_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1071 N_A_4219_613#_M1071_d N_A_4006_599#_M1071_g N_Z_M1071_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1171 N_A_4219_311#_M1171_d N_A_4006_325#_M1171_g N_Z_M1121_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1114 N_A_4219_613#_M1114_d N_A_4006_599#_M1114_g N_Z_M1071_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1243 N_A_4219_311#_M1171_d N_A_4006_325#_M1243_g N_Z_M1243_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1260 N_A_4219_613#_M1114_d N_A_4006_599#_M1260_g N_Z_M1260_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1287 N_A_4219_311#_M1287_d N_A_4006_325#_M1287_g N_Z_M1243_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1313 N_A_4219_613#_M1313_d N_A_4006_599#_M1313_g N_Z_M1260_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1042 N_VPWR_M1042_d N_D[3]_M1042_g N_A_4219_311#_M1042_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1052 N_VPWR_M1052_d N_D[11]_M1052_g N_A_4219_613#_M1052_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1089 N_VPWR_M1089_d N_D[3]_M1089_g N_A_4219_311#_M1042_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1101 N_VPWR_M1101_d N_D[11]_M1101_g N_A_4219_613#_M1052_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1116 N_VPWR_M1089_d N_D[3]_M1116_g N_A_4219_311#_M1116_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1129 N_VPWR_M1101_d N_D[11]_M1129_g N_A_4219_613#_M1129_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1289 N_VPWR_M1289_d N_D[3]_M1289_g N_A_4219_311#_M1116_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1297 N_VPWR_M1297_d N_D[11]_M1297_g N_A_4219_613#_M1129_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1158 N_VPWR_M1158_d N_D[4]_M1158_g N_A_5361_297#_M1158_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_5361_591#_M1006_d N_D[12]_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1194 N_VPWR_M1194_d N_D[4]_M1194_g N_A_5361_297#_M1158_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1165 N_A_5361_591#_M1006_d N_D[12]_M1165_g N_VPWR_M1165_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1265 N_VPWR_M1194_d N_D[4]_M1265_g N_A_5361_297#_M1265_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1203 N_A_5361_591#_M1203_d N_D[12]_M1203_g N_VPWR_M1165_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1319 N_VPWR_M1319_d N_D[4]_M1319_g N_A_5361_297#_M1265_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1277 N_A_5361_591#_M1203_d N_D[12]_M1277_g N_VPWR_M1277_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1050 N_A_5361_297#_M1050_d N_A_5803_265#_M1050_g N_Z_M1050_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1055 N_Z_M1055_d N_A_5803_793#_M1055_g N_A_5361_591#_M1055_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1118 N_A_5361_297#_M1118_d N_A_5803_265#_M1118_g N_Z_M1050_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1119 N_Z_M1055_d N_A_5803_793#_M1119_g N_A_5361_591#_M1119_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1231 N_A_5361_297#_M1118_d N_A_5803_265#_M1231_g N_Z_M1231_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1200 N_Z_M1200_d N_A_5803_793#_M1200_g N_A_5361_591#_M1119_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1295 N_A_5361_297#_M1295_d N_A_5803_265#_M1295_g N_Z_M1231_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1257 N_Z_M1200_d N_A_5803_793#_M1257_g N_A_5361_591#_M1257_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1016 N_VPWR_M1016_d N_S[4]_M1016_g N_A_5803_265#_M1016_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1120 N_VPWR_M1120_d N_S[12]_M1120_g N_A_5803_793#_M1120_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1095 N_VPWR_M1095_d N_S[4]_M1095_g N_A_5803_265#_M1016_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1201 N_VPWR_M1201_d N_S[12]_M1201_g N_A_5803_793#_M1120_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1022 N_A_6674_325#_M1022_d N_S[5]_M1022_g N_VPWR_M1022_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1034 N_VPWR_M1034_d N_S[13]_M1034_g N_A_6674_599#_M1034_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1256 N_A_6674_325#_M1022_d N_S[5]_M1256_g N_VPWR_M1256_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1130 N_VPWR_M1130_d N_S[13]_M1130_g N_A_6674_599#_M1034_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1046 N_Z_M1046_d N_A_6674_325#_M1046_g N_A_6887_311#_M1046_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1092 N_Z_M1092_d N_A_6674_599#_M1092_g N_A_6887_613#_M1092_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1094 N_Z_M1046_d N_A_6674_325#_M1094_g N_A_6887_311#_M1094_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1117 N_Z_M1092_d N_A_6674_599#_M1117_g N_A_6887_613#_M1117_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1261 N_Z_M1261_d N_A_6674_325#_M1261_g N_A_6887_311#_M1094_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1196 N_Z_M1196_d N_A_6674_599#_M1196_g N_A_6887_613#_M1117_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1292 N_Z_M1261_d N_A_6674_325#_M1292_g N_A_6887_311#_M1292_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1238 N_Z_M1196_d N_A_6674_599#_M1238_g N_A_6887_613#_M1238_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1088 N_VPWR_M1088_d N_D[5]_M1088_g N_A_6887_311#_M1088_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1102 N_VPWR_M1102_d N_D[13]_M1102_g N_A_6887_613#_M1102_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1183 N_VPWR_M1183_d N_D[5]_M1183_g N_A_6887_311#_M1088_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1186 N_VPWR_M1186_d N_D[13]_M1186_g N_A_6887_613#_M1102_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1217 N_VPWR_M1183_d N_D[5]_M1217_g N_A_6887_311#_M1217_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1224 N_VPWR_M1186_d N_D[13]_M1224_g N_A_6887_613#_M1224_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1255 N_VPWR_M1255_d N_D[5]_M1255_g N_A_6887_311#_M1217_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1264 N_VPWR_M1264_d N_D[13]_M1264_g N_A_6887_613#_M1224_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1099 N_VPWR_M1099_d N_D[6]_M1099_g N_A_7937_297#_M1099_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1109 N_VPWR_M1109_d N_D[14]_M1109_g N_A_7937_591#_M1109_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1176 N_VPWR_M1176_d N_D[6]_M1176_g N_A_7937_297#_M1099_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1184 N_VPWR_M1184_d N_D[14]_M1184_g N_A_7937_591#_M1109_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1246 N_VPWR_M1176_d N_D[6]_M1246_g N_A_7937_297#_M1246_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1251 N_VPWR_M1184_d N_D[14]_M1251_g N_A_7937_591#_M1251_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1282 N_VPWR_M1282_d N_D[6]_M1282_g N_A_7937_297#_M1246_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1293 N_VPWR_M1293_d N_D[14]_M1293_g N_A_7937_591#_M1251_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1081 N_A_7937_297#_M1081_d N_A_8379_265#_M1081_g N_Z_M1081_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1025 N_A_7937_591#_M1025_d N_A_8379_793#_M1025_g N_Z_M1025_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1168 N_A_7937_297#_M1168_d N_A_8379_265#_M1168_g N_Z_M1081_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1077 N_A_7937_591#_M1077_d N_A_8379_793#_M1077_g N_Z_M1025_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1206 N_A_7937_297#_M1168_d N_A_8379_265#_M1206_g N_Z_M1206_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1227 N_A_7937_591#_M1077_d N_A_8379_793#_M1227_g N_Z_M1227_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1248 N_A_7937_297#_M1248_d N_A_8379_265#_M1248_g N_Z_M1206_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1314 N_A_7937_591#_M1314_d N_A_8379_793#_M1314_g N_Z_M1227_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1015 N_VPWR_M1015_d N_S[6]_M1015_g N_A_8379_265#_M1015_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1124 N_VPWR_M1124_d N_S[14]_M1124_g N_A_8379_793#_M1124_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1063 N_VPWR_M1063_d N_S[6]_M1063_g N_A_8379_265#_M1015_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1170 N_VPWR_M1170_d N_S[14]_M1170_g N_A_8379_793#_M1124_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1142 N_VPWR_M1142_d N_S[7]_M1142_g N_A_9250_325#_M1142_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1233 N_VPWR_M1233_d N_S[15]_M1233_g N_A_9250_599#_M1233_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1185 N_VPWR_M1185_d N_S[7]_M1185_g N_A_9250_325#_M1142_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1279 N_VPWR_M1279_d N_S[15]_M1279_g N_A_9250_599#_M1233_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1013 N_Z_M1013_d N_A_9250_325#_M1013_g N_A_9463_311#_M1013_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1166 N_Z_M1166_d N_A_9250_599#_M1166_g N_A_9463_613#_M1166_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1058 N_Z_M1013_d N_A_9250_325#_M1058_g N_A_9463_311#_M1058_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1204 N_Z_M1166_d N_A_9250_599#_M1204_g N_A_9463_613#_M1204_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1153 N_Z_M1153_d N_A_9250_325#_M1153_g N_A_9463_311#_M1058_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1286 N_Z_M1286_d N_A_9250_599#_M1286_g N_A_9463_613#_M1204_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1163 N_Z_M1153_d N_A_9250_325#_M1163_g N_A_9463_311#_M1163_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1303 N_Z_M1286_d N_A_9250_599#_M1303_g N_A_9463_613#_M1303_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1040 N_VPWR_M1040_d N_D[7]_M1040_g N_A_9463_311#_M1040_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1056 N_VPWR_M1056_d N_D[15]_M1056_g N_A_9463_613#_M1056_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1087 N_VPWR_M1087_d N_D[7]_M1087_g N_A_9463_311#_M1040_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1103 N_VPWR_M1103_d N_D[15]_M1103_g N_A_9463_613#_M1056_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1131 N_VPWR_M1087_d N_D[7]_M1131_g N_A_9463_311#_M1131_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1145 N_VPWR_M1103_d N_D[15]_M1145_g N_A_9463_613#_M1145_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1151 N_VPWR_M1151_d N_D[7]_M1151_g N_A_9463_311#_M1131_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1156 N_VPWR_M1156_d N_D[15]_M1156_g N_A_9463_613#_M1145_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX320_noxref VNB VPB NWDIODE A=148.179 P=110.38
*
.include "sky130_fd_sc_hdll__muxb16to1_4.pxi.spice"
*
.ends
*
*
