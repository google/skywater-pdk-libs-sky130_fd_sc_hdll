* File: sky130_fd_sc_hdll__sdlclkp_2.pex.spice
* Created: Wed Sep  2 08:52:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%SCE 2 3 5 8 10 11 19
c29 3 0 1.61703e-19 $X=0.495 $Y=1.77
r30 18 19 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r31 15 18 43.7153 $w=3.3e-07 $l=2.5e-07 $layer=POLY_cond $X=0.245 $Y=1.16
+ $X2=0.495 $Y2=1.16
r32 10 11 17.4042 $w=2.43e-07 $l=3.7e-07 $layer=LI1_cond $X=0.207 $Y=1.16
+ $X2=0.207 $Y2=1.53
r33 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r34 6 19 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.16
r35 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.445
r36 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r37 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.67 $X2=0.495
+ $Y2=1.77
r38 1 18 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.16
r39 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.495 $Y=1.325
+ $X2=0.495 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GATE 2 3 5 8 10 11 15 16
c41 16 0 1.90185e-19 $X=0.975 $Y=1.16
c42 15 0 8.05567e-20 $X=0.975 $Y=1.16
c43 2 0 1.52835e-19 $X=0.905 $Y=1.67
r44 15 18 39.5599 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.957 $Y=1.16
+ $X2=0.957 $Y2=1.325
r45 15 17 47.9606 $w=3.05e-07 $l=1.65e-07 $layer=POLY_cond $X=0.957 $Y=1.16
+ $X2=0.957 $Y2=0.995
r46 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.975
+ $Y=1.16 $X2=0.975 $Y2=1.16
r47 10 11 9.67483 $w=4.03e-07 $l=3.4e-07 $layer=LI1_cond $X=1.092 $Y=1.53
+ $X2=1.092 $Y2=1.87
r48 10 16 10.5285 $w=4.03e-07 $l=3.7e-07 $layer=LI1_cond $X=1.092 $Y=1.53
+ $X2=1.092 $Y2=1.16
r49 8 17 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.945 $Y=0.445
+ $X2=0.945 $Y2=0.995
r50 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.905 $Y=1.77
+ $X2=0.905 $Y2=2.165
r51 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.905 $Y=1.67 $X2=0.905
+ $Y2=1.77
r52 2 18 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=0.905 $Y=1.67
+ $X2=0.905 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_269_21# 1 2 9 11 13 14 17 20 25 26 28
+ 34 36 39 41 43 45 47 52 53 56 59
c174 52 0 1.44161e-19 $X=4.44 $Y=1.53
c175 45 0 3.5877e-19 $X=1.712 $Y=1.452
c176 25 0 2.99785e-20 $X=1.55 $Y=0.87
c177 9 0 2.2455e-20 $X=1.42 $Y=0.415
r178 67 68 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.875
+ $Y=1.74 $X2=1.875 $Y2=1.74
r179 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.585 $Y=1.53
+ $X2=4.585 $Y2=1.53
r180 56 68 5.07427 $w=4.93e-07 $l=2.1e-07 $layer=LI1_cond $X=1.712 $Y=1.53
+ $X2=1.712 $Y2=1.74
r181 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.71 $Y=1.53
+ $X2=1.71 $Y2=1.53
r182 53 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.855 $Y=1.53
+ $X2=1.71 $Y2=1.53
r183 52 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.44 $Y=1.53
+ $X2=4.585 $Y2=1.53
r184 52 53 3.19925 $w=1.4e-07 $l=2.585e-06 $layer=MET1_cond $X=4.44 $Y=1.53
+ $X2=1.855 $Y2=1.53
r185 45 56 1.88473 $w=4.93e-07 $l=7.8e-08 $layer=LI1_cond $X=1.712 $Y=1.452
+ $X2=1.712 $Y2=1.53
r186 45 46 7.22426 $w=4.93e-07 $l=2.47e-07 $layer=LI1_cond $X=1.712 $Y=1.452
+ $X2=1.712 $Y2=1.205
r187 41 43 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=4.96 $Y=0.615
+ $X2=4.96 $Y2=0.465
r188 37 60 3.79964 $w=2.5e-07 $l=1.53e-07 $layer=LI1_cond $X=4.67 $Y=1.62
+ $X2=4.517 $Y2=1.62
r189 37 39 17.5171 $w=2.48e-07 $l=3.8e-07 $layer=LI1_cond $X=4.67 $Y=1.62
+ $X2=5.05 $Y2=1.62
r190 36 47 3.17288 $w=2.97e-07 $l=8.89101e-08 $layer=LI1_cond $X=4.525 $Y=1.105
+ $X2=4.517 $Y2=1.19
r191 35 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.525 $Y=0.7
+ $X2=4.96 $Y2=0.7
r192 35 36 12.7166 $w=2.88e-07 $l=3.2e-07 $layer=LI1_cond $X=4.525 $Y=0.785
+ $X2=4.525 $Y2=1.105
r193 34 60 3.10428 $w=3.05e-07 $l=1.25e-07 $layer=LI1_cond $X=4.517 $Y=1.495
+ $X2=4.517 $Y2=1.62
r194 33 47 3.17288 $w=2.97e-07 $l=8.5e-08 $layer=LI1_cond $X=4.517 $Y=1.275
+ $X2=4.517 $Y2=1.19
r195 33 34 8.3127 $w=3.03e-07 $l=2.2e-07 $layer=LI1_cond $X=4.517 $Y=1.275
+ $X2=4.517 $Y2=1.495
r196 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.24
+ $Y=1.19 $X2=4.24 $Y2=1.19
r197 28 47 3.41642 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=4.365 $Y=1.19
+ $X2=4.517 $Y2=1.19
r198 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.365 $Y=1.19
+ $X2=4.24 $Y2=1.19
r199 26 62 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=1.55 $Y=0.87
+ $X2=1.42 $Y2=0.87
r200 25 46 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=1.632 $Y=0.87
+ $X2=1.632 $Y2=1.205
r201 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.55
+ $Y=0.87 $X2=1.55 $Y2=0.87
r202 18 31 34.1407 $w=3.26e-07 $l=1.46969e-07 $layer=POLY_cond $X=4.24 $Y=1.055
+ $X2=4.265 $Y2=1.19
r203 18 20 312.787 $w=1.5e-07 $l=6.1e-07 $layer=POLY_cond $X=4.24 $Y=1.055
+ $X2=4.24 $Y2=0.445
r204 14 31 46.5577 $w=3.26e-07 $l=2.73861e-07 $layer=POLY_cond $X=4.215 $Y=1.44
+ $X2=4.265 $Y2=1.19
r205 14 17 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.215 $Y=1.44
+ $X2=4.215 $Y2=1.835
r206 11 67 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.96 $Y=1.99
+ $X2=1.9 $Y2=1.74
r207 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.96 $Y=1.99
+ $X2=1.96 $Y2=2.275
r208 7 62 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=1.42 $Y=0.735
+ $X2=1.42 $Y2=0.87
r209 7 9 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.42 $Y=0.735
+ $X2=1.42 $Y2=0.415
r210 2 39 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.905
+ $Y=1.515 $X2=5.05 $Y2=1.66
r211 1 43 182 $w=1.7e-07 $l=2.89741e-07 $layer=licon1_NDIFF $count=1 $X=4.785
+ $Y=0.235 $X2=4.92 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_266_243# 1 2 8 9 11 12 13 16 18 21 24
+ 28 30 31 37 38 41 42 43
c124 42 0 2.2455e-20 $X=2.06 $Y=0.87
c125 41 0 2.82989e-19 $X=2.06 $Y=0.87
c126 37 0 5.69068e-21 $X=4.075 $Y=0.85
c127 28 0 1.17835e-19 $X=3.98 $Y=1.66
c128 18 0 2.84822e-20 $X=2.022 $Y=1.215
c129 8 0 3.15944e-20 $X=1.43 $Y=1.89
r130 41 44 38.5487 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.082 $Y=0.87
+ $X2=2.082 $Y2=1.035
r131 41 43 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.082 $Y=0.87
+ $X2=2.082 $Y2=0.705
r132 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.06
+ $Y=0.87 $X2=2.06 $Y2=0.87
r133 38 50 6.59116 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.947 $Y=0.85
+ $X2=3.947 $Y2=0.935
r134 38 49 2.91128 $w=4.23e-07 $l=8.5e-08 $layer=LI1_cond $X=3.947 $Y=0.85
+ $X2=3.947 $Y2=0.765
r135 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.075 $Y=0.85
+ $X2=4.075 $Y2=0.85
r136 33 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.22 $Y=0.85
+ $X2=2.22 $Y2=0.85
r137 31 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.365 $Y=0.85
+ $X2=2.22 $Y2=0.85
r138 30 37 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.93 $Y=0.85
+ $X2=4.075 $Y2=0.85
r139 30 31 1.93688 $w=1.4e-07 $l=1.565e-06 $layer=MET1_cond $X=3.93 $Y=0.85
+ $X2=2.365 $Y2=0.85
r140 25 28 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.82 $Y=1.66
+ $X2=3.98 $Y2=1.66
r141 24 25 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.82 $Y=1.575
+ $X2=3.82 $Y2=1.66
r142 24 50 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.82 $Y=1.575
+ $X2=3.82 $Y2=0.935
r143 21 49 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=3.9 $Y=0.465 $X2=3.9
+ $Y2=0.765
r144 18 44 61.2142 $w=1.95e-07 $l=1.8e-07 $layer=POLY_cond $X=2.022 $Y=1.215
+ $X2=2.022 $Y2=1.035
r145 16 43 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2 $Y=0.415 $X2=2
+ $Y2=0.705
r146 12 18 27.531 $w=1.5e-07 $l=1.29167e-07 $layer=POLY_cond $X=1.925 $Y=1.29
+ $X2=2.022 $Y2=1.215
r147 12 13 202.543 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=1.925 $Y=1.29
+ $X2=1.53 $Y2=1.29
r148 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.43 $Y=1.99
+ $X2=1.43 $Y2=2.275
r149 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.43 $Y=1.89 $X2=1.43
+ $Y2=1.99
r150 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=1.43 $Y=1.365
+ $X2=1.53 $Y2=1.29
r151 7 8 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=1.43 $Y=1.365 $X2=1.43
+ $Y2=1.89
r152 2 28 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=3.855
+ $Y=1.515 $X2=3.98 $Y2=1.66
r153 1 21 182 $w=1.7e-07 $l=2.85745e-07 $layer=licon1_NDIFF $count=1 $X=3.855
+ $Y=0.235 $X2=3.98 $Y2=0.465
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_484_315# 1 2 7 9 12 15 16 18 21 23 27
+ 31 33 37 44 45 50
c132 37 0 1.05178e-19 $X=5.63 $Y=1.16
c133 33 0 5.88603e-20 $X=5.405 $Y=2
c134 12 0 1.25378e-19 $X=2.655 $Y=0.445
r135 49 50 4.37153 $w=3.3e-07 $l=2.5e-08 $layer=POLY_cond $X=5.825 $Y=1.16
+ $X2=5.85 $Y2=1.16
r136 41 44 4.25649 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=2.555 $Y=1.74
+ $X2=2.665 $Y2=1.74
r137 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.555
+ $Y=1.74 $X2=2.555 $Y2=1.74
r138 38 49 34.0979 $w=3.3e-07 $l=1.95e-07 $layer=POLY_cond $X=5.63 $Y=1.16
+ $X2=5.825 $Y2=1.16
r139 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.63
+ $Y=1.16 $X2=5.63 $Y2=1.16
r140 35 37 24.8598 $w=3.48e-07 $l=7.55e-07 $layer=LI1_cond $X=5.58 $Y=1.915
+ $X2=5.58 $Y2=1.16
r141 34 45 2.69039 $w=1.7e-07 $l=1.87083e-07 $layer=LI1_cond $X=3.545 $Y=2
+ $X2=3.435 $Y2=1.86
r142 33 35 7.93686 $w=1.7e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.405 $Y=2
+ $X2=5.58 $Y2=1.915
r143 33 34 121.348 $w=1.68e-07 $l=1.86e-06 $layer=LI1_cond $X=5.405 $Y=2
+ $X2=3.545 $Y2=2
r144 29 45 3.42573 $w=1.7e-07 $l=2.37171e-07 $layer=LI1_cond $X=3.46 $Y=1.635
+ $X2=3.435 $Y2=1.86
r145 29 31 79.2674 $w=1.68e-07 $l=1.215e-06 $layer=LI1_cond $X=3.46 $Y=1.635
+ $X2=3.46 $Y2=0.42
r146 25 45 3.42573 $w=2.2e-07 $l=2.25e-07 $layer=LI1_cond $X=3.435 $Y=2.085
+ $X2=3.435 $Y2=1.86
r147 25 27 6.28605 $w=2.18e-07 $l=1.2e-07 $layer=LI1_cond $X=3.435 $Y=2.085
+ $X2=3.435 $Y2=2.205
r148 23 45 2.69039 $w=2.7e-07 $l=1.48324e-07 $layer=LI1_cond $X=3.325 $Y=1.77
+ $X2=3.435 $Y2=1.86
r149 23 44 28.1708 $w=2.68e-07 $l=6.6e-07 $layer=LI1_cond $X=3.325 $Y=1.77
+ $X2=2.665 $Y2=1.77
r150 19 50 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.85 $Y=0.995
+ $X2=5.85 $Y2=1.16
r151 19 21 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=5.85 $Y=0.995
+ $X2=5.85 $Y2=0.445
r152 16 18 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=5.825 $Y=1.77
+ $X2=5.825 $Y2=2.165
r153 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.825 $Y=1.67 $X2=5.825
+ $Y2=1.77
r154 14 49 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.16
r155 14 15 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=5.825 $Y=1.325
+ $X2=5.825 $Y2=1.67
r156 10 42 38.6443 $w=2.87e-07 $l=2.0106e-07 $layer=POLY_cond $X=2.655 $Y=1.575
+ $X2=2.575 $Y2=1.74
r157 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=2.655 $Y=1.575
+ $X2=2.655 $Y2=0.445
r158 7 42 48.651 $w=2.87e-07 $l=2.76134e-07 $layer=POLY_cond $X=2.52 $Y=1.99
+ $X2=2.575 $Y2=1.74
r159 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.52 $Y=1.99
+ $X2=2.52 $Y2=2.275
r160 2 27 600 $w=1.7e-07 $l=7.89177e-07 $layer=licon1_PDIFF $count=1 $X=3.315
+ $Y=1.485 $X2=3.46 $Y2=2.205
r161 1 31 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=3.325
+ $Y=0.235 $X2=3.46 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_299_47# 1 2 7 9 10 12 13 17 22 23 24
+ 26 29 32
c102 32 0 1.38828e-19 $X=2.56 $Y=1.185
c103 26 0 2.99785e-20 $X=2.56 $Y=0.995
c104 24 0 3.15944e-20 $X=2.3 $Y=1.29
r105 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.12
+ $Y=1.16 $X2=3.12 $Y2=1.16
r106 27 32 3.40559 $w=2.75e-07 $l=8.5e-08 $layer=LI1_cond $X=2.645 $Y=1.185
+ $X2=2.56 $Y2=1.185
r107 27 29 14.4055 $w=3.78e-07 $l=4.75e-07 $layer=LI1_cond $X=2.645 $Y=1.185
+ $X2=3.12 $Y2=1.185
r108 26 32 3.11956 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.56 $Y=0.995
+ $X2=2.56 $Y2=1.185
r109 25 26 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.56 $Y=0.535
+ $X2=2.56 $Y2=0.995
r110 23 32 3.40559 $w=2.75e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.475 $Y=1.29
+ $X2=2.56 $Y2=1.185
r111 23 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.475 $Y=1.29
+ $X2=2.3 $Y2=1.29
r112 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.215 $Y=1.375
+ $X2=2.3 $Y2=1.29
r113 21 22 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=2.215 $Y=1.375
+ $X2=2.215 $Y2=2.125
r114 17 22 7.85115 $w=3.4e-07 $l=2.08207e-07 $layer=LI1_cond $X=2.13 $Y=2.295
+ $X2=2.215 $Y2=2.125
r115 17 19 14.7445 $w=3.38e-07 $l=4.35e-07 $layer=LI1_cond $X=2.13 $Y=2.295
+ $X2=1.695 $Y2=2.295
r116 13 25 7.36005 $w=2.8e-07 $l=1.77482e-07 $layer=LI1_cond $X=2.475 $Y=0.395
+ $X2=2.56 $Y2=0.535
r117 13 15 30.6632 $w=2.78e-07 $l=7.45e-07 $layer=LI1_cond $X=2.475 $Y=0.395
+ $X2=1.73 $Y2=0.395
r118 10 30 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.155 $Y2=1.16
r119 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.25 $Y=0.995
+ $X2=3.25 $Y2=0.56
r120 7 30 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.155 $Y2=1.16
r121 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.225 $Y=1.41
+ $X2=3.225 $Y2=1.985
r122 2 19 600 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=1.52 $Y=2.065
+ $X2=1.695 $Y2=2.29
r123 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=1.495
+ $Y=0.235 $X2=1.73 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%CLK 1 3 4 7 10 13 14 16 18 19 21 24 28
+ 30 31 45
c104 30 0 7.91502e-20 $X=6.27 $Y=1.16
c105 28 0 1.33709e-19 $X=5.05 $Y=1.16
c106 14 0 1.64039e-19 $X=6.295 $Y=1.77
c107 7 0 1.17835e-19 $X=4.815 $Y=1.835
c108 4 0 5.69068e-21 $X=4.815 $Y=1.44
r109 30 32 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.16
+ $X2=6.295 $Y2=0.995
r110 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.27
+ $Y=1.16 $X2=6.27 $Y2=1.16
r111 28 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.095 $Y=1.19
+ $X2=5.095 $Y2=1.19
r112 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.05
+ $Y=1.16 $X2=5.05 $Y2=1.16
r113 24 45 0.0128321 $w=2.3e-07 $l=2e-08 $layer=MET1_cond $X=5.055 $Y=1.19
+ $X2=5.075 $Y2=1.19
r114 22 31 6.46067 $w=3.28e-07 $l=1.85e-07 $layer=LI1_cond $X=6.085 $Y=1.16
+ $X2=6.27 $Y2=1.16
r115 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.085 $Y=1.19
+ $X2=6.085 $Y2=1.19
r116 19 45 0.128299 $w=2.3e-07 $l=1.65e-07 $layer=MET1_cond $X=5.24 $Y=1.19
+ $X2=5.075 $Y2=1.19
r117 18 21 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.94 $Y=1.19
+ $X2=6.085 $Y2=1.19
r118 18 19 0.866335 $w=1.4e-07 $l=7e-07 $layer=MET1_cond $X=5.94 $Y=1.19
+ $X2=5.24 $Y2=1.19
r119 14 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.295 $Y=1.77
+ $X2=6.295 $Y2=2.165
r120 13 14 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.295 $Y=1.67 $X2=6.295
+ $Y2=1.77
r121 12 30 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=6.295 $Y=1.325
+ $X2=6.295 $Y2=1.16
r122 12 13 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=6.295 $Y=1.325
+ $X2=6.295 $Y2=1.67
r123 10 32 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=6.21 $Y=0.445
+ $X2=6.21 $Y2=0.995
r124 4 27 47.9649 $w=4.43e-07 $l=3.24037e-07 $layer=POLY_cond $X=4.815 $Y=1.44
+ $X2=4.91 $Y2=1.16
r125 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.815 $Y=1.44
+ $X2=4.815 $Y2=1.835
r126 1 27 69.3486 $w=4.43e-07 $l=5.20481e-07 $layer=POLY_cond $X=4.71 $Y=0.73
+ $X2=4.91 $Y2=1.16
r127 1 3 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.71 $Y=0.73 $X2=4.71
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_1093_47# 1 2 9 11 13 16 18 20 23 25 26
+ 27 31 33 34 40 42 46
c111 46 0 1.64127e-19 $X=7.265 $Y=1.217
c112 42 0 5.46563e-20 $X=6.665 $Y=1.185
c113 33 0 7.91502e-20 $X=6.665 $Y=1.495
r114 46 47 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=7.265 $Y=1.217
+ $X2=7.29 $Y2=1.217
r115 43 44 3.56509 $w=3.38e-07 $l=2.5e-08 $layer=POLY_cond $X=6.795 $Y=1.217
+ $X2=6.82 $Y2=1.217
r116 38 40 12.2649 $w=5.88e-07 $l=6.05e-07 $layer=LI1_cond $X=6.06 $Y=1.79
+ $X2=6.665 $Y2=1.79
r117 37 46 54.1894 $w=3.38e-07 $l=3.8e-07 $layer=POLY_cond $X=6.885 $Y=1.217
+ $X2=7.265 $Y2=1.217
r118 37 44 9.26923 $w=3.38e-07 $l=6.5e-08 $layer=POLY_cond $X=6.885 $Y=1.217
+ $X2=6.82 $Y2=1.217
r119 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.885
+ $Y=1.16 $X2=6.885 $Y2=1.16
r120 34 42 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.75 $Y=1.185
+ $X2=6.665 $Y2=1.185
r121 34 36 6.33462 $w=2.6e-07 $l=1.35e-07 $layer=LI1_cond $X=6.75 $Y=1.185
+ $X2=6.885 $Y2=1.185
r122 33 40 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.665 $Y=1.495
+ $X2=6.665 $Y2=1.79
r123 32 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.665 $Y=1.315
+ $X2=6.665 $Y2=1.185
r124 32 33 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.665 $Y=1.315
+ $X2=6.665 $Y2=1.495
r125 31 42 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.665 $Y=1.055
+ $X2=6.665 $Y2=1.185
r126 30 31 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=6.665 $Y=0.785
+ $X2=6.665 $Y2=1.055
r127 27 38 8.20854 $w=1.7e-07 $l=2.95e-07 $layer=LI1_cond $X=6.06 $Y=2.085
+ $X2=6.06 $Y2=1.79
r128 27 29 2.87059 $w=1.7e-07 $l=4e-08 $layer=LI1_cond $X=6.06 $Y=2.085 $X2=6.06
+ $Y2=2.125
r129 25 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.58 $Y=0.7
+ $X2=6.665 $Y2=0.785
r130 25 26 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=6.58 $Y=0.7
+ $X2=5.675 $Y2=0.7
r131 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.59 $Y=0.615
+ $X2=5.675 $Y2=0.7
r132 21 23 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=5.59 $Y=0.615
+ $X2=5.59 $Y2=0.46
r133 18 47 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.29 $Y=1.41
+ $X2=7.29 $Y2=1.217
r134 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.29 $Y=1.41
+ $X2=7.29 $Y2=1.985
r135 14 46 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.265 $Y=1.025
+ $X2=7.265 $Y2=1.217
r136 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.265 $Y=1.025
+ $X2=7.265 $Y2=0.56
r137 11 44 17.4907 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.82 $Y=1.41
+ $X2=6.82 $Y2=1.217
r138 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.82 $Y=1.41
+ $X2=6.82 $Y2=1.985
r139 7 43 21.7938 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.795 $Y=1.025
+ $X2=6.795 $Y2=1.217
r140 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.795 $Y=1.025
+ $X2=6.795 $Y2=0.56
r141 2 29 600 $w=1.7e-07 $l=3.44964e-07 $layer=licon1_PDIFF $count=1 $X=5.915
+ $Y=1.845 $X2=6.06 $Y2=2.125
r142 1 23 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=5.465
+ $Y=0.235 $X2=5.59 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VPWR 1 2 3 4 5 6 19 21 27 29 31 34 37 39
+ 40 41 48 60 70 76 80 83
r102 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r103 78 80 6.78742 $w=5.48e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=2.53
+ $X2=3.885 $Y2=2.53
r104 78 79 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r105 76 80 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=3.105 $Y=2.72
+ $X2=3.885 $Y2=2.72
r106 75 79 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r107 74 76 10.1774 $w=7.28e-07 $l=1.15e-07 $layer=LI1_cond $X=2.99 $Y=2.44
+ $X2=3.105 $Y2=2.44
r108 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 72 74 1.72039 $w=7.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.885 $Y=2.44
+ $X2=2.99 $Y2=2.44
r110 69 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.99 $Y2=2.72
r111 68 72 5.81655 $w=7.28e-07 $l=3.55e-07 $layer=LI1_cond $X=2.53 $Y=2.44
+ $X2=2.885 $Y2=2.44
r112 68 70 8.45698 $w=7.28e-07 $l=1e-08 $layer=LI1_cond $X=2.53 $Y=2.44 $X2=2.52
+ $Y2=2.44
r113 68 69 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r114 63 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r115 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r116 60 82 3.99177 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.44 $Y=2.72
+ $X2=7.63 $Y2=2.72
r117 60 62 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=7.44 $Y=2.72
+ $X2=7.13 $Y2=2.72
r118 59 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r119 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 56 59 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r121 55 56 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r122 53 55 16.8538 $w=5.48e-07 $l=7.75e-07 $layer=LI1_cond $X=4.515 $Y=2.53
+ $X2=5.29 $Y2=2.53
r123 51 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=5.29 $Y2=2.72
r124 51 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r125 50 53 3.1533 $w=5.48e-07 $l=1.45e-07 $layer=LI1_cond $X=4.37 $Y=2.53
+ $X2=4.515 $Y2=2.53
r126 50 51 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r127 48 78 5.43672 $w=5.48e-07 $l=2.5e-07 $layer=LI1_cond $X=4.16 $Y=2.53
+ $X2=3.91 $Y2=2.53
r128 48 50 4.56684 $w=5.48e-07 $l=2.1e-07 $layer=LI1_cond $X=4.16 $Y=2.53
+ $X2=4.37 $Y2=2.53
r129 47 69 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r130 46 70 119.39 $w=1.68e-07 $l=1.83e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.52 $Y2=2.72
r131 46 47 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r132 44 65 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r133 44 46 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r134 41 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 41 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r136 39 58 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=6.21 $Y2=2.72
r137 39 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.395 $Y=2.72
+ $X2=6.56 $Y2=2.72
r138 38 62 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=6.725 $Y=2.72
+ $X2=7.13 $Y2=2.72
r139 38 40 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.725 $Y=2.72
+ $X2=6.56 $Y2=2.72
r140 37 58 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=5.755 $Y=2.72
+ $X2=6.21 $Y2=2.72
r141 36 37 9.83198 $w=5.48e-07 $l=1.65e-07 $layer=LI1_cond $X=5.59 $Y=2.53
+ $X2=5.755 $Y2=2.53
r142 34 55 4.13191 $w=5.48e-07 $l=1.9e-07 $layer=LI1_cond $X=5.48 $Y=2.53
+ $X2=5.29 $Y2=2.53
r143 34 36 2.39216 $w=5.48e-07 $l=1.1e-07 $layer=LI1_cond $X=5.48 $Y=2.53
+ $X2=5.59 $Y2=2.53
r144 29 82 3.1514 $w=2.5e-07 $l=1.12916e-07 $layer=LI1_cond $X=7.565 $Y=2.635
+ $X2=7.63 $Y2=2.72
r145 29 31 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=7.565 $Y=2.635
+ $X2=7.565 $Y2=2
r146 25 40 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.56 $Y=2.635
+ $X2=6.56 $Y2=2.72
r147 25 27 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=6.56 $Y=2.635
+ $X2=6.56 $Y2=2.36
r148 19 65 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r149 19 21 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=2
r150 6 31 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.38
+ $Y=1.485 $X2=7.525 $Y2=2
r151 5 27 600 $w=1.7e-07 $l=5.96112e-07 $layer=licon1_PDIFF $count=1 $X=6.385
+ $Y=1.845 $X2=6.56 $Y2=2.36
r152 4 36 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=5.445
+ $Y=1.845 $X2=5.59 $Y2=2.36
r153 3 53 600 $w=1.7e-07 $l=9.24054e-07 $layer=licon1_PDIFF $count=1 $X=4.305
+ $Y=1.515 $X2=4.515 $Y2=2.34
r154 2 72 600 $w=1.7e-07 $l=4.10061e-07 $layer=licon1_PDIFF $count=1 $X=2.61
+ $Y=2.065 $X2=2.885 $Y2=2.36
r155 1 21 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%A_27_47# 1 2 3 12 15 16 17 18 20 24
c53 24 0 1.74968e-19 $X=1.2 $Y=0.42
r54 22 24 12.0152 $w=1.78e-07 $l=1.95e-07 $layer=LI1_cond $X=1.205 $Y=0.615
+ $X2=1.205 $Y2=0.42
r55 18 20 16.1003 $w=3.38e-07 $l=4.75e-07 $layer=LI1_cond $X=0.72 $Y=2.295
+ $X2=1.195 $Y2=2.295
r56 16 22 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=1.205 $Y2=0.615
r57 16 17 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=1.115 $Y=0.7
+ $X2=0.72 $Y2=0.7
r58 15 18 7.37505 $w=3.4e-07 $l=2.1543e-07 $layer=LI1_cond $X=0.617 $Y=2.125
+ $X2=0.72 $Y2=2.295
r59 14 17 6.71979 $w=1.68e-07 $l=1.03e-07 $layer=LI1_cond $X=0.617 $Y=0.7
+ $X2=0.72 $Y2=0.7
r60 14 15 72.4967 $w=2.03e-07 $l=1.34e-06 $layer=LI1_cond $X=0.617 $Y=0.785
+ $X2=0.617 $Y2=2.125
r61 10 14 26.2267 $w=1.68e-07 $l=4.02e-07 $layer=LI1_cond $X=0.215 $Y=0.7
+ $X2=0.617 $Y2=0.7
r62 10 12 8.20008 $w=2.58e-07 $l=1.85e-07 $layer=LI1_cond $X=0.215 $Y=0.615
+ $X2=0.215 $Y2=0.43
r63 3 20 600 $w=1.7e-07 $l=5.35747e-07 $layer=licon1_PDIFF $count=1 $X=0.995
+ $Y=1.845 $X2=1.195 $Y2=2.29
r64 2 24 182 $w=1.7e-07 $l=2.59856e-07 $layer=licon1_NDIFF $count=1 $X=1.02
+ $Y=0.235 $X2=1.2 $Y2=0.42
r65 1 12 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%GCLK 1 2 8 9 10 11 12 14 20 21 22
c46 14 0 1.64127e-19 $X=7.005 $Y=0.36
r47 20 21 18.2086 $w=2.48e-07 $l=3.95e-07 $layer=LI1_cond $X=7.095 $Y=1.815
+ $X2=7.095 $Y2=2.21
r48 19 22 17.6855 $w=1.83e-07 $l=2.95e-07 $layer=LI1_cond $X=7.582 $Y=1.485
+ $X2=7.582 $Y2=1.19
r49 18 22 18.285 $w=1.83e-07 $l=3.05e-07 $layer=LI1_cond $X=7.582 $Y=0.885
+ $X2=7.582 $Y2=1.19
r50 17 20 7.37564 $w=2.48e-07 $l=1.6e-07 $layer=LI1_cond $X=7.095 $Y=1.655
+ $X2=7.095 $Y2=1.815
r51 12 17 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=7.22 $Y=1.57
+ $X2=7.095 $Y2=1.655
r52 11 19 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.49 $Y=1.57
+ $X2=7.582 $Y2=1.485
r53 11 12 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=7.49 $Y=1.57 $X2=7.22
+ $Y2=1.57
r54 9 18 6.83233 $w=1.7e-07 $l=1.27609e-07 $layer=LI1_cond $X=7.49 $Y=0.8
+ $X2=7.582 $Y2=0.885
r55 9 10 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=7.49 $Y=0.8 $X2=7.17
+ $Y2=0.8
r56 8 10 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=7.07 $Y=0.715
+ $X2=7.17 $Y2=0.8
r57 7 14 0.40127 $w=2e-07 $l=1.23288e-07 $layer=LI1_cond $X=7.07 $Y=0.445
+ $X2=7.005 $Y2=0.35
r58 7 8 14.9727 $w=1.98e-07 $l=2.7e-07 $layer=LI1_cond $X=7.07 $Y=0.445 $X2=7.07
+ $Y2=0.715
r59 2 20 300 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=2 $X=6.91
+ $Y=1.485 $X2=7.055 $Y2=1.815
r60 1 14 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=6.87
+ $Y=0.235 $X2=7.005 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDLCLKP_2%VGND 1 2 3 4 5 18 22 26 30 33 34 35 37
+ 42 47 59 65 71 74 78 79
r116 78 79 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r117 76 78 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.475 $Y=0
+ $X2=7.59 $Y2=0
r118 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r119 71 72 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r120 65 68 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.36
r121 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r122 62 79 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r123 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r124 59 76 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=7.39 $Y=0 $X2=7.475
+ $Y2=0
r125 59 61 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.39 $Y=0 $X2=7.13
+ $Y2=0
r126 58 62 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r127 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r128 55 58 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=6.21 $Y2=0
r129 55 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=4.37
+ $Y2=0
r130 54 57 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=0 $X2=6.21
+ $Y2=0
r131 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r132 52 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.615 $Y=0 $X2=4.45
+ $Y2=0
r133 52 54 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=4.615 $Y=0
+ $X2=4.83 $Y2=0
r134 51 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r135 51 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=2.99
+ $Y2=0
r136 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r137 48 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.995
+ $Y2=0
r138 48 50 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.91
+ $Y2=0
r139 47 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.285 $Y=0 $X2=4.45
+ $Y2=0
r140 47 50 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=4.285 $Y=0
+ $X2=3.91 $Y2=0
r141 46 72 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r142 46 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r143 45 46 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r144 43 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r145 43 45 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r146 42 71 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.91 $Y=0 $X2=2.995
+ $Y2=0
r147 42 45 114.824 $w=1.68e-07 $l=1.76e-06 $layer=LI1_cond $X=2.91 $Y=0 $X2=1.15
+ $Y2=0
r148 37 65 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r149 37 39 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r150 35 66 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r151 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r152 33 57 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.21 $Y2=0
r153 33 34 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=6.335 $Y=0
+ $X2=6.502 $Y2=0
r154 32 61 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=7.13
+ $Y2=0
r155 32 34 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=6.67 $Y=0 $X2=6.502
+ $Y2=0
r156 28 76 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0
r157 28 30 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.475 $Y=0.085
+ $X2=7.475 $Y2=0.38
r158 24 34 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=6.502 $Y=0.085
+ $X2=6.502 $Y2=0
r159 24 26 9.46035 $w=3.33e-07 $l=2.75e-07 $layer=LI1_cond $X=6.502 $Y=0.085
+ $X2=6.502 $Y2=0.36
r160 20 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0
r161 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.45 $Y=0.085
+ $X2=4.45 $Y2=0.36
r162 16 71 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0
r163 16 18 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=2.995 $Y=0.085
+ $X2=2.995 $Y2=0.51
r164 5 30 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.34
+ $Y=0.235 $X2=7.475 $Y2=0.38
r165 4 26 182 $w=1.7e-07 $l=2.755e-07 $layer=licon1_NDIFF $count=1 $X=6.285
+ $Y=0.235 $X2=6.505 $Y2=0.36
r166 3 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=4.315
+ $Y=0.235 $X2=4.45 $Y2=0.36
r167 2 18 182 $w=1.7e-07 $l=3.85357e-07 $layer=licon1_NDIFF $count=1 $X=2.73
+ $Y=0.235 $X2=2.995 $Y2=0.51
r168 1 68 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.36
.ends

