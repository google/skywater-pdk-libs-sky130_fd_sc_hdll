* File: sky130_fd_sc_hdll__muxb16to1_2.spice
* Created: Thu Aug 27 19:11:31 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb16to1_2.pex.spice"
.subckt sky130_fd_sc_hdll__muxb16to1_2  VNB VPB D[0] D[8] S[0] S[8] S[1] S[9]
+ D[1] D[9] D[2] D[10] S[2] S[10] S[3] S[11] D[3] D[11] D[4] D[12] S[4] S[12]
+ S[5] S[13] D[5] D[13] D[6] D[14] S[6] S[14] S[7] S[15] D[7] D[15] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[15]	D[15]
* D[7]	D[7]
* S[15]	S[15]
* S[7]	S[7]
* S[14]	S[14]
* S[6]	S[6]
* D[14]	D[14]
* D[6]	D[6]
* D[13]	D[13]
* D[5]	D[5]
* S[13]	S[13]
* S[5]	S[5]
* S[12]	S[12]
* S[4]	S[4]
* D[12]	D[12]
* D[4]	D[4]
* D[11]	D[11]
* D[3]	D[3]
* S[11]	S[11]
* S[3]	S[3]
* S[10]	S[10]
* S[2]	S[2]
* D[10]	D[10]
* D[2]	D[2]
* D[9]	D[9]
* D[1]	D[1]
* S[9]	S[9]
* S[1]	S[1]
* S[8]	S[8]
* S[0]	S[0]
* D[8]	D[8]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1042 N_A_27_47#_M1042_d N_D[0]_M1042_g N_VGND_M1042_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1047 N_VGND_M1047_d N_D[8]_M1047_g N_A_27_911#_M1047_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1108 N_A_27_47#_M1108_d N_D[0]_M1108_g N_VGND_M1042_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1118 N_VGND_M1047_d N_D[8]_M1118_g N_A_27_911#_M1118_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1032 N_A_27_47#_M1108_d N_S[0]_M1032_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1020 N_A_27_911#_M1118_s N_S[8]_M1020_g N_Z_M1020_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1041 N_A_27_47#_M1041_d N_S[0]_M1041_g N_Z_M1032_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1104 N_A_27_911#_M1104_d N_S[8]_M1104_g N_Z_M1020_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1081 N_VGND_M1081_d N_S[0]_M1081_g N_A_278_265#_M1081_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1115 N_VGND_M1115_d N_S[8]_M1115_g N_A_278_793#_M1115_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1072 N_A_701_47#_M1072_d N_S[1]_M1072_g N_VGND_M1081_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1039 N_A_701_937#_M1039_d N_S[9]_M1039_g N_VGND_M1115_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1028 N_A_845_69#_M1028_d N_S[1]_M1028_g N_Z_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1048 N_Z_M1048_d N_S[9]_M1048_g N_A_845_915#_M1048_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1037 N_A_845_69#_M1037_d N_S[1]_M1037_g N_Z_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1130 N_Z_M1048_d N_S[9]_M1130_g N_A_845_915#_M1130_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1074 N_VGND_M1074_d N_D[1]_M1074_g N_A_845_69#_M1037_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1026 N_VGND_M1026_d N_D[9]_M1026_g N_A_845_915#_M1130_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1105 N_VGND_M1074_d N_D[1]_M1105_g N_A_845_69#_M1105_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1059 N_VGND_M1026_d N_D[9]_M1059_g N_A_845_915#_M1059_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1117 N_A_1315_47#_M1117_d N_D[2]_M1117_g N_VGND_M1117_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1035 N_A_1315_911#_M1035_d N_D[10]_M1035_g N_VGND_M1035_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1127 N_A_1315_47#_M1127_d N_D[2]_M1127_g N_VGND_M1117_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1109 N_A_1315_911#_M1109_d N_D[10]_M1109_g N_VGND_M1035_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1116 N_Z_M1116_d N_S[2]_M1116_g N_A_1315_47#_M1127_d VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1015 N_Z_M1015_d N_S[10]_M1015_g N_A_1315_911#_M1109_d VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1
+ R=3.46667 SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1151 N_Z_M1116_d N_S[2]_M1151_g N_A_1315_47#_M1151_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1043 N_Z_M1015_d N_S[10]_M1043_g N_A_1315_911#_M1043_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1150 N_VGND_M1150_d N_S[2]_M1150_g N_A_1566_265#_M1150_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1033 N_VGND_M1033_d N_S[10]_M1033_g N_A_1566_793#_M1033_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1019 N_A_1989_47#_M1019_d N_S[3]_M1019_g N_VGND_M1150_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1071 N_A_1989_937#_M1071_d N_S[11]_M1071_g N_VGND_M1033_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1102 N_Z_M1102_d N_S[3]_M1102_g N_A_2133_69#_M1102_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1029 N_Z_M1029_d N_S[11]_M1029_g N_A_2133_915#_M1029_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1125 N_Z_M1102_d N_S[3]_M1125_g N_A_2133_69#_M1125_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1067 N_Z_M1029_d N_S[11]_M1067_g N_A_2133_915#_M1067_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1
+ R=3.46667 SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1025 N_A_2133_69#_M1125_s N_D[3]_M1025_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1011 N_A_2133_915#_M1067_s N_D[11]_M1011_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1156 N_A_2133_69#_M1156_d N_D[3]_M1156_g N_VGND_M1025_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1136 N_A_2133_915#_M1136_d N_D[11]_M1136_g N_VGND_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1057 N_VGND_M1057_d N_D[4]_M1057_g N_A_2603_47#_M1057_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1073 N_VGND_M1073_d N_D[12]_M1073_g N_A_2603_911#_M1073_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1094 N_VGND_M1057_d N_D[4]_M1094_g N_A_2603_47#_M1094_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1103 N_VGND_M1073_d N_D[12]_M1103_g N_A_2603_911#_M1103_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1046 N_Z_M1046_d N_S[4]_M1046_g N_A_2603_47#_M1094_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1000 N_A_2603_911#_M1103_s N_S[12]_M1000_g N_Z_M1000_s VNB NSHORT L=0.15
+ W=0.52 AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1
+ R=3.46667 SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1086 N_Z_M1046_d N_S[4]_M1086_g N_A_2603_47#_M1086_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1128 N_A_2603_911#_M1128_d N_S[12]_M1128_g N_Z_M1000_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1064 N_VGND_M1064_d N_S[4]_M1064_g N_A_2854_265#_M1064_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1063 N_VGND_M1063_d N_S[12]_M1063_g N_A_2854_793#_M1063_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1098 N_A_3277_47#_M1098_d N_S[5]_M1098_g N_VGND_M1064_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1096 N_A_3277_937#_M1096_d N_S[13]_M1096_g N_VGND_M1063_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1022 N_Z_M1022_d N_S[5]_M1022_g N_A_3421_69#_M1022_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1016 N_A_3421_915#_M1016_d N_S[13]_M1016_g N_Z_M1016_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1054 N_Z_M1022_d N_S[5]_M1054_g N_A_3421_69#_M1054_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1146 N_A_3421_915#_M1146_d N_S[13]_M1146_g N_Z_M1016_s VNB NSHORT L=0.15
+ W=0.52 AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1
+ R=3.46667 SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1090 N_VGND_M1090_d N_D[5]_M1090_g N_A_3421_69#_M1054_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1100 N_VGND_M1100_d N_D[13]_M1100_g N_A_3421_915#_M1146_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1110 N_VGND_M1090_d N_D[5]_M1110_g N_A_3421_69#_M1110_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1121 N_VGND_M1100_d N_D[13]_M1121_g N_A_3421_915#_M1121_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1139 N_VGND_M1139_d N_D[6]_M1139_g N_A_3891_47#_M1139_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_D[14]_M1018_g N_A_3891_911#_M1018_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1155 N_VGND_M1139_d N_D[6]_M1155_g N_A_3891_47#_M1155_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1119 N_VGND_M1018_d N_D[14]_M1119_g N_A_3891_911#_M1119_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1112 N_Z_M1112_d N_S[6]_M1112_g N_A_3891_47#_M1155_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1021 N_A_3891_911#_M1119_s N_S[14]_M1021_g N_Z_M1021_s VNB NSHORT L=0.15
+ W=0.52 AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1
+ R=3.46667 SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1145 N_Z_M1112_d N_S[6]_M1145_g N_A_3891_47#_M1145_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1153 N_A_3891_911#_M1153_d N_S[14]_M1153_g N_Z_M1021_s VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75001.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1144 N_VGND_M1144_d N_S[6]_M1144_g N_A_4142_265#_M1144_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1012 N_VGND_M1012_d N_S[14]_M1012_g N_A_4142_793#_M1012_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1017 N_A_4565_47#_M1017_d N_S[7]_M1017_g N_VGND_M1144_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1040 N_A_4565_937#_M1040_d N_S[15]_M1040_g N_VGND_M1012_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1107 N_Z_M1107_d N_S[7]_M1107_g N_A_4709_69#_M1107_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1106 N_Z_M1106_d N_S[15]_M1106_g N_A_4709_915#_M1106_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75001.6 A=0.078 P=1.34 MULT=1
MM1138 N_Z_M1107_d N_S[7]_M1138_g N_A_4709_69#_M1138_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1131 N_Z_M1106_d N_S[15]_M1131_g N_A_4709_915#_M1131_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1
+ R=3.46667 SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1024 N_A_4709_69#_M1138_s N_D[7]_M1024_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1147 N_A_4709_915#_M1131_s N_D[15]_M1147_g N_VGND_M1147_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1050 N_A_4709_69#_M1050_d N_D[7]_M1050_g N_VGND_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1154 N_A_4709_915#_M1154_d N_D[15]_M1154_g N_VGND_M1147_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_27_297#_M1010_d N_D[0]_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1014 N_A_27_591#_M1014_d N_D[8]_M1014_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1075 N_A_27_297#_M1075_d N_D[0]_M1075_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1078 N_A_27_591#_M1078_d N_D[8]_M1078_g N_VPWR_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1013 N_A_27_297#_M1075_d N_A_278_265#_M1013_g N_Z_M1013_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1099 N_A_27_591#_M1078_d N_A_278_793#_M1099_g N_Z_M1099_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1031 N_A_27_297#_M1031_d N_A_278_265#_M1031_g N_Z_M1013_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1111 N_A_27_591#_M1111_d N_A_278_793#_M1111_g N_Z_M1099_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1023 N_VPWR_M1023_d N_S[0]_M1023_g N_A_278_265#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1027 N_VPWR_M1027_d N_S[8]_M1027_g N_A_278_793#_M1027_s VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1089 N_A_701_47#_M1089_d N_S[1]_M1089_g N_VPWR_M1023_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1092 N_A_701_937#_M1092_d N_S[9]_M1092_g N_VPWR_M1027_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1084 N_A_824_333#_M1084_d N_A_701_47#_M1084_g N_Z_M1084_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1036 N_Z_M1036_d N_A_701_937#_M1036_g N_A_824_591#_M1036_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1113 N_A_824_333#_M1113_d N_A_701_47#_M1113_g N_Z_M1084_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1157 N_Z_M1036_d N_A_701_937#_M1157_g N_A_824_591#_M1157_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1052 N_A_824_333#_M1113_d N_D[1]_M1052_g N_VPWR_M1052_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1056 N_A_824_591#_M1157_s N_D[9]_M1056_g N_VPWR_M1056_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1097 N_A_824_333#_M1097_d N_D[1]_M1097_g N_VPWR_M1052_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1101 N_A_824_591#_M1101_d N_D[9]_M1101_g N_VPWR_M1056_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_D[2]_M1003_g N_A_1315_297#_M1003_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_D[10]_M1009_g N_A_1315_591#_M1009_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1120 N_VPWR_M1003_d N_D[2]_M1120_g N_A_1315_297#_M1120_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1126 N_VPWR_M1009_d N_D[10]_M1126_g N_A_1315_591#_M1126_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1005 N_Z_M1005_d N_A_1566_265#_M1005_g N_A_1315_297#_M1120_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1044 N_A_1315_591#_M1126_s N_A_1566_793#_M1044_g N_Z_M1044_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1124 N_Z_M1005_d N_A_1566_265#_M1124_g N_A_1315_297#_M1124_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1095 N_A_1315_591#_M1095_d N_A_1566_793#_M1095_g N_Z_M1044_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1133 N_VPWR_M1133_d N_S[2]_M1133_g N_A_1566_265#_M1133_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1137 N_VPWR_M1137_d N_S[10]_M1137_g N_A_1566_793#_M1137_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1053 N_A_1989_47#_M1053_d N_S[3]_M1053_g N_VPWR_M1133_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1060 N_A_1989_937#_M1060_d N_S[11]_M1060_g N_VPWR_M1137_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_1989_47#_M1004_g N_A_2112_333#_M1004_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1045 N_A_2112_591#_M1045_d N_A_1989_937#_M1045_g N_Z_M1045_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1123 N_Z_M1004_d N_A_1989_47#_M1123_g N_A_2112_333#_M1123_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1093 N_A_2112_591#_M1093_d N_A_1989_937#_M1093_g N_Z_M1045_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1002 N_VPWR_M1002_d N_D[3]_M1002_g N_A_2112_333#_M1123_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_D[11]_M1008_g N_A_2112_591#_M1093_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1135 N_VPWR_M1002_d N_D[3]_M1135_g N_A_2112_333#_M1135_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1141 N_VPWR_M1008_d N_D[11]_M1141_g N_A_2112_591#_M1141_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1030 N_A_2603_297#_M1030_d N_D[4]_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1038 N_A_2603_591#_M1038_d N_D[12]_M1038_g N_VPWR_M1038_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1080 N_A_2603_297#_M1080_d N_D[4]_M1080_g N_VPWR_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1088 N_A_2603_591#_M1088_d N_D[12]_M1088_g N_VPWR_M1038_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1034 N_A_2603_297#_M1080_d N_A_2854_265#_M1034_g N_Z_M1034_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1114 N_A_2603_591#_M1088_d N_A_2854_793#_M1114_g N_Z_M1114_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1083 N_A_2603_297#_M1083_d N_A_2854_265#_M1083_g N_Z_M1034_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1159 N_A_2603_591#_M1159_d N_A_2854_793#_M1159_g N_Z_M1114_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1001 N_VPWR_M1001_d N_S[4]_M1001_g N_A_2854_265#_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_S[12]_M1007_g N_A_2854_793#_M1007_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1065 N_A_3277_47#_M1065_d N_S[5]_M1065_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1070 N_A_3277_937#_M1070_d N_S[13]_M1070_g N_VPWR_M1007_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1055 N_A_3400_333#_M1055_d N_A_3277_47#_M1055_g N_Z_M1055_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1134 N_A_3400_591#_M1134_d N_A_3277_937#_M1134_g N_Z_M1134_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1082 N_A_3400_333#_M1082_d N_A_3277_47#_M1082_g N_Z_M1055_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1158 N_A_3400_591#_M1158_d N_A_3277_937#_M1158_g N_Z_M1134_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1051 N_A_3400_333#_M1082_d N_D[5]_M1051_g N_VPWR_M1051_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1058 N_A_3400_591#_M1158_d N_D[13]_M1058_g N_VPWR_M1058_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1079 N_A_3400_333#_M1079_d N_D[5]_M1079_g N_VPWR_M1051_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1087 N_A_3400_591#_M1087_d N_D[13]_M1087_g N_VPWR_M1058_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1062 N_A_3891_297#_M1062_d N_D[6]_M1062_g N_VPWR_M1062_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1069 N_A_3891_591#_M1069_d N_D[14]_M1069_g N_VPWR_M1069_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1143 N_A_3891_297#_M1143_d N_D[6]_M1143_g N_VPWR_M1062_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1152 N_A_3891_591#_M1152_d N_D[14]_M1152_g N_VPWR_M1069_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1066 N_A_3891_297#_M1143_d N_A_4142_265#_M1066_g N_Z_M1066_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1006 N_Z_M1006_d N_A_4142_793#_M1006_g N_A_3891_591#_M1152_d VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1091 N_A_3891_297#_M1091_d N_A_4142_265#_M1091_g N_Z_M1066_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1140 N_Z_M1006_d N_A_4142_793#_M1140_g N_A_3891_591#_M1140_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1077 N_VPWR_M1077_d N_S[6]_M1077_g N_A_4142_265#_M1077_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1085 N_VPWR_M1085_d N_S[14]_M1085_g N_A_4142_793#_M1085_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1129 N_A_4565_47#_M1129_d N_S[7]_M1129_g N_VPWR_M1077_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1132 N_A_4565_937#_M1132_d N_S[15]_M1132_g N_VPWR_M1085_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1122 N_A_4688_333#_M1122_d N_A_4565_47#_M1122_g N_Z_M1122_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1049 N_A_4688_591#_M1049_d N_A_4565_937#_M1049_g N_Z_M1049_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1148 N_A_4688_333#_M1148_d N_A_4565_47#_M1148_g N_Z_M1122_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1076 N_A_4688_591#_M1076_d N_A_4565_937#_M1076_g N_Z_M1049_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182
+ M=1 R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1061 N_A_4688_333#_M1148_d N_D[7]_M1061_g N_VPWR_M1061_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1068 N_A_4688_591#_M1076_d N_D[15]_M1068_g N_VPWR_M1068_s VPB PHIGHVT L=0.18
+ W=1 AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1142 N_A_4688_333#_M1142_d N_D[7]_M1142_g N_VPWR_M1061_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1149 N_A_4688_591#_M1149_d N_D[15]_M1149_g N_VPWR_M1068_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX160_noxref VNB VPB NWDIODE A=73.9762 P=57.94
c_495 VNB 0 0.00218386f $X=25.445 $Y=5.355
*
.include "sky130_fd_sc_hdll__muxb16to1_2.pxi.spice"
*
.ends
*
*
