* File: sky130_fd_sc_hdll__sdfxtp_1.spice
* Created: Wed Sep  2 08:52:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__sdfxtp_1.pex.spice"
.subckt sky130_fd_sc_hdll__sdfxtp_1  VNB VPB CLK SCE D SCD VPWR Q VGND
* 
* VGND	VGND
* Q	Q
* VPWR	VPWR
* SCD	SCD
* D	D
* SCE	SCE
* CLK	CLK
* VPB	VPB
* VNB	VNB
MM1028 N_VGND_M1028_d N_CLK_M1028_g N_A_27_47#_M1028_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1092 PD=0.74 PS=1.36 NRD=12.852 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1007 N_A_203_47#_M1007_d N_A_27_47#_M1007_g N_VGND_M1028_d VNB NSHORT L=0.15
+ W=0.42 AD=0.1302 AS=0.0672 PD=1.46 PS=0.74 NRD=12.852 NRS=0 M=1 R=2.8
+ SA=75000.7 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1013 N_VGND_M1013_d N_SCE_M1013_g N_A_319_47#_M1013_s VNB NSHORT L=0.15 W=0.42
+ AD=0.063 AS=0.1428 PD=0.72 PS=1.52 NRD=4.284 NRS=15.708 M=1 R=2.8 SA=75000.3
+ SB=75002.2 A=0.063 P=1.14 MULT=1
MM1021 A_507_47# N_A_319_47#_M1021_g N_VGND_M1013_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0819 AS=0.063 PD=0.81 PS=0.72 NRD=39.996 NRS=1.428 M=1 R=2.8 SA=75000.7
+ SB=75001.7 A=0.063 P=1.14 MULT=1
MM1003 N_A_608_369#_M1003_d N_D_M1003_g A_507_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.0819 PD=0.8 PS=0.81 NRD=14.28 NRS=39.996 M=1 R=2.8 SA=75001.3
+ SB=75001.2 A=0.063 P=1.14 MULT=1
MM1029 A_721_47# N_SCE_M1029_g N_A_608_369#_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0483 AS=0.0798 PD=0.65 PS=0.8 NRD=17.136 NRS=14.28 M=1 R=2.8 SA=75001.8
+ SB=75000.7 A=0.063 P=1.14 MULT=1
MM1020 N_VGND_M1020_d N_SCD_M1020_g A_721_47# VNB NSHORT L=0.15 W=0.42 AD=0.1512
+ AS=0.0483 PD=1.56 PS=0.65 NRD=21.42 NRS=17.136 M=1 R=2.8 SA=75002.2 SB=75000.3
+ A=0.063 P=1.14 MULT=1
MM1026 N_A_1011_47#_M1026_d N_A_27_47#_M1026_g N_A_608_369#_M1026_s VNB NSHORT
+ L=0.15 W=0.36 AD=0.0684 AS=0.1008 PD=0.74 PS=1.28 NRD=34.992 NRS=4.992 M=1
+ R=2.4 SA=75000.2 SB=75003.7 A=0.054 P=1.02 MULT=1
MM1023 A_1117_47# N_A_203_47#_M1023_g N_A_1011_47#_M1026_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0667385 AS=0.0684 PD=0.72 PS=0.74 NRD=43.452 NRS=0 M=1 R=2.4
+ SA=75000.7 SB=75003.1 A=0.054 P=1.02 MULT=1
MM1005 N_VGND_M1005_d N_A_1189_21#_M1005_g A_1117_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.12386 AS=0.0778615 PD=0.978679 PS=0.84 NRD=69.996 NRS=37.248 M=1 R=2.8
+ SA=75001.1 SB=75002.4 A=0.063 P=1.14 MULT=1
MM1012 N_A_1189_21#_M1012_d N_A_1011_47#_M1012_g N_VGND_M1005_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.134656 AS=0.18874 PD=1.3184 PS=1.49132 NRD=21.552
+ NRS=13.116 M=1 R=4.26667 SA=75001.3 SB=75001.1 A=0.096 P=1.58 MULT=1
MM1018 N_A_1474_413#_M1018_d N_A_203_47#_M1018_g N_A_1189_21#_M1012_d VNB NSHORT
+ L=0.15 W=0.36 AD=0.0675 AS=0.075744 PD=0.735 PS=0.7416 NRD=33.324 NRS=0 M=1
+ R=2.4 SA=75002.5 SB=75001.4 A=0.054 P=1.02 MULT=1
MM1027 A_1581_47# N_A_27_47#_M1027_g N_A_1474_413#_M1018_d VNB NSHORT L=0.15
+ W=0.36 AD=0.0617538 AS=0.0675 PD=0.692308 PS=0.735 NRD=38.844 NRS=0 M=1 R=2.4
+ SA=75003.1 SB=75000.8 A=0.054 P=1.02 MULT=1
MM1008 N_VGND_M1008_d N_A_1647_21#_M1008_g A_1581_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1785 AS=0.0720462 PD=1.69 PS=0.807692 NRD=45.708 NRS=33.288 M=1 R=2.8
+ SA=75003.1 SB=75000.3 A=0.063 P=1.14 MULT=1
MM1001 N_VGND_M1001_d N_A_1474_413#_M1001_g N_A_1647_21#_M1001_s VNB NSHORT
+ L=0.15 W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1
+ R=4.33333 SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1031 N_Q_M1031_d N_A_1647_21#_M1031_g N_VGND_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_CLK_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1017 N_A_203_47#_M1017_d N_A_27_47#_M1017_g N_VPWR_M1002_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1009 N_VPWR_M1009_d N_SCE_M1009_g N_A_319_47#_M1009_s VPB PHIGHVT L=0.18
+ W=0.64 AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90002.2 A=0.1152 P=1.64 MULT=1
MM1006 A_504_369# N_SCE_M1006_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1088 AS=0.0928 PD=0.98 PS=0.93 NRD=35.3812 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90001.7 A=0.1152 P=1.64 MULT=1
MM1030 N_A_608_369#_M1030_d N_D_M1030_g A_504_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1088 PD=0.93 PS=0.98 NRD=1.5366 NRS=35.3812 M=1 R=3.55556
+ SA=90001.2 SB=90001.2 A=0.1152 P=1.64 MULT=1
MM1022 A_702_369# N_A_319_47#_M1022_g N_A_608_369#_M1030_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1072 AS=0.0928 PD=0.975 PS=0.93 NRD=34.6129 NRS=1.5366 M=1
+ R=3.55556 SA=90001.6 SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1019 N_VPWR_M1019_d N_SCD_M1019_g A_702_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1888 AS=0.1072 PD=1.87 PS=0.975 NRD=9.2196 NRS=34.6129 M=1 R=3.55556
+ SA=90002.2 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1014 N_A_1011_47#_M1014_d N_A_203_47#_M1014_g N_A_608_369#_M1014_s VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.07035 AS=0.1344 PD=0.755 PS=1.48 NRD=14.0658 NRS=25.7873
+ M=1 R=2.33333 SA=90000.2 SB=90003.6 A=0.0756 P=1.2 MULT=1
MM1011 A_1121_413# N_A_27_47#_M1011_g N_A_1011_47#_M1014_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.0735 AS=0.07035 PD=0.77 PS=0.755 NRD=56.2829 NRS=11.7215 M=1
+ R=2.33333 SA=90000.7 SB=90003.1 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A_1189_21#_M1000_g A_1121_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.128585 AS=0.0735 PD=0.908205 PS=0.77 NRD=99.6623 NRS=56.2829 M=1
+ R=2.33333 SA=90001.3 SB=90002.6 A=0.0756 P=1.2 MULT=1
MM1025 N_A_1189_21#_M1025_d N_A_1011_47#_M1025_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.75 AD=0.155096 AS=0.229615 PD=1.42308 PS=1.62179 NRD=1.3002
+ NRS=6.5601 M=1 R=4.16667 SA=90001.3 SB=90001.1 A=0.135 P=1.86 MULT=1
MM1004 N_A_1474_413#_M1004_d N_A_27_47#_M1004_g N_A_1189_21#_M1025_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.063 AS=0.0868538 PD=0.72 PS=0.796923 NRD=2.3443 NRS=35.1645
+ M=1 R=2.33333 SA=90002.5 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1015 A_1570_413# N_A_203_47#_M1015_g N_A_1474_413#_M1004_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.08295 AS=0.063 PD=0.815 PS=0.72 NRD=66.8224 NRS=7.0329 M=1
+ R=2.33333 SA=90003 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1010 N_VPWR_M1010_d N_A_1647_21#_M1010_g A_1570_413# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1617 AS=0.08295 PD=1.61 PS=0.815 NRD=53.9386 NRS=66.8224 M=1 R=2.33333
+ SA=90003.6 SB=90000.3 A=0.0756 P=1.2 MULT=1
MM1024 N_VPWR_M1024_d N_A_1474_413#_M1024_g N_A_1647_21#_M1024_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.2 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1016 N_Q_M1016_d N_A_1647_21#_M1016_g N_VPWR_M1024_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=17.5908 P=25.13
c_193 VPB 0 3.04607e-19 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__sdfxtp_1.pxi.spice"
*
.ends
*
*
