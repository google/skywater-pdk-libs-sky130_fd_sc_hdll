* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdfbbp_1 CLK D RESET_B SCD SCE SET_B VGND VNB VPB VPWR
+ Q Q_N
X0 a_1469_329# a_1525_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X1 a_1353_47# a_1003_47# a_1197_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X2 a_1769_47# a_211_363# a_1864_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X3 VGND a_2845_47# Q VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1525_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X5 VPWR SCD a_409_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X6 a_1864_47# a_211_363# a_1968_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X7 VGND SET_B a_1353_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X9 a_1710_329# a_27_47# a_1864_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 a_453_315# SCE VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X11 a_453_315# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 a_1105_413# a_1197_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X13 a_1121_47# a_1197_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 a_1992_47# a_2058_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X15 VPWR a_2845_47# Q VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VGND SCD a_411_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 a_483_47# a_211_363# a_1003_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X18 VPWR SET_B a_1197_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X19 VGND a_27_47# a_211_363# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X20 a_824_47# D a_483_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1197_21# a_1003_47# a_1469_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X22 a_1968_413# a_2058_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X23 a_1003_47# a_211_363# a_1121_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X24 a_2845_47# a_2058_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X25 a_810_413# D a_483_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X26 a_1525_21# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X27 a_27_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X28 a_2845_47# a_2058_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X29 VPWR a_2058_21# Q_N VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X30 a_2058_21# a_1525_21# a_2216_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X31 a_2216_47# a_1864_47# a_2058_21# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X32 VPWR a_27_47# a_211_363# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X33 a_2320_329# a_1525_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X34 a_1864_47# a_27_47# a_1992_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X35 a_1003_47# a_27_47# a_1105_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X36 VPWR SET_B a_2058_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X37 a_409_363# a_453_315# a_483_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X38 VPWR SCE a_810_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X39 VGND a_1197_21# a_1769_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X40 VGND a_453_315# a_824_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X41 a_1197_21# a_1525_21# a_1353_47# VNB sky130_fd_pr__nfet_01v8 w=640000u l=150000u
X42 a_411_47# SCE a_483_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X43 a_483_47# a_27_47# a_1003_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X44 a_2058_21# a_1864_47# a_2320_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X45 VGND a_2058_21# Q_N VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 VPWR a_1197_21# a_1710_329# VPB sky130_fd_pr__pfet_01v8_hvt w=840000u l=180000u
X47 VGND SET_B a_2216_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
