* NGSPICE file created from sky130_fd_sc_hdll__clkinv_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__clkinv_2 A VGND VNB VPB VPWR Y
M1000 VGND A Y VNB nshort w=420000u l=150000u
+  ad=2.415e+11p pd=2.83e+06u as=1.386e+11p ps=1.5e+06u
M1001 Y A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.9e+11p pd=5.18e+06u as=5.75e+11p ps=5.15e+06u
M1002 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1003 Y A VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VPWR A Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

