* File: sky130_fd_sc_hdll__o22a_1.pex.spice
* Created: Thu Aug 27 19:20:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22A_1%A_83_21# 1 2 7 9 10 12 16 19 20 21 22 24 27
+ 28
c66 27 0 8.11014e-20 $X=1.64 $Y=0.73
c67 16 0 1.4405e-19 $X=0.62 $Y=1.16
r68 27 28 10.1417 $w=2.48e-07 $l=2e-07 $layer=LI1_cond $X=1.64 $Y=0.77 $X2=1.44
+ $Y2=0.77
r69 22 31 2.53261 $w=4.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.04 $Y=1.705
+ $X2=2.04 $Y2=1.6
r70 22 24 15.1418 $w=4.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.04 $Y=1.705
+ $X2=2.04 $Y2=2.3
r71 20 31 5.66822 $w=2.1e-07 $l=2.35e-07 $layer=LI1_cond $X=1.805 $Y=1.6
+ $X2=2.04 $Y2=1.6
r72 20 21 49.9091 $w=2.08e-07 $l=9.45e-07 $layer=LI1_cond $X=1.805 $Y=1.6
+ $X2=0.86 $Y2=1.6
r73 19 28 35.7374 $w=1.78e-07 $l=5.8e-07 $layer=LI1_cond $X=0.86 $Y=0.805
+ $X2=1.44 $Y2=0.805
r74 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r75 14 21 7.23431 $w=2.1e-07 $l=2.09007e-07 $layer=LI1_cond $X=0.697 $Y=1.495
+ $X2=0.86 $Y2=1.6
r76 14 16 11.879 $w=3.23e-07 $l=3.35e-07 $layer=LI1_cond $X=0.697 $Y=1.495
+ $X2=0.697 $Y2=1.16
r77 13 19 7.57412 $w=1.8e-07 $l=2.03074e-07 $layer=LI1_cond $X=0.697 $Y=0.895
+ $X2=0.86 $Y2=0.805
r78 13 16 9.39684 $w=3.23e-07 $l=2.65e-07 $layer=LI1_cond $X=0.697 $Y=0.895
+ $X2=0.697 $Y2=1.16
r79 10 17 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.585 $Y2=1.16
r80 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r81 7 17 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.585 $Y2=1.16
r82 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
r83 2 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.485 $X2=2.11 $Y2=1.62
r84 2 24 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.965
+ $Y=1.485 $X2=2.11 $Y2=2.3
r85 1 27 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=1.505
+ $Y=0.235 $X2=1.64 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%B1 1 3 4 6 7 15
r29 7 15 2.0744 $w=2.48e-07 $l=4.5e-08 $layer=LI1_cond $X=1.37 $Y=1.2 $X2=1.415
+ $Y2=1.2
r30 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r31 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.37 $Y2=1.16
r32 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
r33 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.405 $Y=1.41
+ $X2=1.37 $Y2=1.16
r34 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.405 $Y=1.41
+ $X2=1.405 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%B2 1 3 4 6 7
r33 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.91
+ $Y=1.16 $X2=1.91 $Y2=1.16
r34 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.875 $Y=1.41
+ $X2=1.91 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.875 $Y=1.41
+ $X2=1.875 $Y2=1.985
r36 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.85 $Y=0.995
+ $X2=1.91 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.85 $Y=0.995 $X2=1.85
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%A2 1 3 4 6 9 13
c39 1 0 8.11014e-20 $X=2.44 $Y=0.995
r40 12 13 28.5492 $w=2.18e-07 $l=5.45e-07 $layer=LI1_cond $X=2.555 $Y=1.325
+ $X2=2.555 $Y2=1.87
r41 9 12 7.04571 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=2.5 $Y=1.16 $X2=2.5
+ $Y2=1.325
r42 9 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.5 $Y=1.16
+ $X2=2.5 $Y2=1.16
r43 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.465 $Y=1.41
+ $X2=2.5 $Y2=1.16
r44 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.465 $Y=1.41
+ $X2=2.465 $Y2=1.985
r45 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=2.44 $Y=0.995
+ $X2=2.5 $Y2=1.16
r46 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.44 $Y=0.995 $X2=2.44
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%A1 1 3 4 6 7 15
r22 7 15 4.71364 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3 $Y=1.175 $X2=3.085
+ $Y2=1.175
r23 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r24 4 10 49.9093 $w=2.71e-07 $l=2.7157e-07 $layer=POLY_cond $X=2.945 $Y=1.41
+ $X2=2.99 $Y2=1.16
r25 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.945 $Y=1.41
+ $X2=2.945 $Y2=1.985
r26 1 10 38.8824 $w=2.71e-07 $l=1.96914e-07 $layer=POLY_cond $X=2.92 $Y=0.995
+ $X2=2.99 $Y2=1.16
r27 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.92 $Y=0.995 $X2=2.92
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%X 1 2 7 10
r14 10 13 42.1876 $w=2.78e-07 $l=1.025e-06 $layer=LI1_cond $X=0.225 $Y=0.595
+ $X2=0.225 $Y2=1.62
r15 7 17 3.70428 $w=2.78e-07 $l=9e-08 $layer=LI1_cond $X=0.225 $Y=2.21 $X2=0.225
+ $Y2=2.3
r16 7 13 24.2836 $w=2.78e-07 $l=5.9e-07 $layer=LI1_cond $X=0.225 $Y=2.21
+ $X2=0.225 $Y2=1.62
r17 2 17 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
r18 2 13 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r19 1 10 182 $w=1.7e-07 $l=4.17852e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.595
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%VPWR 1 2 9 11 13 17 19 24 30 34
c42 1 0 1.4405e-19 $X=0.605 $Y=1.485
r43 34 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r44 33 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 33 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 28 36 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r48 28 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r49 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r50 25 30 14.2108 $w=1.7e-07 $l=3.78e-07 $layer=LI1_cond $X=1.36 $Y=2.72
+ $X2=0.982 $Y2=2.72
r51 25 27 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=1.36 $Y=2.72
+ $X2=1.61 $Y2=2.72
r52 24 33 6.69489 $w=1.7e-07 $l=3.47e-07 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=3.332 $Y2=2.72
r53 24 27 89.7059 $w=1.68e-07 $l=1.375e-06 $layer=LI1_cond $X=2.985 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 19 30 14.2108 $w=1.7e-07 $l=3.77e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.982 $Y2=2.72
r55 19 21 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=0.605 $Y=2.72
+ $X2=0.23 $Y2=2.72
r56 17 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r57 17 21 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 13 16 14.6547 $w=5.53e-07 $l=6.8e-07 $layer=LI1_cond $X=3.262 $Y=1.66
+ $X2=3.262 $Y2=2.34
r59 11 33 2.99051 $w=5.55e-07 $l=1.14782e-07 $layer=LI1_cond $X=3.262 $Y=2.635
+ $X2=3.332 $Y2=2.72
r60 11 16 6.35753 $w=5.53e-07 $l=2.95e-07 $layer=LI1_cond $X=3.262 $Y=2.635
+ $X2=3.262 $Y2=2.34
r61 7 30 3.01793 $w=7.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.982 $Y=2.635
+ $X2=0.982 $Y2=2.72
r62 7 9 10.6934 $w=7.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.982 $Y=2.635
+ $X2=0.982 $Y2=1.96
r63 2 16 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.485 $X2=3.18 $Y2=2.34
r64 2 13 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.035
+ $Y=1.485 $X2=3.18 $Y2=1.66
r65 1 9 150 $w=1.7e-07 $l=7.19305e-07 $layer=licon1_PDIFF $count=4 $X=0.605
+ $Y=1.485 $X2=1.125 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%VGND 1 2 11 15 18 19 20 30 31 34
r50 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r51 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r52 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r53 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r54 25 28 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r55 25 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r56 24 27 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.53
+ $Y2=0
r57 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r58 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.785 $Y=0 $X2=0.7
+ $Y2=0
r59 22 24 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.785 $Y=0 $X2=1.15
+ $Y2=0
r60 20 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r61 18 27 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.53
+ $Y2=0
r62 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.625 $Y=0 $X2=2.71
+ $Y2=0
r63 17 30 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=2.795 $Y=0 $X2=3.45
+ $Y2=0
r64 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0 $X2=2.71
+ $Y2=0
r65 13 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0
r66 13 15 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0.36
r67 9 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r68 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0.38
r69 2 15 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.71 $Y2=0.36
r70 1 11 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.565
+ $Y=0.235 $X2=0.7 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_1%A_219_47# 1 2 3 10 14 15 16 20
r45 18 20 9.0127 $w=3.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.16 $Y=0.695
+ $X2=3.16 $Y2=0.39
r46 17 25 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.395 $Y=0.78
+ $X2=2.23 $Y2=0.78
r47 16 18 8.28377 $w=1.7e-07 $l=2.33666e-07 $layer=LI1_cond $X=2.965 $Y=0.78
+ $X2=3.16 $Y2=0.695
r48 16 17 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=2.965 $Y=0.78
+ $X2=2.395 $Y2=0.78
r49 15 25 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.23 $Y=0.695 $X2=2.23
+ $Y2=0.78
r50 14 23 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=2.23 $Y=0.475 $X2=2.23
+ $Y2=0.385
r51 14 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=2.23 $Y=0.475
+ $X2=2.23 $Y2=0.695
r52 10 23 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=0.385
+ $X2=2.23 $Y2=0.385
r53 10 12 52.0657 $w=1.78e-07 $l=8.45e-07 $layer=LI1_cond $X=2.065 $Y=0.385
+ $X2=1.22 $Y2=0.385
r54 3 20 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=2.995
+ $Y=0.235 $X2=3.18 $Y2=0.39
r55 2 25 182 $w=1.7e-07 $l=6.29285e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.23 $Y2=0.73
r56 2 23 182 $w=1.7e-07 $l=3.74566e-07 $layer=licon1_NDIFF $count=1 $X=1.925
+ $Y=0.235 $X2=2.23 $Y2=0.39
r57 1 12 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.095
+ $Y=0.235 $X2=1.22 $Y2=0.39
.ends

