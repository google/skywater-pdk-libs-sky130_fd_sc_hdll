* File: sky130_fd_sc_hdll__o21bai_4.pxi.spice
* Created: Wed Sep  2 08:44:23 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%B1_N N_B1_N_c_107_n N_B1_N_M1008_g
+ N_B1_N_c_108_n N_B1_N_M1009_g B1_N B1_N PM_SKY130_FD_SC_HDLL__O21BAI_4%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%A_33_297# N_A_33_297#_M1009_d
+ N_A_33_297#_M1008_s N_A_33_297#_c_143_n N_A_33_297#_M1001_g
+ N_A_33_297#_c_144_n N_A_33_297#_M1011_g N_A_33_297#_c_133_n
+ N_A_33_297#_M1006_g N_A_33_297#_c_145_n N_A_33_297#_M1014_g
+ N_A_33_297#_c_134_n N_A_33_297#_M1013_g N_A_33_297#_c_146_n
+ N_A_33_297#_M1021_g N_A_33_297#_c_135_n N_A_33_297#_M1019_g
+ N_A_33_297#_c_136_n N_A_33_297#_M1024_g N_A_33_297#_c_147_n
+ N_A_33_297#_c_148_n N_A_33_297#_c_149_n N_A_33_297#_c_137_n
+ N_A_33_297#_c_138_n N_A_33_297#_c_139_n N_A_33_297#_c_190_p
+ N_A_33_297#_c_140_n N_A_33_297#_c_141_n N_A_33_297#_c_142_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_4%A_33_297#
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%A2 N_A2_c_231_n N_A2_M1004_g N_A2_c_237_n
+ N_A2_M1002_g N_A2_c_232_n N_A2_M1010_g N_A2_c_238_n N_A2_M1012_g N_A2_c_233_n
+ N_A2_M1017_g N_A2_c_239_n N_A2_M1016_g N_A2_c_240_n N_A2_M1025_g N_A2_c_234_n
+ N_A2_M1018_g A2 N_A2_c_235_n N_A2_c_236_n A2 PM_SKY130_FD_SC_HDLL__O21BAI_4%A2
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%A1 N_A1_c_317_n N_A1_M1005_g N_A1_c_323_n
+ N_A1_M1000_g N_A1_c_318_n N_A1_M1007_g N_A1_c_324_n N_A1_M1003_g N_A1_c_319_n
+ N_A1_M1020_g N_A1_c_325_n N_A1_M1015_g N_A1_c_326_n N_A1_M1022_g N_A1_c_320_n
+ N_A1_M1023_g A1 A1 N_A1_c_322_n A1 PM_SKY130_FD_SC_HDLL__O21BAI_4%A1
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%VPWR N_VPWR_M1008_d N_VPWR_M1011_s
+ N_VPWR_M1021_s N_VPWR_M1000_s N_VPWR_M1015_s N_VPWR_c_393_n N_VPWR_c_394_n
+ N_VPWR_c_395_n N_VPWR_c_396_n N_VPWR_c_397_n N_VPWR_c_398_n N_VPWR_c_399_n
+ N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n N_VPWR_c_403_n N_VPWR_c_404_n
+ N_VPWR_c_405_n N_VPWR_c_406_n VPWR N_VPWR_c_407_n N_VPWR_c_392_n
+ N_VPWR_c_409_n PM_SKY130_FD_SC_HDLL__O21BAI_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%Y N_Y_M1006_s N_Y_M1019_s N_Y_M1001_d
+ N_Y_M1014_d N_Y_M1002_d N_Y_M1016_d N_Y_c_494_n N_Y_c_502_n N_Y_c_495_n
+ N_Y_c_513_n N_Y_c_551_n N_Y_c_575_p N_Y_c_496_n N_Y_c_497_n N_Y_c_498_n
+ N_Y_c_499_n N_Y_c_500_n Y N_Y_c_493_n PM_SKY130_FD_SC_HDLL__O21BAI_4%Y
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%A_621_297# N_A_621_297#_M1002_s
+ N_A_621_297#_M1012_s N_A_621_297#_M1025_s N_A_621_297#_M1003_d
+ N_A_621_297#_M1022_d N_A_621_297#_c_580_n N_A_621_297#_c_588_n
+ N_A_621_297#_c_581_n N_A_621_297#_c_639_n N_A_621_297#_c_590_n
+ N_A_621_297#_c_582_n N_A_621_297#_c_618_n N_A_621_297#_c_583_n
+ N_A_621_297#_c_622_n N_A_621_297#_c_584_n N_A_621_297#_c_585_n
+ N_A_621_297#_c_626_n N_A_621_297#_c_628_n N_A_621_297#_c_586_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_4%A_621_297#
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%VGND N_VGND_M1009_s N_VGND_M1004_s
+ N_VGND_M1017_s N_VGND_M1005_d N_VGND_M1020_d N_VGND_c_645_n N_VGND_c_646_n
+ N_VGND_c_647_n N_VGND_c_648_n N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n
+ N_VGND_c_652_n N_VGND_c_653_n N_VGND_c_654_n N_VGND_c_655_n N_VGND_c_656_n
+ N_VGND_c_657_n N_VGND_c_658_n VGND N_VGND_c_659_n N_VGND_c_660_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_4%VGND
x_PM_SKY130_FD_SC_HDLL__O21BAI_4%A_245_47# N_A_245_47#_M1006_d
+ N_A_245_47#_M1013_d N_A_245_47#_M1024_d N_A_245_47#_M1010_d
+ N_A_245_47#_M1018_d N_A_245_47#_M1007_s N_A_245_47#_M1023_s
+ N_A_245_47#_c_750_n N_A_245_47#_c_767_n N_A_245_47#_c_751_n
+ N_A_245_47#_c_752_n N_A_245_47#_c_775_n N_A_245_47#_c_753_n
+ N_A_245_47#_c_783_n N_A_245_47#_c_754_n N_A_245_47#_c_797_n
+ N_A_245_47#_c_755_n N_A_245_47#_c_756_n N_A_245_47#_c_757_n
+ N_A_245_47#_c_758_n N_A_245_47#_c_759_n
+ PM_SKY130_FD_SC_HDLL__O21BAI_4%A_245_47#
cc_1 VNB N_B1_N_c_107_n 0.0415843f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.41
cc_2 VNB N_B1_N_c_108_n 0.0249175f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.995
cc_3 VNB B1_N 0.0151212f $X=-0.19 $Y=-0.24 $X2=0.375 $Y2=1.19
cc_4 VNB N_A_33_297#_c_133_n 0.020602f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VNB N_A_33_297#_c_134_n 0.016968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_33_297#_c_135_n 0.0169283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_33_297#_c_136_n 0.0166801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_33_297#_c_137_n 0.005897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_33_297#_c_138_n 0.00315117f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_33_297#_c_139_n 3.44862e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_33_297#_c_140_n 0.00319326f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_33_297#_c_141_n 0.00384754f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_33_297#_c_142_n 0.116193f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_231_n 0.0164874f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.41
cc_15 VNB N_A2_c_232_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_16 VNB N_A2_c_233_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A2_c_234_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A2_c_235_n 0.00255635f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_236_n 0.0733814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A1_c_317_n 0.0164927f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.41
cc_21 VNB N_A1_c_318_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_22 VNB N_A1_c_319_n 0.0172028f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_c_320_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB A1 0.026556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A1_c_322_n 0.0801709f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VPWR_c_392_n 0.30769f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB Y 0.00282199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_Y_c_493_n 0.00200357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_645_n 0.012648f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_646_n 0.00618788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_647_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_648_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_649_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_650_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_651_n 0.0794043f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_652_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_653_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_654_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_655_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_656_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_657_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_658_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_659_n 0.02183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_660_n 0.370167f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_245_47#_c_750_n 0.00254893f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_245_47#_c_751_n 0.003225f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_245_47#_c_752_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_245_47#_c_753_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_245_47#_c_754_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_245_47#_c_755_n 0.0132268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_245_47#_c_756_n 0.0187437f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_245_47#_c_757_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_245_47#_c_758_n 0.00384439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_245_47#_c_759_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VPB N_B1_N_c_107_n 0.036326f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.41
cc_56 VPB N_A_33_297#_c_143_n 0.0162716f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_57 VPB N_A_33_297#_c_144_n 0.0159554f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_58 VPB N_A_33_297#_c_145_n 0.015974f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_33_297#_c_146_n 0.0192137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_33_297#_c_147_n 0.00924758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_33_297#_c_148_n 0.0308647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_33_297#_c_149_n 7.41046e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_33_297#_c_139_n 0.00270647f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_33_297#_c_142_n 0.0625916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A2_c_237_n 0.0192297f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=0.995
cc_66 VPB N_A2_c_238_n 0.0158906f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_67 VPB N_A2_c_239_n 0.0158911f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A2_c_240_n 0.0164196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A2_c_236_n 0.0463124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A1_c_323_n 0.0161059f $X=-0.19 $Y=1.305 $X2=0.57 $Y2=0.995
cc_71 VPB N_A1_c_324_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.345 $Y2=1.16
cc_72 VPB N_A1_c_325_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A1_c_326_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_A1_c_322_n 0.048391f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_393_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_394_n 0.0198475f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_395_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_396_n 0.00518f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_397_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_398_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_399_n 0.0213496f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_400_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_401_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_402_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_403_n 0.0635591f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_404_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_405_n 0.0195604f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_406_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_407_n 0.0225629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_392_n 0.0623712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_409_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_Y_c_494_n 0.0016295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_Y_c_495_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_Y_c_496_n 0.00282553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_Y_c_497_n 0.00192868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_Y_c_498_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_Y_c_499_n 0.0014926f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_Y_c_500_n 0.00188018f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB Y 0.0166889f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_621_297#_c_580_n 0.00612452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_621_297#_c_581_n 0.00248232f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_A_621_297#_c_582_n 0.00362897f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_A_621_297#_c_583_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_A_621_297#_c_584_n 0.00196267f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_A_621_297#_c_585_n 0.00366598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_A_621_297#_c_586_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 N_B1_N_c_107_n N_A_33_297#_c_143_n 0.0200302f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_108 N_B1_N_c_107_n N_A_33_297#_c_147_n 0.00721448f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_109 B1_N N_A_33_297#_c_147_n 0.027158f $X=0.375 $Y=1.19 $X2=0 $Y2=0
cc_110 N_B1_N_c_107_n N_A_33_297#_c_148_n 0.0107663f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_111 N_B1_N_c_107_n N_A_33_297#_c_149_n 0.0161433f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_112 B1_N N_A_33_297#_c_149_n 0.00237761f $X=0.375 $Y=1.19 $X2=0 $Y2=0
cc_113 N_B1_N_c_108_n N_A_33_297#_c_137_n 0.00672357f $X=0.57 $Y=0.995 $X2=0
+ $Y2=0
cc_114 N_B1_N_c_108_n N_A_33_297#_c_138_n 0.00633394f $X=0.57 $Y=0.995 $X2=0
+ $Y2=0
cc_115 N_B1_N_c_107_n N_A_33_297#_c_139_n 0.00417188f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_116 N_B1_N_c_108_n N_A_33_297#_c_140_n 0.00491195f $X=0.57 $Y=0.995 $X2=0
+ $Y2=0
cc_117 N_B1_N_c_107_n N_A_33_297#_c_141_n 0.00202946f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_118 B1_N N_A_33_297#_c_141_n 0.0179337f $X=0.375 $Y=1.19 $X2=0 $Y2=0
cc_119 N_B1_N_c_107_n N_A_33_297#_c_142_n 0.0182723f $X=0.545 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_B1_N_c_107_n N_VPWR_c_393_n 0.0058284f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B1_N_c_107_n N_VPWR_c_399_n 0.00674404f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B1_N_c_107_n N_VPWR_c_392_n 0.0128249f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B1_N_c_107_n N_Y_c_502_n 6.60746e-19 $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_N_c_107_n N_VGND_c_646_n 0.00429275f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B1_N_c_108_n N_VGND_c_646_n 0.00671047f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_126 B1_N N_VGND_c_646_n 0.0131644f $X=0.375 $Y=1.19 $X2=0 $Y2=0
cc_127 N_B1_N_c_108_n N_VGND_c_651_n 0.0046926f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_128 N_B1_N_c_108_n N_VGND_c_660_n 0.0101446f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_129 N_A_33_297#_c_136_n N_A2_c_231_n 0.0143687f $X=3.02 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_130 N_A_33_297#_c_142_n N_A2_c_235_n 2.06878e-19 $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_131 N_A_33_297#_c_142_n N_A2_c_236_n 0.0143687f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_33_297#_c_149_n N_VPWR_M1008_d 0.00319401f $X=0.68 $Y=1.54 $X2=-0.19
+ $Y2=-0.24
cc_133 N_A_33_297#_c_143_n N_VPWR_c_393_n 0.00486097f $X=1.015 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A_33_297#_c_148_n N_VPWR_c_393_n 0.0387469f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_135 N_A_33_297#_c_149_n N_VPWR_c_393_n 0.0138849f $X=0.68 $Y=1.54 $X2=0 $Y2=0
cc_136 N_A_33_297#_c_141_n N_VPWR_c_393_n 5.82871e-19 $X=0.812 $Y=1.18 $X2=0
+ $Y2=0
cc_137 N_A_33_297#_c_143_n N_VPWR_c_394_n 0.00597712f $X=1.015 $Y=1.41 $X2=0
+ $Y2=0
cc_138 N_A_33_297#_c_144_n N_VPWR_c_394_n 0.00702461f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_139 N_A_33_297#_c_144_n N_VPWR_c_395_n 0.00300743f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_140 N_A_33_297#_c_145_n N_VPWR_c_395_n 0.00300743f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_33_297#_c_146_n N_VPWR_c_396_n 0.00479105f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_33_297#_c_142_n N_VPWR_c_396_n 5.95839e-19 $X=2.55 $Y=1.202 $X2=0
+ $Y2=0
cc_143 N_A_33_297#_c_148_n N_VPWR_c_399_n 0.0176517f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_144 N_A_33_297#_c_145_n N_VPWR_c_401_n 0.00702461f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_145 N_A_33_297#_c_146_n N_VPWR_c_401_n 0.00702461f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_146 N_A_33_297#_M1008_s N_VPWR_c_392_n 0.00235527f $X=0.165 $Y=1.485 $X2=0
+ $Y2=0
cc_147 N_A_33_297#_c_143_n N_VPWR_c_392_n 0.0100198f $X=1.015 $Y=1.41 $X2=0
+ $Y2=0
cc_148 N_A_33_297#_c_144_n N_VPWR_c_392_n 0.0124092f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_149 N_A_33_297#_c_145_n N_VPWR_c_392_n 0.0124092f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_150 N_A_33_297#_c_146_n N_VPWR_c_392_n 0.0136915f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_A_33_297#_c_148_n N_VPWR_c_392_n 0.0122874f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_152 N_A_33_297#_c_143_n N_Y_c_494_n 0.00379574f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_153 N_A_33_297#_c_149_n N_Y_c_494_n 0.0140017f $X=0.68 $Y=1.54 $X2=0 $Y2=0
cc_154 N_A_33_297#_c_190_p N_Y_c_494_n 0.027498f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_155 N_A_33_297#_c_142_n N_Y_c_494_n 0.00664071f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_156 N_A_33_297#_c_143_n N_Y_c_502_n 0.0136295f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A_33_297#_c_148_n N_Y_c_502_n 0.00476769f $X=0.31 $Y=2.3 $X2=0 $Y2=0
cc_158 N_A_33_297#_c_144_n N_Y_c_495_n 0.0156273f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_33_297#_c_145_n N_Y_c_495_n 0.0156202f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_33_297#_c_190_p N_Y_c_495_n 0.0486996f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_161 N_A_33_297#_c_142_n N_Y_c_495_n 0.00878951f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_162 N_A_33_297#_c_133_n N_Y_c_513_n 0.00930809f $X=1.61 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_33_297#_c_134_n N_Y_c_513_n 0.00917588f $X=2.08 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_33_297#_c_135_n N_Y_c_513_n 0.00999491f $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_165 N_A_33_297#_c_190_p N_Y_c_513_n 0.0443969f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_166 N_A_33_297#_c_142_n N_Y_c_513_n 0.00690047f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_167 N_A_33_297#_c_190_p N_Y_c_498_n 0.0204509f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_33_297#_c_142_n N_Y_c_498_n 0.00685366f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_33_297#_c_146_n Y 0.0191827f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_33_297#_c_190_p Y 0.0316614f $X=2.25 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_33_297#_c_142_n Y 0.0385826f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_172 N_A_33_297#_c_135_n N_Y_c_493_n 0.00421061f $X=2.55 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_33_297#_c_136_n N_Y_c_493_n 0.00260235f $X=3.02 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_33_297#_c_142_n N_Y_c_493_n 0.0095102f $X=2.55 $Y=1.202 $X2=0 $Y2=0
cc_175 N_A_33_297#_c_142_n N_A_621_297#_c_580_n 2.80671e-19 $X=2.55 $Y=1.202
+ $X2=0 $Y2=0
cc_176 N_A_33_297#_c_137_n N_VGND_c_646_n 0.0451414f $X=0.78 $Y=0.39 $X2=0 $Y2=0
cc_177 N_A_33_297#_c_133_n N_VGND_c_651_n 0.00368123f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_178 N_A_33_297#_c_134_n N_VGND_c_651_n 0.00368123f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_179 N_A_33_297#_c_135_n N_VGND_c_651_n 0.00368123f $X=2.55 $Y=0.995 $X2=0
+ $Y2=0
cc_180 N_A_33_297#_c_136_n N_VGND_c_651_n 0.00368123f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_33_297#_c_137_n N_VGND_c_651_n 0.0199288f $X=0.78 $Y=0.39 $X2=0 $Y2=0
cc_182 N_A_33_297#_M1009_d N_VGND_c_660_n 0.00211145f $X=0.645 $Y=0.235 $X2=0
+ $Y2=0
cc_183 N_A_33_297#_c_133_n N_VGND_c_660_n 0.00670426f $X=1.61 $Y=0.995 $X2=0
+ $Y2=0
cc_184 N_A_33_297#_c_134_n N_VGND_c_660_n 0.00550516f $X=2.08 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_33_297#_c_135_n N_VGND_c_660_n 0.00550516f $X=2.55 $Y=0.995 $X2=0
+ $Y2=0
cc_186 N_A_33_297#_c_136_n N_VGND_c_660_n 0.0054054f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_187 N_A_33_297#_c_137_n N_VGND_c_660_n 0.0138528f $X=0.78 $Y=0.39 $X2=0 $Y2=0
cc_188 N_A_33_297#_c_133_n N_A_245_47#_c_750_n 0.00825287f $X=1.61 $Y=0.995
+ $X2=0 $Y2=0
cc_189 N_A_33_297#_c_134_n N_A_245_47#_c_750_n 0.00825287f $X=2.08 $Y=0.995
+ $X2=0 $Y2=0
cc_190 N_A_33_297#_c_135_n N_A_245_47#_c_750_n 0.00825287f $X=2.55 $Y=0.995
+ $X2=0 $Y2=0
cc_191 N_A_33_297#_c_136_n N_A_245_47#_c_750_n 0.0102764f $X=3.02 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A_33_297#_c_137_n N_A_245_47#_c_750_n 0.0119612f $X=0.78 $Y=0.39 $X2=0
+ $Y2=0
cc_193 N_A_33_297#_c_190_p N_A_245_47#_c_750_n 0.00847565f $X=2.25 $Y=1.16 $X2=0
+ $Y2=0
cc_194 N_A_33_297#_c_142_n N_A_245_47#_c_750_n 0.00665065f $X=2.55 $Y=1.202
+ $X2=0 $Y2=0
cc_195 N_A2_c_234_n N_A1_c_317_n 0.0175841f $X=4.9 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_196 N_A2_c_240_n N_A1_c_323_n 0.00966468f $X=4.875 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A2_c_235_n A1 0.0176526f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_198 N_A2_c_236_n A1 0.00106988f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A2_c_235_n N_A1_c_322_n 2.06428e-19 $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A2_c_236_n N_A1_c_322_n 0.0175841f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_201 N_A2_c_237_n N_VPWR_c_396_n 0.00196069f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A2_c_237_n N_VPWR_c_403_n 0.00429453f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A2_c_238_n N_VPWR_c_403_n 0.00429453f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_c_239_n N_VPWR_c_403_n 0.00429453f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A2_c_240_n N_VPWR_c_403_n 0.00429453f $X=4.875 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_237_n N_VPWR_c_392_n 0.00734734f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_238_n N_VPWR_c_392_n 0.00606499f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_239_n N_VPWR_c_392_n 0.00606499f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_240_n N_VPWR_c_392_n 0.00609021f $X=4.875 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_237_n N_Y_c_496_n 0.0143265f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A2_c_235_n N_Y_c_496_n 0.0145519f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A2_c_236_n N_Y_c_496_n 8.96166e-19 $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_213 N_A2_c_238_n N_Y_c_497_n 0.0133055f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A2_c_239_n N_Y_c_497_n 0.0132328f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A2_c_235_n N_Y_c_497_n 0.0487345f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A2_c_236_n N_Y_c_497_n 0.00876269f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A2_c_235_n N_Y_c_499_n 0.020385f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_218 N_A2_c_236_n N_Y_c_499_n 0.00663436f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_219 N_A2_c_240_n N_Y_c_500_n 6.32035e-19 $X=4.875 $Y=1.41 $X2=0 $Y2=0
cc_220 N_A2_c_235_n N_Y_c_500_n 0.020385f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A2_c_236_n N_Y_c_500_n 0.00642616f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_222 N_A2_c_237_n Y 0.0022548f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A2_c_235_n Y 0.0171514f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_224 N_A2_c_236_n Y 0.00552541f $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_225 N_A2_c_236_n N_Y_c_493_n 4.27419e-19 $X=4.875 $Y=1.202 $X2=0 $Y2=0
cc_226 N_A2_c_237_n N_A_621_297#_c_588_n 0.01161f $X=3.465 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A2_c_238_n N_A_621_297#_c_588_n 0.01161f $X=3.935 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A2_c_239_n N_A_621_297#_c_590_n 0.01161f $X=4.405 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A2_c_240_n N_A_621_297#_c_590_n 0.0143578f $X=4.875 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A2_c_240_n N_A_621_297#_c_582_n 2.98195e-19 $X=4.875 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A2_c_231_n N_VGND_c_647_n 0.00456563f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A2_c_232_n N_VGND_c_647_n 0.00276126f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A2_c_233_n N_VGND_c_648_n 0.00385467f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A2_c_234_n N_VGND_c_648_n 0.00365402f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A2_c_231_n N_VGND_c_651_n 0.00423866f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A2_c_232_n N_VGND_c_653_n 0.00423334f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_237 N_A2_c_233_n N_VGND_c_653_n 0.00423334f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A2_c_234_n N_VGND_c_655_n 0.00396605f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_239 N_A2_c_231_n N_VGND_c_660_n 0.00600634f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A2_c_232_n N_VGND_c_660_n 0.00597024f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A2_c_233_n N_VGND_c_660_n 0.00620835f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A2_c_234_n N_VGND_c_660_n 0.00583042f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_243 N_A2_c_231_n N_A_245_47#_c_767_n 0.00230607f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_244 N_A2_c_231_n N_A_245_47#_c_751_n 0.00513756f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A2_c_232_n N_A_245_47#_c_751_n 4.74935e-19 $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A2_c_235_n N_A_245_47#_c_751_n 0.00228728f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_247 N_A2_c_231_n N_A_245_47#_c_752_n 0.00901745f $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A2_c_232_n N_A_245_47#_c_752_n 0.00895898f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_249 N_A2_c_235_n N_A_245_47#_c_752_n 0.0397461f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A2_c_236_n N_A_245_47#_c_752_n 0.00345541f $X=4.875 $Y=1.202 $X2=0
+ $Y2=0
cc_251 N_A2_c_231_n N_A_245_47#_c_775_n 5.24597e-19 $X=3.44 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A2_c_232_n N_A_245_47#_c_775_n 0.00651696f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_253 N_A2_c_233_n N_A_245_47#_c_775_n 0.00693563f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_254 N_A2_c_234_n N_A_245_47#_c_775_n 5.34196e-19 $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A2_c_233_n N_A_245_47#_c_753_n 0.00929182f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A2_c_234_n N_A_245_47#_c_753_n 0.00650032f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A2_c_235_n N_A_245_47#_c_753_n 0.0399344f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_258 N_A2_c_236_n N_A_245_47#_c_753_n 0.00468948f $X=4.875 $Y=1.202 $X2=0
+ $Y2=0
cc_259 N_A2_c_233_n N_A_245_47#_c_783_n 5.69266e-19 $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A2_c_234_n N_A_245_47#_c_783_n 0.00857123f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A2_c_232_n N_A_245_47#_c_757_n 0.00116636f $X=3.91 $Y=0.995 $X2=0 $Y2=0
cc_262 N_A2_c_233_n N_A_245_47#_c_757_n 0.00116636f $X=4.38 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A2_c_235_n N_A_245_47#_c_757_n 0.0306016f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A2_c_236_n N_A_245_47#_c_757_n 0.00358305f $X=4.875 $Y=1.202 $X2=0
+ $Y2=0
cc_265 N_A2_c_234_n N_A_245_47#_c_758_n 0.00269873f $X=4.9 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A2_c_235_n N_A_245_47#_c_758_n 0.00614022f $X=4.7 $Y=1.16 $X2=0 $Y2=0
cc_267 N_A1_c_323_n N_VPWR_c_397_n 0.00300743f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A1_c_324_n N_VPWR_c_397_n 0.00300743f $X=5.815 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A1_c_325_n N_VPWR_c_398_n 0.00300743f $X=6.285 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A1_c_326_n N_VPWR_c_398_n 0.00300743f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A1_c_323_n N_VPWR_c_403_n 0.00702461f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A1_c_324_n N_VPWR_c_405_n 0.00702461f $X=5.815 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A1_c_325_n N_VPWR_c_405_n 0.00702461f $X=6.285 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A1_c_326_n N_VPWR_c_407_n 0.00702461f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A1_c_323_n N_VPWR_c_392_n 0.0124344f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A1_c_324_n N_VPWR_c_392_n 0.0124092f $X=5.815 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A1_c_325_n N_VPWR_c_392_n 0.0124092f $X=6.285 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A1_c_326_n N_VPWR_c_392_n 0.013408f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_279 A1 N_A_621_297#_c_582_n 0.00771248f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_280 N_A1_c_323_n N_A_621_297#_c_583_n 0.0155666f $X=5.345 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A1_c_324_n N_A_621_297#_c_583_n 0.0156273f $X=5.815 $Y=1.41 $X2=0 $Y2=0
cc_282 A1 N_A_621_297#_c_583_n 0.0487385f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_283 N_A1_c_322_n N_A_621_297#_c_583_n 0.00837544f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_284 N_A1_c_325_n N_A_621_297#_c_584_n 0.0156273f $X=6.285 $Y=1.41 $X2=0 $Y2=0
cc_285 N_A1_c_326_n N_A_621_297#_c_584_n 0.0158328f $X=6.755 $Y=1.41 $X2=0 $Y2=0
cc_286 A1 N_A_621_297#_c_584_n 0.0487385f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_287 N_A1_c_322_n N_A_621_297#_c_584_n 0.00816971f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_288 A1 N_A_621_297#_c_585_n 0.0214236f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_289 A1 N_A_621_297#_c_586_n 0.0204509f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_290 N_A1_c_322_n N_A_621_297#_c_586_n 0.00656533f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_291 N_A1_c_317_n N_VGND_c_649_n 0.00379224f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_292 N_A1_c_318_n N_VGND_c_649_n 0.00276126f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_293 N_A1_c_319_n N_VGND_c_650_n 0.00385467f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_294 N_A1_c_320_n N_VGND_c_650_n 0.00365402f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_295 N_A1_c_317_n N_VGND_c_655_n 0.00423334f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_296 N_A1_c_318_n N_VGND_c_657_n 0.00423334f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_297 N_A1_c_319_n N_VGND_c_657_n 0.00423334f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_298 N_A1_c_320_n N_VGND_c_659_n 0.00396605f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_299 N_A1_c_317_n N_VGND_c_660_n 0.00599324f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_300 N_A1_c_318_n N_VGND_c_660_n 0.00597024f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_301 N_A1_c_319_n N_VGND_c_660_n 0.00620835f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_302 N_A1_c_320_n N_VGND_c_660_n 0.00684747f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_303 N_A1_c_317_n N_A_245_47#_c_783_n 0.00686626f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_304 N_A1_c_318_n N_A_245_47#_c_783_n 5.45498e-19 $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A1_c_317_n N_A_245_47#_c_754_n 0.00901745f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A1_c_318_n N_A_245_47#_c_754_n 0.00901745f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_307 A1 N_A_245_47#_c_754_n 0.0398926f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_308 N_A1_c_322_n N_A_245_47#_c_754_n 0.00345541f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_309 N_A1_c_317_n N_A_245_47#_c_797_n 5.24597e-19 $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_310 N_A1_c_318_n N_A_245_47#_c_797_n 0.00651696f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_311 N_A1_c_319_n N_A_245_47#_c_797_n 0.00693563f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_312 N_A1_c_320_n N_A_245_47#_c_797_n 5.34196e-19 $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_313 N_A1_c_319_n N_A_245_47#_c_755_n 0.00929182f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A1_c_320_n N_A_245_47#_c_755_n 0.00936658f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_315 A1 N_A_245_47#_c_755_n 0.071856f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_316 N_A1_c_322_n N_A_245_47#_c_755_n 0.00468948f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_317 N_A1_c_319_n N_A_245_47#_c_756_n 5.69266e-19 $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A1_c_320_n N_A_245_47#_c_756_n 0.00857123f $X=6.78 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A1_c_317_n N_A_245_47#_c_758_n 0.00112787f $X=5.32 $Y=0.995 $X2=0 $Y2=0
cc_320 A1 N_A_245_47#_c_758_n 0.0108485f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_321 N_A1_c_318_n N_A_245_47#_c_759_n 0.00116636f $X=5.79 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A1_c_319_n N_A_245_47#_c_759_n 0.00116636f $X=6.26 $Y=0.995 $X2=0 $Y2=0
cc_323 A1 N_A_245_47#_c_759_n 0.0307014f $X=6.775 $Y=1.105 $X2=0 $Y2=0
cc_324 N_A1_c_322_n N_A_245_47#_c_759_n 0.00358305f $X=6.755 $Y=1.202 $X2=0
+ $Y2=0
cc_325 N_VPWR_c_392_n N_Y_M1001_d 0.00300692f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_326 N_VPWR_c_392_n N_Y_M1014_d 0.00370124f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_392_n N_Y_M1002_d 0.00232895f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_c_392_n N_Y_M1016_d 0.00232895f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_329 N_VPWR_c_393_n N_Y_c_502_n 0.0495854f $X=0.78 $Y=1.96 $X2=0 $Y2=0
cc_330 N_VPWR_c_394_n N_Y_c_502_n 0.0203479f $X=1.595 $Y=2.72 $X2=0 $Y2=0
cc_331 N_VPWR_c_392_n N_Y_c_502_n 0.012629f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_332 N_VPWR_M1011_s N_Y_c_495_n 0.00187091f $X=1.575 $Y=1.485 $X2=0 $Y2=0
cc_333 N_VPWR_c_395_n N_Y_c_495_n 0.0143191f $X=1.72 $Y=1.96 $X2=0 $Y2=0
cc_334 N_VPWR_c_401_n N_Y_c_551_n 0.0149311f $X=2.535 $Y=2.72 $X2=0 $Y2=0
cc_335 N_VPWR_c_392_n N_Y_c_551_n 0.00955092f $X=7.13 $Y=2.72 $X2=0 $Y2=0
cc_336 N_VPWR_M1021_s Y 0.00359918f $X=2.515 $Y=1.485 $X2=0 $Y2=0
cc_337 N_VPWR_c_396_n Y 0.0179413f $X=2.66 $Y=1.96 $X2=0 $Y2=0
cc_338 N_VPWR_c_392_n N_A_621_297#_M1002_s 0.00217519f $X=7.13 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_339 N_VPWR_c_392_n N_A_621_297#_M1012_s 0.00231264f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_340 N_VPWR_c_392_n N_A_621_297#_M1025_s 0.00297222f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_341 N_VPWR_c_392_n N_A_621_297#_M1003_d 0.00370124f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_342 N_VPWR_c_392_n N_A_621_297#_M1022_d 0.00376247f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_343 N_VPWR_c_396_n N_A_621_297#_c_580_n 0.0312508f $X=2.66 $Y=1.96 $X2=0
+ $Y2=0
cc_344 N_VPWR_c_403_n N_A_621_297#_c_588_n 0.0386815f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_345 N_VPWR_c_392_n N_A_621_297#_c_588_n 0.0239144f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_346 N_VPWR_c_396_n N_A_621_297#_c_581_n 0.0113145f $X=2.66 $Y=1.96 $X2=0
+ $Y2=0
cc_347 N_VPWR_c_403_n N_A_621_297#_c_581_n 0.0219693f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_348 N_VPWR_c_392_n N_A_621_297#_c_581_n 0.0126987f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_349 N_VPWR_c_403_n N_A_621_297#_c_590_n 0.0386815f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_350 N_VPWR_c_392_n N_A_621_297#_c_590_n 0.0239144f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_351 N_VPWR_c_403_n N_A_621_297#_c_618_n 0.015002f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_352 N_VPWR_c_392_n N_A_621_297#_c_618_n 0.00962794f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_353 N_VPWR_M1000_s N_A_621_297#_c_583_n 0.00187091f $X=5.435 $Y=1.485 $X2=0
+ $Y2=0
cc_354 N_VPWR_c_397_n N_A_621_297#_c_583_n 0.0143191f $X=5.58 $Y=1.96 $X2=0
+ $Y2=0
cc_355 N_VPWR_c_405_n N_A_621_297#_c_622_n 0.0149311f $X=6.395 $Y=2.72 $X2=0
+ $Y2=0
cc_356 N_VPWR_c_392_n N_A_621_297#_c_622_n 0.00955092f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_357 N_VPWR_M1015_s N_A_621_297#_c_584_n 0.00187091f $X=6.375 $Y=1.485 $X2=0
+ $Y2=0
cc_358 N_VPWR_c_398_n N_A_621_297#_c_584_n 0.0143191f $X=6.52 $Y=1.96 $X2=0
+ $Y2=0
cc_359 N_VPWR_c_407_n N_A_621_297#_c_626_n 0.0161853f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_360 N_VPWR_c_392_n N_A_621_297#_c_626_n 0.00955092f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_361 N_VPWR_c_403_n N_A_621_297#_c_628_n 0.0149886f $X=5.455 $Y=2.72 $X2=0
+ $Y2=0
cc_362 N_VPWR_c_392_n N_A_621_297#_c_628_n 0.00962421f $X=7.13 $Y=2.72 $X2=0
+ $Y2=0
cc_363 N_Y_c_496_n N_A_621_297#_M1002_s 0.00169948f $X=3.575 $Y=1.535 $X2=-0.19
+ $Y2=-0.24
cc_364 Y N_A_621_297#_M1002_s 0.00190672f $X=2.695 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_365 N_Y_c_497_n N_A_621_297#_M1012_s 0.00187422f $X=4.515 $Y=1.535 $X2=0
+ $Y2=0
cc_366 N_Y_c_496_n N_A_621_297#_c_580_n 0.0100336f $X=3.575 $Y=1.535 $X2=0 $Y2=0
cc_367 Y N_A_621_297#_c_580_n 0.0151689f $X=2.695 $Y=1.445 $X2=0 $Y2=0
cc_368 N_Y_M1002_d N_A_621_297#_c_588_n 0.00352392f $X=3.555 $Y=1.485 $X2=0
+ $Y2=0
cc_369 N_Y_c_496_n N_A_621_297#_c_588_n 0.00387236f $X=3.575 $Y=1.535 $X2=0
+ $Y2=0
cc_370 N_Y_c_497_n N_A_621_297#_c_588_n 0.00387236f $X=4.515 $Y=1.535 $X2=0
+ $Y2=0
cc_371 N_Y_c_499_n N_A_621_297#_c_588_n 0.0134104f $X=3.7 $Y=1.62 $X2=0 $Y2=0
cc_372 N_Y_c_497_n N_A_621_297#_c_639_n 0.0143571f $X=4.515 $Y=1.535 $X2=0 $Y2=0
cc_373 N_Y_M1016_d N_A_621_297#_c_590_n 0.00352392f $X=4.495 $Y=1.485 $X2=0
+ $Y2=0
cc_374 N_Y_c_497_n N_A_621_297#_c_590_n 0.00387236f $X=4.515 $Y=1.535 $X2=0
+ $Y2=0
cc_375 N_Y_c_500_n N_A_621_297#_c_590_n 0.0134104f $X=4.64 $Y=1.62 $X2=0 $Y2=0
cc_376 N_Y_c_500_n N_A_621_297#_c_582_n 0.00226124f $X=4.64 $Y=1.62 $X2=0 $Y2=0
cc_377 N_Y_M1006_s N_VGND_c_660_n 0.00261035f $X=1.685 $Y=0.235 $X2=0 $Y2=0
cc_378 N_Y_M1019_s N_VGND_c_660_n 0.00261035f $X=2.625 $Y=0.235 $X2=0 $Y2=0
cc_379 N_Y_c_513_n N_A_245_47#_M1013_d 0.00436017f $X=2.695 $Y=0.73 $X2=0 $Y2=0
cc_380 N_Y_M1006_s N_A_245_47#_c_750_n 0.00418804f $X=1.685 $Y=0.235 $X2=0 $Y2=0
cc_381 N_Y_M1019_s N_A_245_47#_c_750_n 0.00417299f $X=2.625 $Y=0.235 $X2=0 $Y2=0
cc_382 N_Y_c_513_n N_A_245_47#_c_750_n 0.0581171f $X=2.695 $Y=0.73 $X2=0 $Y2=0
cc_383 N_Y_c_575_p N_A_245_47#_c_750_n 0.0148563f $X=2.81 $Y=0.815 $X2=0 $Y2=0
cc_384 Y N_A_245_47#_c_750_n 0.00515509f $X=2.695 $Y=1.445 $X2=0 $Y2=0
cc_385 N_Y_c_496_n N_A_245_47#_c_751_n 0.00638629f $X=3.575 $Y=1.535 $X2=0 $Y2=0
cc_386 Y N_A_245_47#_c_751_n 0.00447631f $X=2.695 $Y=1.445 $X2=0 $Y2=0
cc_387 N_Y_c_493_n N_A_245_47#_c_751_n 0.00136495f $X=2.945 $Y=1.075 $X2=0 $Y2=0
cc_388 N_A_621_297#_c_582_n N_A_245_47#_c_758_n 0.00658191f $X=5.11 $Y=1.625
+ $X2=0 $Y2=0
cc_389 N_VGND_c_660_n N_A_245_47#_M1006_d 0.00254247f $X=7.13 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_390 N_VGND_c_660_n N_A_245_47#_M1013_d 0.00259403f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_391 N_VGND_c_660_n N_A_245_47#_M1024_d 0.00218529f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_392 N_VGND_c_660_n N_A_245_47#_M1010_d 0.0025535f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_393 N_VGND_c_660_n N_A_245_47#_M1018_d 0.00215201f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_394 N_VGND_c_660_n N_A_245_47#_M1007_s 0.0025535f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_395 N_VGND_c_660_n N_A_245_47#_M1023_s 0.00209319f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_396 N_VGND_c_651_n N_A_245_47#_c_750_n 0.0841928f $X=3.615 $Y=0 $X2=0 $Y2=0
cc_397 N_VGND_c_660_n N_A_245_47#_c_750_n 0.0678713f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_398 N_VGND_c_647_n N_A_245_47#_c_767_n 0.0109395f $X=3.7 $Y=0.39 $X2=0 $Y2=0
cc_399 N_VGND_c_651_n N_A_245_47#_c_767_n 0.0114777f $X=3.615 $Y=0 $X2=0 $Y2=0
cc_400 N_VGND_c_660_n N_A_245_47#_c_767_n 0.00913984f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_401 N_VGND_c_647_n N_A_245_47#_c_751_n 0.00471242f $X=3.7 $Y=0.39 $X2=0 $Y2=0
cc_402 N_VGND_M1004_s N_A_245_47#_c_752_n 0.00251047f $X=3.515 $Y=0.235 $X2=0
+ $Y2=0
cc_403 N_VGND_c_647_n N_A_245_47#_c_752_n 0.0127273f $X=3.7 $Y=0.39 $X2=0 $Y2=0
cc_404 N_VGND_c_651_n N_A_245_47#_c_752_n 0.00266636f $X=3.615 $Y=0 $X2=0 $Y2=0
cc_405 N_VGND_c_653_n N_A_245_47#_c_752_n 0.00198695f $X=4.555 $Y=0 $X2=0 $Y2=0
cc_406 N_VGND_c_660_n N_A_245_47#_c_752_n 0.00972452f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_407 N_VGND_c_648_n N_A_245_47#_c_775_n 0.0183628f $X=4.64 $Y=0.39 $X2=0 $Y2=0
cc_408 N_VGND_c_653_n N_A_245_47#_c_775_n 0.0223596f $X=4.555 $Y=0 $X2=0 $Y2=0
cc_409 N_VGND_c_660_n N_A_245_47#_c_775_n 0.0141302f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_410 N_VGND_M1017_s N_A_245_47#_c_753_n 0.00348805f $X=4.455 $Y=0.235 $X2=0
+ $Y2=0
cc_411 N_VGND_c_648_n N_A_245_47#_c_753_n 0.0131987f $X=4.64 $Y=0.39 $X2=0 $Y2=0
cc_412 N_VGND_c_653_n N_A_245_47#_c_753_n 0.00266636f $X=4.555 $Y=0 $X2=0 $Y2=0
cc_413 N_VGND_c_655_n N_A_245_47#_c_753_n 0.00199443f $X=5.495 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_660_n N_A_245_47#_c_753_n 0.0100158f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_648_n N_A_245_47#_c_783_n 0.0223967f $X=4.64 $Y=0.39 $X2=0 $Y2=0
cc_416 N_VGND_c_649_n N_A_245_47#_c_783_n 0.0183628f $X=5.58 $Y=0.39 $X2=0 $Y2=0
cc_417 N_VGND_c_655_n N_A_245_47#_c_783_n 0.0222529f $X=5.495 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_660_n N_A_245_47#_c_783_n 0.0139016f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_M1005_d N_A_245_47#_c_754_n 0.00251047f $X=5.395 $Y=0.235 $X2=0
+ $Y2=0
cc_420 N_VGND_c_649_n N_A_245_47#_c_754_n 0.0127273f $X=5.58 $Y=0.39 $X2=0 $Y2=0
cc_421 N_VGND_c_655_n N_A_245_47#_c_754_n 0.00266636f $X=5.495 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_657_n N_A_245_47#_c_754_n 0.00198695f $X=6.435 $Y=0 $X2=0 $Y2=0
cc_423 N_VGND_c_660_n N_A_245_47#_c_754_n 0.00972452f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_424 N_VGND_c_650_n N_A_245_47#_c_797_n 0.0183628f $X=6.52 $Y=0.39 $X2=0 $Y2=0
cc_425 N_VGND_c_657_n N_A_245_47#_c_797_n 0.0223596f $X=6.435 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_660_n N_A_245_47#_c_797_n 0.0141302f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_M1020_d N_A_245_47#_c_755_n 0.00348805f $X=6.335 $Y=0.235 $X2=0
+ $Y2=0
cc_428 N_VGND_c_650_n N_A_245_47#_c_755_n 0.0131987f $X=6.52 $Y=0.39 $X2=0 $Y2=0
cc_429 N_VGND_c_657_n N_A_245_47#_c_755_n 0.00266636f $X=6.435 $Y=0 $X2=0 $Y2=0
cc_430 N_VGND_c_659_n N_A_245_47#_c_755_n 0.00199443f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_660_n N_A_245_47#_c_755_n 0.0100158f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_c_650_n N_A_245_47#_c_756_n 0.0223967f $X=6.52 $Y=0.39 $X2=0 $Y2=0
cc_433 N_VGND_c_659_n N_A_245_47#_c_756_n 0.024373f $X=7.13 $Y=0 $X2=0 $Y2=0
cc_434 N_VGND_c_660_n N_A_245_47#_c_756_n 0.0141066f $X=7.13 $Y=0 $X2=0 $Y2=0
