# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o2bb2a_2
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A1_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.315000 1.075000 1.835000 1.275000 ;
    END
  END A1_N
  PIN A2_N
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.520000 0.380000 1.885000 0.735000 ;
        RECT 1.520000 0.735000 2.225000 0.905000 ;
        RECT 2.005000 0.905000 2.225000 1.100000 ;
    END
  END A2_N
  PIN B1
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.000000 1.075000 4.465000 1.645000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.220000 1.075000 3.825000 1.325000 ;
        RECT 3.655000 1.325000 3.825000 1.915000 ;
        RECT 3.655000 1.915000 3.995000 2.425000 ;
    END
  END B2
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.498000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.920000 0.825000 ;
        RECT 0.535000 0.825000 0.755000 1.795000 ;
        RECT 0.535000 1.795000 0.840000 2.465000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.110000  0.085000 0.365000 0.910000 ;
      RECT 0.110000  1.410000 0.365000 2.635000 ;
      RECT 0.925000  0.995000 1.145000 1.445000 ;
      RECT 0.925000  1.445000 1.370000 1.615000 ;
      RECT 1.010000  2.235000 1.390000 2.635000 ;
      RECT 1.135000  0.085000 1.305000 0.750000 ;
      RECT 1.200000  1.615000 1.370000 1.885000 ;
      RECT 1.200000  1.885000 3.435000 2.055000 ;
      RECT 1.540000  1.495000 2.660000 1.715000 ;
      RECT 2.055000  0.395000 2.565000 0.565000 ;
      RECT 2.360000  2.235000 2.765000 2.635000 ;
      RECT 2.395000  0.565000 2.565000 1.355000 ;
      RECT 2.395000  1.355000 2.660000 1.495000 ;
      RECT 2.735000  0.320000 2.980000 0.690000 ;
      RECT 2.810000  0.690000 2.980000 1.075000 ;
      RECT 2.810000  1.075000 3.000000 1.245000 ;
      RECT 2.830000  1.245000 3.000000 1.495000 ;
      RECT 2.830000  1.495000 3.435000 1.885000 ;
      RECT 3.035000  2.055000 3.435000 2.425000 ;
      RECT 3.205000  0.320000 3.435000 0.725000 ;
      RECT 3.205000  0.725000 4.405000 0.905000 ;
      RECT 3.675000  0.085000 3.845000 0.555000 ;
      RECT 4.015000  0.320000 4.405000 0.725000 ;
      RECT 4.165000  1.815000 4.480000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o2bb2a_2
END LIBRARY
