* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
X0 VGND a_216_93# a_336_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_426_413# a_27_410# a_532_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND B a_336_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X3 VGND D_N a_216_93# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 a_336_413# a_216_93# a_426_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 X a_336_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 X a_336_413# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_336_413# a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 a_27_410# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X9 VPWR D_N a_216_93# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X10 a_336_413# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 a_27_410# C_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X12 VPWR a_336_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VGND a_336_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_532_297# B a_614_297# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X15 a_614_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
