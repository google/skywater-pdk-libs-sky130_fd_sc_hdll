* File: sky130_fd_sc_hdll__o22ai_2.spice
* Created: Thu Aug 27 19:21:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o22ai_2  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_Y_M1006_d N_B1_M1006_g N_A_27_47#_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.182 PD=1.02 PS=1.86 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75004.1 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1006_d N_B1_M1013_g N_A_27_47#_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75003.6 A=0.0975 P=1.6 MULT=1
MM1007 N_A_27_47#_M1013_s N_B2_M1007_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.1
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1012 N_A_27_47#_M1012_d N_B2_M1012_g N_Y_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26975 AS=0.12025 PD=1.48 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.7
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_47#_M1012_d N_A2_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.26975 AS=0.12025 PD=1.48 PS=1.02 NRD=0 NRS=17.532 M=1 R=4.33333
+ SA=75002.6 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1009 N_A_27_47#_M1009_d N_A2_M1009_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=0 M=1 R=4.33333 SA=75003.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A1_M1004_g N_A_27_47#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1014 N_VGND_M1004_d N_A1_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_B1_M1001_g N_A_27_297#_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1001_d N_B1_M1011_g N_A_27_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1003 N_A_27_297#_M1011_s N_B2_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_A_27_297#_M1005_d N_B2_M1005_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g N_A_515_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1000_d N_A2_M1015_g N_A_515_297#_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1008 N_A_515_297#_M1015_s N_A1_M1008_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1010 N_A_515_297#_M1010_d N_A1_M1010_g N_VPWR_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX17_noxref noxref_13 B2 B2 PROBETYPE=1
pX18_noxref noxref_14 A2 A2 PROBETYPE=1
pX19_noxref noxref_15 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o22ai_2.pxi.spice"
*
.ends
*
*
