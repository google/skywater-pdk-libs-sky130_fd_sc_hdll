* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__or3_2 A B C VGND VNB VPB VPWR X
M1000 VGND a_30_53# X VNB nshort w=650000u l=150000u
+  ad=6.469e+11p pd=5.71e+06u as=2.405e+11p ps=2.04e+06u
M1001 a_120_297# C a_30_53# VPB phighvt w=420000u l=180000u
+  ad=9.66e+10p pd=1.3e+06u as=1.134e+11p ps=1.38e+06u
M1002 VGND A a_30_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=2.646e+11p ps=2.94e+06u
M1003 VPWR a_30_53# X VPB phighvt w=1e+06u l=180000u
+  ad=8.257e+11p pd=5.75e+06u as=2.9e+11p ps=2.58e+06u
M1004 a_30_53# B VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_30_53# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VPWR A a_202_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=1.47e+11p ps=1.54e+06u
M1007 X a_30_53# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 VGND C a_30_53# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_202_297# B a_120_297# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
