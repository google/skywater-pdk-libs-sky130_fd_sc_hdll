# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdfbbp_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfbbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  15.64000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.975000 0.435000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.155000 1.325000 4.475000 2.375000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.439000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 15.260000 0.255000 15.545000 0.825000 ;
        RECT 15.260000 1.605000 15.545000 2.465000 ;
        RECT 15.310000 0.825000 15.545000 1.605000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.595750 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 13.715000 0.255000 14.115000 0.715000 ;
        RECT 13.715000 1.630000 14.095000 2.465000 ;
        RECT 13.820000 0.715000 14.115000 1.520000 ;
        RECT 13.820000 1.520000 14.095000 1.630000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.515000 1.095000 13.090000 1.325000 ;
    END
  END RESET_B
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.490000 1.025000 1.765000 1.685000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.935000 0.760000 2.255000 0.765000 ;
        RECT 1.935000 0.765000 2.605000 1.015000 ;
        RECT 1.935000 1.015000 2.255000 1.695000 ;
        RECT 1.975000 0.345000 2.255000 0.760000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.277200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT  6.525000 0.735000  6.815000 0.780000 ;
        RECT  6.525000 0.780000 10.945000 0.920000 ;
        RECT  6.525000 0.920000  6.815000 0.965000 ;
        RECT 10.655000 0.735000 10.945000 0.780000 ;
        RECT 10.655000 0.920000 10.945000 0.965000 ;
    END
  END SET_B
  PIN VGND
    ANTENNADIFFAREA  1.524700 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 15.640000 0.085000 ;
        RECT  0.515000  0.085000  0.895000 0.465000 ;
        RECT  1.555000  0.085000  1.805000 0.635000 ;
        RECT  3.620000  0.085000  3.950000 0.445000 ;
        RECT  6.385000  0.085000  6.555000 0.525000 ;
        RECT  8.290000  0.085000  8.675000 0.465000 ;
        RECT 10.410000  0.085000 10.720000 0.525000 ;
        RECT 13.100000  0.085000 13.430000 0.805000 ;
        RECT 14.750000  0.085000 15.040000 0.545000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
        RECT 14.865000 -0.085000 15.035000 0.085000 ;
        RECT 15.325000 -0.085000 15.495000 0.085000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 15.640000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  2.152000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 15.640000 2.805000 ;
        RECT  0.515000 2.135000  0.895000 2.635000 ;
        RECT  1.555000 1.885000  1.885000 2.635000 ;
        RECT  3.510000 2.215000  3.890000 2.635000 ;
        RECT  6.205000 2.205000  6.585000 2.635000 ;
        RECT  7.825000 1.915000  8.155000 2.635000 ;
        RECT 10.520000 2.255000 10.900000 2.635000 ;
        RECT 11.940000 2.255000 13.430000 2.635000 ;
        RECT 14.745000 1.765000 15.040000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
        RECT 14.405000 2.635000 14.575000 2.805000 ;
        RECT 14.865000 2.635000 15.035000 2.805000 ;
        RECT 15.325000 2.635000 15.495000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 15.640000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.170000 0.345000  0.345000 0.635000 ;
      RECT  0.170000 0.635000  0.885000 0.805000 ;
      RECT  0.170000 1.795000  0.885000 1.965000 ;
      RECT  0.170000 1.965000  0.345000 2.465000 ;
      RECT  0.655000 0.805000  0.885000 1.795000 ;
      RECT  1.115000 0.345000  1.320000 2.465000 ;
      RECT  2.385000 1.875000  2.765000 2.385000 ;
      RECT  2.550000 0.265000  2.955000 0.595000 ;
      RECT  2.550000 1.185000  3.275000 1.365000 ;
      RECT  2.550000 1.365000  2.765000 1.875000 ;
      RECT  2.785000 0.595000  2.955000 1.075000 ;
      RECT  2.785000 1.075000  3.275000 1.185000 ;
      RECT  2.945000 1.575000  3.895000 1.745000 ;
      RECT  2.945000 1.745000  3.265000 1.905000 ;
      RECT  3.095000 1.905000  3.265000 2.465000 ;
      RECT  3.125000 0.305000  3.325000 0.625000 ;
      RECT  3.125000 0.625000  3.895000 0.765000 ;
      RECT  3.125000 0.765000  4.070000 0.795000 ;
      RECT  3.725000 0.795000  4.070000 1.095000 ;
      RECT  3.725000 1.095000  3.895000 1.575000 ;
      RECT  4.645000 0.305000  4.815000 2.465000 ;
      RECT  4.985000 0.705000  5.245000 1.575000 ;
      RECT  4.985000 1.575000  5.575000 1.955000 ;
      RECT  5.035000 2.250000  5.915000 2.420000 ;
      RECT  5.100000 0.265000  6.215000 0.465000 ;
      RECT  5.425000 0.645000  5.825000 1.015000 ;
      RECT  5.745000 1.195000  6.215000 1.235000 ;
      RECT  5.745000 1.235000  7.195000 1.405000 ;
      RECT  5.745000 1.405000  5.915000 2.250000 ;
      RECT  5.995000 0.465000  6.215000 1.195000 ;
      RECT  6.085000 1.575000  6.385000 1.785000 ;
      RECT  6.085000 1.785000  7.585000 2.035000 ;
      RECT  6.385000 0.735000  6.795000 1.065000 ;
      RECT  6.775000 0.255000  8.045000 0.425000 ;
      RECT  6.775000 0.425000  7.105000 0.465000 ;
      RECT  6.935000 2.035000  7.105000 2.375000 ;
      RECT  6.945000 1.405000  7.195000 1.485000 ;
      RECT  6.975000 1.155000  7.195000 1.235000 ;
      RECT  7.275000 0.595000  7.655000 0.765000 ;
      RECT  7.415000 0.765000  7.655000 0.895000 ;
      RECT  7.415000 0.895000  8.875000 1.065000 ;
      RECT  7.415000 1.065000  7.585000 1.785000 ;
      RECT  7.805000 1.235000  8.135000 1.415000 ;
      RECT  7.805000 1.415000  8.910000 1.655000 ;
      RECT  7.850000 0.425000  8.045000 0.715000 ;
      RECT  8.445000 1.065000  8.875000 1.235000 ;
      RECT  9.110000 1.575000  9.345000 1.985000 ;
      RECT  9.170000 0.705000  9.510000 1.125000 ;
      RECT  9.170000 1.125000  9.890000 1.305000 ;
      RECT  9.300000 2.250000 10.230000 2.420000 ;
      RECT  9.415000 0.265000 10.230000 0.465000 ;
      RECT  9.635000 1.305000  9.890000 1.905000 ;
      RECT 10.060000 0.465000 10.230000 1.235000 ;
      RECT 10.060000 1.235000 11.510000 1.405000 ;
      RECT 10.060000 1.405000 10.230000 2.250000 ;
      RECT 10.400000 1.575000 10.700000 1.915000 ;
      RECT 10.400000 1.915000 13.430000 2.085000 ;
      RECT 10.655000 0.735000 11.080000 1.065000 ;
      RECT 10.980000 0.255000 12.300000 0.425000 ;
      RECT 10.980000 0.425000 11.380000 0.465000 ;
      RECT 11.190000 2.085000 11.360000 2.375000 ;
      RECT 11.290000 1.075000 11.510000 1.235000 ;
      RECT 11.535000 0.645000 11.915000 0.815000 ;
      RECT 11.730000 0.815000 11.915000 1.915000 ;
      RECT 12.125000 0.425000 12.300000 0.585000 ;
      RECT 12.130000 0.755000 12.815000 0.925000 ;
      RECT 12.130000 0.925000 12.345000 1.575000 ;
      RECT 12.130000 1.575000 12.905000 1.745000 ;
      RECT 12.615000 0.265000 12.815000 0.755000 ;
      RECT 13.260000 0.995000 13.525000 1.325000 ;
      RECT 13.260000 1.325000 13.430000 1.915000 ;
      RECT 14.265000 1.725000 14.520000 2.415000 ;
      RECT 14.315000 0.255000 14.520000 0.995000 ;
      RECT 14.315000 0.995000 15.090000 1.325000 ;
      RECT 14.315000 1.325000 14.520000 1.725000 ;
    LAYER mcon ;
      RECT  0.655000 1.785000  0.825000 1.955000 ;
      RECT  1.150000 0.765000  1.320000 0.935000 ;
      RECT  3.105000 1.105000  3.275000 1.275000 ;
      RECT  4.645000 1.105000  4.815000 1.275000 ;
      RECT  5.145000 1.785000  5.315000 1.955000 ;
      RECT  5.655000 0.765000  5.825000 0.935000 ;
      RECT  6.585000 0.765000  6.755000 0.935000 ;
      RECT  8.715000 1.445000  8.885000 1.615000 ;
      RECT  9.175000 1.105000  9.345000 1.275000 ;
      RECT  9.175000 1.785000  9.345000 1.955000 ;
      RECT 10.715000 0.765000 10.885000 0.935000 ;
      RECT 12.165000 1.445000 12.335000 1.615000 ;
    LAYER met1 ;
      RECT  0.595000 1.755000  0.885000 1.800000 ;
      RECT  0.595000 1.800000  9.405000 1.940000 ;
      RECT  0.595000 1.940000  0.885000 1.985000 ;
      RECT  1.090000 0.735000  1.380000 0.780000 ;
      RECT  1.090000 0.780000  5.885000 0.920000 ;
      RECT  1.090000 0.920000  1.380000 0.965000 ;
      RECT  3.045000 1.075000  3.335000 1.120000 ;
      RECT  3.045000 1.120000  4.875000 1.260000 ;
      RECT  3.045000 1.260000  3.335000 1.305000 ;
      RECT  4.585000 1.075000  4.875000 1.120000 ;
      RECT  4.585000 1.260000  4.875000 1.305000 ;
      RECT  5.085000 1.755000  5.375000 1.800000 ;
      RECT  5.085000 1.940000  5.375000 1.985000 ;
      RECT  5.595000 0.735000  5.885000 0.780000 ;
      RECT  5.595000 0.920000  5.885000 0.965000 ;
      RECT  5.670000 0.965000  5.885000 1.120000 ;
      RECT  5.670000 1.120000  9.405000 1.260000 ;
      RECT  8.655000 1.415000  8.945000 1.460000 ;
      RECT  8.655000 1.460000 12.395000 1.600000 ;
      RECT  8.655000 1.600000  8.945000 1.645000 ;
      RECT  9.115000 1.075000  9.405000 1.120000 ;
      RECT  9.115000 1.260000  9.405000 1.305000 ;
      RECT  9.115000 1.755000  9.405000 1.800000 ;
      RECT  9.115000 1.940000  9.405000 1.985000 ;
      RECT 12.105000 1.415000 12.395000 1.460000 ;
      RECT 12.105000 1.600000 12.395000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfbbp_1
END LIBRARY
