* File: sky130_fd_sc_hdll__o2bb2a_1.spice
* Created: Thu Aug 27 19:21:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o2bb2a_1.pex.spice"
.subckt sky130_fd_sc_hdll__o2bb2a_1  VNB VPB A1_N A2_N B2 B1 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* B1	B1
* B2	B2
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1009 N_VGND_M1009_d N_A_76_199#_M1009_g N_X_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.132582 AS=0.2015 PD=1.2514 PS=1.92 NRD=3.684 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1001 A_225_47# N_A1_N_M1001_g N_VGND_M1009_d VNB NSHORT L=0.15 W=0.42
+ AD=0.06615 AS=0.0856682 PD=0.735 PS=0.808598 NRD=29.28 NRS=22.848 M=1 R=2.8
+ SA=75000.8 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1004 N_A_224_369#_M1004_d N_A2_N_M1004_g A_225_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.06615 PD=1.46 PS=0.735 NRD=12.852 NRS=29.28 M=1 R=2.8
+ SA=75001.2 SB=75000.2 A=0.063 P=1.14 MULT=1
MM1010 N_A_529_47#_M1010_d N_A_224_369#_M1010_g N_A_76_199#_M1010_s VNB NSHORT
+ L=0.15 W=0.42 AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.3 A=0.063 P=1.14 MULT=1
MM1003 N_VGND_M1003_d N_B2_M1003_g N_A_529_47#_M1010_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0903 AS=0.0672 PD=0.85 PS=0.74 NRD=17.136 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75000.8 A=0.063 P=1.14 MULT=1
MM1008 N_A_529_47#_M1008_d N_B1_M1008_g N_VGND_M1003_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.0903 PD=1.46 PS=0.85 NRD=12.852 NRS=25.704 M=1 R=2.8 SA=75001.3
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_A_76_199#_M1002_g N_X_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.215282 AS=0.27 PD=1.90845 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1006 N_A_224_369#_M1006_d N_A1_N_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1332 AS=0.0904183 PD=1.2 PS=0.801549 NRD=122.948 NRS=35.1645 M=1
+ R=2.33333 SA=90000.7 SB=90002.8 A=0.0756 P=1.2 MULT=1
MM1000 N_VPWR_M1000_d N_A2_N_M1000_g N_A_224_369#_M1006_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.21035 AS=0.1332 PD=1.355 PS=1.2 NRD=98.4803 NRS=122.948 M=1
+ R=2.33333 SA=90001.3 SB=90002.2 A=0.0756 P=1.2 MULT=1
MM1011 N_A_76_199#_M1011_d N_A_224_369#_M1011_g N_VPWR_M1000_d VPB PHIGHVT
+ L=0.18 W=0.42 AD=0.0735 AS=0.21035 PD=0.77 PS=1.355 NRD=0 NRS=209.116 M=1
+ R=2.33333 SA=90002.2 SB=90001.3 A=0.0756 P=1.2 MULT=1
MM1005 A_633_369# N_B2_M1005_g N_A_76_199#_M1011_d VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0819 AS=0.0735 PD=0.81 PS=0.77 NRD=65.6601 NRS=25.7873 M=1 R=2.33333
+ SA=90002.8 SB=90000.7 A=0.0756 P=1.2 MULT=1
MM1007 N_VPWR_M1007_d N_B1_M1007_g A_633_369# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.1134 AS=0.0819 PD=1.38 PS=0.81 NRD=2.3443 NRS=65.6601 M=1 R=2.33333
+ SA=90003.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_15 B2 B2 PROBETYPE=1
pX14_noxref noxref_16 B1 B1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o2bb2a_1.pxi.spice"
*
.ends
*
*
