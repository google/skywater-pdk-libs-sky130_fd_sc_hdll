* File: sky130_fd_sc_hdll__nand4b_4.pxi.spice
* Created: Thu Aug 27 19:14:54 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%A_N N_A_N_c_134_n N_A_N_M1011_g N_A_N_M1023_g
+ A_N N_A_N_c_133_n PM_SKY130_FD_SC_HDLL__NAND4B_4%A_N
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%A_27_47# N_A_27_47#_M1023_s N_A_27_47#_M1011_s
+ N_A_27_47#_c_174_n N_A_27_47#_M1006_g N_A_27_47#_M1009_g N_A_27_47#_c_175_n
+ N_A_27_47#_M1014_g N_A_27_47#_M1010_g N_A_27_47#_c_176_n N_A_27_47#_M1020_g
+ N_A_27_47#_M1013_g N_A_27_47#_c_177_n N_A_27_47#_M1030_g N_A_27_47#_M1026_g
+ N_A_27_47#_c_165_n N_A_27_47#_c_178_n N_A_27_47#_c_179_n N_A_27_47#_c_166_n
+ N_A_27_47#_c_167_n N_A_27_47#_c_180_n N_A_27_47#_c_168_n N_A_27_47#_c_169_n
+ N_A_27_47#_c_170_n N_A_27_47#_c_171_n N_A_27_47#_c_172_n N_A_27_47#_c_173_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%B N_B_c_297_n N_B_M1004_g N_B_M1000_g
+ N_B_c_298_n N_B_M1019_g N_B_M1003_g N_B_c_299_n N_B_M1025_g N_B_M1022_g
+ N_B_c_300_n N_B_M1033_g N_B_M1027_g B B B B N_B_c_295_n B B B B
+ PM_SKY130_FD_SC_HDLL__NAND4B_4%B
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%C N_C_c_378_n N_C_M1001_g N_C_M1016_g
+ N_C_c_379_n N_C_M1015_g N_C_M1018_g N_C_c_380_n N_C_M1021_g N_C_M1029_g
+ N_C_c_381_n N_C_M1031_g N_C_M1032_g C C C C N_C_c_375_n N_C_c_376_n
+ N_C_c_377_n C C C C PM_SKY130_FD_SC_HDLL__NAND4B_4%C
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%D N_D_M1002_g N_D_c_458_n N_D_M1005_g
+ N_D_M1012_g N_D_c_459_n N_D_M1007_g N_D_M1024_g N_D_c_460_n N_D_M1008_g
+ N_D_M1028_g N_D_c_461_n N_D_M1017_g D D D D N_D_c_455_n N_D_c_456_n D D D D
+ PM_SKY130_FD_SC_HDLL__NAND4B_4%D
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%VPWR N_VPWR_M1011_d N_VPWR_M1006_d
+ N_VPWR_M1014_d N_VPWR_M1030_d N_VPWR_M1019_s N_VPWR_M1033_s N_VPWR_M1015_s
+ N_VPWR_M1031_s N_VPWR_M1007_d N_VPWR_M1017_d N_VPWR_c_540_n N_VPWR_c_541_n
+ N_VPWR_c_542_n N_VPWR_c_543_n N_VPWR_c_544_n N_VPWR_c_545_n N_VPWR_c_546_n
+ N_VPWR_c_547_n N_VPWR_c_548_n N_VPWR_c_549_n N_VPWR_c_550_n N_VPWR_c_551_n
+ N_VPWR_c_552_n N_VPWR_c_553_n N_VPWR_c_554_n N_VPWR_c_555_n N_VPWR_c_556_n
+ N_VPWR_c_557_n N_VPWR_c_558_n N_VPWR_c_559_n N_VPWR_c_560_n N_VPWR_c_561_n
+ N_VPWR_c_562_n N_VPWR_c_563_n VPWR N_VPWR_c_564_n N_VPWR_c_565_n
+ N_VPWR_c_566_n N_VPWR_c_567_n N_VPWR_c_539_n
+ PM_SKY130_FD_SC_HDLL__NAND4B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%Y N_Y_M1009_s N_Y_M1013_s N_Y_M1006_s
+ N_Y_M1020_s N_Y_M1004_d N_Y_M1025_d N_Y_M1001_d N_Y_M1021_d N_Y_M1005_s
+ N_Y_M1008_s N_Y_c_691_n N_Y_c_693_n N_Y_c_717_n N_Y_c_694_n N_Y_c_724_n
+ N_Y_c_727_n N_Y_c_695_n N_Y_c_749_n N_Y_c_696_n N_Y_c_772_n N_Y_c_697_n
+ N_Y_c_779_n N_Y_c_698_n N_Y_c_785_n N_Y_c_699_n N_Y_c_700_n N_Y_c_808_n
+ N_Y_c_701_n N_Y_c_702_n N_Y_c_703_n N_Y_c_704_n N_Y_c_705_n N_Y_c_706_n Y Y Y
+ N_Y_c_739_n PM_SKY130_FD_SC_HDLL__NAND4B_4%Y
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%VGND N_VGND_M1023_d N_VGND_M1002_d
+ N_VGND_M1024_d N_VGND_c_883_n N_VGND_c_884_n N_VGND_c_885_n N_VGND_c_886_n
+ N_VGND_c_887_n N_VGND_c_888_n N_VGND_c_889_n VGND N_VGND_c_890_n
+ N_VGND_c_891_n N_VGND_c_892_n PM_SKY130_FD_SC_HDLL__NAND4B_4%VGND
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%A_225_47# N_A_225_47#_M1009_d
+ N_A_225_47#_M1010_d N_A_225_47#_M1026_d N_A_225_47#_M1003_d
+ N_A_225_47#_M1027_d N_A_225_47#_c_986_n N_A_225_47#_c_987_n
+ N_A_225_47#_c_988_n PM_SKY130_FD_SC_HDLL__NAND4B_4%A_225_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%A_693_47# N_A_693_47#_M1000_s
+ N_A_693_47#_M1022_s N_A_693_47#_M1016_s N_A_693_47#_M1029_s
+ N_A_693_47#_c_1030_n PM_SKY130_FD_SC_HDLL__NAND4B_4%A_693_47#
x_PM_SKY130_FD_SC_HDLL__NAND4B_4%A_1081_47# N_A_1081_47#_M1016_d
+ N_A_1081_47#_M1018_d N_A_1081_47#_M1032_d N_A_1081_47#_M1012_s
+ N_A_1081_47#_M1028_s N_A_1081_47#_c_1063_n N_A_1081_47#_c_1073_n
+ N_A_1081_47#_c_1074_n N_A_1081_47#_c_1064_n N_A_1081_47#_c_1065_n
+ N_A_1081_47#_c_1081_n N_A_1081_47#_c_1066_n N_A_1081_47#_c_1067_n
+ N_A_1081_47#_c_1068_n PM_SKY130_FD_SC_HDLL__NAND4B_4%A_1081_47#
cc_1 VNB N_A_N_M1023_g 0.0265299f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB A_N 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_133_n 0.0406212f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_4 VNB N_A_27_47#_M1009_g 0.022257f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.212
cc_5 VNB N_A_27_47#_M1010_g 0.0183542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_27_47#_M1013_g 0.0178704f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_47#_M1026_g 0.0187975f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_47#_c_165_n 0.0189842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_166_n 0.0025002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_27_47#_c_167_n 0.00939234f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_47#_c_168_n 0.00420118f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_c_169_n 7.99113e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_c_170_n 0.00934767f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_171_n 0.00267593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_172_n 0.0330574f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_173_n 0.086168f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_B_M1000_g 0.0187461f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_18 VNB N_B_M1003_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_19 VNB N_B_M1022_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_B_M1027_g 0.023617f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_B_c_295_n 0.101123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB B 0.00350438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_C_M1016_g 0.0242928f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_24 VNB N_C_M1018_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.212
cc_25 VNB N_C_M1029_g 0.0183897f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_C_M1032_g 0.0183319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_C_c_375_n 0.0331062f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_C_c_376_n 0.00184776f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_C_c_377_n 0.0846646f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_D_M1002_g 0.0180932f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_31 VNB N_D_M1012_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.212
cc_32 VNB N_D_M1024_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_D_M1028_g 0.0235985f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_D_c_455_n 0.0847647f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_D_c_456_n 0.0291228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB D 0.00946594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VPWR_c_539_n 0.402575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_691_n 0.00597884f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB Y 0.00120246f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_883_n 0.00869034f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.212
cc_41 VNB N_VGND_c_884_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_885_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_886_n 0.15691f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_887_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_888_n 0.0192031f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_889_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_890_n 0.021812f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_891_n 0.463538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_892_n 0.0235067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_225_47#_c_986_n 0.00217944f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_225_47#_c_987_n 0.00651087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_225_47#_c_988_n 0.00256809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_693_47#_c_1030_n 0.0277237f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_1081_47#_c_1063_n 0.00245677f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_1081_47#_c_1064_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_1081_47#_c_1065_n 0.00355458f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_A_1081_47#_c_1066_n 0.0118443f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_A_1081_47#_c_1067_n 0.0192914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_A_1081_47#_c_1068_n 0.00253093f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VPB N_A_N_c_134_n 0.0239744f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_61 VPB N_A_N_c_133_n 0.017029f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_62 VPB N_A_27_47#_c_174_n 0.0195378f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_175_n 0.0158656f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_176_n 0.0157312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_177_n 0.0158458f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_178_n 0.00765454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_179_n 0.0314532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_180_n 0.00131456f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_169_n 0.00467396f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_47#_c_173_n 0.0262074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_B_c_297_n 0.0159794f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_72 VPB N_B_c_298_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_73 VPB N_B_c_299_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_B_c_300_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_B_c_295_n 0.0325788f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_C_c_378_n 0.0201049f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_77 VPB N_C_c_379_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_78 VPB N_C_c_380_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_C_c_381_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_C_c_377_n 0.0287129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_D_c_458_n 0.0160015f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_82 VPB N_D_c_459_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_83 VPB N_D_c_460_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_D_c_461_n 0.0198539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_D_c_455_n 0.0289993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_D_c_456_n 0.00976317f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_540_n 0.0106419f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_541_n 0.00474491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_542_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_543_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_544_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_545_n 0.00760606f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_546_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_547_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_VPWR_c_548_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_549_n 0.0134596f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_550_n 0.0463636f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_551_n 0.00644865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_552_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_553_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_554_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_555_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_556_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_557_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_558_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_559_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_560_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_561_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_562_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_563_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_564_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_565_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_566_n 0.0326527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_567_n 0.0132428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_539_n 0.0486981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_Y_c_693_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_Y_c_694_n 0.0022967f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_695_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_696_n 0.00728445f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_Y_c_697_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_Y_c_698_n 0.00528316f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_Y_c_699_n 0.00173134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_Y_c_700_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_Y_c_701_n 0.00730119f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_Y_c_702_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_Y_c_703_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_Y_c_704_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_Y_c_705_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_Y_c_706_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 N_A_N_c_134_n N_A_27_47#_c_178_n 6.2e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 A_N N_A_27_47#_c_178_n 0.0184539f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_N_c_133_n N_A_27_47#_c_178_n 0.006079f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_133 N_A_N_c_134_n N_A_27_47#_c_179_n 0.0115942f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_N_M1023_g N_A_27_47#_c_166_n 0.0137691f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_135 A_N N_A_27_47#_c_166_n 0.00104802f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_N_c_133_n N_A_27_47#_c_166_n 5.86657e-19 $X=0.495 $Y=1.212 $X2=0
+ $Y2=0
cc_137 A_N N_A_27_47#_c_167_n 0.0255857f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_138 N_A_N_c_133_n N_A_27_47#_c_167_n 0.0077859f $X=0.495 $Y=1.212 $X2=0 $Y2=0
cc_139 N_A_N_c_134_n N_A_27_47#_c_180_n 0.0168914f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_140 A_N N_A_27_47#_c_180_n 8.10212e-19 $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_141 N_A_N_M1023_g N_A_27_47#_c_168_n 0.00609467f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_142 N_A_N_c_134_n N_A_27_47#_c_169_n 0.0033081f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_N_c_133_n N_A_27_47#_c_169_n 0.00523181f $X=0.495 $Y=1.212 $X2=0
+ $Y2=0
cc_144 A_N N_A_27_47#_c_171_n 0.0138154f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_N_c_133_n N_A_27_47#_c_171_n 0.00264337f $X=0.495 $Y=1.212 $X2=0
+ $Y2=0
cc_146 N_A_N_c_133_n N_A_27_47#_c_172_n 0.00570182f $X=0.495 $Y=1.212 $X2=0
+ $Y2=0
cc_147 N_A_N_c_134_n N_VPWR_c_541_n 0.00329148f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_N_c_134_n N_VPWR_c_551_n 0.00824863f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_N_c_134_n N_VPWR_c_566_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_N_c_134_n N_VPWR_c_539_n 0.0140376f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_N_M1023_g N_VGND_c_883_n 0.0044954f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_N_M1023_g N_VGND_c_891_n 0.00823623f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_N_M1023_g N_VGND_c_892_n 0.00439206f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A_N_M1023_g N_A_225_47#_c_987_n 0.00359645f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_27_47#_c_177_n N_B_c_297_n 0.0229862f $X=2.895 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_156 N_A_27_47#_M1026_g N_B_M1000_g 0.0223757f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_173_n N_B_c_295_n 0.0245486f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_158 N_A_27_47#_c_173_n B 0.00180429f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_180_n N_VPWR_M1011_d 0.00520922f $X=0.66 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_160 N_A_27_47#_c_169_n N_VPWR_M1011_d 3.02568e-19 $X=0.757 $Y=1.495 $X2=-0.19
+ $Y2=-0.24
cc_161 N_A_27_47#_c_174_n N_VPWR_c_541_n 0.0086715f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_179_n N_VPWR_c_541_n 0.00496819f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_180_n N_VPWR_c_541_n 0.0134641f $X=0.66 $Y=1.58 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_170_n N_VPWR_c_541_n 0.0190248f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_172_n N_VPWR_c_541_n 0.00624109f $X=1.485 $Y=1.217 $X2=0
+ $Y2=0
cc_166 N_A_27_47#_c_175_n N_VPWR_c_542_n 0.0052072f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_176_n N_VPWR_c_542_n 0.004751f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_27_47#_c_177_n N_VPWR_c_543_n 0.0052072f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_179_n N_VPWR_c_551_n 0.0425456f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_180_n N_VPWR_c_551_n 0.0185488f $X=0.66 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_170_n N_VPWR_c_551_n 0.00706024f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_174_n N_VPWR_c_552_n 0.00597712f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_173 N_A_27_47#_c_175_n N_VPWR_c_552_n 0.00673617f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_176_n N_VPWR_c_554_n 0.00597712f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_177_n N_VPWR_c_554_n 0.00673617f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_179_n N_VPWR_c_566_n 0.021418f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_177 N_A_27_47#_M1011_s N_VPWR_c_539_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_174_n N_VPWR_c_539_n 0.0112769f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_27_47#_c_175_n N_VPWR_c_539_n 0.0118438f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_176_n N_VPWR_c_539_n 0.00999457f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_177_n N_VPWR_c_539_n 0.011869f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A_27_47#_c_179_n N_VPWR_c_539_n 0.0126651f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1009_g N_Y_c_691_n 0.00630077f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_184 N_A_27_47#_M1010_g N_Y_c_691_n 0.0126025f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_185 N_A_27_47#_M1013_g N_Y_c_691_n 0.0057546f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_186 N_A_27_47#_c_170_n N_Y_c_691_n 0.034711f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_187 N_A_27_47#_c_173_n N_Y_c_691_n 0.00711941f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_188 N_A_27_47#_c_174_n N_Y_c_693_n 0.0052648f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_27_47#_c_175_n N_Y_c_693_n 0.00116723f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_27_47#_c_169_n N_Y_c_693_n 0.00141131f $X=0.757 $Y=1.495 $X2=0 $Y2=0
cc_191 N_A_27_47#_c_170_n N_Y_c_693_n 0.0305808f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_173_n N_Y_c_693_n 0.0074788f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_193 N_A_27_47#_c_174_n N_Y_c_717_n 0.0121679f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_175_n N_Y_c_717_n 0.0106251f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_27_47#_c_176_n N_Y_c_717_n 6.24674e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_175_n N_Y_c_694_n 0.0161811f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_27_47#_c_176_n N_Y_c_694_n 0.00943113f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_170_n N_Y_c_694_n 0.00626555f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_27_47#_c_173_n N_Y_c_694_n 0.00849036f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_175_n N_Y_c_724_n 6.48386e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_176_n N_Y_c_724_n 0.0130707f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_27_47#_c_177_n N_Y_c_724_n 0.0106251f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_177_n N_Y_c_727_n 6.48386e-19 $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_177_n N_Y_c_701_n 0.018707f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_27_47#_c_173_n N_Y_c_701_n 4.93319e-19 $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1010_g Y 6.69312e-19 $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_176_n Y 0.00124952f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_27_47#_M1013_g Y 0.00444494f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_209 N_A_27_47#_c_177_n Y 0.00107825f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_27_47#_M1026_g Y 0.00368424f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_170_n Y 0.00751579f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_173_n Y 0.0416946f $X=2.895 $Y=1.217 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_176_n Y 0.0044033f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_177_n Y 0.00191486f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_27_47#_M1013_g N_Y_c_739_n 0.00475315f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_216 N_A_27_47#_M1026_g N_Y_c_739_n 3.43088e-19 $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_166_n N_VGND_M1023_d 0.00466472f $X=0.66 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_218 N_A_27_47#_M1009_g N_VGND_c_883_n 0.00211277f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_166_n N_VGND_c_883_n 0.015871f $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_170_n N_VGND_c_883_n 0.00148402f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1009_g N_VGND_c_886_n 0.00357877f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_27_47#_M1010_g N_VGND_c_886_n 0.00357877f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_223 N_A_27_47#_M1013_g N_VGND_c_886_n 0.00357877f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1026_g N_VGND_c_886_n 0.00357877f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1023_s N_VGND_c_891_n 0.00259235f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_226 N_A_27_47#_M1009_g N_VGND_c_891_n 0.00668309f $X=1.51 $Y=0.56 $X2=0 $Y2=0
cc_227 N_A_27_47#_M1010_g N_VGND_c_891_n 0.00548399f $X=1.98 $Y=0.56 $X2=0 $Y2=0
cc_228 N_A_27_47#_M1013_g N_VGND_c_891_n 0.00548399f $X=2.45 $Y=0.56 $X2=0 $Y2=0
cc_229 N_A_27_47#_M1026_g N_VGND_c_891_n 0.00550244f $X=2.92 $Y=0.56 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_165_n N_VGND_c_891_n 0.0128092f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_166_n N_VGND_c_891_n 0.00585608f $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_232 N_A_27_47#_c_165_n N_VGND_c_892_n 0.0221535f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_166_n N_VGND_c_892_n 0.00248202f $X=0.66 $Y=0.82 $X2=0 $Y2=0
cc_234 N_A_27_47#_M1009_g N_A_225_47#_c_987_n 0.00459803f $X=1.51 $Y=0.56 $X2=0
+ $Y2=0
cc_235 N_A_27_47#_c_166_n N_A_225_47#_c_987_n 0.0116449f $X=0.66 $Y=0.82 $X2=0
+ $Y2=0
cc_236 N_A_27_47#_c_170_n N_A_225_47#_c_987_n 0.0201437f $X=1.72 $Y=1.16 $X2=0
+ $Y2=0
cc_237 N_A_27_47#_c_172_n N_A_225_47#_c_987_n 0.00588114f $X=1.485 $Y=1.217
+ $X2=0 $Y2=0
cc_238 N_A_27_47#_M1009_g N_A_225_47#_c_988_n 0.00999874f $X=1.51 $Y=0.56 $X2=0
+ $Y2=0
cc_239 N_A_27_47#_M1010_g N_A_225_47#_c_988_n 0.00903374f $X=1.98 $Y=0.56 $X2=0
+ $Y2=0
cc_240 N_A_27_47#_M1013_g N_A_225_47#_c_988_n 0.00902896f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_241 N_A_27_47#_M1026_g N_A_225_47#_c_988_n 0.0137288f $X=2.92 $Y=0.56 $X2=0
+ $Y2=0
cc_242 N_A_27_47#_c_170_n N_A_225_47#_c_988_n 0.00348133f $X=1.72 $Y=1.16 $X2=0
+ $Y2=0
cc_243 N_A_27_47#_c_172_n N_A_225_47#_c_988_n 0.00156368f $X=1.485 $Y=1.217
+ $X2=0 $Y2=0
cc_244 N_A_27_47#_c_173_n N_A_225_47#_c_988_n 4.47034e-19 $X=2.895 $Y=1.217
+ $X2=0 $Y2=0
cc_245 N_A_27_47#_M1026_g N_A_693_47#_c_1030_n 8.91337e-19 $X=2.92 $Y=0.56 $X2=0
+ $Y2=0
cc_246 N_B_c_295_n N_C_M1016_g 2.26972e-19 $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_247 N_B_c_295_n N_C_c_375_n 0.0171123f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_248 B N_C_c_375_n 2.32928e-19 $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_249 N_B_c_295_n N_C_c_376_n 7.96599e-19 $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_250 B N_C_c_376_n 0.0156078f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_251 N_B_c_295_n N_C_c_377_n 2.65226e-19 $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_252 N_B_c_297_n N_VPWR_c_543_n 0.004751f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_298_n N_VPWR_c_544_n 0.0052072f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_299_n N_VPWR_c_544_n 0.004751f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_300_n N_VPWR_c_545_n 0.021146f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_297_n N_VPWR_c_556_n 0.00597712f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_298_n N_VPWR_c_556_n 0.00673617f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_299_n N_VPWR_c_564_n 0.00597712f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_259 N_B_c_300_n N_VPWR_c_564_n 0.00673617f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_260 N_B_c_297_n N_VPWR_c_539_n 0.0100198f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B_c_298_n N_VPWR_c_539_n 0.0118438f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B_c_299_n N_VPWR_c_539_n 0.00999457f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B_c_300_n N_VPWR_c_539_n 0.0132531f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B_c_297_n N_Y_c_724_n 6.24674e-19 $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B_c_297_n N_Y_c_727_n 0.0130707f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_298_n N_Y_c_727_n 0.0106251f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_267 N_B_c_299_n N_Y_c_727_n 6.24674e-19 $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_268 N_B_c_298_n N_Y_c_695_n 0.0153933f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B_c_299_n N_Y_c_695_n 0.0113962f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B_c_295_n N_Y_c_695_n 0.00725062f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_271 B N_Y_c_695_n 0.040258f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_272 N_B_c_298_n N_Y_c_749_n 6.48386e-19 $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B_c_299_n N_Y_c_749_n 0.0130707f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_300_n N_Y_c_749_n 0.0153658f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_275 N_B_c_300_n N_Y_c_696_n 0.0179883f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_276 N_B_c_295_n N_Y_c_696_n 0.00406635f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_277 B N_Y_c_696_n 0.0240956f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_278 N_B_c_297_n N_Y_c_701_n 0.0113403f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_295_n N_Y_c_701_n 0.00160364f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_280 B N_Y_c_701_n 0.0147812f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_281 N_B_c_297_n N_Y_c_702_n 0.00292783f $X=3.365 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B_c_298_n N_Y_c_702_n 0.00116723f $X=3.835 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B_c_295_n N_Y_c_702_n 0.0074788f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_284 B N_Y_c_702_n 0.0305808f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_285 N_B_c_299_n N_Y_c_703_n 0.00292783f $X=4.305 $Y=1.41 $X2=0 $Y2=0
cc_286 N_B_c_300_n N_Y_c_703_n 0.00116723f $X=4.775 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B_c_295_n N_Y_c_703_n 0.0074788f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_288 B N_Y_c_703_n 0.0305808f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_289 N_B_c_295_n Y 0.00113076f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_290 B Y 0.010142f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_291 N_B_M1000_g N_VGND_c_886_n 0.00357877f $X=3.39 $Y=0.56 $X2=0 $Y2=0
cc_292 N_B_M1003_g N_VGND_c_886_n 0.00357877f $X=3.86 $Y=0.56 $X2=0 $Y2=0
cc_293 N_B_M1022_g N_VGND_c_886_n 0.00357877f $X=4.33 $Y=0.56 $X2=0 $Y2=0
cc_294 N_B_M1027_g N_VGND_c_886_n 0.00357877f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_295 N_B_M1000_g N_VGND_c_891_n 0.00550244f $X=3.39 $Y=0.56 $X2=0 $Y2=0
cc_296 N_B_M1003_g N_VGND_c_891_n 0.00548399f $X=3.86 $Y=0.56 $X2=0 $Y2=0
cc_297 N_B_M1022_g N_VGND_c_891_n 0.00548399f $X=4.33 $Y=0.56 $X2=0 $Y2=0
cc_298 N_B_M1027_g N_VGND_c_891_n 0.00668309f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_299 N_B_M1000_g N_A_225_47#_c_988_n 0.00999874f $X=3.39 $Y=0.56 $X2=0 $Y2=0
cc_300 N_B_M1003_g N_A_225_47#_c_988_n 0.00903374f $X=3.86 $Y=0.56 $X2=0 $Y2=0
cc_301 N_B_M1022_g N_A_225_47#_c_988_n 0.00903374f $X=4.33 $Y=0.56 $X2=0 $Y2=0
cc_302 N_B_M1027_g N_A_225_47#_c_988_n 0.00903374f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_303 N_B_c_295_n N_A_225_47#_c_988_n 0.00174447f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_304 B N_A_225_47#_c_988_n 0.00452933f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_305 N_B_M1000_g N_A_693_47#_c_1030_n 0.0082344f $X=3.39 $Y=0.56 $X2=0 $Y2=0
cc_306 N_B_M1003_g N_A_693_47#_c_1030_n 0.0117281f $X=3.86 $Y=0.56 $X2=0 $Y2=0
cc_307 N_B_M1022_g N_A_693_47#_c_1030_n 0.0117281f $X=4.33 $Y=0.56 $X2=0 $Y2=0
cc_308 N_B_M1027_g N_A_693_47#_c_1030_n 0.0146104f $X=4.8 $Y=0.56 $X2=0 $Y2=0
cc_309 N_B_c_295_n N_A_693_47#_c_1030_n 0.0136147f $X=4.8 $Y=1.212 $X2=0 $Y2=0
cc_310 B N_A_693_47#_c_1030_n 0.122218f $X=4.84 $Y=1.19 $X2=0 $Y2=0
cc_311 N_C_M1032_g N_D_M1002_g 0.0178323f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_312 N_C_c_381_n N_D_c_458_n 0.0231619f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_313 N_C_c_376_n N_D_c_455_n 7.08716e-19 $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_314 N_C_c_377_n N_D_c_455_n 0.0178323f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_315 N_C_c_376_n D 0.00629771f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_316 N_C_c_377_n D 7.7315e-19 $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_317 N_C_c_378_n N_VPWR_c_545_n 0.0205167f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_318 N_C_c_379_n N_VPWR_c_546_n 0.0052072f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_319 N_C_c_380_n N_VPWR_c_546_n 0.004751f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_320 N_C_c_381_n N_VPWR_c_547_n 0.0052072f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_321 N_C_c_378_n N_VPWR_c_558_n 0.00597712f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_322 N_C_c_379_n N_VPWR_c_558_n 0.00673617f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_323 N_C_c_380_n N_VPWR_c_560_n 0.00597712f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_324 N_C_c_381_n N_VPWR_c_560_n 0.00673617f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_325 N_C_c_378_n N_VPWR_c_539_n 0.0114039f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_326 N_C_c_379_n N_VPWR_c_539_n 0.0118438f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_327 N_C_c_380_n N_VPWR_c_539_n 0.00999457f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_328 N_C_c_381_n N_VPWR_c_539_n 0.011869f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_329 N_C_c_378_n N_Y_c_696_n 0.0139912f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_330 N_C_c_375_n N_Y_c_696_n 0.00873655f $X=5.665 $Y=1.16 $X2=0 $Y2=0
cc_331 N_C_c_376_n N_Y_c_696_n 0.0398863f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_332 N_C_c_377_n N_Y_c_696_n 2.73568e-19 $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_333 N_C_c_378_n N_Y_c_772_n 0.0178402f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_334 N_C_c_379_n N_Y_c_772_n 0.0106251f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_335 N_C_c_380_n N_Y_c_772_n 6.24674e-19 $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_336 N_C_c_379_n N_Y_c_697_n 0.0153933f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_337 N_C_c_380_n N_Y_c_697_n 0.0113962f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_338 N_C_c_376_n N_Y_c_697_n 0.040258f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_339 N_C_c_377_n N_Y_c_697_n 0.00725062f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_340 N_C_c_379_n N_Y_c_779_n 6.48386e-19 $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_341 N_C_c_380_n N_Y_c_779_n 0.0130707f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_342 N_C_c_381_n N_Y_c_779_n 0.0106251f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_343 N_C_c_381_n N_Y_c_698_n 0.0201997f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_344 N_C_c_376_n N_Y_c_698_n 3.14784e-19 $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_345 N_C_c_377_n N_Y_c_698_n 4.93319e-19 $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_346 N_C_c_381_n N_Y_c_785_n 6.48386e-19 $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_347 N_C_c_378_n N_Y_c_704_n 0.00292783f $X=5.765 $Y=1.41 $X2=0 $Y2=0
cc_348 N_C_c_379_n N_Y_c_704_n 0.00116723f $X=6.235 $Y=1.41 $X2=0 $Y2=0
cc_349 N_C_c_376_n N_Y_c_704_n 0.0305808f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_350 N_C_c_377_n N_Y_c_704_n 0.0074788f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_351 N_C_c_380_n N_Y_c_705_n 0.00292783f $X=6.705 $Y=1.41 $X2=0 $Y2=0
cc_352 N_C_c_381_n N_Y_c_705_n 0.00116723f $X=7.175 $Y=1.41 $X2=0 $Y2=0
cc_353 N_C_c_376_n N_Y_c_705_n 0.0305808f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_354 N_C_c_377_n N_Y_c_705_n 0.0074788f $X=7.175 $Y=1.217 $X2=0 $Y2=0
cc_355 N_C_M1016_g N_VGND_c_886_n 0.00357877f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_356 N_C_M1018_g N_VGND_c_886_n 0.00357877f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_357 N_C_M1029_g N_VGND_c_886_n 0.00357877f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_358 N_C_M1032_g N_VGND_c_886_n 0.00357877f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_359 N_C_M1016_g N_VGND_c_891_n 0.00668309f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_360 N_C_M1018_g N_VGND_c_891_n 0.00548399f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_361 N_C_M1029_g N_VGND_c_891_n 0.00548399f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_362 N_C_M1032_g N_VGND_c_891_n 0.00538422f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_363 N_C_M1016_g N_A_693_47#_c_1030_n 0.0146104f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_364 N_C_M1018_g N_A_693_47#_c_1030_n 0.0117281f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_365 N_C_M1029_g N_A_693_47#_c_1030_n 0.0116916f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_366 N_C_c_375_n N_A_693_47#_c_1030_n 0.0104802f $X=5.665 $Y=1.16 $X2=0 $Y2=0
cc_367 N_C_c_376_n N_A_693_47#_c_1030_n 0.138391f $X=6.945 $Y=1.16 $X2=0 $Y2=0
cc_368 N_C_c_377_n N_A_693_47#_c_1030_n 0.00970138f $X=7.175 $Y=1.217 $X2=0
+ $Y2=0
cc_369 N_C_M1016_g N_A_1081_47#_c_1063_n 0.00903374f $X=5.79 $Y=0.56 $X2=0 $Y2=0
cc_370 N_C_M1018_g N_A_1081_47#_c_1063_n 0.00903374f $X=6.26 $Y=0.56 $X2=0 $Y2=0
cc_371 N_C_M1029_g N_A_1081_47#_c_1063_n 0.00903374f $X=6.73 $Y=0.56 $X2=0 $Y2=0
cc_372 N_C_M1032_g N_A_1081_47#_c_1063_n 0.0137288f $X=7.2 $Y=0.56 $X2=0 $Y2=0
cc_373 N_D_c_458_n N_VPWR_c_547_n 0.004751f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_374 N_D_c_459_n N_VPWR_c_548_n 0.0052072f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_375 N_D_c_460_n N_VPWR_c_548_n 0.004751f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_376 N_D_c_461_n N_VPWR_c_550_n 0.00952555f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_377 N_D_c_456_n N_VPWR_c_550_n 0.00595724f $X=9.32 $Y=1.16 $X2=0 $Y2=0
cc_378 D N_VPWR_c_550_n 0.0206302f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_379 N_D_c_458_n N_VPWR_c_562_n 0.00597712f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_380 N_D_c_459_n N_VPWR_c_562_n 0.00673617f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_381 N_D_c_460_n N_VPWR_c_565_n 0.00597712f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_382 N_D_c_461_n N_VPWR_c_565_n 0.00673617f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_383 N_D_c_458_n N_VPWR_c_539_n 0.0100198f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_384 N_D_c_459_n N_VPWR_c_539_n 0.0118438f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_385 N_D_c_460_n N_VPWR_c_539_n 0.00999457f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_386 N_D_c_461_n N_VPWR_c_539_n 0.0128426f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_387 N_D_c_458_n N_Y_c_779_n 6.24674e-19 $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_388 N_D_c_458_n N_Y_c_698_n 0.0126784f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_389 N_D_c_455_n N_Y_c_698_n 3.62694e-19 $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_390 N_D_c_458_n N_Y_c_785_n 0.0130707f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_391 N_D_c_459_n N_Y_c_785_n 0.0106251f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_392 N_D_c_460_n N_Y_c_785_n 6.24674e-19 $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_393 N_D_c_459_n N_Y_c_699_n 0.0153933f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_394 N_D_c_460_n N_Y_c_699_n 0.0113962f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_395 N_D_c_455_n N_Y_c_699_n 0.00725062f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_396 D N_Y_c_699_n 0.040258f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_397 N_D_c_460_n N_Y_c_700_n 0.00292783f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_398 N_D_c_461_n N_Y_c_700_n 0.00349846f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_399 N_D_c_455_n N_Y_c_700_n 0.0074788f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_400 D N_Y_c_700_n 0.0305808f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_401 N_D_c_459_n N_Y_c_808_n 6.48386e-19 $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_402 N_D_c_460_n N_Y_c_808_n 0.0130707f $X=8.585 $Y=1.41 $X2=0 $Y2=0
cc_403 N_D_c_461_n N_Y_c_808_n 0.0100147f $X=9.055 $Y=1.41 $X2=0 $Y2=0
cc_404 N_D_c_458_n N_Y_c_706_n 0.00292783f $X=7.645 $Y=1.41 $X2=0 $Y2=0
cc_405 N_D_c_459_n N_Y_c_706_n 0.00116723f $X=8.115 $Y=1.41 $X2=0 $Y2=0
cc_406 N_D_c_455_n N_Y_c_706_n 0.0074788f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_407 D N_Y_c_706_n 0.0305808f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_408 N_D_M1002_g N_VGND_c_884_n 0.00375751f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_409 N_D_M1012_g N_VGND_c_884_n 0.00276126f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_410 N_D_M1024_g N_VGND_c_885_n 0.00376026f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_411 N_D_M1028_g N_VGND_c_885_n 0.00276126f $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_412 N_D_M1002_g N_VGND_c_886_n 0.00422898f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_413 N_D_M1012_g N_VGND_c_888_n 0.00424416f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_414 N_D_M1024_g N_VGND_c_888_n 0.00424416f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_415 N_D_M1028_g N_VGND_c_890_n 0.00424416f $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_416 N_D_M1002_g N_VGND_c_891_n 0.00602209f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_417 N_D_M1012_g N_VGND_c_891_n 0.00599001f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_418 N_D_M1024_g N_VGND_c_891_n 0.00611278f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_419 N_D_M1028_g N_VGND_c_891_n 0.00693927f $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_420 N_D_M1002_g N_A_1081_47#_c_1073_n 0.00271016f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_421 N_D_M1002_g N_A_1081_47#_c_1074_n 0.0044152f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_422 N_D_M1012_g N_A_1081_47#_c_1074_n 5.3593e-19 $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_423 N_D_M1002_g N_A_1081_47#_c_1064_n 0.00987731f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_424 N_D_M1012_g N_A_1081_47#_c_1064_n 0.00874287f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_425 N_D_c_455_n N_A_1081_47#_c_1064_n 0.0031956f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_426 D N_A_1081_47#_c_1064_n 0.0334265f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_427 N_D_M1002_g N_A_1081_47#_c_1065_n 0.00140666f $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_428 N_D_M1002_g N_A_1081_47#_c_1081_n 5.82865e-19 $X=7.62 $Y=0.56 $X2=0 $Y2=0
cc_429 N_D_M1012_g N_A_1081_47#_c_1081_n 0.00678142f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_430 N_D_M1024_g N_A_1081_47#_c_1081_n 0.00711907f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_431 N_D_M1028_g N_A_1081_47#_c_1081_n 6.0307e-19 $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_432 N_D_M1024_g N_A_1081_47#_c_1066_n 0.00879805f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_433 N_D_M1028_g N_A_1081_47#_c_1066_n 0.0100812f $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_434 N_D_c_455_n N_A_1081_47#_c_1066_n 0.0120263f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_435 D N_A_1081_47#_c_1066_n 0.0706725f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_436 N_D_M1024_g N_A_1081_47#_c_1067_n 5.82794e-19 $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_437 N_D_M1028_g N_A_1081_47#_c_1067_n 0.00678142f $X=9.03 $Y=0.56 $X2=0 $Y2=0
cc_438 N_D_M1012_g N_A_1081_47#_c_1068_n 0.00113905f $X=8.09 $Y=0.56 $X2=0 $Y2=0
cc_439 N_D_M1024_g N_A_1081_47#_c_1068_n 0.00113905f $X=8.56 $Y=0.56 $X2=0 $Y2=0
cc_440 N_D_c_455_n N_A_1081_47#_c_1068_n 0.00332f $X=9.155 $Y=1.16 $X2=0 $Y2=0
cc_441 D N_A_1081_47#_c_1068_n 0.030602f $X=9.39 $Y=1.19 $X2=0 $Y2=0
cc_442 N_VPWR_c_539_n N_Y_M1006_s 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_443 N_VPWR_c_539_n N_Y_M1020_s 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_444 N_VPWR_c_539_n N_Y_M1004_d 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_445 N_VPWR_c_539_n N_Y_M1025_d 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_446 N_VPWR_c_539_n N_Y_M1001_d 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_447 N_VPWR_c_539_n N_Y_M1021_d 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_448 N_VPWR_c_539_n N_Y_M1005_s 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_449 N_VPWR_c_539_n N_Y_M1008_s 0.00231261f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_450 N_VPWR_c_541_n N_Y_c_693_n 0.0138777f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_451 N_VPWR_c_541_n N_Y_c_717_n 0.065436f $X=1.25 $Y=1.66 $X2=0 $Y2=0
cc_452 N_VPWR_c_542_n N_Y_c_717_n 0.0385613f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_453 N_VPWR_c_552_n N_Y_c_717_n 0.0223557f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_454 N_VPWR_c_539_n N_Y_c_717_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_455 N_VPWR_M1014_d N_Y_c_694_n 0.00180012f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_456 N_VPWR_c_542_n N_Y_c_694_n 0.0139097f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_457 N_VPWR_c_542_n N_Y_c_724_n 0.0470327f $X=2.19 $Y=2 $X2=0 $Y2=0
cc_458 N_VPWR_c_543_n N_Y_c_724_n 0.0385613f $X=3.13 $Y=2 $X2=0 $Y2=0
cc_459 N_VPWR_c_554_n N_Y_c_724_n 0.0223557f $X=3.045 $Y=2.72 $X2=0 $Y2=0
cc_460 N_VPWR_c_539_n N_Y_c_724_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_461 N_VPWR_c_543_n N_Y_c_727_n 0.0470327f $X=3.13 $Y=2 $X2=0 $Y2=0
cc_462 N_VPWR_c_544_n N_Y_c_727_n 0.0385613f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_463 N_VPWR_c_556_n N_Y_c_727_n 0.0223557f $X=3.985 $Y=2.72 $X2=0 $Y2=0
cc_464 N_VPWR_c_539_n N_Y_c_727_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_465 N_VPWR_M1019_s N_Y_c_695_n 0.00180012f $X=3.925 $Y=1.485 $X2=0 $Y2=0
cc_466 N_VPWR_c_544_n N_Y_c_695_n 0.0139097f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_467 N_VPWR_c_544_n N_Y_c_749_n 0.0470327f $X=4.07 $Y=2 $X2=0 $Y2=0
cc_468 N_VPWR_c_545_n N_Y_c_749_n 0.0429581f $X=5.45 $Y=2 $X2=0 $Y2=0
cc_469 N_VPWR_c_564_n N_Y_c_749_n 0.0223557f $X=4.925 $Y=2.72 $X2=0 $Y2=0
cc_470 N_VPWR_c_539_n N_Y_c_749_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_471 N_VPWR_M1033_s N_Y_c_696_n 0.0118304f $X=4.865 $Y=1.485 $X2=0 $Y2=0
cc_472 N_VPWR_c_545_n N_Y_c_696_n 0.0569634f $X=5.45 $Y=2 $X2=0 $Y2=0
cc_473 N_VPWR_c_545_n N_Y_c_772_n 0.0523533f $X=5.45 $Y=2 $X2=0 $Y2=0
cc_474 N_VPWR_c_546_n N_Y_c_772_n 0.0385613f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_475 N_VPWR_c_558_n N_Y_c_772_n 0.0223557f $X=6.385 $Y=2.72 $X2=0 $Y2=0
cc_476 N_VPWR_c_539_n N_Y_c_772_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_477 N_VPWR_M1015_s N_Y_c_697_n 0.00180012f $X=6.325 $Y=1.485 $X2=0 $Y2=0
cc_478 N_VPWR_c_546_n N_Y_c_697_n 0.0139097f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_479 N_VPWR_c_546_n N_Y_c_779_n 0.0470327f $X=6.47 $Y=2 $X2=0 $Y2=0
cc_480 N_VPWR_c_547_n N_Y_c_779_n 0.0385613f $X=7.41 $Y=2 $X2=0 $Y2=0
cc_481 N_VPWR_c_560_n N_Y_c_779_n 0.0223557f $X=7.325 $Y=2.72 $X2=0 $Y2=0
cc_482 N_VPWR_c_539_n N_Y_c_779_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_483 N_VPWR_M1031_s N_Y_c_698_n 0.00180012f $X=7.265 $Y=1.485 $X2=0 $Y2=0
cc_484 N_VPWR_c_547_n N_Y_c_698_n 0.0139097f $X=7.41 $Y=2 $X2=0 $Y2=0
cc_485 N_VPWR_c_547_n N_Y_c_785_n 0.0470327f $X=7.41 $Y=2 $X2=0 $Y2=0
cc_486 N_VPWR_c_548_n N_Y_c_785_n 0.0385613f $X=8.35 $Y=2 $X2=0 $Y2=0
cc_487 N_VPWR_c_562_n N_Y_c_785_n 0.0223557f $X=8.265 $Y=2.72 $X2=0 $Y2=0
cc_488 N_VPWR_c_539_n N_Y_c_785_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_489 N_VPWR_M1007_d N_Y_c_699_n 0.00180012f $X=8.205 $Y=1.485 $X2=0 $Y2=0
cc_490 N_VPWR_c_548_n N_Y_c_699_n 0.0139097f $X=8.35 $Y=2 $X2=0 $Y2=0
cc_491 N_VPWR_c_550_n N_Y_c_700_n 0.0146317f $X=9.29 $Y=1.66 $X2=0 $Y2=0
cc_492 N_VPWR_c_548_n N_Y_c_808_n 0.0470327f $X=8.35 $Y=2 $X2=0 $Y2=0
cc_493 N_VPWR_c_550_n N_Y_c_808_n 0.0504385f $X=9.29 $Y=1.66 $X2=0 $Y2=0
cc_494 N_VPWR_c_565_n N_Y_c_808_n 0.0223557f $X=9.205 $Y=2.72 $X2=0 $Y2=0
cc_495 N_VPWR_c_539_n N_Y_c_808_n 0.0140101f $X=9.43 $Y=2.72 $X2=0 $Y2=0
cc_496 N_VPWR_M1030_d N_Y_c_701_n 0.00180012f $X=2.985 $Y=1.485 $X2=0 $Y2=0
cc_497 N_VPWR_c_543_n N_Y_c_701_n 0.0139097f $X=3.13 $Y=2 $X2=0 $Y2=0
cc_498 N_Y_M1009_s N_VGND_c_891_n 0.00256987f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_499 N_Y_M1013_s N_VGND_c_891_n 0.00256987f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_500 N_Y_c_691_n N_A_225_47#_M1010_d 0.00214196f $X=2.41 $Y=0.77 $X2=0 $Y2=0
cc_501 N_Y_c_691_n N_A_225_47#_c_987_n 0.0216726f $X=2.41 $Y=0.77 $X2=0 $Y2=0
cc_502 N_Y_M1009_s N_A_225_47#_c_988_n 0.00401386f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_503 N_Y_M1013_s N_A_225_47#_c_988_n 0.00400901f $X=2.525 $Y=0.235 $X2=0 $Y2=0
cc_504 N_Y_c_691_n N_A_225_47#_c_988_n 0.0476124f $X=2.41 $Y=0.77 $X2=0 $Y2=0
cc_505 N_Y_c_739_n N_A_225_47#_c_988_n 0.0244305f $X=2.625 $Y=0.905 $X2=0 $Y2=0
cc_506 N_Y_c_696_n N_A_693_47#_c_1030_n 0.00714173f $X=5.785 $Y=1.555 $X2=0
+ $Y2=0
cc_507 N_Y_c_739_n N_A_693_47#_c_1030_n 0.00470114f $X=2.625 $Y=0.905 $X2=0
+ $Y2=0
cc_508 N_Y_c_698_n N_A_1081_47#_c_1064_n 0.00238597f $X=7.665 $Y=1.555 $X2=0
+ $Y2=0
cc_509 N_Y_c_698_n N_A_1081_47#_c_1065_n 0.00936811f $X=7.665 $Y=1.555 $X2=0
+ $Y2=0
cc_510 N_VGND_c_891_n N_A_225_47#_M1009_d 0.00250318f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_511 N_VGND_c_891_n N_A_225_47#_M1010_d 0.00255381f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_512 N_VGND_c_891_n N_A_225_47#_M1026_d 0.00255381f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_513 N_VGND_c_891_n N_A_225_47#_M1003_d 0.00255381f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_514 N_VGND_c_891_n N_A_225_47#_M1027_d 0.00209344f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_515 N_VGND_c_883_n N_A_225_47#_c_986_n 0.0168366f $X=0.73 $Y=0.38 $X2=0 $Y2=0
cc_516 N_VGND_c_886_n N_A_225_47#_c_986_n 0.017577f $X=7.795 $Y=0 $X2=0 $Y2=0
cc_517 N_VGND_c_891_n N_A_225_47#_c_986_n 0.00961661f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_518 N_VGND_c_883_n N_A_225_47#_c_987_n 0.00586971f $X=0.73 $Y=0.38 $X2=0
+ $Y2=0
cc_519 N_VGND_c_886_n N_A_225_47#_c_988_n 0.217929f $X=7.795 $Y=0 $X2=0 $Y2=0
cc_520 N_VGND_c_891_n N_A_225_47#_c_988_n 0.137642f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_521 N_VGND_c_891_n N_A_693_47#_M1000_s 0.00256987f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_522 N_VGND_c_891_n N_A_693_47#_M1022_s 0.00256987f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_523 N_VGND_c_891_n N_A_693_47#_M1016_s 0.00256987f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_524 N_VGND_c_891_n N_A_693_47#_M1029_s 0.00256987f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_525 N_VGND_c_886_n N_A_693_47#_c_1030_n 0.00358979f $X=7.795 $Y=0 $X2=0 $Y2=0
cc_526 N_VGND_c_891_n N_A_693_47#_c_1030_n 0.0126052f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_527 N_VGND_c_891_n N_A_1081_47#_M1016_d 0.00250339f $X=9.43 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_528 N_VGND_c_891_n N_A_1081_47#_M1018_d 0.00255381f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_529 N_VGND_c_891_n N_A_1081_47#_M1032_d 0.00215206f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_530 N_VGND_c_891_n N_A_1081_47#_M1012_s 0.0025535f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_531 N_VGND_c_891_n N_A_1081_47#_M1028_s 0.00250309f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_532 N_VGND_c_886_n N_A_1081_47#_c_1063_n 0.111776f $X=7.795 $Y=0 $X2=0 $Y2=0
cc_533 N_VGND_c_891_n N_A_1081_47#_c_1063_n 0.0703157f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_534 N_VGND_c_884_n N_A_1081_47#_c_1073_n 0.0135136f $X=7.88 $Y=0.38 $X2=0
+ $Y2=0
cc_535 N_VGND_c_886_n N_A_1081_47#_c_1073_n 0.0152108f $X=7.795 $Y=0 $X2=0 $Y2=0
cc_536 N_VGND_c_891_n N_A_1081_47#_c_1073_n 0.00940698f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_537 N_VGND_c_884_n N_A_1081_47#_c_1074_n 0.00471242f $X=7.88 $Y=0.38 $X2=0
+ $Y2=0
cc_538 N_VGND_M1002_d N_A_1081_47#_c_1064_n 0.00259473f $X=7.695 $Y=0.235 $X2=0
+ $Y2=0
cc_539 N_VGND_c_884_n N_A_1081_47#_c_1064_n 0.0115453f $X=7.88 $Y=0.38 $X2=0
+ $Y2=0
cc_540 N_VGND_c_886_n N_A_1081_47#_c_1064_n 0.00260082f $X=7.795 $Y=0 $X2=0
+ $Y2=0
cc_541 N_VGND_c_888_n N_A_1081_47#_c_1064_n 0.00193763f $X=8.735 $Y=0 $X2=0
+ $Y2=0
cc_542 N_VGND_c_891_n N_A_1081_47#_c_1064_n 0.00964063f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_543 N_VGND_c_885_n N_A_1081_47#_c_1081_n 0.0177507f $X=8.82 $Y=0.38 $X2=0
+ $Y2=0
cc_544 N_VGND_c_888_n N_A_1081_47#_c_1081_n 0.0223596f $X=8.735 $Y=0 $X2=0 $Y2=0
cc_545 N_VGND_c_891_n N_A_1081_47#_c_1081_n 0.0141302f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_546 N_VGND_M1024_d N_A_1081_47#_c_1066_n 0.00259473f $X=8.635 $Y=0.235 $X2=0
+ $Y2=0
cc_547 N_VGND_c_885_n N_A_1081_47#_c_1066_n 0.0115453f $X=8.82 $Y=0.38 $X2=0
+ $Y2=0
cc_548 N_VGND_c_888_n N_A_1081_47#_c_1066_n 0.00260082f $X=8.735 $Y=0 $X2=0
+ $Y2=0
cc_549 N_VGND_c_890_n N_A_1081_47#_c_1066_n 0.00193763f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_550 N_VGND_c_891_n N_A_1081_47#_c_1066_n 0.00964063f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_551 N_VGND_c_890_n N_A_1081_47#_c_1067_n 0.0248368f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_552 N_VGND_c_891_n N_A_1081_47#_c_1067_n 0.0145275f $X=9.43 $Y=0 $X2=0 $Y2=0
cc_553 N_A_225_47#_c_988_n N_A_693_47#_M1000_s 0.00401386f $X=5.01 $Y=0.38
+ $X2=-0.19 $Y2=-0.24
cc_554 N_A_225_47#_c_988_n N_A_693_47#_M1022_s 0.00401386f $X=5.01 $Y=0.38 $X2=0
+ $Y2=0
cc_555 N_A_225_47#_M1003_d N_A_693_47#_c_1030_n 0.00214196f $X=3.935 $Y=0.235
+ $X2=0 $Y2=0
cc_556 N_A_225_47#_M1027_d N_A_693_47#_c_1030_n 0.00321334f $X=4.875 $Y=0.235
+ $X2=0 $Y2=0
cc_557 N_A_225_47#_c_988_n N_A_693_47#_c_1030_n 0.0981138f $X=5.01 $Y=0.38 $X2=0
+ $Y2=0
cc_558 N_A_225_47#_c_988_n N_A_1081_47#_c_1063_n 0.0180052f $X=5.01 $Y=0.38
+ $X2=0 $Y2=0
cc_559 N_A_693_47#_c_1030_n N_A_1081_47#_M1016_d 0.00442235f $X=6.94 $Y=0.72
+ $X2=-0.19 $Y2=-0.24
cc_560 N_A_693_47#_c_1030_n N_A_1081_47#_M1018_d 0.00214196f $X=6.94 $Y=0.72
+ $X2=0 $Y2=0
cc_561 N_A_693_47#_M1016_s N_A_1081_47#_c_1063_n 0.00401386f $X=5.865 $Y=0.235
+ $X2=0 $Y2=0
cc_562 N_A_693_47#_M1029_s N_A_1081_47#_c_1063_n 0.00401386f $X=6.805 $Y=0.235
+ $X2=0 $Y2=0
cc_563 N_A_693_47#_c_1030_n N_A_1081_47#_c_1063_n 0.0963535f $X=6.94 $Y=0.72
+ $X2=0 $Y2=0
cc_564 N_A_693_47#_c_1030_n N_A_1081_47#_c_1065_n 0.00140356f $X=6.94 $Y=0.72
+ $X2=0 $Y2=0
