* File: sky130_fd_sc_hdll__dfstp_4.pex.spice
* Created: Thu Aug 27 19:04:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%CLK 4 5 7 8 10 13 19 20 24 26
c41 13 0 2.71124e-20 $X=0.52 $Y=0.805
r42 24 27 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.4
r43 24 26 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.245 $Y=1.235
+ $X2=0.245 $Y2=1.07
r44 19 20 11.1952 $w=3.48e-07 $l=3.4e-07 $layer=LI1_cond $X=0.265 $Y=1.19
+ $X2=0.265 $Y2=1.53
r45 19 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.235 $X2=0.245 $Y2=1.235
r46 11 13 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=0.305 $Y=0.805
+ $X2=0.52 $Y2=0.805
r47 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r48 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r49 5 15 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.495 $Y=1.665
+ $X2=0.305 $Y2=1.665
r50 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r51 4 15 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.665
r52 4 27 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=1.59
+ $X2=0.305 $Y2=1.4
r53 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=0.805
r54 1 26 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.305 $Y=0.88
+ $X2=0.305 $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_27_47# 1 2 8 9 11 14 16 18 19 21 22 24
+ 25 27 30 34 35 36 39 41 45 46 49 50 51 53 54 68 72 73 75 76 77 82 90 96
c262 73 0 3.46126e-20 $X=2.875 $Y=1.825
c263 50 0 1.75333e-19 $X=6.37 $Y=0.81
c264 46 0 9.81997e-20 $X=2.585 $Y=0.87
c265 36 0 1.76957e-19 $X=0.66 $Y=1.88
c266 22 0 1.37207e-19 $X=5.54 $Y=1.99
c267 19 0 2.53929e-20 $X=2.96 $Y=1.99
r268 93 104 7.06336 $w=3.08e-07 $l=1.9e-07 $layer=LI1_cond $X=5.605 $Y=1.81
+ $X2=5.415 $Y2=1.81
r269 92 93 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.605
+ $Y=1.74 $X2=5.605 $Y2=1.74
r270 89 90 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.965
+ $Y=1.74 $X2=2.965 $Y2=1.74
r271 81 82 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.235
+ $X2=0.99 $Y2=1.235
r272 76 93 6.87748 $w=3.08e-07 $l=1.85e-07 $layer=LI1_cond $X=5.79 $Y=1.81
+ $X2=5.605 $Y2=1.81
r273 75 77 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.79 $Y=1.825
+ $X2=5.645 $Y2=1.825
r274 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.79 $Y=1.825
+ $X2=5.79 $Y2=1.825
r275 73 77 3.42821 $w=1.4e-07 $l=2.77e-06 $layer=MET1_cond $X=2.875 $Y=1.87
+ $X2=5.645 $Y2=1.87
r276 71 90 7.12695 $w=3.78e-07 $l=2.35e-07 $layer=LI1_cond $X=2.73 $Y=1.765
+ $X2=2.965 $Y2=1.765
r277 71 99 2.88111 $w=3.78e-07 $l=9.5e-08 $layer=LI1_cond $X=2.73 $Y=1.765
+ $X2=2.635 $Y2=1.765
r278 70 73 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.73 $Y=1.825
+ $X2=2.875 $Y2=1.825
r279 70 72 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.73 $Y=1.825
+ $X2=2.585 $Y2=1.825
r280 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.73 $Y=1.825
+ $X2=2.73 $Y2=1.825
r281 68 72 2.09158 $w=1.4e-07 $l=1.69e-06 $layer=MET1_cond $X=0.895 $Y=1.87
+ $X2=2.585 $Y2=1.87
r282 65 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.75 $Y=1.825
+ $X2=0.895 $Y2=1.825
r283 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.75 $Y=1.825
+ $X2=0.75 $Y2=1.825
r284 58 96 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=6.535 $Y=0.93
+ $X2=6.645 $Y2=0.93
r285 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.535
+ $Y=0.93 $X2=6.535 $Y2=0.93
r286 54 57 3.63929 $w=3.78e-07 $l=1.2e-07 $layer=LI1_cond $X=6.56 $Y=0.81
+ $X2=6.56 $Y2=0.93
r287 50 54 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.37 $Y=0.81
+ $X2=6.56 $Y2=0.81
r288 50 51 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=6.37 $Y=0.81
+ $X2=5.5 $Y2=0.81
r289 49 104 4.25403 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=5.415 $Y=1.655
+ $X2=5.415 $Y2=1.81
r290 48 51 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.415 $Y=0.895
+ $X2=5.5 $Y2=0.81
r291 48 49 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=5.415 $Y=0.895
+ $X2=5.415 $Y2=1.655
r292 46 84 22.732 $w=3.3e-07 $l=1.3e-07 $layer=POLY_cond $X=2.585 $Y=0.87
+ $X2=2.455 $Y2=0.87
r293 45 46 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.585
+ $Y=0.87 $X2=2.585 $Y2=0.87
r294 43 99 2.7393 $w=2.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.635 $Y=1.575
+ $X2=2.635 $Y2=1.765
r295 43 45 30.0916 $w=2.68e-07 $l=7.05e-07 $layer=LI1_cond $X=2.635 $Y=1.575
+ $X2=2.635 $Y2=0.87
r296 42 81 35.5478 $w=2.7e-07 $l=1.6e-07 $layer=POLY_cond $X=0.805 $Y=1.235
+ $X2=0.965 $Y2=1.235
r297 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.805
+ $Y=1.235 $X2=0.805 $Y2=1.235
r298 39 66 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.88
r299 39 41 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.775 $Y=1.795
+ $X2=0.775 $Y2=1.235
r300 38 41 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.775 $Y=0.805
+ $X2=0.775 $Y2=1.235
r301 37 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=1.88
+ $X2=0.26 $Y2=1.88
r302 36 66 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.775 $Y2=1.88
r303 36 37 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=1.88
+ $X2=0.345 $Y2=1.88
r304 34 38 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.775 $Y2=0.805
r305 34 35 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.66 $Y=0.72
+ $X2=0.345 $Y2=0.72
r306 28 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r307 28 30 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r308 25 96 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=6.645 $Y=0.765
+ $X2=6.645 $Y2=0.93
r309 25 27 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=6.645 $Y=0.765
+ $X2=6.645 $Y2=0.445
r310 22 92 46.5577 $w=3.26e-07 $l=2.91548e-07 $layer=POLY_cond $X=5.54 $Y=1.99
+ $X2=5.63 $Y2=1.74
r311 22 24 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.54 $Y=1.99
+ $X2=5.54 $Y2=2.275
r312 19 89 46.5577 $w=3.26e-07 $l=2.64575e-07 $layer=POLY_cond $X=2.96 $Y=1.99
+ $X2=2.99 $Y2=1.74
r313 19 21 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.96 $Y=1.99
+ $X2=2.96 $Y2=2.275
r314 16 84 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=2.455 $Y=0.705
+ $X2=2.455 $Y2=0.87
r315 16 18 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.455 $Y=0.705
+ $X2=2.455 $Y2=0.415
r316 12 82 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=1.235
r317 12 14 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.99 $Y=1.1
+ $X2=0.99 $Y2=0.445
r318 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r319 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.64 $X2=0.965
+ $Y2=1.74
r320 7 81 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.37
+ $X2=0.965 $Y2=1.235
r321 7 8 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.965 $Y=1.37 $X2=0.965
+ $Y2=1.64
r322 2 53 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r323 1 30 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%D 1 3 6 8 9 14
c38 1 0 1.46624e-19 $X=1.955 $Y=1.57
r39 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.955
+ $Y=1.17 $X2=1.955 $Y2=1.17
r40 8 9 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=2.1 $Y=1.19 $X2=2.1
+ $Y2=1.53
r41 8 14 0.520034 $w=4.58e-07 $l=2e-08 $layer=LI1_cond $X=2.1 $Y=1.19 $X2=2.1
+ $Y2=1.17
r42 4 13 38.9026 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.98 $Y=1.005
+ $X2=1.98 $Y2=1.17
r43 4 6 230.745 $w=1.5e-07 $l=4.5e-07 $layer=POLY_cond $X=1.98 $Y=1.005 $X2=1.98
+ $Y2=0.555
r44 1 13 76.7755 $w=2.7e-07 $l=4.12311e-07 $layer=POLY_cond $X=1.955 $Y=1.57
+ $X2=1.98 $Y2=1.17
r45 1 3 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=1.955 $Y=1.57
+ $X2=1.955 $Y2=2.065
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_211_363# 1 2 8 9 11 12 13 16 19 21 24 26
+ 28 29 30 31 34 36 41 43 44 49 50 51 58 63
c199 51 0 1.51904e-19 $X=5.665 $Y=1.195
c200 50 0 4.09811e-20 $X=5.81 $Y=1.195
c201 49 0 2.54518e-19 $X=5.81 $Y=1.195
c202 36 0 2.53929e-20 $X=3.385 $Y=1.19
c203 34 0 9.81997e-20 $X=3.277 $Y=1.12
c204 30 0 1.75333e-19 $X=5.97 $Y=1.125
c205 21 0 1.7977e-19 $X=6.13 $Y=1.89
c206 8 0 4.36039e-20 $X=2.49 $Y=1.89
r207 58 61 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=0.93
+ $X2=3.165 $Y2=1.095
r208 58 60 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.165 $Y=0.93
+ $X2=3.165 $Y2=0.765
r209 50 54 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.815
+ $Y=1.26 $X2=5.815 $Y2=1.26
r210 49 51 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.81 $Y=1.195
+ $X2=5.665 $Y2=1.195
r211 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.81 $Y=1.195
+ $X2=5.81 $Y2=1.195
r212 46 47 0.0440827 $w=2.9e-07 $l=7e-08 $layer=MET1_cond $X=3.24 $Y=0.85
+ $X2=3.24 $Y2=0.92
r213 44 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.165
+ $Y=0.93 $X2=3.165 $Y2=0.93
r214 43 46 0.0220415 $w=2.9e-07 $l=4.5e-08 $layer=MET1_cond $X=3.24 $Y=0.805
+ $X2=3.24 $Y2=0.85
r215 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.24 $Y=0.805
+ $X2=3.24 $Y2=0.805
r216 39 67 59.1587 $w=2.23e-07 $l=1.155e-06 $layer=LI1_cond $X=1.227 $Y=0.805
+ $X2=1.227 $Y2=1.96
r217 39 63 15.1098 $w=2.23e-07 $l=2.95e-07 $layer=LI1_cond $X=1.227 $Y=0.805
+ $X2=1.227 $Y2=0.51
r218 38 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.25 $Y=0.805
+ $X2=1.395 $Y2=0.805
r219 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.25 $Y=0.805
+ $X2=1.25 $Y2=0.805
r220 36 51 2.82178 $w=1.4e-07 $l=2.28e-06 $layer=MET1_cond $X=3.385 $Y=1.19
+ $X2=5.665 $Y2=1.19
r221 34 36 0.0739737 $w=1.4e-07 $l=1.38651e-07 $layer=MET1_cond $X=3.277 $Y=1.12
+ $X2=3.385 $Y2=1.19
r222 34 47 0.142799 $w=2.15e-07 $l=2e-07 $layer=MET1_cond $X=3.277 $Y=1.12
+ $X2=3.277 $Y2=0.92
r223 31 46 0.0513368 $w=1.4e-07 $l=1.45e-07 $layer=MET1_cond $X=3.095 $Y=0.85
+ $X2=3.24 $Y2=0.85
r224 31 41 2.10396 $w=1.4e-07 $l=1.7e-06 $layer=MET1_cond $X=3.095 $Y=0.85
+ $X2=1.395 $Y2=0.85
r225 29 54 34.4369 $w=2.7e-07 $l=1.55e-07 $layer=POLY_cond $X=5.97 $Y=1.26
+ $X2=5.815 $Y2=1.26
r226 29 30 0.63749 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=5.97 $Y=1.26
+ $X2=5.97 $Y2=1.125
r227 26 28 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.13 $Y=1.99
+ $X2=6.13 $Y2=2.275
r228 22 30 28.793 $w=1.75e-07 $l=1.45e-07 $layer=POLY_cond $X=6.115 $Y=1.125
+ $X2=5.97 $Y2=1.125
r229 22 24 348.681 $w=1.5e-07 $l=6.8e-07 $layer=POLY_cond $X=6.115 $Y=1.125
+ $X2=6.115 $Y2=0.445
r230 21 26 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.13 $Y=1.89 $X2=6.13
+ $Y2=1.99
r231 20 30 28.793 $w=1.75e-07 $l=4.02119e-07 $layer=POLY_cond $X=6.13 $Y=1.455
+ $X2=5.97 $Y2=1.125
r232 20 21 144.236 $w=2e-07 $l=4.35e-07 $layer=POLY_cond $X=6.13 $Y=1.455
+ $X2=6.13 $Y2=1.89
r233 19 61 76.9149 $w=1.5e-07 $l=1.5e-07 $layer=POLY_cond $X=3.105 $Y=1.245
+ $X2=3.105 $Y2=1.095
r234 16 60 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.105 $Y=0.415
+ $X2=3.105 $Y2=0.765
r235 12 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.03 $Y=1.32
+ $X2=3.105 $Y2=1.245
r236 12 13 225.617 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=3.03 $Y=1.32
+ $X2=2.59 $Y2=1.32
r237 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.49 $Y=1.99
+ $X2=2.49 $Y2=2.275
r238 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.49 $Y=1.89 $X2=2.49
+ $Y2=1.99
r239 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=2.49 $Y=1.395
+ $X2=2.59 $Y2=1.32
r240 7 8 164.131 $w=2e-07 $l=4.95e-07 $layer=POLY_cond $X=2.49 $Y=1.395 $X2=2.49
+ $Y2=1.89
r241 2 67 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r242 1 63 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_702_21# 1 2 9 11 13 14 18 20 24 27 29 34
+ 36
c108 36 0 2.23858e-19 $X=4.95 $Y=1.065
c109 34 0 2.11834e-19 $X=4.425 $Y=1.96
c110 29 0 1.15651e-19 $X=3.695 $Y=1.74
r111 35 36 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=4.95 $Y=0.725
+ $X2=4.95 $Y2=1.065
r112 29 32 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=3.76 $Y=1.74
+ $X2=3.76 $Y2=1.96
r113 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.695
+ $Y=1.74 $X2=3.695 $Y2=1.74
r114 27 36 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.025 $Y=1.835
+ $X2=5.025 $Y2=1.065
r115 24 35 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=4.875 $Y=0.46
+ $X2=4.875 $Y2=0.725
r116 21 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.51 $Y=1.96
+ $X2=4.425 $Y2=1.96
r117 20 27 7.14316 $w=2.5e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.94 $Y=1.96
+ $X2=5.025 $Y2=1.835
r118 20 21 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.94 $Y=1.96
+ $X2=4.51 $Y2=1.96
r119 16 34 2.76166 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.085
+ $X2=4.425 $Y2=1.96
r120 16 18 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=4.425 $Y=2.085
+ $X2=4.425 $Y2=2.21
r121 15 32 1.80669 $w=2.5e-07 $l=1.5e-07 $layer=LI1_cond $X=3.91 $Y=1.96
+ $X2=3.76 $Y2=1.96
r122 14 34 3.70735 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.34 $Y=1.96
+ $X2=4.425 $Y2=1.96
r123 14 15 19.822 $w=2.48e-07 $l=4.3e-07 $layer=LI1_cond $X=4.34 $Y=1.96
+ $X2=3.91 $Y2=1.96
r124 11 30 46.2237 $w=3.35e-07 $l=2.89396e-07 $layer=POLY_cond $X=3.61 $Y=1.99
+ $X2=3.695 $Y2=1.74
r125 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.61 $Y=1.99
+ $X2=3.61 $Y2=2.275
r126 7 30 38.6365 $w=3.35e-07 $l=2.13014e-07 $layer=POLY_cond $X=3.585 $Y=1.575
+ $X2=3.695 $Y2=1.74
r127 7 9 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=3.585 $Y=1.575
+ $X2=3.585 $Y2=0.445
r128 2 18 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.28
+ $Y=2.065 $X2=4.425 $Y2=2.21
r129 1 24 182 $w=1.7e-07 $l=3.03727e-07 $layer=licon1_NDIFF $count=1 $X=4.69
+ $Y=0.235 $X2=4.875 $Y2=0.46
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%SET_B 2 3 5 8 12 17 18 20 21 22 23 24 26
+ 29 34 37 38 44
c130 44 0 7.40925e-20 $X=4.365 $Y=0.85
c131 26 0 1.71107e-19 $X=7.59 $Y=0.85
c132 24 0 3.91725e-20 $X=4.51 $Y=0.85
c133 23 0 1.86694e-20 $X=7.445 $Y=0.85
c134 8 0 1.90694e-19 $X=4.255 $Y=0.445
c135 3 0 1.15651e-19 $X=4.19 $Y=1.99
r136 37 40 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=0.98
+ $X2=7.45 $Y2=1.145
r137 37 39 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.45 $Y=0.98
+ $X2=7.45 $Y2=0.815
r138 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.425
+ $Y=0.98 $X2=7.425 $Y2=0.98
r139 34 35 10.074 $w=3.11e-07 $l=6.5e-08 $layer=POLY_cond $X=4.19 $Y=0.98
+ $X2=4.255 $Y2=0.98
r140 33 44 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=4.075 $Y=0.9
+ $X2=4.365 $Y2=0.9
r141 32 34 17.8232 $w=3.11e-07 $l=1.15e-07 $layer=POLY_cond $X=4.075 $Y=0.98
+ $X2=4.19 $Y2=0.98
r142 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.075
+ $Y=0.98 $X2=4.075 $Y2=0.98
r143 29 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.365 $Y=0.85
+ $X2=4.365 $Y2=0.85
r144 26 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0.85
+ $X2=7.59 $Y2=0.85
r145 24 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.51 $Y=0.85
+ $X2=4.365 $Y2=0.85
r146 23 26 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.445 $Y=0.85
+ $X2=7.59 $Y2=0.85
r147 23 24 3.63242 $w=1.4e-07 $l=2.935e-06 $layer=MET1_cond $X=7.445 $Y=0.85
+ $X2=4.51 $Y2=0.85
r148 21 22 43.7534 $w=2.2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.52 $Y=1.535
+ $X2=7.52 $Y2=1.685
r149 21 40 129.315 $w=2e-07 $l=3.9e-07 $layer=POLY_cond $X=7.51 $Y=1.535
+ $X2=7.51 $Y2=1.145
r150 18 20 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.53 $Y=1.99
+ $X2=7.53 $Y2=2.275
r151 17 18 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.53 $Y=1.89 $X2=7.53
+ $Y2=1.99
r152 17 22 67.9733 $w=2e-07 $l=2.05e-07 $layer=POLY_cond $X=7.53 $Y=1.89
+ $X2=7.53 $Y2=1.685
r153 12 39 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=7.365 $Y=0.445
+ $X2=7.365 $Y2=0.815
r154 6 35 19.8172 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.255 $Y=0.815
+ $X2=4.255 $Y2=0.98
r155 6 8 189.723 $w=1.5e-07 $l=3.7e-07 $layer=POLY_cond $X=4.255 $Y=0.815
+ $X2=4.255 $Y2=0.445
r156 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.19 $Y=1.99
+ $X2=4.19 $Y2=2.275
r157 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.19 $Y=1.89 $X2=4.19
+ $Y2=1.99
r158 1 34 13.1188 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.19 $Y=1.145
+ $X2=4.19 $Y2=0.98
r159 1 2 247.025 $w=2e-07 $l=7.45e-07 $layer=POLY_cond $X=4.19 $Y=1.145 $X2=4.19
+ $Y2=1.89
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_506_47# 1 2 7 9 11 13 14 16 17 20 21 23
+ 24 26 27 28 32 37 39 40 45 46 56
c160 56 0 1.34022e-19 $X=5.13 $Y=1.4
c161 46 0 3.91725e-20 $X=4.62 $Y=1.32
c162 45 0 4.36039e-20 $X=3.74 $Y=1.317
c163 24 0 3.31643e-20 $X=5.705 $Y=0.735
c164 17 0 1.50733e-19 $X=5.63 $Y=0.825
r165 55 56 82.1848 $w=3.3e-07 $l=4.7e-07 $layer=POLY_cond $X=4.66 $Y=1.4
+ $X2=5.13 $Y2=1.4
r166 54 55 3.49723 $w=3.3e-07 $l=2e-08 $layer=POLY_cond $X=4.64 $Y=1.4 $X2=4.66
+ $Y2=1.4
r167 50 54 0.874306 $w=3.3e-07 $l=5e-09 $layer=POLY_cond $X=4.635 $Y=1.4
+ $X2=4.64 $Y2=1.4
r168 49 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.635
+ $Y=1.4 $X2=4.635 $Y2=1.4
r169 46 49 3.07318 $w=2.98e-07 $l=8e-08 $layer=LI1_cond $X=4.62 $Y=1.32 $X2=4.62
+ $Y2=1.4
r170 40 46 4.061 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=4.47 $Y=1.32 $X2=4.62
+ $Y2=1.32
r171 40 45 47.6257 $w=1.68e-07 $l=7.3e-07 $layer=LI1_cond $X=4.47 $Y=1.32
+ $X2=3.74 $Y2=1.32
r172 39 45 6.97143 $w=1.73e-07 $l=1.1e-07 $layer=LI1_cond $X=3.63 $Y=1.317
+ $X2=3.74 $Y2=1.317
r173 39 42 17.4286 $w=1.73e-07 $l=2.75e-07 $layer=LI1_cond $X=3.63 $Y=1.317
+ $X2=3.355 $Y2=1.317
r174 38 39 40.0736 $w=2.18e-07 $l=7.65e-07 $layer=LI1_cond $X=3.63 $Y=0.465
+ $X2=3.63 $Y2=1.23
r175 36 42 0.89264 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=3.355 $Y=1.405
+ $X2=3.355 $Y2=1.317
r176 36 37 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=3.355 $Y=1.405
+ $X2=3.355 $Y2=2.25
r177 32 38 6.83662 $w=2e-07 $l=1.51987e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=3.63 $Y2=0.465
r178 32 34 40.4818 $w=1.98e-07 $l=7.3e-07 $layer=LI1_cond $X=3.52 $Y=0.365
+ $X2=2.79 $Y2=0.365
r179 28 37 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.27 $Y=2.335
+ $X2=3.355 $Y2=2.25
r180 28 30 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.27 $Y=2.335
+ $X2=2.725 $Y2=2.335
r181 24 26 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.705 $Y=0.735
+ $X2=5.705 $Y2=0.445
r182 21 23 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.13 $Y=1.99
+ $X2=5.13 $Y2=2.275
r183 20 21 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=5.13 $Y=1.89 $X2=5.13
+ $Y2=1.99
r184 19 56 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=5.13 $Y=1.565
+ $X2=5.13 $Y2=1.4
r185 19 20 107.763 $w=2e-07 $l=3.25e-07 $layer=POLY_cond $X=5.13 $Y=1.565
+ $X2=5.13 $Y2=1.89
r186 18 27 4.90422 $w=1.8e-07 $l=1e-07 $layer=POLY_cond $X=4.74 $Y=0.825
+ $X2=4.64 $Y2=0.825
r187 17 24 27.2212 $w=1.8e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.63 $Y=0.825
+ $X2=5.705 $Y2=0.735
r188 17 18 345.952 $w=1.8e-07 $l=8.9e-07 $layer=POLY_cond $X=5.63 $Y=0.825
+ $X2=4.74 $Y2=0.825
r189 14 16 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=4.66 $Y=1.99
+ $X2=4.66 $Y2=2.275
r190 13 14 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.66 $Y=1.89 $X2=4.66
+ $Y2=1.99
r191 12 55 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.66 $Y=1.565
+ $X2=4.66 $Y2=1.4
r192 12 13 107.763 $w=2e-07 $l=3.25e-07 $layer=POLY_cond $X=4.66 $Y=1.565
+ $X2=4.66 $Y2=1.89
r193 11 54 14.4873 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.64 $Y=1.235
+ $X2=4.64 $Y2=1.4
r194 10 27 20.8929 $w=1.75e-07 $l=9e-08 $layer=POLY_cond $X=4.64 $Y=0.915
+ $X2=4.64 $Y2=0.825
r195 10 11 106.105 $w=2e-07 $l=3.2e-07 $layer=POLY_cond $X=4.64 $Y=0.915
+ $X2=4.64 $Y2=1.235
r196 7 27 20.8929 $w=1.75e-07 $l=1.01735e-07 $layer=POLY_cond $X=4.615 $Y=0.735
+ $X2=4.64 $Y2=0.825
r197 7 9 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.615 $Y=0.735
+ $X2=4.615 $Y2=0.445
r198 2 30 600 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=1 $X=2.58
+ $Y=2.065 $X2=2.725 $Y2=2.335
r199 1 34 182 $w=1.7e-07 $l=3.245e-07 $layer=licon1_NDIFF $count=1 $X=2.53
+ $Y=0.235 $X2=2.79 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1288_261# 1 2 7 9 12 21 24 28 31 32
c72 31 0 1.7977e-19 $X=8.21 $Y=1.67
c73 24 0 1.58039e-19 $X=8.445 $Y=1.575
c74 7 0 5.96505e-20 $X=6.54 $Y=1.99
r75 30 32 8.75598 $w=1.88e-07 $l=1.5e-07 $layer=LI1_cond $X=8.295 $Y=1.67
+ $X2=8.445 $Y2=1.67
r76 30 31 5.10991 $w=1.88e-07 $l=8.5e-08 $layer=LI1_cond $X=8.295 $Y=1.67
+ $X2=8.21 $Y2=1.67
r77 26 28 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=8.295 $Y=0.515
+ $X2=8.445 $Y2=0.515
r78 24 32 0.0965754 $w=2.1e-07 $l=9.5e-08 $layer=LI1_cond $X=8.445 $Y=1.575
+ $X2=8.445 $Y2=1.67
r79 23 28 3.38185 $w=2.1e-07 $l=1.65e-07 $layer=LI1_cond $X=8.445 $Y=0.68
+ $X2=8.445 $Y2=0.515
r80 23 24 47.2684 $w=2.08e-07 $l=8.95e-07 $layer=LI1_cond $X=8.445 $Y=0.68
+ $X2=8.445 $Y2=1.575
r81 19 30 1.386 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=8.295 $Y=1.765
+ $X2=8.295 $Y2=1.67
r82 19 21 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=8.295 $Y=1.765
+ $X2=8.295 $Y2=1.87
r83 16 31 103.406 $w=1.68e-07 $l=1.585e-06 $layer=LI1_cond $X=6.625 $Y=1.66
+ $X2=8.21 $Y2=1.66
r84 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.625
+ $Y=1.66 $X2=6.625 $Y2=1.66
r85 10 17 62.9618 $w=3.88e-07 $l=4.61519e-07 $layer=POLY_cond $X=7.005 $Y=1.305
+ $X2=6.76 $Y2=1.66
r86 10 12 440.979 $w=1.5e-07 $l=8.6e-07 $layer=POLY_cond $X=7.005 $Y=1.305
+ $X2=7.005 $Y2=0.445
r87 7 17 54.9609 $w=3.88e-07 $l=4.26028e-07 $layer=POLY_cond $X=6.54 $Y=1.99
+ $X2=6.76 $Y2=1.66
r88 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.54 $Y=1.99 $X2=6.54
+ $Y2=2.275
r89 2 21 300 $w=1.7e-07 $l=2.88531e-07 $layer=licon1_PDIFF $count=2 $X=8.15
+ $Y=1.645 $X2=8.295 $Y2=1.87
r90 1 26 182 $w=1.7e-07 $l=3.40881e-07 $layer=licon1_NDIFF $count=1 $X=8.16
+ $Y=0.235 $X2=8.295 $Y2=0.515
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1126_413# 1 2 3 10 12 15 17 18 20 21 23
+ 26 28 29 34 35 39 40 41 44 49 51 54 56 58
c163 54 0 9.39049e-20 $X=7.005 $Y=1.32
c164 10 0 1.58039e-19 $X=8.06 $Y=1.57
r165 61 62 2.90361 $w=4.15e-07 $l=2.5e-08 $layer=POLY_cond $X=8.06 $Y=1.332
+ $X2=8.085 $Y2=1.332
r166 57 61 12.1952 $w=4.15e-07 $l=1.05e-07 $layer=POLY_cond $X=7.955 $Y=1.332
+ $X2=8.06 $Y2=1.332
r167 56 58 9.07524 $w=2.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.955 $Y=1.29
+ $X2=7.79 $Y2=1.29
r168 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.955
+ $Y=1.26 $X2=7.955 $Y2=1.26
r169 47 49 6.00231 $w=2.38e-07 $l=1.25e-07 $layer=LI1_cond $X=7.26 $Y=2.085
+ $X2=7.26 $Y2=2.21
r170 46 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.09 $Y=1.32
+ $X2=7.005 $Y2=1.32
r171 46 58 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.09 $Y=1.32 $X2=7.79
+ $Y2=1.32
r172 44 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.005 $Y=1.235
+ $X2=7.005 $Y2=1.32
r173 43 44 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=7.005 $Y=0.475
+ $X2=7.005 $Y2=1.235
r174 42 51 2.2496 $w=1.7e-07 $l=1.1e-07 $layer=LI1_cond $X=6.29 $Y=2 $X2=6.18
+ $Y2=2
r175 41 47 7.07814 $w=1.7e-07 $l=1.56844e-07 $layer=LI1_cond $X=7.14 $Y=2
+ $X2=7.26 $Y2=2.085
r176 41 42 55.4545 $w=1.68e-07 $l=8.5e-07 $layer=LI1_cond $X=7.14 $Y=2 $X2=6.29
+ $Y2=2
r177 39 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.92 $Y=1.32
+ $X2=7.005 $Y2=1.32
r178 39 40 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=6.92 $Y=1.32
+ $X2=6.29 $Y2=1.32
r179 35 43 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.92 $Y=0.39
+ $X2=7.005 $Y2=0.475
r180 35 37 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=6.92 $Y=0.39
+ $X2=6.355 $Y2=0.39
r181 34 51 4.45262 $w=2.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.18 $Y=1.915
+ $X2=6.18 $Y2=2
r182 33 40 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.18 $Y=1.405
+ $X2=6.29 $Y2=1.32
r183 33 34 26.7157 $w=2.18e-07 $l=5.1e-07 $layer=LI1_cond $X=6.18 $Y=1.405
+ $X2=6.18 $Y2=1.915
r184 29 51 15.1913 $w=2.18e-07 $l=2.9e-07 $layer=LI1_cond $X=6.18 $Y=2.29
+ $X2=6.18 $Y2=2
r185 29 31 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=6.07 $Y=2.29
+ $X2=5.775 $Y2=2.29
r186 24 28 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=9.075 $Y=1.095
+ $X2=9.05 $Y2=1.26
r187 24 26 333.298 $w=1.5e-07 $l=6.5e-07 $layer=POLY_cond $X=9.075 $Y=1.095
+ $X2=9.075 $Y2=0.445
r188 21 23 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=9.05 $Y=1.77
+ $X2=9.05 $Y2=2.165
r189 20 21 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.05 $Y=1.67 $X2=9.05
+ $Y2=1.77
r190 19 28 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=9.05 $Y=1.425
+ $X2=9.05 $Y2=1.26
r191 19 20 81.2364 $w=2e-07 $l=2.45e-07 $layer=POLY_cond $X=9.05 $Y=1.425
+ $X2=9.05 $Y2=1.67
r192 18 62 10.8699 $w=4.15e-07 $l=1.05e-07 $layer=POLY_cond $X=8.16 $Y=1.26
+ $X2=8.085 $Y2=1.332
r193 17 28 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=8.95 $Y=1.26 $X2=9.05
+ $Y2=1.26
r194 17 18 138.14 $w=3.3e-07 $l=7.9e-07 $layer=POLY_cond $X=8.95 $Y=1.26
+ $X2=8.16 $Y2=1.26
r195 13 62 26.7644 $w=1.5e-07 $l=2.37e-07 $layer=POLY_cond $X=8.085 $Y=1.095
+ $X2=8.085 $Y2=1.332
r196 13 15 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.085 $Y=1.095
+ $X2=8.085 $Y2=0.505
r197 10 61 22.3416 $w=1.8e-07 $l=2.38e-07 $layer=POLY_cond $X=8.06 $Y=1.57
+ $X2=8.06 $Y2=1.332
r198 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.06 $Y=1.57
+ $X2=8.06 $Y2=2.065
r199 3 49 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=7.17
+ $Y=2.065 $X2=7.295 $Y2=2.21
r200 2 31 600 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_PDIFF $count=1 $X=5.63
+ $Y=2.065 $X2=5.775 $Y2=2.33
r201 1 37 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=6.19
+ $Y=0.235 $X2=6.355 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_1738_47# 1 2 9 11 13 16 18 20 23 25 27
+ 30 32 34 35 37 40 46 55 59 60 61 72
r125 72 73 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=11.455 $Y=1.217
+ $X2=11.48 $Y2=1.217
r126 69 70 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=10.96 $Y=1.217
+ $X2=10.985 $Y2=1.217
r127 68 69 65.9969 $w=3.25e-07 $l=4.45e-07 $layer=POLY_cond $X=10.515 $Y=1.217
+ $X2=10.96 $Y2=1.217
r128 67 68 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=10.49 $Y=1.217
+ $X2=10.515 $Y2=1.217
r129 66 67 65.9969 $w=3.25e-07 $l=4.45e-07 $layer=POLY_cond $X=10.045 $Y=1.217
+ $X2=10.49 $Y2=1.217
r130 65 66 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=10.02 $Y=1.217
+ $X2=10.045 $Y2=1.217
r131 62 63 3.70769 $w=3.25e-07 $l=2.5e-08 $layer=POLY_cond $X=9.55 $Y=1.217
+ $X2=9.575 $Y2=1.217
r132 59 60 3.67308 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=8.815 $Y=2
+ $X2=8.815 $Y2=1.915
r133 56 72 37.8185 $w=3.25e-07 $l=2.55e-07 $layer=POLY_cond $X=11.2 $Y=1.217
+ $X2=11.455 $Y2=1.217
r134 56 70 31.8862 $w=3.25e-07 $l=2.15e-07 $layer=POLY_cond $X=11.2 $Y=1.217
+ $X2=10.985 $Y2=1.217
r135 55 56 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=11.2
+ $Y=1.16 $X2=11.2 $Y2=1.16
r136 53 65 56.3569 $w=3.25e-07 $l=3.8e-07 $layer=POLY_cond $X=9.64 $Y=1.217
+ $X2=10.02 $Y2=1.217
r137 53 63 9.64 $w=3.25e-07 $l=6.5e-08 $layer=POLY_cond $X=9.64 $Y=1.217
+ $X2=9.575 $Y2=1.217
r138 52 55 81.7187 $w=2.18e-07 $l=1.56e-06 $layer=LI1_cond $X=9.64 $Y=1.165
+ $X2=11.2 $Y2=1.165
r139 52 53 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=9.64
+ $Y=1.16 $X2=9.64 $Y2=1.16
r140 50 61 1.80668 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=8.98 $Y=1.165
+ $X2=8.855 $Y2=1.165
r141 50 52 34.5733 $w=2.18e-07 $l=6.6e-07 $layer=LI1_cond $X=8.98 $Y=1.165
+ $X2=9.64 $Y2=1.165
r142 48 61 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.855 $Y=1.275
+ $X2=8.855 $Y2=1.165
r143 48 60 29.5025 $w=2.48e-07 $l=6.4e-07 $layer=LI1_cond $X=8.855 $Y=1.275
+ $X2=8.855 $Y2=1.915
r144 44 61 4.63873 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=8.855 $Y=1.055
+ $X2=8.855 $Y2=1.165
r145 44 46 25.1233 $w=2.48e-07 $l=5.45e-07 $layer=LI1_cond $X=8.855 $Y=1.055
+ $X2=8.855 $Y2=0.51
r146 38 73 20.86 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=11.48 $Y=1.025
+ $X2=11.48 $Y2=1.217
r147 38 40 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.48 $Y=1.025
+ $X2=11.48 $Y2=0.56
r148 35 72 16.5763 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.217
r149 35 37 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=11.455 $Y=1.41
+ $X2=11.455 $Y2=1.985
r150 32 70 16.5763 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.217
r151 32 34 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.985 $Y=1.41
+ $X2=10.985 $Y2=1.985
r152 28 69 20.86 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.96 $Y=1.025
+ $X2=10.96 $Y2=1.217
r153 28 30 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.96 $Y=1.025
+ $X2=10.96 $Y2=0.56
r154 25 68 16.5763 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.217
r155 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.515 $Y=1.41
+ $X2=10.515 $Y2=1.985
r156 21 67 20.86 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.49 $Y=1.025
+ $X2=10.49 $Y2=1.217
r157 21 23 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.49 $Y=1.025
+ $X2=10.49 $Y2=0.56
r158 18 66 16.5763 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.045 $Y=1.41
+ $X2=10.045 $Y2=1.217
r159 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.045 $Y=1.41
+ $X2=10.045 $Y2=1.985
r160 14 65 20.86 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.02 $Y=1.025
+ $X2=10.02 $Y2=1.217
r161 14 16 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.02 $Y=1.025
+ $X2=10.02 $Y2=0.56
r162 11 63 16.5763 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.575 $Y=1.41
+ $X2=9.575 $Y2=1.217
r163 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.575 $Y=1.41
+ $X2=9.575 $Y2=1.985
r164 7 62 20.86 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.55 $Y=1.025
+ $X2=9.55 $Y2=1.217
r165 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.55 $Y=1.025
+ $X2=9.55 $Y2=0.56
r166 2 59 300 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_PDIFF $count=2 $X=8.69
+ $Y=1.845 $X2=8.815 $Y2=2
r167 1 46 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=8.69
+ $Y=0.235 $X2=8.815 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 30 32 36 40 44 48
+ 52 55 56 58 59 60 62 64 70 78 83 95 106 112 113 116 119 122 129 136 143 146
c196 1 0 1.76957e-19 $X=0.585 $Y=1.815
r197 146 147 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r198 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r199 139 140 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r200 136 139 9.67042 $w=4.68e-07 $l=3.8e-07 $layer=LI1_cond $X=6.705 $Y=2.34
+ $X2=6.705 $Y2=2.72
r201 132 133 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r202 129 132 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=4.87 $Y=2.34
+ $X2=4.87 $Y2=2.72
r203 125 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r204 122 125 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=3.92 $Y=2.34
+ $X2=3.92 $Y2=2.72
r205 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r206 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.61 $Y2=2.72
r207 116 117 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r208 113 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r209 112 113 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r210 110 146 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.435 $Y=2.72
+ $X2=11.245 $Y2=2.72
r211 110 112 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.435 $Y=2.72
+ $X2=11.73 $Y2=2.72
r212 109 147 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=2.72
+ $X2=11.27 $Y2=2.72
r213 108 109 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r214 106 146 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.055 $Y=2.72
+ $X2=11.245 $Y2=2.72
r215 106 108 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.055 $Y=2.72
+ $X2=10.81 $Y2=2.72
r216 105 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.81 $Y2=2.72
r217 105 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=9.43 $Y2=2.72
r218 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r219 102 143 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=9.545 $Y=2.72
+ $X2=9.367 $Y2=2.72
r220 102 104 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=9.545 $Y=2.72
+ $X2=9.89 $Y2=2.72
r221 101 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.43 $Y2=2.72
r222 100 101 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r223 98 101 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r224 97 100 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r225 97 98 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r226 95 143 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=9.19 $Y=2.72
+ $X2=9.367 $Y2=2.72
r227 95 100 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.19 $Y=2.72
+ $X2=8.97 $Y2=2.72
r228 94 98 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.05 $Y2=2.72
r229 94 140 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r230 93 94 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r231 91 139 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=6.705 $Y2=2.72
r232 91 93 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=6.94 $Y=2.72
+ $X2=7.59 $Y2=2.72
r233 90 140 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r234 89 90 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r235 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r236 87 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.83 $Y2=2.72
r237 86 89 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r238 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r239 84 132 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=4.87 $Y2=2.72
r240 84 86 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=5.06 $Y=2.72
+ $X2=5.29 $Y2=2.72
r241 83 139 6.76998 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=6.47 $Y=2.72
+ $X2=6.705 $Y2=2.72
r242 83 89 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=6.47 $Y=2.72
+ $X2=6.21 $Y2=2.72
r243 82 133 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r244 82 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r245 81 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r246 79 125 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=3.92 $Y2=2.72
r247 79 81 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=4.37 $Y2=2.72
r248 78 132 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.68 $Y=2.72
+ $X2=4.87 $Y2=2.72
r249 78 81 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=4.68 $Y=2.72
+ $X2=4.37 $Y2=2.72
r250 77 126 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r251 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r252 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r253 74 120 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r254 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=3.45 $Y2=2.72
r255 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r256 71 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=1.72 $Y2=2.72
r257 71 73 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=2.72
+ $X2=2.07 $Y2=2.72
r258 70 125 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.92 $Y2=2.72
r259 70 76 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.45 $Y2=2.72
r260 64 116 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r261 62 117 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r262 60 64 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=0.515 $Y2=2.72
r263 60 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r264 58 104 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=10.165 $Y=2.72
+ $X2=9.89 $Y2=2.72
r265 58 59 7.13466 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=10.165 $Y=2.72
+ $X2=10.292 $Y2=2.72
r266 57 108 25.4438 $w=1.68e-07 $l=3.9e-07 $layer=LI1_cond $X=10.42 $Y=2.72
+ $X2=10.81 $Y2=2.72
r267 57 59 7.13466 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=10.42 $Y=2.72
+ $X2=10.292 $Y2=2.72
r268 55 93 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r269 55 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.875 $Y2=2.72
r270 54 97 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=8.05 $Y2=2.72
r271 54 56 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=8.04 $Y=2.72
+ $X2=7.875 $Y2=2.72
r272 50 146 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.245 $Y=2.635
+ $X2=11.245 $Y2=2.72
r273 50 52 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=11.245 $Y=2.635
+ $X2=11.245 $Y2=2.02
r274 46 59 0.067832 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=10.292 $Y=2.635
+ $X2=10.292 $Y2=2.72
r275 46 48 21.4671 $w=2.53e-07 $l=4.75e-07 $layer=LI1_cond $X=10.292 $Y=2.635
+ $X2=10.292 $Y2=2.16
r276 42 143 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=9.367 $Y=2.635
+ $X2=9.367 $Y2=2.72
r277 42 44 20.6141 $w=3.53e-07 $l=6.35e-07 $layer=LI1_cond $X=9.367 $Y=2.635
+ $X2=9.367 $Y2=2
r278 38 56 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.72
r279 38 40 14.8421 $w=3.28e-07 $l=4.25e-07 $layer=LI1_cond $X=7.875 $Y=2.635
+ $X2=7.875 $Y2=2.21
r280 34 119 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.72
r281 34 36 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=1.72 $Y=2.635
+ $X2=1.72 $Y2=2.22
r282 33 116 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r283 32 119 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=1.72 $Y2=2.72
r284 32 33 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=2.72
+ $X2=0.895 $Y2=2.72
r285 28 116 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r286 28 30 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.22
r287 9 52 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=11.075
+ $Y=1.485 $X2=11.22 $Y2=2.02
r288 8 48 600 $w=1.7e-07 $l=7.43976e-07 $layer=licon1_PDIFF $count=1 $X=10.135
+ $Y=1.485 $X2=10.28 $Y2=2.16
r289 7 44 300 $w=1.7e-07 $l=2.66458e-07 $layer=licon1_PDIFF $count=2 $X=9.14
+ $Y=1.845 $X2=9.34 $Y2=2
r290 6 40 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=7.62
+ $Y=2.065 $X2=7.825 $Y2=2.21
r291 5 136 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=6.63
+ $Y=2.065 $X2=6.775 $Y2=2.34
r292 4 129 600 $w=1.7e-07 $l=3.39853e-07 $layer=licon1_PDIFF $count=1 $X=4.75
+ $Y=2.065 $X2=4.895 $Y2=2.34
r293 3 122 600 $w=1.7e-07 $l=3.59514e-07 $layer=licon1_PDIFF $count=1 $X=3.7
+ $Y=2.065 $X2=3.895 $Y2=2.34
r294 2 36 600 $w=1.7e-07 $l=6.34429e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.645 $X2=1.72 $Y2=2.22
r295 1 30 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%A_409_329# 1 2 8 9 10 11 12 15 20
c59 20 0 1.81236e-19 $X=2.19 $Y=1.96
r60 13 15 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.19 $Y=0.635
+ $X2=2.19 $Y2=0.47
r61 11 20 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=1.88
+ $X2=2.19 $Y2=1.88
r62 11 12 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=2.105 $Y=1.88
+ $X2=1.7 $Y2=1.88
r63 9 13 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=2.105 $Y=0.73
+ $X2=2.19 $Y2=0.635
r64 9 10 23.6411 $w=1.88e-07 $l=4.05e-07 $layer=LI1_cond $X=2.105 $Y=0.73
+ $X2=1.7 $Y2=0.73
r65 8 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.615 $Y=1.795
+ $X2=1.7 $Y2=1.88
r66 7 10 6.84389 $w=1.9e-07 $l=1.30767e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.7 $Y2=0.73
r67 7 8 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=1.615 $Y=0.825
+ $X2=1.615 $Y2=1.795
r68 2 20 300 $w=1.7e-07 $l=3.80657e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.645 $X2=2.19 $Y2=1.96
r69 1 15 182 $w=1.7e-07 $l=2.94873e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%Q 1 2 3 4 5 6 19 20 21 22 23 28 30 32 36
+ 37 38 39 40 41 42 43 44 45 46
r90 69 74 3.84148 $w=2.53e-07 $l=8.5e-08 $layer=LI1_cond $X=11.732 $Y=0.715
+ $X2=11.732 $Y2=0.63
r91 45 46 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=11.732 $Y=1.82
+ $X2=11.732 $Y2=2.21
r92 45 81 8.13489 $w=2.53e-07 $l=1.8e-07 $layer=LI1_cond $X=11.732 $Y=1.82
+ $X2=11.732 $Y2=1.64
r93 44 76 3.67481 $w=2.52e-07 $l=8.6487e-08 $layer=LI1_cond $X=11.732 $Y=1.555
+ $X2=11.735 $Y2=1.47
r94 44 81 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=11.732 $Y=1.555
+ $X2=11.732 $Y2=1.64
r95 44 76 0.59927 $w=2.48e-07 $l=1.3e-08 $layer=LI1_cond $X=11.735 $Y=1.457
+ $X2=11.735 $Y2=1.47
r96 43 44 12.3081 $w=2.48e-07 $l=2.67e-07 $layer=LI1_cond $X=11.735 $Y=1.19
+ $X2=11.735 $Y2=1.457
r97 42 69 3.67481 $w=2.52e-07 $l=8.5e-08 $layer=LI1_cond $X=11.732 $Y=0.8
+ $X2=11.732 $Y2=0.715
r98 42 75 3.67481 $w=2.52e-07 $l=8.6487e-08 $layer=LI1_cond $X=11.732 $Y=0.8
+ $X2=11.735 $Y2=0.885
r99 42 43 12.9074 $w=2.48e-07 $l=2.8e-07 $layer=LI1_cond $X=11.735 $Y=0.91
+ $X2=11.735 $Y2=1.19
r100 42 75 1.15244 $w=2.48e-07 $l=2.5e-08 $layer=LI1_cond $X=11.735 $Y=0.91
+ $X2=11.735 $Y2=0.885
r101 41 74 5.42326 $w=2.53e-07 $l=1.2e-07 $layer=LI1_cond $X=11.732 $Y=0.51
+ $X2=11.732 $Y2=0.63
r102 39 40 16.6464 $w=2.68e-07 $l=3.9e-07 $layer=LI1_cond $X=9.86 $Y=1.82
+ $X2=9.86 $Y2=2.21
r103 38 62 4.60977 $w=2.98e-07 $l=1.2e-07 $layer=LI1_cond $X=9.875 $Y=0.51
+ $X2=9.875 $Y2=0.63
r104 35 39 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=9.86 $Y=1.64
+ $X2=9.86 $Y2=1.82
r105 34 62 3.26526 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=9.875 $Y=0.715
+ $X2=9.875 $Y2=0.63
r106 33 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.835 $Y=1.555
+ $X2=10.75 $Y2=1.555
r107 32 44 2.79892 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.605 $Y=1.555
+ $X2=11.732 $Y2=1.555
r108 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=11.605 $Y=1.555
+ $X2=10.835 $Y2=1.555
r109 31 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.835 $Y=0.8
+ $X2=10.75 $Y2=0.8
r110 30 42 2.79892 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=11.605 $Y=0.8
+ $X2=11.732 $Y2=0.8
r111 30 31 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=11.605 $Y=0.8
+ $X2=10.835 $Y2=0.8
r112 26 37 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=1.64
+ $X2=10.75 $Y2=1.555
r113 26 28 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.75 $Y=1.64
+ $X2=10.75 $Y2=1.82
r114 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.715
+ $X2=10.75 $Y2=0.8
r115 23 25 6.1 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.75 $Y=0.715 $X2=10.75
+ $Y2=0.63
r116 22 34 7.51767 $w=1.7e-07 $l=1.8775e-07 $layer=LI1_cond $X=10.025 $Y=0.8
+ $X2=9.875 $Y2=0.715
r117 21 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.665 $Y=0.8
+ $X2=10.75 $Y2=0.8
r118 21 22 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=10.665 $Y=0.8
+ $X2=10.025 $Y2=0.8
r119 20 35 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=9.995 $Y=1.555
+ $X2=9.86 $Y2=1.64
r120 19 37 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.665 $Y=1.555
+ $X2=10.75 $Y2=1.555
r121 19 20 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=10.665 $Y=1.555
+ $X2=9.995 $Y2=1.555
r122 6 45 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=11.545
+ $Y=1.485 $X2=11.69 $Y2=1.82
r123 5 28 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=10.605
+ $Y=1.485 $X2=10.75 $Y2=1.82
r124 4 39 300 $w=1.7e-07 $l=4.00999e-07 $layer=licon1_PDIFF $count=2 $X=9.665
+ $Y=1.485 $X2=9.81 $Y2=1.82
r125 3 74 182 $w=1.7e-07 $l=4.57548e-07 $layer=licon1_NDIFF $count=1 $X=11.555
+ $Y=0.235 $X2=11.69 $Y2=0.63
r126 2 25 182 $w=1.7e-07 $l=4.78644e-07 $layer=licon1_NDIFF $count=1 $X=10.565
+ $Y=0.235 $X2=10.75 $Y2=0.63
r127 1 62 182 $w=1.7e-07 $l=4.78644e-07 $layer=licon1_NDIFF $count=1 $X=9.625
+ $Y=0.235 $X2=9.81 $Y2=0.63
.ends

.subckt PM_SKY130_FD_SC_HDLL__DFSTP_4%VGND 1 2 3 4 5 6 7 8 25 29 33 37 41 45 48
+ 49 50 52 54 60 65 85 89 96 97 101 107 110 117 122 125 127 130
c192 122 0 3.3422e-20 $X=7.32 $Y=0.24
c193 97 0 2.71124e-20 $X=11.73 $Y=0
c194 5 0 1.71107e-19 $X=7.44 $Y=0.235
r195 130 131 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r196 127 128 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r197 124 125 13.0581 $w=6.48e-07 $l=3.05e-07 $layer=LI1_cond $X=7.725 $Y=0.24
+ $X2=8.03 $Y2=0.24
r198 120 124 2.48416 $w=6.48e-07 $l=1.35e-07 $layer=LI1_cond $X=7.59 $Y=0.24
+ $X2=7.725 $Y2=0.24
r199 120 122 12.4141 $w=6.48e-07 $l=2.7e-07 $layer=LI1_cond $X=7.59 $Y=0.24
+ $X2=7.32 $Y2=0.24
r200 120 121 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r201 117 118 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r202 110 114 9.36061 $w=4.58e-07 $l=3.6e-07 $layer=LI1_cond $X=4.14 $Y=0
+ $X2=4.14 $Y2=0.36
r203 110 111 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r204 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0
+ $X2=1.61 $Y2=0
r205 102 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=1.61 $Y2=0
r206 101 104 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r207 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r208 97 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r209 96 97 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r210 94 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.435 $Y=0
+ $X2=11.245 $Y2=0
r211 94 96 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=11.435 $Y=0
+ $X2=11.73 $Y2=0
r212 93 131 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r213 93 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=10.35 $Y2=0
r214 92 93 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r215 90 127 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.345 $Y2=0
r216 90 92 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.495 $Y=0
+ $X2=10.81 $Y2=0
r217 89 130 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=11.245 $Y2=0
r218 89 92 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=11.055 $Y=0
+ $X2=10.81 $Y2=0
r219 88 128 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.35 $Y2=0
r220 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r221 85 127 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=10.345 $Y2=0
r222 85 87 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=10.195 $Y=0
+ $X2=9.89 $Y2=0
r223 84 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r224 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r225 81 84 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r226 81 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.05 $Y=0
+ $X2=7.59 $Y2=0
r227 80 83 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r228 80 125 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.03
+ $Y2=0
r229 80 81 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r230 77 121 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=7.59 $Y2=0
r231 76 122 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=7.13 $Y=0 $X2=7.32
+ $Y2=0
r232 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r233 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=7.13 $Y2=0
r234 74 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=5.29 $Y2=0
r235 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=5.75 $Y=0 $X2=7.13
+ $Y2=0
r236 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r237 71 117 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.335
+ $Y2=0
r238 71 73 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=5.53 $Y=0 $X2=5.75
+ $Y2=0
r239 69 118 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.29 $Y2=0
r240 69 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=3.91 $Y2=0
r241 68 69 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r242 66 110 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.14
+ $Y2=0
r243 66 68 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=4.83
+ $Y2=0
r244 65 117 9.6488 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=5.335
+ $Y2=0
r245 65 68 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.14 $Y=0 $X2=4.83
+ $Y2=0
r246 64 111 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=3.91 $Y2=0
r247 64 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=1.61 $Y2=0
r248 63 64 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r249 61 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=1.72 $Y2=0
r250 61 63 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=0
+ $X2=2.07 $Y2=0
r251 60 110 6.6364 $w=1.7e-07 $l=2.3e-07 $layer=LI1_cond $X=3.91 $Y=0 $X2=4.14
+ $Y2=0
r252 60 63 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.91 $Y=0 $X2=2.07
+ $Y2=0
r253 54 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.705 $Y2=0
r254 52 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r255 50 54 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.515 $Y2=0
r256 50 52 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r257 48 83 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=9.19 $Y=0 $X2=8.97
+ $Y2=0
r258 48 49 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=9.19 $Y=0 $X2=9.332
+ $Y2=0
r259 47 87 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.475 $Y=0
+ $X2=9.89 $Y2=0
r260 47 49 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=9.475 $Y=0
+ $X2=9.332 $Y2=0
r261 43 130 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.245 $Y=0.085
+ $X2=11.245 $Y2=0
r262 43 45 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=11.245 $Y=0.085
+ $X2=11.245 $Y2=0.38
r263 39 127 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0
r264 39 41 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=10.345 $Y=0.085
+ $X2=10.345 $Y2=0.38
r265 35 49 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=9.332 $Y=0.085
+ $X2=9.332 $Y2=0
r266 35 37 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=9.332 $Y=0.085
+ $X2=9.332 $Y2=0.38
r267 31 117 1.39532 $w=3.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.335 $Y=0.085
+ $X2=5.335 $Y2=0
r268 31 33 8.7172 $w=3.88e-07 $l=2.95e-07 $layer=LI1_cond $X=5.335 $Y=0.085
+ $X2=5.335 $Y2=0.38
r269 27 107 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0
r270 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.72 $Y=0.085
+ $X2=1.72 $Y2=0.38
r271 26 101 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=0.705 $Y2=0
r272 25 107 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=1.72 $Y2=0
r273 25 26 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.555 $Y=0
+ $X2=0.895 $Y2=0
r274 8 45 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=11.035
+ $Y=0.235 $X2=11.22 $Y2=0.38
r275 7 41 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=10.095
+ $Y=0.235 $X2=10.28 $Y2=0.38
r276 6 37 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=9.15
+ $Y=0.235 $X2=9.34 $Y2=0.38
r277 5 124 182 $w=1.7e-07 $l=3.88652e-07 $layer=licon1_NDIFF $count=1 $X=7.44
+ $Y=0.235 $X2=7.725 $Y2=0.48
r278 4 33 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.32
+ $Y=0.235 $X2=5.445 $Y2=0.38
r279 3 114 182 $w=1.7e-07 $l=3.92556e-07 $layer=licon1_NDIFF $count=1 $X=3.66
+ $Y=0.235 $X2=3.995 $Y2=0.36
r280 2 29 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.72 $Y2=0.38
r281 1 104 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

