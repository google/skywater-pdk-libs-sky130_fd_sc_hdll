* File: sky130_fd_sc_hdll__or4_2.pex.spice
* Created: Thu Aug 27 19:24:55 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR4_2%D 1 3 6 8 9 15
c28 8 0 1.35736e-19 $X=0.235 $Y=0.85
r29 15 16 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r30 13 15 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r31 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r32 8 9 10.2074 $w=3.48e-07 $l=3.1e-07 $layer=LI1_cond $X=0.26 $Y=0.85 $X2=0.26
+ $Y2=1.16
r33 4 16 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r34 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.475
r35 1 15 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r36 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%C 1 3 6 8 9 10 11 20 27
r35 18 27 4.14769 $w=6.18e-07 $l=2.15e-07 $layer=LI1_cond $X=0.94 $Y=1.305
+ $X2=1.155 $Y2=1.305
r36 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.94
+ $Y=1.16 $X2=0.94 $Y2=1.16
r37 10 11 0.578748 $w=6.18e-07 $l=3e-08 $layer=LI1_cond $X=1.16 $Y=1.305
+ $X2=1.19 $Y2=1.305
r38 10 27 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=1.16 $Y=1.305
+ $X2=1.155 $Y2=1.305
r39 9 18 3.76186 $w=6.18e-07 $l=1.95e-07 $layer=LI1_cond $X=0.745 $Y=1.305
+ $X2=0.94 $Y2=1.305
r40 8 9 0.675206 $w=6.18e-07 $l=3.5e-08 $layer=LI1_cond $X=0.71 $Y=1.305
+ $X2=0.745 $Y2=1.305
r41 8 20 0.289374 $w=6.18e-07 $l=1.5e-08 $layer=LI1_cond $X=0.71 $Y=1.305
+ $X2=0.695 $Y2=1.305
r42 4 17 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=1.05 $Y=0.995
+ $X2=0.965 $Y2=1.16
r43 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.05 $Y=0.995 $X2=1.05
+ $Y2=0.475
r44 1 17 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=0.965 $Y2=1.16
r45 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.025 $Y=1.41
+ $X2=1.025 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%B 2 3 4 6 9 10 11 12 13 14 15 27 30
c44 11 0 6.13246e-20 $X=1.465 $Y=0.91
c45 4 0 1.73735e-19 $X=1.435 $Y=2.035
c46 2 0 8.49032e-20 $X=1.435 $Y=1.31
r47 15 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.52
+ $Y=2.28 $X2=1.52 $Y2=2.28
r48 14 15 13.9088 $w=2.88e-07 $l=3.5e-07 $layer=LI1_cond $X=1.17 $Y=2.27
+ $X2=1.52 $Y2=2.27
r49 14 30 0.198697 $w=2.88e-07 $l=5e-09 $layer=LI1_cond $X=1.17 $Y=2.27
+ $X2=1.165 $Y2=2.27
r50 13 30 17.8827 $w=2.88e-07 $l=4.5e-07 $layer=LI1_cond $X=0.715 $Y=2.27
+ $X2=1.165 $Y2=2.27
r51 13 27 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=0.715 $Y=2.27
+ $X2=0.695 $Y2=2.27
r52 12 27 18.2801 $w=2.88e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=2.27
+ $X2=0.695 $Y2=2.27
r53 10 11 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=1.465 $Y=0.76
+ $X2=1.465 $Y2=0.91
r54 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.52 $Y=0.475 $X2=1.52
+ $Y2=0.76
r55 4 21 46.6963 $w=3.06e-07 $l=2.8e-07 $layer=POLY_cond $X=1.435 $Y=2.035
+ $X2=1.51 $Y2=2.28
r56 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.435 $Y=2.035
+ $X2=1.435 $Y2=1.695
r57 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.695
r58 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.435 $Y=1.31 $X2=1.435
+ $Y2=1.41
r59 2 11 132.631 $w=2e-07 $l=4e-07 $layer=POLY_cond $X=1.435 $Y=1.31 $X2=1.435
+ $Y2=0.91
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%A 1 3 6 8 12 14
r41 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.925
+ $Y=1.16 $X2=1.925 $Y2=1.16
r42 8 12 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.925 $Y2=1.16
r43 8 14 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=1.765 $Y=1.16
+ $X2=1.615 $Y2=1.16
r44 4 11 38.578 $w=2.95e-07 $l=1.83916e-07 $layer=POLY_cond $X=1.99 $Y=0.995
+ $X2=1.95 $Y2=1.16
r45 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.99 $Y=0.995 $X2=1.99
+ $Y2=0.475
r46 1 11 48.1208 $w=2.95e-07 $l=2.57391e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.95 $Y2=1.16
r47 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.965 $Y=1.41
+ $X2=1.965 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%A_27_297# 1 2 3 10 12 13 15 16 18 19 21 23
+ 24 25 26 30 32 33 36 38 40 43 45 47 51 52 59
c122 52 0 1.73735e-19 $X=1.745 $Y=1.58
c123 45 0 1.07404e-19 $X=2.35 $Y=1.495
r124 59 60 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.615
+ $Y=1.16 $X2=2.615 $Y2=1.16
r125 56 59 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.35 $Y=1.16
+ $X2=2.615 $Y2=1.16
r126 52 54 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=1.745 $Y=1.58
+ $X2=1.745 $Y2=1.87
r127 47 49 6.56006 $w=3.23e-07 $l=1.85e-07 $layer=LI1_cond $X=0.247 $Y=1.685
+ $X2=0.247 $Y2=1.87
r128 44 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=1.325
+ $X2=2.35 $Y2=1.16
r129 44 45 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.35 $Y=1.325
+ $X2=2.35 $Y2=1.495
r130 43 56 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.35 $Y=0.995
+ $X2=2.35 $Y2=1.16
r131 42 43 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.35 $Y=0.825
+ $X2=2.35 $Y2=0.995
r132 41 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.83 $Y=1.58
+ $X2=1.745 $Y2=1.58
r133 40 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=1.58
+ $X2=2.35 $Y2=1.495
r134 40 41 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=2.265 $Y=1.58
+ $X2=1.83 $Y2=1.58
r135 39 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.815 $Y=0.74
+ $X2=1.73 $Y2=0.74
r136 38 42 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.265 $Y=0.74
+ $X2=2.35 $Y2=0.825
r137 38 39 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.265 $Y=0.74
+ $X2=1.815 $Y2=0.74
r138 34 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.73 $Y=0.655
+ $X2=1.73 $Y2=0.74
r139 34 36 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.73 $Y=0.655
+ $X2=1.73 $Y2=0.47
r140 32 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.74
+ $X2=1.73 $Y2=0.74
r141 32 33 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.645 $Y=0.74
+ $X2=0.845 $Y2=0.74
r142 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.845 $Y2=0.74
r143 28 30 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.76 $Y=0.655
+ $X2=0.76 $Y2=0.47
r144 27 49 4.53325 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=0.41 $Y=1.87
+ $X2=0.247 $Y2=1.87
r145 26 54 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=1.745 $Y2=1.87
r146 26 27 81.5508 $w=1.68e-07 $l=1.25e-06 $layer=LI1_cond $X=1.66 $Y=1.87
+ $X2=0.41 $Y2=1.87
r147 24 60 74.316 $w=3.3e-07 $l=4.25e-07 $layer=POLY_cond $X=3.04 $Y=1.16
+ $X2=2.615 $Y2=1.16
r148 24 25 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.04 $Y=1.16
+ $X2=3.14 $Y2=1.202
r149 22 60 1.74861 $w=3.3e-07 $l=1e-08 $layer=POLY_cond $X=2.605 $Y=1.16
+ $X2=2.615 $Y2=1.16
r150 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=2.605 $Y=1.16
+ $X2=2.505 $Y2=1.202
r151 19 25 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=3.165 $Y=0.995
+ $X2=3.14 $Y2=1.202
r152 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.165 $Y=0.995
+ $X2=3.165 $Y2=0.56
r153 16 25 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=3.14 $Y=1.41
+ $X2=3.14 $Y2=1.202
r154 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.14 $Y=1.41
+ $X2=3.14 $Y2=1.985
r155 13 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.202
r156 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.505 $Y=1.41
+ $X2=2.505 $Y2=1.985
r157 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.505 $Y2=1.202
r158 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.48 $Y=0.995
+ $X2=2.48 $Y2=0.56
r159 3 47 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.685
r160 2 36 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.265 $X2=1.73 $Y2=0.47
r161 1 30 182 $w=1.7e-07 $l=2.75409e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.265 $X2=0.76 $Y2=0.47
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%VPWR 1 2 9 11 13 18 19 20 29 35
c31 1 0 1.07404e-19 $X=2.055 $Y=1.485
r32 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r33 32 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r34 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r35 29 34 3.73837 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=3.497 $Y2=2.72
r36 29 31 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=2.72
+ $X2=2.99 $Y2=2.72
r37 28 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r38 27 28 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 23 27 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 20 28 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r41 20 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r42 18 27 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 18 19 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.115 $Y=2.72
+ $X2=2.255 $Y2=2.72
r44 17 31 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 17 19 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.395 $Y=2.72
+ $X2=2.255 $Y2=2.72
r46 13 16 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=3.425 $Y=1.66
+ $X2=3.425 $Y2=2.34
r47 11 34 3.22486 $w=2.2e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.425 $Y=2.635
+ $X2=3.497 $Y2=2.72
r48 11 16 15.4532 $w=2.18e-07 $l=2.95e-07 $layer=LI1_cond $X=3.425 $Y=2.635
+ $X2=3.425 $Y2=2.34
r49 7 19 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2.72
r50 7 9 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.255 $Y=2.635
+ $X2=2.255 $Y2=2
r51 2 16 400 $w=1.7e-07 $l=9.36149e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.4 $Y2=2.34
r52 2 13 400 $w=1.7e-07 $l=2.45713e-07 $layer=licon1_PDIFF $count=1 $X=3.23
+ $Y=1.485 $X2=3.4 $Y2=1.66
r53 1 9 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.055
+ $Y=1.485 $X2=2.265 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%X 1 2 10 13 14 15
r31 13 15 7.48143 $w=3.03e-07 $l=1.98e-07 $layer=LI1_cond $X=2.972 $Y=1.647
+ $X2=2.972 $Y2=1.845
r32 13 14 6.38002 $w=3.03e-07 $l=1.52e-07 $layer=LI1_cond $X=2.972 $Y=1.647
+ $X2=2.972 $Y2=1.495
r33 12 14 36.0445 $w=2.33e-07 $l=7.35e-07 $layer=LI1_cond $X=3.007 $Y=0.76
+ $X2=3.007 $Y2=1.495
r34 10 12 7.06015 $w=3.03e-07 $l=1.7e-07 $layer=LI1_cond $X=2.972 $Y=0.59
+ $X2=2.972 $Y2=0.76
r35 2 15 300 $w=1.7e-07 $l=4.91121e-07 $layer=licon1_PDIFF $count=2 $X=2.595
+ $Y=1.485 $X2=2.905 $Y2=1.845
r36 1 10 182 $w=1.7e-07 $l=5.00275e-07 $layer=licon1_NDIFF $count=1 $X=2.555
+ $Y=0.235 $X2=2.905 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR4_2%VGND 1 2 3 4 13 15 19 21 23 25 27 32 37 46
+ 50 57
c59 32 0 6.13246e-20 $X=1.985 $Y=0
c60 27 0 1.35736e-19 $X=1.045 $Y=0
r61 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r62 50 53 10.7204 $w=4.28e-07 $l=4e-07 $layer=LI1_cond $X=2.2 $Y=0 $X2=2.2
+ $Y2=0.4
r63 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r64 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r65 41 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r66 41 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.07
+ $Y2=0
r67 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r68 38 50 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.2
+ $Y2=0
r69 38 40 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=2.415 $Y=0 $X2=2.99
+ $Y2=0
r70 37 56 3.73837 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=3.497
+ $Y2=0
r71 37 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=3.315 $Y=0 $X2=2.99
+ $Y2=0
r72 36 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r73 36 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r74 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r75 33 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.235
+ $Y2=0
r76 33 35 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.425 $Y=0 $X2=1.61
+ $Y2=0
r77 32 50 6.22023 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=2.2
+ $Y2=0
r78 32 35 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.985 $Y=0 $X2=1.61
+ $Y2=0
r79 31 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r80 30 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r81 28 43 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r82 28 30 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r83 27 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=1.235
+ $Y2=0
r84 27 30 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.045 $Y=0 $X2=0.69
+ $Y2=0
r85 25 31 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r86 25 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r87 21 56 3.22486 $w=2.2e-07 $l=1.15521e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.497 $Y2=0
r88 21 23 16.5009 $w=2.18e-07 $l=3.15e-07 $layer=LI1_cond $X=3.425 $Y=0.085
+ $X2=3.425 $Y2=0.4
r89 17 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r90 17 19 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.4
r91 13 43 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.212 $Y2=0
r92 13 15 14.2765 $w=3.33e-07 $l=4.15e-07 $layer=LI1_cond $X=0.257 $Y=0.085
+ $X2=0.257 $Y2=0.5
r93 4 23 91 $w=1.7e-07 $l=2.31571e-07 $layer=licon1_NDIFF $count=2 $X=3.24
+ $Y=0.235 $X2=3.4 $Y2=0.4
r94 3 53 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.065
+ $Y=0.265 $X2=2.25 $Y2=0.4
r95 2 19 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.265 $X2=1.26 $Y2=0.4
r96 1 15 182 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.265 $X2=0.26 $Y2=0.5
.ends

