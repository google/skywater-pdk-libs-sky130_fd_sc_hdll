* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__isobufsrc_16 A SLEEP VGND VNB VPB VPWR X
X0 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR A a_151_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR A a_151_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 VGND A a_151_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_151_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VGND A a_151_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X40 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X41 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X42 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X43 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 a_151_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X46 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X47 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X49 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 a_151_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X52 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X53 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X54 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X55 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X56 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X58 a_585_297# SLEEP X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X59 a_151_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X60 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X61 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X62 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X63 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X64 X SLEEP a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 X a_151_297# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X66 a_585_297# a_151_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X67 VGND a_151_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X68 VGND SLEEP X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X69 X SLEEP VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X70 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X71 VPWR a_151_297# a_585_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
