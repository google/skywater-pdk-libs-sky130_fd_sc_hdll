* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
X0 a_601_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR A1 a_1369_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 Y B2 a_601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 Y B2 a_601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_601_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A2 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 a_1369_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_511_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 a_27_47# B2 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND A1 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 Y C1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_511_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND A2 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_511_47# B1 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 a_601_297# B2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_511_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND A1 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 VPWR B1 a_601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_601_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 a_511_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 Y A2 a_1369_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X25 a_27_47# C1 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 a_1369_297# A2 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_1369_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X28 a_511_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X29 a_27_47# B1 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 VPWR C1 Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X31 VPWR B1 a_601_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 Y A2 a_1369_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_511_47# B2 a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_511_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X35 a_1369_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_27_47# B1 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 a_27_47# B2 a_511_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X38 Y C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 VPWR A1 a_1369_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
