* NGSPICE file created from sky130_fd_sc_hdll__conb_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__conb_1 VGND VNB VPB VPWR HI LO
R0 VGND LO short w=480000u l=45000u
R1 HI VPWR short w=480000u l=45000u
.ends

