* File: sky130_fd_sc_hdll__muxb8to1_2.pex.spice
* Created: Wed Sep  2 08:36:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[0] 3 7 11 15 17 27 29
r47 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.16
+ $X2=0.965 $Y2=1.16
r48 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.75 $Y=1.16 $X2=0.94
+ $Y2=1.16
r49 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.75
+ $Y=1.16 $X2=0.75 $Y2=1.16
r50 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=0.52 $Y=1.16 $X2=0.75
+ $Y2=1.16
r51 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.16
+ $X2=0.52 $Y2=1.16
r52 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=0.41 $Y=1.19
+ $X2=0.75 $Y2=1.19
r53 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=0.41 $Y=1.16
+ $X2=0.495 $Y2=1.16
r54 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.41
+ $Y=1.16 $X2=0.41 $Y2=1.16
r55 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=0.23 $Y=1.19
+ $X2=0.41 $Y2=1.19
r56 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.16
r57 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.965 $Y=1.295
+ $X2=0.965 $Y2=1.985
r58 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.16
r59 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r60 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=1.16
r61 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.52 $Y=1.025
+ $X2=0.52 $Y2=0.56
r62 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.16
r63 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=0.495 $Y=1.295
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_278_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c77 9 0 1.30521e-19 $X=1.49 $Y=2.075
r78 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=2.43 $Y=1.42
+ $X2=2.715 $Y2=1.63
r79 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=2.265 $Y=1.34
+ $X2=1.96 $Y2=1.34
r80 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=2.265 $Y=1.42
+ $X2=2.43 $Y2=1.42
r81 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.265
+ $Y=1.34 $X2=2.265 $Y2=1.34
r82 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=2.715 $Y=2.31
+ $X2=2.715 $Y2=1.635
r83 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=2.43 $Y=1.205
+ $X2=2.43 $Y2=1.42
r84 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.8 $Y2=0.457
r85 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=2.43 $Y=0.755
+ $X2=2.43 $Y2=1.205
r86 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=1.96 $Y=1.475
+ $X2=1.96 $Y2=1.34
r87 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.96 $Y=1.475 $X2=1.96
+ $Y2=2.075
r88 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=1.87 $Y=1.4
+ $X2=1.96 $Y2=1.34
r89 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=1.4 $X2=1.58
+ $Y2=1.4
r90 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=1.49 $Y=1.475
+ $X2=1.58 $Y2=1.4
r91 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=1.49 $Y=1.475 $X2=1.49
+ $Y2=2.075
r92 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=1.63
r93 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=2.59
+ $Y=1.485 $X2=2.715 $Y2=2.31
r94 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=2.675
+ $Y=0.235 $X2=2.8 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[0] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=2.955 $Y=0.92
+ $X2=2.955 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=2.955 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.01 $Y=0.845
+ $X2=3.01 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.955 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.95 $Y=1.41
+ $X2=2.95 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.955 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=2.82 $Y=0.92
+ $X2=2.44 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.365 $Y=0.845
+ $X2=2.44 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=2.365 $Y=0.255
+ $X2=2.365 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.955 $Y=0.18
+ $X2=1.88 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=2.365 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=2.29 $Y=0.18
+ $X2=1.955 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.88 $Y=0.255
+ $X2=1.88 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.88 $Y=0.255 $X2=1.88
+ $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.88 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=1.805 $Y=0.18
+ $X2=1.535 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.46 $Y=0.255
+ $X2=1.535 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=1.46 $Y=0.255 $X2=1.46
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[1] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=3.485 $Y=0.92
+ $X2=3.485 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.485
+ $Y=1.16 $X2=3.485 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.98 $Y=0.255
+ $X2=4.98 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.635 $Y=0.18
+ $X2=4.56 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.98 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=4.905 $Y=0.18
+ $X2=4.635 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=4.56 $Y=0.255
+ $X2=4.56 $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.56 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=4.485 $Y=0.18
+ $X2=4.15 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.15 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=4.075 $Y=0.255
+ $X2=4.075 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=3.62 $Y=0.92
+ $X2=3.485 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4 $Y=0.92
+ $X2=4.075 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=4 $Y=0.92 $X2=3.62
+ $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.49 $Y=1.41
+ $X2=3.485 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.49 $Y=1.41 $X2=3.49
+ $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=3.43 $Y=0.845
+ $X2=3.485 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=3.43 $Y=0.845 $X2=3.43
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_701_47# 1 2 9 11 12 15 19 22 24 28
c74 15 0 1.69024e-19 $X=4.95 $Y=2.075
c75 11 0 1.93373e-19 $X=4.86 $Y=1.4
r76 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=4.175 $Y=1.34
+ $X2=4.48 $Y2=1.34
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.175
+ $Y=1.34 $X2=4.175 $Y2=1.34
r78 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=4.01 $Y=1.42
+ $X2=4.175 $Y2=1.42
r79 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=3.725 $Y=1.63
+ $X2=4.01 $Y2=1.42
r80 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=4.01 $Y=1.205
+ $X2=4.01 $Y2=1.42
r81 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=3.64 $Y2=0.457
r82 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=4.01 $Y=0.755
+ $X2=4.01 $Y2=1.205
r83 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=3.725 $Y=2.31
+ $X2=3.725 $Y2=1.635
r84 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.95 $Y=1.475 $X2=4.95
+ $Y2=2.075
r85 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=4.57 $Y=1.4
+ $X2=4.48 $Y2=1.34
r86 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=4.86 $Y=1.4
+ $X2=4.95 $Y2=1.475
r87 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=4.86 $Y=1.4 $X2=4.57
+ $Y2=1.4
r88 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=4.48 $Y=1.475
+ $X2=4.48 $Y2=1.34
r89 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=4.48 $Y=1.475 $X2=4.48
+ $Y2=2.075
r90 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=1.63
r91 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.58
+ $Y=1.485 $X2=3.725 $Y2=2.31
r92 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.505
+ $Y=0.235 $X2=3.64 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[1] 3 7 11 15 17 28
c53 17 0 1.17966e-19 $X=6.21 $Y=1.19
c54 15 0 1.17966e-19 $X=5.945 $Y=1.985
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.03
+ $Y=1.16 $X2=6.03 $Y2=1.16
r56 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=5.945 $Y=1.16
+ $X2=6.03 $Y2=1.16
r57 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.92 $Y=1.16
+ $X2=5.945 $Y2=1.16
r58 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=5.69 $Y=1.19
+ $X2=6.03 $Y2=1.19
r59 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=5.69 $Y=1.16 $X2=5.92
+ $Y2=1.16
r60 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.69
+ $Y=1.16 $X2=5.69 $Y2=1.16
r61 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=5.5 $Y=1.16 $X2=5.69
+ $Y2=1.16
r62 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.5 $Y2=1.16
r63 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.21 $Y=1.19
+ $X2=6.03 $Y2=1.19
r64 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.16
r65 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.945 $Y=1.295
+ $X2=5.945 $Y2=1.985
r66 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=1.16
r67 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.92 $Y=1.025
+ $X2=5.92 $Y2=0.56
r68 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=1.16
r69 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.5 $Y=1.025 $X2=5.5
+ $Y2=0.56
r70 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.16
r71 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=5.475 $Y=1.295
+ $X2=5.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[2] 3 7 11 15 17 27 29
c54 27 0 1.17966e-19 $X=7.19 $Y=1.16
c55 3 0 1.17966e-19 $X=6.935 $Y=1.985
r56 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=7.38 $Y=1.16
+ $X2=7.405 $Y2=1.16
r57 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=7.19 $Y=1.16 $X2=7.38
+ $Y2=1.16
r58 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.19
+ $Y=1.16 $X2=7.19 $Y2=1.16
r59 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=6.96 $Y=1.16 $X2=7.19
+ $Y2=1.16
r60 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=6.935 $Y=1.16
+ $X2=6.96 $Y2=1.16
r61 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=6.85 $Y=1.19
+ $X2=7.19 $Y2=1.19
r62 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=6.85 $Y=1.16
+ $X2=6.935 $Y2=1.16
r63 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.85
+ $Y=1.16 $X2=6.85 $Y2=1.16
r64 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=6.67 $Y=1.19
+ $X2=6.85 $Y2=1.19
r65 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.16
r66 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=7.405 $Y=1.295
+ $X2=7.405 $Y2=1.985
r67 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=1.16
r68 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.38 $Y=1.025
+ $X2=7.38 $Y2=0.56
r69 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=1.16
r70 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.96 $Y=1.025
+ $X2=6.96 $Y2=0.56
r71 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.16
r72 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=6.935 $Y=1.295
+ $X2=6.935 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1566_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c78 12 0 1.93373e-19 $X=8.02 $Y=1.4
c79 9 0 1.69024e-19 $X=7.93 $Y=2.075
r80 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=8.87 $Y=1.42
+ $X2=9.155 $Y2=1.63
r81 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=8.705 $Y=1.34
+ $X2=8.4 $Y2=1.34
r82 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=8.705 $Y=1.42
+ $X2=8.87 $Y2=1.42
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.705
+ $Y=1.34 $X2=8.705 $Y2=1.34
r84 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=9.155 $Y=2.31
+ $X2=9.155 $Y2=1.635
r85 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=8.87 $Y=1.205
+ $X2=8.87 $Y2=1.42
r86 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=9.24 $Y2=0.457
r87 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=8.87 $Y=0.755
+ $X2=8.87 $Y2=1.205
r88 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=8.4 $Y=1.475
+ $X2=8.4 $Y2=1.34
r89 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=8.4 $Y=1.475 $X2=8.4
+ $Y2=2.075
r90 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=8.31 $Y=1.4
+ $X2=8.4 $Y2=1.34
r91 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=8.31 $Y=1.4 $X2=8.02
+ $Y2=1.4
r92 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=7.93 $Y=1.475
+ $X2=8.02 $Y2=1.4
r93 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=7.93 $Y=1.475 $X2=7.93
+ $Y2=2.075
r94 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=1.63
r95 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=9.03
+ $Y=1.485 $X2=9.155 $Y2=2.31
r96 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=9.115
+ $Y=0.235 $X2=9.24 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[2] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.395 $Y=0.92
+ $X2=9.395 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.395
+ $Y=1.16 $X2=9.395 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.395 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.45 $Y=0.845
+ $X2=9.45 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.395 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.39 $Y=1.41
+ $X2=9.39 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=9.395 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=9.26 $Y=0.92
+ $X2=8.88 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.805 $Y=0.845
+ $X2=8.88 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=8.805 $Y=0.255
+ $X2=8.805 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.395 $Y=0.18
+ $X2=8.32 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.805 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=8.73 $Y=0.18
+ $X2=8.395 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.32 $Y=0.255
+ $X2=8.32 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=8.32 $Y=0.255 $X2=8.32
+ $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=8.32 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=8.245 $Y=0.18
+ $X2=7.975 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.9 $Y=0.255
+ $X2=7.975 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=7.9 $Y=0.255 $X2=7.9
+ $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[3] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=9.925 $Y=0.92
+ $X2=9.925 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.925
+ $Y=1.16 $X2=9.925 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11.42 $Y=0.255
+ $X2=11.42 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11.075 $Y=0.18
+ $X2=11 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.42 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=11.345 $Y=0.18
+ $X2=11.075 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=11 $Y=0.255 $X2=11
+ $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=11 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=10.925 $Y=0.18
+ $X2=10.59 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.59 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=10.515 $Y=0.255
+ $X2=10.515 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=10.06 $Y=0.92
+ $X2=9.925 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.515 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=10.44 $Y=0.92
+ $X2=10.06 $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=9.93 $Y=1.41
+ $X2=9.925 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.93 $Y=1.41 $X2=9.93
+ $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=9.87 $Y=0.845
+ $X2=9.925 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=9.87 $Y=0.845 $X2=9.87
+ $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1989_47# 1 2 9 11 12 15 19 22 24 28
c74 15 0 1.69024e-19 $X=11.39 $Y=2.075
c75 11 0 1.93373e-19 $X=11.3 $Y=1.4
r76 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=10.615 $Y=1.34
+ $X2=10.92 $Y2=1.34
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.615
+ $Y=1.34 $X2=10.615 $Y2=1.34
r78 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=10.45 $Y=1.42
+ $X2=10.615 $Y2=1.42
r79 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=10.165 $Y=1.63
+ $X2=10.45 $Y2=1.42
r80 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=10.45 $Y=1.205
+ $X2=10.45 $Y2=1.42
r81 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.08 $Y2=0.457
r82 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=10.45 $Y=0.755
+ $X2=10.45 $Y2=1.205
r83 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=10.165 $Y=2.31
+ $X2=10.165 $Y2=1.635
r84 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=11.39 $Y=1.475
+ $X2=11.39 $Y2=2.075
r85 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=11.01 $Y=1.4
+ $X2=10.92 $Y2=1.34
r86 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.39 $Y2=1.475
r87 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=11.3 $Y=1.4
+ $X2=11.01 $Y2=1.4
r88 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=10.92 $Y=1.475
+ $X2=10.92 $Y2=1.34
r89 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=10.92 $Y=1.475 $X2=10.92
+ $Y2=2.075
r90 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=1.63
r91 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.02
+ $Y=1.485 $X2=10.165 $Y2=2.31
r92 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.945
+ $Y=0.235 $X2=10.08 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[3] 3 7 11 15 17 28
c53 17 0 1.17966e-19 $X=12.65 $Y=1.19
c54 15 0 1.17966e-19 $X=12.385 $Y=1.985
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.47
+ $Y=1.16 $X2=12.47 $Y2=1.16
r56 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=12.385 $Y=1.16
+ $X2=12.47 $Y2=1.16
r57 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=12.36 $Y=1.16
+ $X2=12.385 $Y2=1.16
r58 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=12.13 $Y=1.19
+ $X2=12.47 $Y2=1.19
r59 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=12.13 $Y=1.16 $X2=12.36
+ $Y2=1.16
r60 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=12.13
+ $Y=1.16 $X2=12.13 $Y2=1.16
r61 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=11.94 $Y=1.16
+ $X2=12.13 $Y2=1.16
r62 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=11.915 $Y=1.16
+ $X2=11.94 $Y2=1.16
r63 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=12.65 $Y=1.19
+ $X2=12.47 $Y2=1.19
r64 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.16
r65 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=12.385 $Y=1.295
+ $X2=12.385 $Y2=1.985
r66 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=1.16
r67 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=12.36 $Y=1.025
+ $X2=12.36 $Y2=0.56
r68 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=1.16
r69 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=11.94 $Y=1.025
+ $X2=11.94 $Y2=0.56
r70 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.16
r71 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=11.915 $Y=1.295
+ $X2=11.915 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[4] 3 7 11 15 17 27 29
c54 27 0 1.17966e-19 $X=13.63 $Y=1.16
c55 3 0 1.17966e-19 $X=13.375 $Y=1.985
r56 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.82 $Y=1.16
+ $X2=13.845 $Y2=1.16
r57 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=13.63 $Y=1.16
+ $X2=13.82 $Y2=1.16
r58 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.63
+ $Y=1.16 $X2=13.63 $Y2=1.16
r59 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=13.4 $Y=1.16 $X2=13.63
+ $Y2=1.16
r60 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=13.375 $Y=1.16
+ $X2=13.4 $Y2=1.16
r61 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=13.29 $Y=1.19
+ $X2=13.63 $Y2=1.19
r62 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=13.29 $Y=1.16
+ $X2=13.375 $Y2=1.16
r63 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.29
+ $Y=1.16 $X2=13.29 $Y2=1.16
r64 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=13.11 $Y=1.19
+ $X2=13.29 $Y2=1.19
r65 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.16
r66 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.845 $Y=1.295
+ $X2=13.845 $Y2=1.985
r67 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=1.16
r68 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.82 $Y=1.025
+ $X2=13.82 $Y2=0.56
r69 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=1.16
r70 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=13.4 $Y=1.025
+ $X2=13.4 $Y2=0.56
r71 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.16
r72 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=13.375 $Y=1.295
+ $X2=13.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2854_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c78 12 0 1.93373e-19 $X=14.46 $Y=1.4
c79 9 0 1.69024e-19 $X=14.37 $Y=2.075
r80 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=15.31 $Y=1.42
+ $X2=15.595 $Y2=1.63
r81 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=15.145 $Y=1.34
+ $X2=14.84 $Y2=1.34
r82 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=15.145 $Y=1.42
+ $X2=15.31 $Y2=1.42
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.145
+ $Y=1.34 $X2=15.145 $Y2=1.34
r84 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=15.595 $Y=2.31
+ $X2=15.595 $Y2=1.635
r85 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=15.31 $Y=1.205
+ $X2=15.31 $Y2=1.42
r86 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=15.31 $Y=0.755
+ $X2=15.68 $Y2=0.457
r87 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=15.31 $Y=0.755
+ $X2=15.31 $Y2=1.205
r88 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=14.84 $Y=1.475
+ $X2=14.84 $Y2=1.34
r89 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.84 $Y=1.475
+ $X2=14.84 $Y2=2.075
r90 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=14.75 $Y=1.4
+ $X2=14.84 $Y2=1.34
r91 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=14.75 $Y=1.4
+ $X2=14.46 $Y2=1.4
r92 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=14.37 $Y=1.475
+ $X2=14.46 $Y2=1.4
r93 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=14.37 $Y=1.475 $X2=14.37
+ $Y2=2.075
r94 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=1.485 $X2=15.595 $Y2=1.63
r95 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=15.47
+ $Y=1.485 $X2=15.595 $Y2=2.31
r96 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=15.555
+ $Y=0.235 $X2=15.68 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[4] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=15.835 $Y=0.92
+ $X2=15.835 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=15.835
+ $Y=1.16 $X2=15.835 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=15.89 $Y=0.845
+ $X2=15.835 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=15.89 $Y=0.845
+ $X2=15.89 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=15.83 $Y=1.41
+ $X2=15.835 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=15.83 $Y=1.41
+ $X2=15.83 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=15.7 $Y=0.92
+ $X2=15.835 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=15.7 $Y=0.92
+ $X2=15.32 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.245 $Y=0.845
+ $X2=15.32 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=15.245 $Y=0.255
+ $X2=15.245 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.835 $Y=0.18
+ $X2=14.76 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=15.17 $Y=0.18
+ $X2=15.245 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=15.17 $Y=0.18
+ $X2=14.835 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.76 $Y=0.255
+ $X2=14.76 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.76 $Y=0.255
+ $X2=14.76 $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=14.685 $Y=0.18
+ $X2=14.76 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=14.685 $Y=0.18
+ $X2=14.415 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=14.34 $Y=0.255
+ $X2=14.415 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=14.34 $Y=0.255
+ $X2=14.34 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[5] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=16.365 $Y=0.92
+ $X2=16.365 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=16.365
+ $Y=1.16 $X2=16.365 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.86 $Y=0.255
+ $X2=17.86 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.515 $Y=0.18
+ $X2=17.44 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=17.785 $Y=0.18
+ $X2=17.86 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=17.785 $Y=0.18
+ $X2=17.515 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.44 $Y=0.255
+ $X2=17.44 $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=17.44 $Y=0.255
+ $X2=17.44 $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=17.365 $Y=0.18
+ $X2=17.44 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=17.365 $Y=0.18
+ $X2=17.03 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.955 $Y=0.255
+ $X2=17.03 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=16.955 $Y=0.255
+ $X2=16.955 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=16.5 $Y=0.92
+ $X2=16.365 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=16.88 $Y=0.92
+ $X2=16.955 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=16.88 $Y=0.92 $X2=16.5
+ $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=16.37 $Y=1.41
+ $X2=16.365 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=16.37 $Y=1.41
+ $X2=16.37 $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=16.31 $Y=0.845
+ $X2=16.365 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=16.31 $Y=0.845
+ $X2=16.31 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3277_47# 1 2 9 11 12 15 19 22 24 28
c74 15 0 1.69024e-19 $X=17.83 $Y=2.075
c75 11 0 1.93373e-19 $X=17.74 $Y=1.4
r76 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=17.055 $Y=1.34
+ $X2=17.36 $Y2=1.34
r77 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=17.055
+ $Y=1.34 $X2=17.055 $Y2=1.34
r78 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=16.89 $Y=1.42
+ $X2=17.055 $Y2=1.42
r79 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=16.605 $Y=1.63
+ $X2=16.89 $Y2=1.42
r80 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=16.89 $Y=1.205
+ $X2=16.89 $Y2=1.42
r81 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=16.89 $Y=0.755
+ $X2=16.52 $Y2=0.457
r82 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=16.89 $Y=0.755
+ $X2=16.89 $Y2=1.205
r83 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=16.605 $Y=2.31
+ $X2=16.605 $Y2=1.635
r84 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.83 $Y=1.475
+ $X2=17.83 $Y2=2.075
r85 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=17.45 $Y=1.4
+ $X2=17.36 $Y2=1.34
r86 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=17.74 $Y=1.4
+ $X2=17.83 $Y2=1.475
r87 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=17.74 $Y=1.4
+ $X2=17.45 $Y2=1.4
r88 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=17.36 $Y=1.475
+ $X2=17.36 $Y2=1.34
r89 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=17.36 $Y=1.475 $X2=17.36
+ $Y2=2.075
r90 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=1.485 $X2=16.605 $Y2=1.63
r91 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=16.46
+ $Y=1.485 $X2=16.605 $Y2=2.31
r92 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=16.385
+ $Y=0.235 $X2=16.52 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[5] 3 7 11 15 17 28
c53 17 0 1.17966e-19 $X=19.09 $Y=1.19
c54 15 0 1.17966e-19 $X=18.825 $Y=1.985
r55 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.91
+ $Y=1.16 $X2=18.91 $Y2=1.16
r56 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=18.825 $Y=1.16
+ $X2=18.91 $Y2=1.16
r57 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.8 $Y=1.16
+ $X2=18.825 $Y2=1.16
r58 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=18.57 $Y=1.19
+ $X2=18.91 $Y2=1.19
r59 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=18.57 $Y=1.16 $X2=18.8
+ $Y2=1.16
r60 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=18.57
+ $Y=1.16 $X2=18.57 $Y2=1.16
r61 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=18.38 $Y=1.16
+ $X2=18.57 $Y2=1.16
r62 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=18.355 $Y=1.16
+ $X2=18.38 $Y2=1.16
r63 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.09 $Y=1.19
+ $X2=18.91 $Y2=1.19
r64 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.825 $Y=1.295
+ $X2=18.825 $Y2=1.16
r65 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.825 $Y=1.295
+ $X2=18.825 $Y2=1.985
r66 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.8 $Y=1.025
+ $X2=18.8 $Y2=1.16
r67 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.8 $Y=1.025
+ $X2=18.8 $Y2=0.56
r68 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=18.38 $Y=1.025
+ $X2=18.38 $Y2=1.16
r69 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=18.38 $Y=1.025
+ $X2=18.38 $Y2=0.56
r70 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=18.355 $Y=1.295
+ $X2=18.355 $Y2=1.16
r71 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=18.355 $Y=1.295
+ $X2=18.355 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[6] 3 7 11 15 17 27 29
c54 27 0 1.17966e-19 $X=20.07 $Y=1.16
c55 3 0 1.17966e-19 $X=19.815 $Y=1.985
r56 28 29 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=20.26 $Y=1.16
+ $X2=20.285 $Y2=1.16
r57 26 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=20.07 $Y=1.16
+ $X2=20.26 $Y2=1.16
r58 26 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=20.07
+ $Y=1.16 $X2=20.07 $Y2=1.16
r59 24 26 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=19.84 $Y=1.16 $X2=20.07
+ $Y2=1.16
r60 23 24 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=19.815 $Y=1.16
+ $X2=19.84 $Y2=1.16
r61 21 27 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=19.73 $Y=1.19
+ $X2=20.07 $Y2=1.19
r62 20 23 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=19.73 $Y=1.16
+ $X2=19.815 $Y2=1.16
r63 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=19.73
+ $Y=1.16 $X2=19.73 $Y2=1.16
r64 17 21 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=19.55 $Y=1.19
+ $X2=19.73 $Y2=1.19
r65 13 29 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=20.285 $Y=1.295
+ $X2=20.285 $Y2=1.16
r66 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=20.285 $Y=1.295
+ $X2=20.285 $Y2=1.985
r67 9 28 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=20.26 $Y=1.025
+ $X2=20.26 $Y2=1.16
r68 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=20.26 $Y=1.025
+ $X2=20.26 $Y2=0.56
r69 5 24 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=19.84 $Y=1.025
+ $X2=19.84 $Y2=1.16
r70 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=19.84 $Y=1.025
+ $X2=19.84 $Y2=0.56
r71 1 23 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=19.815 $Y=1.295
+ $X2=19.815 $Y2=1.16
r72 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=19.815 $Y=1.295
+ $X2=19.815 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4142_265# 1 2 9 11 12 15 17 18 21 28
+ 32
c78 12 0 1.93373e-19 $X=20.9 $Y=1.4
c79 9 0 1.69024e-19 $X=20.81 $Y=2.075
r80 26 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=21.75 $Y=1.42
+ $X2=22.035 $Y2=1.63
r81 25 32 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=21.585 $Y=1.34
+ $X2=21.28 $Y2=1.34
r82 24 26 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=21.585 $Y=1.42
+ $X2=21.75 $Y2=1.42
r83 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=21.585
+ $Y=1.34 $X2=21.585 $Y2=1.34
r84 21 28 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=22.035 $Y=2.31
+ $X2=22.035 $Y2=1.635
r85 18 26 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=21.75 $Y=1.205
+ $X2=21.75 $Y2=1.42
r86 17 31 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=21.75 $Y=0.755
+ $X2=22.12 $Y2=0.457
r87 17 18 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=21.75 $Y=0.755
+ $X2=21.75 $Y2=1.205
r88 13 32 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=21.28 $Y=1.475
+ $X2=21.28 $Y2=1.34
r89 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=21.28 $Y=1.475
+ $X2=21.28 $Y2=2.075
r90 11 32 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=21.19 $Y=1.4
+ $X2=21.28 $Y2=1.34
r91 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=21.19 $Y=1.4
+ $X2=20.9 $Y2=1.4
r92 7 12 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=20.81 $Y=1.475
+ $X2=20.9 $Y2=1.4
r93 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=20.81 $Y=1.475 $X2=20.81
+ $Y2=2.075
r94 2 28 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=1.485 $X2=22.035 $Y2=1.63
r95 2 21 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=21.91
+ $Y=1.485 $X2=22.035 $Y2=2.31
r96 1 31 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=21.995
+ $Y=0.235 $X2=22.12 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[6] 1 3 4 5 6 8 9 12 13 14 15 17 18 20
+ 21 22
r65 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.275 $Y=0.92
+ $X2=22.275 $Y2=1.16
r66 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.275
+ $Y=1.16 $X2=22.275 $Y2=1.16
r67 18 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.33 $Y=0.845
+ $X2=22.275 $Y2=0.92
r68 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.33 $Y=0.845
+ $X2=22.33 $Y2=0.495
r69 15 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.27 $Y=1.41
+ $X2=22.275 $Y2=1.16
r70 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.27 $Y=1.41
+ $X2=22.27 $Y2=1.985
r71 13 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.14 $Y=0.92
+ $X2=22.275 $Y2=0.92
r72 13 14 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=22.14 $Y=0.92
+ $X2=21.76 $Y2=0.92
r73 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.685 $Y=0.845
+ $X2=21.76 $Y2=0.92
r74 11 12 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=21.685 $Y=0.255
+ $X2=21.685 $Y2=0.845
r75 10 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.275 $Y=0.18
+ $X2=21.2 $Y2=0.18
r76 9 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=21.61 $Y=0.18
+ $X2=21.685 $Y2=0.255
r77 9 10 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=21.61 $Y=0.18
+ $X2=21.275 $Y2=0.18
r78 6 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.2 $Y=0.255
+ $X2=21.2 $Y2=0.18
r79 6 8 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=21.2 $Y=0.255 $X2=21.2
+ $Y2=0.605
r80 4 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=21.125 $Y=0.18
+ $X2=21.2 $Y2=0.18
r81 4 5 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=21.125 $Y=0.18
+ $X2=20.855 $Y2=0.18
r82 1 5 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=20.78 $Y=0.255
+ $X2=20.855 $Y2=0.18
r83 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=20.78 $Y=0.255
+ $X2=20.78 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%S[7] 1 3 4 6 7 10 11 12 13 15 16 18 20
+ 21 22
r62 24 26 44.8372 $w=2.58e-07 $l=2.4e-07 $layer=POLY_cond $X=22.805 $Y=0.92
+ $X2=22.805 $Y2=1.16
r63 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=22.805
+ $Y=1.16 $X2=22.805 $Y2=1.16
r64 18 20 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=24.3 $Y=0.255
+ $X2=24.3 $Y2=0.605
r65 17 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.955 $Y=0.18
+ $X2=23.88 $Y2=0.18
r66 16 18 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=24.225 $Y=0.18
+ $X2=24.3 $Y2=0.255
r67 16 17 138.447 $w=1.5e-07 $l=2.7e-07 $layer=POLY_cond $X=24.225 $Y=0.18
+ $X2=23.955 $Y2=0.18
r68 13 21 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.88 $Y=0.255
+ $X2=23.88 $Y2=0.18
r69 13 15 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=23.88 $Y=0.255
+ $X2=23.88 $Y2=0.605
r70 11 21 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=23.805 $Y=0.18
+ $X2=23.88 $Y2=0.18
r71 11 12 171.777 $w=1.5e-07 $l=3.35e-07 $layer=POLY_cond $X=23.805 $Y=0.18
+ $X2=23.47 $Y2=0.18
r72 9 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.395 $Y=0.255
+ $X2=23.47 $Y2=0.18
r73 9 10 302.532 $w=1.5e-07 $l=5.9e-07 $layer=POLY_cond $X=23.395 $Y=0.255
+ $X2=23.395 $Y2=0.845
r74 8 24 15.449 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=22.94 $Y=0.92
+ $X2=22.805 $Y2=0.92
r75 7 10 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=23.32 $Y=0.92
+ $X2=23.395 $Y2=0.845
r76 7 8 194.851 $w=1.5e-07 $l=3.8e-07 $layer=POLY_cond $X=23.32 $Y=0.92
+ $X2=22.94 $Y2=0.92
r77 4 26 51.1626 $w=2.58e-07 $l=2.52488e-07 $layer=POLY_cond $X=22.81 $Y=1.41
+ $X2=22.805 $Y2=1.16
r78 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=22.81 $Y=1.41
+ $X2=22.81 $Y2=1.985
r79 1 24 22.3869 $w=2.58e-07 $l=9.87421e-08 $layer=POLY_cond $X=22.75 $Y=0.845
+ $X2=22.805 $Y2=0.92
r80 1 3 112.467 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=22.75 $Y=0.845
+ $X2=22.75 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4565_47# 1 2 9 11 12 15 19 22 24 28
c73 15 0 1.30521e-19 $X=24.27 $Y=2.075
r74 31 33 66.8227 $w=2.2e-07 $l=3.05e-07 $layer=POLY_cond $X=23.495 $Y=1.34
+ $X2=23.8 $Y2=1.34
r75 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=23.495
+ $Y=1.34 $X2=23.495 $Y2=1.34
r76 28 30 7.80233 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=23.33 $Y=1.42
+ $X2=23.495 $Y2=1.42
r77 27 28 13.4767 $w=2.58e-07 $l=3.756e-07 $layer=LI1_cond $X=23.045 $Y=1.63
+ $X2=23.33 $Y2=1.42
r78 22 28 3.17874 $w=1.7e-07 $l=2.15e-07 $layer=LI1_cond $X=23.33 $Y=1.205
+ $X2=23.33 $Y2=1.42
r79 21 24 16.1792 $w=2.79e-07 $l=4.97152e-07 $layer=LI1_cond $X=23.33 $Y=0.755
+ $X2=22.96 $Y2=0.457
r80 21 22 29.3583 $w=1.68e-07 $l=4.5e-07 $layer=LI1_cond $X=23.33 $Y=0.755
+ $X2=23.33 $Y2=1.205
r81 19 27 23.5727 $w=3.28e-07 $l=6.75e-07 $layer=LI1_cond $X=23.045 $Y=2.31
+ $X2=23.045 $Y2=1.635
r82 13 15 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=24.27 $Y=1.475
+ $X2=24.27 $Y2=2.075
r83 12 33 24.6297 $w=2.2e-07 $l=1.16189e-07 $layer=POLY_cond $X=23.89 $Y=1.4
+ $X2=23.8 $Y2=1.34
r84 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=24.18 $Y=1.4
+ $X2=24.27 $Y2=1.475
r85 11 12 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=24.18 $Y=1.4
+ $X2=23.89 $Y2=1.4
r86 7 33 7.56431 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=23.8 $Y=1.475
+ $X2=23.8 $Y2=1.34
r87 7 9 233.226 $w=1.8e-07 $l=6e-07 $layer=POLY_cond $X=23.8 $Y=1.475 $X2=23.8
+ $Y2=2.075
r88 2 27 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=1.485 $X2=23.045 $Y2=1.63
r89 2 19 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=22.9
+ $Y=1.485 $X2=23.045 $Y2=2.31
r90 1 24 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.825
+ $Y=0.235 $X2=22.96 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%D[7] 3 7 11 15 17 28
r46 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.35
+ $Y=1.16 $X2=25.35 $Y2=1.16
r47 26 28 18.8848 $w=2.7e-07 $l=8.5e-08 $layer=POLY_cond $X=25.265 $Y=1.16
+ $X2=25.35 $Y2=1.16
r48 25 26 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=25.24 $Y=1.16
+ $X2=25.265 $Y2=1.16
r49 24 29 14.5122 $w=2.68e-07 $l=3.4e-07 $layer=LI1_cond $X=25.01 $Y=1.19
+ $X2=25.35 $Y2=1.19
r50 23 25 51.1 $w=2.7e-07 $l=2.3e-07 $layer=POLY_cond $X=25.01 $Y=1.16 $X2=25.24
+ $Y2=1.16
r51 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=25.01
+ $Y=1.16 $X2=25.01 $Y2=1.16
r52 21 23 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=24.82 $Y=1.16
+ $X2=25.01 $Y2=1.16
r53 19 21 5.55434 $w=2.7e-07 $l=2.5e-08 $layer=POLY_cond $X=24.795 $Y=1.16
+ $X2=24.82 $Y2=1.16
r54 17 29 7.68295 $w=2.68e-07 $l=1.8e-07 $layer=LI1_cond $X=25.53 $Y=1.19
+ $X2=25.35 $Y2=1.19
r55 13 26 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.16
r56 13 15 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=25.265 $Y=1.295
+ $X2=25.265 $Y2=1.985
r57 9 25 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=1.16
r58 9 11 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=25.24 $Y=1.025
+ $X2=25.24 $Y2=0.56
r59 5 21 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=1.16
r60 5 7 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=24.82 $Y=1.025
+ $X2=24.82 $Y2=0.56
r61 1 19 12.2893 $w=1.8e-07 $l=1.35e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.16
r62 1 3 268.21 $w=1.8e-07 $l=6.9e-07 $layer=POLY_cond $X=24.795 $Y=1.295
+ $X2=24.795 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_297# 1 2 3 10 12 17 18 19 22 27 28
r47 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=0.26 $Y=2.34
+ $X2=0.26 $Y2=2.21
r48 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=2.195 $Y=2.295
+ $X2=2.195 $Y2=1.81
r49 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.11 $Y=2.38
+ $X2=2.195 $Y2=2.295
r50 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=2.11 $Y=2.38
+ $X2=1.285 $Y2=2.38
r51 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.285 $Y2=2.38
r52 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=1.78
r53 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=1.2 $Y=1.665
+ $X2=1.2 $Y2=1.78
r54 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.395 $Y=1.58
+ $X2=0.245 $Y2=1.58
r55 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=1.2 $Y2=1.665
r56 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=1.115 $Y=1.58
+ $X2=0.395 $Y2=1.58
r57 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=1.58
r58 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=0.245 $Y=1.665
+ $X2=0.245 $Y2=2.21
r59 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.665 $X2=2.195 $Y2=1.81
r60 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.78
r61 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r62 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 40 43
+ 50 54 57 64 68 71 78 82 85 92 94 98 99 101 105 109 110 112 116 120 121 123 127
+ 131 132 134 137 138 139 140 141 142 143 144 153 165 172 184 191 203 210 222
+ 231 235 238 241 244 247 250 253 256
c368 134 0 1.30521e-19 $X=25.03 $Y=1.94
c369 127 0 1.69024e-19 $X=20.05 $Y=1.94
c370 123 0 1.69024e-19 $X=18.59 $Y=1.94
c371 116 0 1.69024e-19 $X=13.61 $Y=1.94
c372 112 0 1.69024e-19 $X=12.15 $Y=1.94
c373 105 0 1.69024e-19 $X=7.17 $Y=1.94
c374 101 0 1.69024e-19 $X=5.71 $Y=1.94
c375 94 0 1.30521e-19 $X=0.73 $Y=1.94
r376 256 257 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.07 $Y=2.72
+ $X2=25.07 $Y2=2.72
r377 253 254 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.01 $Y=2.72
+ $X2=20.01 $Y2=2.72
r378 250 251 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=18.63 $Y=2.72
+ $X2=18.63 $Y2=2.72
r379 247 248 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r380 244 245 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=12.19 $Y=2.72
+ $X2=12.19 $Y2=2.72
r381 241 242 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r382 238 239 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r383 235 236 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r384 229 256 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=25.165 $Y=2.72
+ $X2=25.015 $Y2=2.72
r385 229 231 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=25.165 $Y=2.72
+ $X2=25.53 $Y2=2.72
r386 228 257 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=24.61 $Y=2.72
+ $X2=25.07 $Y2=2.72
r387 227 228 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=24.61 $Y=2.72
+ $X2=24.61 $Y2=2.72
r388 225 228 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=22.77 $Y=2.72
+ $X2=24.61 $Y2=2.72
r389 224 227 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=22.77 $Y=2.72
+ $X2=24.61 $Y2=2.72
r390 224 225 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.77 $Y=2.72
+ $X2=22.77 $Y2=2.72
r391 222 256 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=24.865 $Y=2.72
+ $X2=25.015 $Y2=2.72
r392 222 227 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=24.865 $Y=2.72
+ $X2=24.61 $Y2=2.72
r393 221 225 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=22.31 $Y=2.72
+ $X2=22.77 $Y2=2.72
r394 220 221 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.31 $Y=2.72
+ $X2=22.31 $Y2=2.72
r395 218 221 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=22.31 $Y2=2.72
r396 218 254 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=2.72
+ $X2=20.01 $Y2=2.72
r397 217 220 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=20.47 $Y=2.72
+ $X2=22.31 $Y2=2.72
r398 217 218 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=20.47 $Y=2.72
+ $X2=20.47 $Y2=2.72
r399 215 253 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=20.215 $Y=2.72
+ $X2=20.065 $Y2=2.72
r400 215 217 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=20.215 $Y=2.72
+ $X2=20.47 $Y2=2.72
r401 211 250 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.725 $Y=2.72
+ $X2=18.575 $Y2=2.72
r402 211 213 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=18.725 $Y=2.72
+ $X2=19.55 $Y2=2.72
r403 210 253 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.915 $Y=2.72
+ $X2=20.065 $Y2=2.72
r404 210 213 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=19.915 $Y=2.72
+ $X2=19.55 $Y2=2.72
r405 209 251 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=2.72
+ $X2=18.63 $Y2=2.72
r406 208 209 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18.17 $Y=2.72
+ $X2=18.17 $Y2=2.72
r407 206 209 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=16.33 $Y=2.72
+ $X2=18.17 $Y2=2.72
r408 205 208 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=16.33 $Y=2.72
+ $X2=18.17 $Y2=2.72
r409 205 206 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.33 $Y=2.72
+ $X2=16.33 $Y2=2.72
r410 203 250 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.425 $Y=2.72
+ $X2=18.575 $Y2=2.72
r411 203 208 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=18.425 $Y=2.72
+ $X2=18.17 $Y2=2.72
r412 202 206 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=2.72
+ $X2=16.33 $Y2=2.72
r413 201 202 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.87 $Y=2.72
+ $X2=15.87 $Y2=2.72
r414 199 202 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=15.87 $Y2=2.72
r415 199 248 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=2.72
+ $X2=13.57 $Y2=2.72
r416 198 201 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=14.03 $Y=2.72
+ $X2=15.87 $Y2=2.72
r417 198 199 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=14.03 $Y=2.72
+ $X2=14.03 $Y2=2.72
r418 196 247 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.775 $Y=2.72
+ $X2=13.625 $Y2=2.72
r419 196 198 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=13.775 $Y=2.72
+ $X2=14.03 $Y2=2.72
r420 192 244 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=12.135 $Y2=2.72
r421 192 194 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=12.285 $Y=2.72
+ $X2=13.11 $Y2=2.72
r422 191 247 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.475 $Y=2.72
+ $X2=13.625 $Y2=2.72
r423 191 194 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=13.475 $Y=2.72
+ $X2=13.11 $Y2=2.72
r424 190 245 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.19 $Y2=2.72
r425 189 190 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r426 187 190 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=11.73 $Y2=2.72
r427 186 189 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=2.72
+ $X2=11.73 $Y2=2.72
r428 186 187 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r429 184 244 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=12.135 $Y2=2.72
r430 184 189 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=11.985 $Y=2.72
+ $X2=11.73 $Y2=2.72
r431 183 187 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r432 182 183 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r433 180 183 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r434 180 242 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=7.13 $Y2=2.72
r435 179 182 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=2.72
+ $X2=9.43 $Y2=2.72
r436 179 180 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r437 177 241 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.185 $Y2=2.72
r438 177 179 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.335 $Y=2.72
+ $X2=7.59 $Y2=2.72
r439 173 238 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=5.695 $Y2=2.72
r440 173 175 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.845 $Y=2.72
+ $X2=6.67 $Y2=2.72
r441 172 241 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=7.185 $Y2=2.72
r442 172 175 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=7.035 $Y=2.72
+ $X2=6.67 $Y2=2.72
r443 171 239 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r444 170 171 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r445 168 171 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=5.29 $Y2=2.72
r446 167 170 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=5.29 $Y2=2.72
r447 167 168 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r448 165 238 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.695 $Y2=2.72
r449 165 170 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.545 $Y=2.72
+ $X2=5.29 $Y2=2.72
r450 164 168 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r451 163 164 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r452 161 164 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r453 161 236 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r454 160 163 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r455 160 161 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r456 158 235 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.745 $Y2=2.72
r457 158 160 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r458 153 235 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.745 $Y2=2.72
r459 153 155 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=0.595 $Y=2.72
+ $X2=0.23 $Y2=2.72
r460 144 257 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=25.53 $Y=2.72
+ $X2=25.07 $Y2=2.72
r461 144 231 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=25.53 $Y=2.72
+ $X2=25.53 $Y2=2.72
r462 143 254 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.55 $Y=2.72
+ $X2=20.01 $Y2=2.72
r463 143 213 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=19.55 $Y=2.72
+ $X2=19.55 $Y2=2.72
r464 142 143 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=2.72
+ $X2=19.55 $Y2=2.72
r465 142 251 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=2.72
+ $X2=18.63 $Y2=2.72
r466 141 248 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=2.72
+ $X2=13.57 $Y2=2.72
r467 141 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.11 $Y=2.72
+ $X2=13.11 $Y2=2.72
r468 140 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=13.11 $Y2=2.72
r469 140 245 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=2.72
+ $X2=12.19 $Y2=2.72
r470 139 242 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.13 $Y2=2.72
r471 139 175 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r472 138 139 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r473 138 239 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r474 137 236 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r475 137 155 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r476 134 136 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=25.03 $Y=1.94
+ $X2=25.03 $Y2=2.105
r477 131 220 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=22.375 $Y=2.72
+ $X2=22.31 $Y2=2.72
r478 131 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.375 $Y=2.72
+ $X2=22.54 $Y2=2.72
r479 130 224 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=22.705 $Y=2.72
+ $X2=22.77 $Y2=2.72
r480 130 132 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=22.705 $Y=2.72
+ $X2=22.54 $Y2=2.72
r481 127 129 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=20.05 $Y=1.94
+ $X2=20.05 $Y2=2.105
r482 123 125 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=18.59 $Y=1.94
+ $X2=18.59 $Y2=2.105
r483 120 201 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=15.935 $Y=2.72
+ $X2=15.87 $Y2=2.72
r484 120 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=15.935 $Y=2.72
+ $X2=16.1 $Y2=2.72
r485 119 205 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=16.265 $Y=2.72
+ $X2=16.33 $Y2=2.72
r486 119 121 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=16.265 $Y=2.72
+ $X2=16.1 $Y2=2.72
r487 116 118 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.61 $Y=1.94
+ $X2=13.61 $Y2=2.105
r488 112 114 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=12.15 $Y=1.94
+ $X2=12.15 $Y2=2.105
r489 109 182 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.43 $Y2=2.72
r490 109 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.495 $Y=2.72
+ $X2=9.66 $Y2=2.72
r491 108 186 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.89 $Y2=2.72
r492 108 110 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.825 $Y=2.72
+ $X2=9.66 $Y2=2.72
r493 105 107 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=7.17 $Y=1.94
+ $X2=7.17 $Y2=2.105
r494 101 103 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=5.71 $Y=1.94
+ $X2=5.71 $Y2=2.105
r495 98 163 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=2.99 $Y2=2.72
r496 98 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.055 $Y=2.72
+ $X2=3.22 $Y2=2.72
r497 97 167 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.45 $Y2=2.72
r498 97 99 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.385 $Y=2.72
+ $X2=3.22 $Y2=2.72
r499 94 96 5.8804 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=1.94
+ $X2=0.73 $Y2=2.105
r500 92 136 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=25.015 $Y=2.34
+ $X2=25.015 $Y2=2.105
r501 90 256 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.015 $Y=2.635
+ $X2=25.015 $Y2=2.72
r502 90 92 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=25.015 $Y=2.635
+ $X2=25.015 $Y2=2.34
r503 85 88 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=22.54 $Y=1.63
+ $X2=22.54 $Y2=2.31
r504 83 132 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=2.635
+ $X2=22.54 $Y2=2.72
r505 83 88 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=22.54 $Y=2.635
+ $X2=22.54 $Y2=2.31
r506 82 129 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=20.065 $Y=2.34
+ $X2=20.065 $Y2=2.105
r507 80 253 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=20.065 $Y=2.635
+ $X2=20.065 $Y2=2.72
r508 80 82 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=20.065 $Y=2.635
+ $X2=20.065 $Y2=2.34
r509 78 125 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=18.575 $Y=2.34
+ $X2=18.575 $Y2=2.105
r510 76 250 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=18.575 $Y=2.635
+ $X2=18.575 $Y2=2.72
r511 76 78 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=18.575 $Y=2.635
+ $X2=18.575 $Y2=2.34
r512 71 74 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=16.1 $Y=1.63
+ $X2=16.1 $Y2=2.31
r513 69 121 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=2.635
+ $X2=16.1 $Y2=2.72
r514 69 74 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=16.1 $Y=2.635
+ $X2=16.1 $Y2=2.31
r515 68 118 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=13.625 $Y=2.34
+ $X2=13.625 $Y2=2.105
r516 66 247 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.625 $Y=2.635
+ $X2=13.625 $Y2=2.72
r517 66 68 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=13.625 $Y=2.635
+ $X2=13.625 $Y2=2.34
r518 64 114 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=12.135 $Y=2.34
+ $X2=12.135 $Y2=2.105
r519 62 244 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.72
r520 62 64 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=12.135 $Y=2.635
+ $X2=12.135 $Y2=2.34
r521 57 60 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=9.66 $Y=1.63
+ $X2=9.66 $Y2=2.31
r522 55 110 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r523 55 60 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.31
r524 54 107 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=7.185 $Y=2.34
+ $X2=7.185 $Y2=2.105
r525 52 241 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.72
r526 52 54 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=7.185 $Y=2.635
+ $X2=7.185 $Y2=2.34
r527 50 103 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.695 $Y=2.34
+ $X2=5.695 $Y2=2.105
r528 48 238 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.72
r529 48 50 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.695 $Y=2.635
+ $X2=5.695 $Y2=2.34
r530 43 46 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=3.22 $Y=1.63
+ $X2=3.22 $Y2=2.31
r531 41 99 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.72
r532 41 46 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=3.22 $Y=2.635
+ $X2=3.22 $Y2=2.31
r533 40 96 9.02747 $w=2.98e-07 $l=2.35e-07 $layer=LI1_cond $X=0.745 $Y=2.34
+ $X2=0.745 $Y2=2.105
r534 38 235 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.72
r535 38 40 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.745 $Y=2.635
+ $X2=0.745 $Y2=2.34
r536 12 134 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=1.94
r537 12 92 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=24.885
+ $Y=1.485 $X2=25.03 $Y2=2.34
r538 11 88 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=1.485 $X2=22.54 $Y2=2.31
r539 11 85 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=22.36
+ $Y=1.485 $X2=22.54 $Y2=1.63
r540 10 127 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=19.905
+ $Y=1.485 $X2=20.05 $Y2=1.94
r541 10 82 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=19.905
+ $Y=1.485 $X2=20.05 $Y2=2.34
r542 9 123 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=18.445
+ $Y=1.485 $X2=18.59 $Y2=1.94
r543 9 78 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=18.445
+ $Y=1.485 $X2=18.59 $Y2=2.34
r544 8 74 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=1.485 $X2=16.1 $Y2=2.31
r545 8 71 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=15.92
+ $Y=1.485 $X2=16.1 $Y2=1.63
r546 7 116 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=1.94
r547 7 68 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=13.465
+ $Y=1.485 $X2=13.61 $Y2=2.34
r548 6 112 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=1.94
r549 6 64 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.005
+ $Y=1.485 $X2=12.15 $Y2=2.34
r550 5 60 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=2.31
r551 5 57 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=9.48
+ $Y=1.485 $X2=9.66 $Y2=1.63
r552 4 105 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=1.94
r553 4 54 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.025
+ $Y=1.485 $X2=7.17 $Y2=2.34
r554 3 101 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=1.94
r555 3 50 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.565
+ $Y=1.485 $X2=5.71 $Y2=2.34
r556 2 46 400 $w=1.7e-07 $l=9.10563e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=2.31
r557 2 43 400 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.485 $X2=3.22 $Y2=1.63
r558 1 94 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.94
r559 1 40 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%Z 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15
+ 16 66 69 72 75 78 81 84 87 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 120 122 126 128 132 134 138 140 144 146 150 152
+ 156 158 162 164
c482 99 0 6.32252e-19 $X=20.785 $Y=1.87
c483 95 0 6.32252e-19 $X=14.345 $Y=1.87
c484 91 0 6.32252e-19 $X=7.905 $Y=1.87
r485 162 164 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=24.08 $Y=1.87
+ $X2=24.08 $Y2=1.755
r486 156 158 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=21 $Y=1.87
+ $X2=21 $Y2=1.755
r487 150 152 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=17.64 $Y=1.87
+ $X2=17.64 $Y2=1.755
r488 144 146 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=14.56 $Y=1.87
+ $X2=14.56 $Y2=1.755
r489 138 140 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=11.2 $Y=1.87
+ $X2=11.2 $Y2=1.755
r490 132 134 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=8.12 $Y=1.87
+ $X2=8.12 $Y2=1.755
r491 126 128 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=4.76 $Y=1.87
+ $X2=4.76 $Y2=1.755
r492 120 122 7.44484 $w=4.28e-07 $l=1.15e-07 $layer=LI1_cond $X=1.68 $Y=1.87
+ $X2=1.68 $Y2=1.755
r493 110 162 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=24.15 $Y=1.87
+ $X2=24.15 $Y2=1.87
r494 109 156 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=20.93 $Y=1.87
+ $X2=20.93 $Y2=1.87
r495 108 150 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=17.71 $Y=1.87
+ $X2=17.71 $Y2=1.87
r496 107 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.49 $Y=1.87
+ $X2=14.49 $Y2=1.87
r497 106 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=1.87
+ $X2=11.27 $Y2=1.87
r498 105 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.05 $Y=1.87
+ $X2=8.05 $Y2=1.87
r499 104 126 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=1.87
+ $X2=4.83 $Y2=1.87
r500 103 120 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=1.87
+ $X2=1.61 $Y2=1.87
r501 102 109 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=21.075 $Y=1.87
+ $X2=20.93 $Y2=1.87
r502 101 110 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=24.005 $Y=1.87
+ $X2=24.15 $Y2=1.87
r503 101 102 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=24.005 $Y=1.87
+ $X2=21.075 $Y2=1.87
r504 100 108 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.855 $Y=1.87
+ $X2=17.71 $Y2=1.87
r505 99 109 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=20.785 $Y=1.87
+ $X2=20.93 $Y2=1.87
r506 99 100 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=20.785 $Y=1.87
+ $X2=17.855 $Y2=1.87
r507 98 107 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.635 $Y=1.87
+ $X2=14.49 $Y2=1.87
r508 97 108 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=17.565 $Y=1.87
+ $X2=17.71 $Y2=1.87
r509 97 98 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=17.565 $Y=1.87
+ $X2=14.635 $Y2=1.87
r510 96 106 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.415 $Y=1.87
+ $X2=11.27 $Y2=1.87
r511 95 107 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=14.345 $Y=1.87
+ $X2=14.49 $Y2=1.87
r512 95 96 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=14.345 $Y=1.87
+ $X2=11.415 $Y2=1.87
r513 94 105 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.195 $Y=1.87
+ $X2=8.05 $Y2=1.87
r514 93 106 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=11.27 $Y2=1.87
r515 93 94 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=11.125 $Y=1.87
+ $X2=8.195 $Y2=1.87
r516 92 104 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.975 $Y=1.87
+ $X2=4.83 $Y2=1.87
r517 91 105 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=8.05 $Y2=1.87
r518 91 92 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=7.905 $Y=1.87
+ $X2=4.975 $Y2=1.87
r519 90 103 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.755 $Y=1.87
+ $X2=1.61 $Y2=1.87
r520 89 104 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=4.83 $Y2=1.87
r521 89 90 3.62623 $w=1.4e-07 $l=2.93e-06 $layer=MET1_cond $X=4.685 $Y=1.87
+ $X2=1.755 $Y2=1.87
r522 63 87 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=24.09 $Y=0.885
+ $X2=24.09 $Y2=0.68
r523 63 164 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=24.09 $Y=0.885
+ $X2=24.09 $Y2=1.755
r524 61 84 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=20.99 $Y=0.885
+ $X2=20.99 $Y2=0.68
r525 61 158 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=20.99 $Y=0.885
+ $X2=20.99 $Y2=1.755
r526 59 81 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=17.65 $Y=0.885
+ $X2=17.65 $Y2=0.68
r527 59 152 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=17.65 $Y=0.885
+ $X2=17.65 $Y2=1.755
r528 57 78 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=14.55 $Y=0.885
+ $X2=14.55 $Y2=0.68
r529 57 146 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=14.55 $Y=0.885
+ $X2=14.55 $Y2=1.755
r530 55 75 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=0.68
r531 55 140 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=11.21 $Y=0.885
+ $X2=11.21 $Y2=1.755
r532 53 72 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=0.68
r533 53 134 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=8.11 $Y=0.885
+ $X2=8.11 $Y2=1.755
r534 51 69 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=0.68
r535 51 128 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=4.77 $Y=0.885
+ $X2=4.77 $Y2=1.755
r536 49 66 9.85908 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=0.68
r537 49 122 56.7594 $w=1.68e-07 $l=8.7e-07 $layer=LI1_cond $X=1.67 $Y=0.885
+ $X2=1.67 $Y2=1.755
r538 16 162 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=23.89
+ $Y=1.665 $X2=24.035 $Y2=2.02
r539 15 156 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=20.9
+ $Y=1.665 $X2=21.045 $Y2=2.02
r540 14 150 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=17.45
+ $Y=1.665 $X2=17.595 $Y2=2.02
r541 13 144 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=14.46
+ $Y=1.665 $X2=14.605 $Y2=2.02
r542 12 138 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=11.01
+ $Y=1.665 $X2=11.155 $Y2=2.02
r543 11 132 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=8.02
+ $Y=1.665 $X2=8.165 $Y2=2.02
r544 10 126 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=4.57
+ $Y=1.665 $X2=4.715 $Y2=2.02
r545 9 120 600 $w=1.7e-07 $l=4.21307e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.665 $X2=1.725 $Y2=2.02
r546 8 87 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=23.955
+ $Y=0.345 $X2=24.09 $Y2=0.68
r547 7 84 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=20.855
+ $Y=0.345 $X2=20.99 $Y2=0.68
r548 6 81 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=17.515
+ $Y=0.345 $X2=17.65 $Y2=0.68
r549 5 78 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=14.415
+ $Y=0.345 $X2=14.55 $Y2=0.68
r550 4 75 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=11.075
+ $Y=0.345 $X2=11.21 $Y2=0.68
r551 3 72 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=7.975
+ $Y=0.345 $X2=8.11 $Y2=0.68
r552 2 69 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=4.635
+ $Y=0.345 $X2=4.77 $Y2=0.68
r553 1 66 182 $w=1.7e-07 $l=3.968e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.345 $X2=1.67 $Y2=0.68
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_824_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
c59 3 0 1.22753e-19 $X=6.035 $Y=1.485
r60 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.18 $Y=2.34
+ $X2=6.18 $Y2=2.21
r61 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=1.58
r62 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.195 $Y=1.665
+ $X2=6.195 $Y2=2.21
r63 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=6.195 $Y2=1.58
r64 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=6.045 $Y=1.58
+ $X2=5.325 $Y2=1.58
r65 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.24 $Y=2.295
+ $X2=5.24 $Y2=1.78
r66 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.24 $Y=1.665
+ $X2=5.325 $Y2=1.58
r67 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=5.24 $Y=1.665
+ $X2=5.24 $Y2=1.78
r68 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.155 $Y=2.38
+ $X2=5.24 $Y2=2.295
r69 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=5.155 $Y=2.38
+ $X2=4.33 $Y2=2.38
r70 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.245 $Y=2.295
+ $X2=4.33 $Y2=2.38
r71 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=4.245 $Y=2.295
+ $X2=4.245 $Y2=1.81
r72 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.66
r73 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=2.34
r74 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=5.04
+ $Y=1.665 $X2=5.24 $Y2=1.78
r75 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.12
+ $Y=1.665 $X2=4.245 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_297# 1 2 3 10 12 17 18 19 22 27
+ 28
c57 1 0 1.22753e-19 $X=6.575 $Y=1.485
r58 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=6.7 $Y=2.34 $X2=6.7
+ $Y2=2.21
r59 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=8.635 $Y=2.295
+ $X2=8.635 $Y2=1.81
r60 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.55 $Y=2.38
+ $X2=8.635 $Y2=2.295
r61 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=8.55 $Y=2.38
+ $X2=7.725 $Y2=2.38
r62 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.64 $Y=2.295
+ $X2=7.725 $Y2=2.38
r63 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=7.64 $Y=2.295
+ $X2=7.64 $Y2=1.78
r64 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=7.64 $Y=1.665
+ $X2=7.64 $Y2=1.78
r65 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=6.835 $Y=1.58
+ $X2=6.685 $Y2=1.58
r66 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=7.64 $Y2=1.665
r67 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=7.555 $Y=1.58
+ $X2=6.835 $Y2=1.58
r68 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=1.58
r69 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.685 $Y=1.665
+ $X2=6.685 $Y2=2.21
r70 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=8.49
+ $Y=1.665 $X2=8.635 $Y2=1.81
r71 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=7.495
+ $Y=1.485 $X2=7.64 $Y2=1.78
r72 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=2.34
r73 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=6.575
+ $Y=1.485 $X2=6.7 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2112_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
c59 3 0 1.22753e-19 $X=12.475 $Y=1.485
r60 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=12.62 $Y=2.34
+ $X2=12.62 $Y2=2.21
r61 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=1.58
r62 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=12.635 $Y=1.665
+ $X2=12.635 $Y2=2.21
r63 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=12.635 $Y2=1.58
r64 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=12.485 $Y=1.58
+ $X2=11.765 $Y2=1.58
r65 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=11.68 $Y=2.295
+ $X2=11.68 $Y2=1.78
r66 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.68 $Y=1.665
+ $X2=11.765 $Y2=1.58
r67 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=11.68 $Y=1.665
+ $X2=11.68 $Y2=1.78
r68 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=11.595 $Y=2.38
+ $X2=11.68 $Y2=2.295
r69 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=11.595 $Y=2.38
+ $X2=10.77 $Y2=2.38
r70 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.685 $Y=2.295
+ $X2=10.77 $Y2=2.38
r71 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=10.685 $Y=2.295
+ $X2=10.685 $Y2=1.81
r72 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=1.66
r73 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=12.475
+ $Y=1.485 $X2=12.62 $Y2=2.34
r74 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=11.48
+ $Y=1.665 $X2=11.68 $Y2=1.78
r75 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=10.56
+ $Y=1.665 $X2=10.685 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_297# 1 2 3 10 12 17 18 19 22 27
+ 28
c57 1 0 1.22753e-19 $X=13.015 $Y=1.485
r58 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=13.14 $Y=2.34
+ $X2=13.14 $Y2=2.21
r59 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=15.075 $Y=2.295
+ $X2=15.075 $Y2=1.81
r60 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.99 $Y=2.38
+ $X2=15.075 $Y2=2.295
r61 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=14.99 $Y=2.38
+ $X2=14.165 $Y2=2.38
r62 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.08 $Y=2.295
+ $X2=14.165 $Y2=2.38
r63 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=14.08 $Y=2.295
+ $X2=14.08 $Y2=1.78
r64 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=14.08 $Y=1.665
+ $X2=14.08 $Y2=1.78
r65 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=13.275 $Y=1.58
+ $X2=13.125 $Y2=1.58
r66 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=13.995 $Y=1.58
+ $X2=14.08 $Y2=1.665
r67 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=13.995 $Y=1.58
+ $X2=13.275 $Y2=1.58
r68 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=13.125 $Y=1.665
+ $X2=13.125 $Y2=1.58
r69 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=13.125 $Y=1.665
+ $X2=13.125 $Y2=2.21
r70 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=14.93
+ $Y=1.665 $X2=15.075 $Y2=1.81
r71 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=13.935
+ $Y=1.485 $X2=14.08 $Y2=1.78
r72 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=2.34
r73 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=13.015
+ $Y=1.485 $X2=13.14 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3400_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
c59 3 0 1.22753e-19 $X=18.915 $Y=1.485
r60 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=19.06 $Y=2.34
+ $X2=19.06 $Y2=2.21
r61 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.075 $Y=1.665
+ $X2=19.075 $Y2=1.58
r62 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=19.075 $Y=1.665
+ $X2=19.075 $Y2=2.21
r63 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=18.925 $Y=1.58
+ $X2=19.075 $Y2=1.58
r64 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=18.925 $Y=1.58
+ $X2=18.205 $Y2=1.58
r65 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=18.12 $Y=2.295
+ $X2=18.12 $Y2=1.78
r66 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=18.12 $Y=1.665
+ $X2=18.205 $Y2=1.58
r67 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=18.12 $Y=1.665
+ $X2=18.12 $Y2=1.78
r68 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=18.035 $Y=2.38
+ $X2=18.12 $Y2=2.295
r69 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=18.035 $Y=2.38
+ $X2=17.21 $Y2=2.38
r70 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.125 $Y=2.295
+ $X2=17.21 $Y2=2.38
r71 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=17.125 $Y=2.295
+ $X2=17.125 $Y2=1.81
r72 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=18.915
+ $Y=1.485 $X2=19.06 $Y2=1.66
r73 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=18.915
+ $Y=1.485 $X2=19.06 $Y2=2.34
r74 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=17.92
+ $Y=1.665 $X2=18.12 $Y2=1.78
r75 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=17
+ $Y=1.665 $X2=17.125 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_297# 1 2 3 10 12 17 18 19 22 27
+ 28
c57 1 0 1.22753e-19 $X=19.455 $Y=1.485
r58 27 28 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=19.58 $Y=2.34
+ $X2=19.58 $Y2=2.21
r59 20 22 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=21.515 $Y=2.295
+ $X2=21.515 $Y2=1.81
r60 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=21.43 $Y=2.38
+ $X2=21.515 $Y2=2.295
r61 18 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=21.43 $Y=2.38
+ $X2=20.605 $Y2=2.38
r62 15 19 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=20.52 $Y=2.295
+ $X2=20.605 $Y2=2.38
r63 15 17 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=20.52 $Y=2.295
+ $X2=20.52 $Y2=1.78
r64 14 17 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=20.52 $Y=1.665
+ $X2=20.52 $Y2=1.78
r65 13 25 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=19.715 $Y=1.58
+ $X2=19.565 $Y2=1.58
r66 12 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=20.435 $Y=1.58
+ $X2=20.52 $Y2=1.665
r67 12 13 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=20.435 $Y=1.58
+ $X2=19.715 $Y2=1.58
r68 10 25 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=19.565 $Y=1.665
+ $X2=19.565 $Y2=1.58
r69 10 28 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=19.565 $Y=1.665
+ $X2=19.565 $Y2=2.21
r70 3 22 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=21.37
+ $Y=1.665 $X2=21.515 $Y2=1.81
r71 2 17 300 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_PDIFF $count=2 $X=20.375
+ $Y=1.485 $X2=20.52 $Y2=1.78
r72 1 27 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=19.455
+ $Y=1.485 $X2=19.58 $Y2=2.34
r73 1 25 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=19.455
+ $Y=1.485 $X2=19.58 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4688_333# 1 2 3 12 14 15 19 20 21 22
+ 25 26
r49 25 26 4.65811 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=25.5 $Y=2.34
+ $X2=25.5 $Y2=2.21
r50 22 29 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=25.515 $Y=1.665
+ $X2=25.515 $Y2=1.58
r51 22 26 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=25.515 $Y=1.665
+ $X2=25.515 $Y2=2.21
r52 20 29 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=25.365 $Y=1.58
+ $X2=25.515 $Y2=1.58
r53 20 21 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=25.365 $Y=1.58
+ $X2=24.645 $Y2=1.58
r54 17 19 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=24.56 $Y=2.295
+ $X2=24.56 $Y2=1.78
r55 16 21 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=24.56 $Y=1.665
+ $X2=24.645 $Y2=1.58
r56 16 19 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=24.56 $Y=1.665
+ $X2=24.56 $Y2=1.78
r57 14 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=24.475 $Y=2.38
+ $X2=24.56 $Y2=2.295
r58 14 15 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=24.475 $Y=2.38
+ $X2=23.65 $Y2=2.38
r59 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=23.565 $Y=2.295
+ $X2=23.65 $Y2=2.38
r60 10 12 31.6417 $w=1.68e-07 $l=4.85e-07 $layer=LI1_cond $X=23.565 $Y=2.295
+ $X2=23.565 $Y2=1.81
r61 3 29 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=1.66
r62 3 25 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=25.355
+ $Y=1.485 $X2=25.5 $Y2=2.34
r63 2 19 300 $w=1.7e-07 $l=2.50998e-07 $layer=licon1_PDIFF $count=2 $X=24.36
+ $Y=1.665 $X2=24.56 $Y2=1.78
r64 1 12 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=23.44
+ $Y=1.665 $X2=23.565 $Y2=1.81
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_27_47# 1 2 3 12 14 15 16 18 22
c42 16 0 1.81988e-19 $X=1.182 $Y=0.425
r43 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=2.09 $Y=0.425
+ $X2=2.09 $Y2=0.605
r44 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=1.335 $Y=0.34
+ $X2=1.182 $Y2=0.34
r45 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=2.09 $Y2=0.425
r46 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=2.005 $Y=0.34
+ $X2=1.335 $Y2=0.34
r47 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.34
r48 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=1.182 $Y=0.425
+ $X2=1.182 $Y2=0.715
r49 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=1.182 $Y2=0.715
r50 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=1.03 $Y=0.8
+ $X2=0.475 $Y2=0.8
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.475 $Y2=0.8
r52 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.31 $Y=0.715
+ $X2=0.31 $Y2=0.38
r53 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.345 $X2=2.09 $Y2=0.605
r54 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=1.015
+ $Y=0.235 $X2=1.175 $Y2=0.42
r55 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.31 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%VGND 1 2 3 4 5 6 7 8 9 10 11 12 41 45
+ 49 51 55 59 63 65 69 73 77 79 83 87 91 94 95 97 98 100 101 103 104 106 107 108
+ 109 110 111 112 113 114 115 131 145 159 180 184 187 190 193 196 199 202
r285 202 203 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=20.01 $Y=0
+ $X2=20.01 $Y2=0
r286 199 200 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=18.63 $Y=0
+ $X2=18.63 $Y2=0
r287 196 197 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r288 193 194 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=12.19 $Y=0
+ $X2=12.19 $Y2=0
r289 190 191 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0
+ $X2=7.13 $Y2=0
r290 187 188 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r291 184 185 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r292 177 178 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=24.61 $Y=0
+ $X2=24.61 $Y2=0
r293 175 178 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=22.77 $Y=0
+ $X2=24.61 $Y2=0
r294 174 177 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=22.77 $Y=0
+ $X2=24.61 $Y2=0
r295 174 175 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.77 $Y=0
+ $X2=22.77 $Y2=0
r296 172 175 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=22.31 $Y=0
+ $X2=22.77 $Y2=0
r297 171 172 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=22.31 $Y=0
+ $X2=22.31 $Y2=0
r298 169 172 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=22.31 $Y2=0
r299 169 203 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=20.47 $Y=0
+ $X2=20.01 $Y2=0
r300 168 171 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=20.47 $Y=0
+ $X2=22.31 $Y2=0
r301 168 169 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=20.47 $Y=0
+ $X2=20.47 $Y2=0
r302 166 202 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=20.18 $Y=0
+ $X2=20.072 $Y2=0
r303 166 168 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=20.18 $Y=0
+ $X2=20.47 $Y2=0
r304 165 200 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=18.17 $Y=0
+ $X2=18.63 $Y2=0
r305 164 165 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=18.17 $Y=0
+ $X2=18.17 $Y2=0
r306 162 165 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=16.33 $Y=0
+ $X2=18.17 $Y2=0
r307 161 164 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=16.33 $Y=0
+ $X2=18.17 $Y2=0
r308 161 162 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=16.33 $Y=0
+ $X2=16.33 $Y2=0
r309 159 199 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=18.46 $Y=0
+ $X2=18.567 $Y2=0
r310 159 164 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=18.46 $Y=0
+ $X2=18.17 $Y2=0
r311 158 162 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=15.87 $Y=0
+ $X2=16.33 $Y2=0
r312 157 158 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=15.87 $Y=0
+ $X2=15.87 $Y2=0
r313 155 158 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=15.87 $Y2=0
r314 155 197 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.03 $Y=0
+ $X2=13.57 $Y2=0
r315 154 157 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=14.03 $Y=0
+ $X2=15.87 $Y2=0
r316 154 155 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=14.03 $Y=0
+ $X2=14.03 $Y2=0
r317 152 196 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=13.74 $Y=0
+ $X2=13.632 $Y2=0
r318 152 154 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=13.74 $Y=0
+ $X2=14.03 $Y2=0
r319 151 194 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.19 $Y2=0
r320 150 151 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r321 148 151 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r322 147 150 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=9.89 $Y=0
+ $X2=11.73 $Y2=0
r323 147 148 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r324 145 193 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=12.127 $Y2=0
r325 145 150 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=12.02 $Y=0
+ $X2=11.73 $Y2=0
r326 144 148 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r327 143 144 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r328 141 144 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r329 141 191 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=7.13 $Y2=0
r330 140 143 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=7.59 $Y=0
+ $X2=9.43 $Y2=0
r331 140 141 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r332 138 190 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=7.3 $Y=0
+ $X2=7.192 $Y2=0
r333 138 140 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=7.3 $Y=0 $X2=7.59
+ $Y2=0
r334 137 188 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0
+ $X2=5.75 $Y2=0
r335 136 137 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=5.29 $Y=0
+ $X2=5.29 $Y2=0
r336 134 137 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r337 133 136 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=3.45 $Y=0
+ $X2=5.29 $Y2=0
r338 133 134 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=3.45 $Y=0
+ $X2=3.45 $Y2=0
r339 131 187 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=5.58 $Y=0
+ $X2=5.687 $Y2=0
r340 131 136 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=5.58 $Y=0
+ $X2=5.29 $Y2=0
r341 130 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.45 $Y2=0
r342 129 130 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r343 127 130 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r344 127 185 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=0.69 $Y2=0
r345 126 129 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=1.15 $Y=0
+ $X2=2.99 $Y2=0
r346 126 127 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r347 124 184 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=0.86 $Y=0
+ $X2=0.752 $Y2=0
r348 124 126 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.86 $Y=0
+ $X2=1.15 $Y2=0
r349 115 178 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=25.53 $Y=0
+ $X2=24.61 $Y2=0
r350 115 180 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=25.53 $Y=0
+ $X2=25.53 $Y2=0
r351 114 203 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.55 $Y=0
+ $X2=20.01 $Y2=0
r352 113 114 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=0
+ $X2=19.55 $Y2=0
r353 113 200 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=19.09 $Y=0
+ $X2=18.63 $Y2=0
r354 112 197 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=13.11 $Y=0
+ $X2=13.57 $Y2=0
r355 111 112 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=13.11 $Y2=0
r356 111 194 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=12.65 $Y=0
+ $X2=12.19 $Y2=0
r357 110 191 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.13 $Y2=0
r358 109 110 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=6.67 $Y2=0
r359 109 188 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0
+ $X2=5.75 $Y2=0
r360 108 185 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r361 106 177 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=24.9 $Y=0
+ $X2=24.61 $Y2=0
r362 106 107 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=24.9 $Y=0
+ $X2=25.007 $Y2=0
r363 105 180 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=25.115 $Y=0
+ $X2=25.53 $Y2=0
r364 105 107 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=25.115 $Y=0
+ $X2=25.007 $Y2=0
r365 103 171 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.415 $Y=0
+ $X2=22.31 $Y2=0
r366 103 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.415 $Y=0
+ $X2=22.54 $Y2=0
r367 102 174 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=22.665 $Y=0
+ $X2=22.77 $Y2=0
r368 102 104 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=22.665 $Y=0
+ $X2=22.54 $Y2=0
r369 100 157 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=15.975 $Y=0
+ $X2=15.87 $Y2=0
r370 100 101 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=15.975 $Y=0
+ $X2=16.1 $Y2=0
r371 99 161 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=16.225 $Y=0
+ $X2=16.33 $Y2=0
r372 99 101 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=16.225 $Y=0
+ $X2=16.1 $Y2=0
r373 97 143 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.535 $Y=0
+ $X2=9.43 $Y2=0
r374 97 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.535 $Y=0 $X2=9.66
+ $Y2=0
r375 96 147 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=9.785 $Y=0
+ $X2=9.89 $Y2=0
r376 96 98 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=9.785 $Y=0 $X2=9.66
+ $Y2=0
r377 94 129 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.095 $Y=0
+ $X2=2.99 $Y2=0
r378 94 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.095 $Y=0 $X2=3.22
+ $Y2=0
r379 93 133 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=3.345 $Y=0
+ $X2=3.45 $Y2=0
r380 93 95 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.345 $Y=0 $X2=3.22
+ $Y2=0
r381 89 107 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=25.007 $Y=0.085
+ $X2=25.007 $Y2=0
r382 89 91 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=25.007 $Y=0.085
+ $X2=25.007 $Y2=0.38
r383 85 104 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=22.54 $Y=0.085
+ $X2=22.54 $Y2=0
r384 85 87 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=22.54 $Y=0.085
+ $X2=22.54 $Y2=0.495
r385 81 202 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=20.072 $Y=0.085
+ $X2=20.072 $Y2=0
r386 81 83 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=20.072 $Y=0.085
+ $X2=20.072 $Y2=0.38
r387 80 199 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=18.675 $Y=0
+ $X2=18.567 $Y2=0
r388 79 202 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=19.965 $Y=0
+ $X2=20.072 $Y2=0
r389 79 80 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=19.965 $Y=0
+ $X2=18.675 $Y2=0
r390 75 199 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=18.567 $Y=0.085
+ $X2=18.567 $Y2=0
r391 75 77 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=18.567 $Y=0.085
+ $X2=18.567 $Y2=0.38
r392 71 101 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=16.1 $Y=0.085
+ $X2=16.1 $Y2=0
r393 71 73 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=16.1 $Y=0.085
+ $X2=16.1 $Y2=0.495
r394 67 196 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=13.632 $Y=0.085
+ $X2=13.632 $Y2=0
r395 67 69 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=13.632 $Y=0.085
+ $X2=13.632 $Y2=0.38
r396 66 193 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=12.235 $Y=0
+ $X2=12.127 $Y2=0
r397 65 196 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=13.525 $Y=0
+ $X2=13.632 $Y2=0
r398 65 66 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=13.525 $Y=0
+ $X2=12.235 $Y2=0
r399 61 193 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0
r400 61 63 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=12.127 $Y=0.085
+ $X2=12.127 $Y2=0.38
r401 57 98 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0
r402 57 59 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0.495
r403 53 190 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0
r404 53 55 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=7.192 $Y=0.085
+ $X2=7.192 $Y2=0.38
r405 52 187 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=5.795 $Y=0
+ $X2=5.687 $Y2=0
r406 51 190 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=7.192 $Y2=0
r407 51 52 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=7.085 $Y=0
+ $X2=5.795 $Y2=0
r408 47 187 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0
r409 47 49 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=5.687 $Y=0.085
+ $X2=5.687 $Y2=0.38
r410 43 95 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0
r411 43 45 18.9001 $w=2.48e-07 $l=4.1e-07 $layer=LI1_cond $X=3.22 $Y=0.085
+ $X2=3.22 $Y2=0.495
r412 39 184 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0
r413 39 41 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=0.752 $Y=0.085
+ $X2=0.752 $Y2=0.38
r414 12 91 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=24.895
+ $Y=0.235 $X2=25.03 $Y2=0.38
r415 11 87 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=22.405
+ $Y=0.235 $X2=22.54 $Y2=0.495
r416 10 83 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=19.915
+ $Y=0.235 $X2=20.05 $Y2=0.38
r417 9 77 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=18.455
+ $Y=0.235 $X2=18.59 $Y2=0.38
r418 8 73 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=15.965
+ $Y=0.235 $X2=16.1 $Y2=0.495
r419 7 69 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=13.475
+ $Y=0.235 $X2=13.61 $Y2=0.38
r420 6 63 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=12.015
+ $Y=0.235 $X2=12.15 $Y2=0.38
r421 5 59 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=9.525
+ $Y=0.235 $X2=9.66 $Y2=0.495
r422 4 55 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=7.035
+ $Y=0.235 $X2=7.17 $Y2=0.38
r423 3 49 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=5.575
+ $Y=0.235 $X2=5.71 $Y2=0.38
r424 2 45 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.22 $Y2=0.495
r425 1 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_845_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=5.257 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.13 $Y=0.715
+ $X2=6.13 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=6.13 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=5.965 $Y=0.8
+ $X2=5.41 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=5.257 $Y=0.715
+ $X2=5.41 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=5.257 $Y=0.425
+ $X2=5.257 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=5.257 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.105 $Y=0.34
+ $X2=4.435 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.435 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=4.35 $Y=0.425
+ $X2=4.35 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.995
+ $Y=0.235 $X2=6.13 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=5.055
+ $Y=0.345 $X2=5.265 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=4.225
+ $Y=0.345 $X2=4.35 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_1315_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=7.622 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=8.53 $Y=0.425
+ $X2=8.53 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=7.775 $Y=0.34
+ $X2=7.622 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=8.53 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=8.445 $Y=0.34
+ $X2=7.775 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=7.622 $Y=0.425
+ $X2=7.622 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=7.622 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=7.47 $Y=0.8
+ $X2=6.915 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.915 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=6.75 $Y=0.715
+ $X2=6.75 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=8.395
+ $Y=0.345 $X2=8.53 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=7.455
+ $Y=0.235 $X2=7.615 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=6.575
+ $Y=0.235 $X2=6.75 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2133_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=11.697 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=12.57 $Y=0.715
+ $X2=12.57 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=12.57 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=12.405 $Y=0.8
+ $X2=11.85 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=11.697 $Y=0.715
+ $X2=11.85 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=11.697 $Y=0.425
+ $X2=11.697 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=11.697 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=11.545 $Y=0.34
+ $X2=10.875 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.875 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=10.79 $Y=0.425
+ $X2=10.79 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=12.435
+ $Y=0.235 $X2=12.57 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=11.495
+ $Y=0.345 $X2=11.705 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=10.665
+ $Y=0.345 $X2=10.79 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_2603_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=14.062 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=14.97 $Y=0.425
+ $X2=14.97 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=14.215 $Y=0.34
+ $X2=14.062 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=14.885 $Y=0.34
+ $X2=14.97 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=14.885 $Y=0.34
+ $X2=14.215 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=14.062 $Y=0.425
+ $X2=14.062 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=14.062 $Y=0.425
+ $X2=14.062 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=13.91 $Y=0.8
+ $X2=14.062 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=13.91 $Y=0.8
+ $X2=13.355 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=13.19 $Y=0.715
+ $X2=13.355 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=13.19 $Y=0.715
+ $X2=13.19 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=14.835
+ $Y=0.345 $X2=14.97 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=13.895
+ $Y=0.235 $X2=14.055 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=13.015
+ $Y=0.235 $X2=13.19 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3421_69# 1 2 3 12 14 15 16 18 19 22
c48 16 0 1.81988e-19 $X=18.137 $Y=0.425
r49 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=19.01 $Y=0.715
+ $X2=19.01 $Y2=0.38
r50 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=18.845 $Y=0.8
+ $X2=19.01 $Y2=0.715
r51 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=18.845 $Y=0.8
+ $X2=18.29 $Y2=0.8
r52 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=18.137 $Y=0.715
+ $X2=18.29 $Y2=0.8
r53 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=18.137 $Y=0.425
+ $X2=18.137 $Y2=0.34
r54 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=18.137 $Y=0.425
+ $X2=18.137 $Y2=0.715
r55 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=17.985 $Y=0.34
+ $X2=18.137 $Y2=0.34
r56 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=17.985 $Y=0.34
+ $X2=17.315 $Y2=0.34
r57 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=17.23 $Y=0.425
+ $X2=17.315 $Y2=0.34
r58 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=17.23 $Y=0.425
+ $X2=17.23 $Y2=0.605
r59 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=18.875
+ $Y=0.235 $X2=19.01 $Y2=0.38
r60 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=17.935
+ $Y=0.345 $X2=18.145 $Y2=0.42
r61 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=17.105
+ $Y=0.345 $X2=17.23 $Y2=0.605
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_3891_47# 1 2 3 12 14 15 16 18 22
c44 16 0 1.81988e-19 $X=20.502 $Y=0.425
r45 20 22 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=21.41 $Y=0.425
+ $X2=21.41 $Y2=0.605
r46 19 25 4.85887 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=20.655 $Y=0.34
+ $X2=20.502 $Y2=0.34
r47 18 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=21.325 $Y=0.34
+ $X2=21.41 $Y2=0.425
r48 18 19 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=21.325 $Y=0.34
+ $X2=20.655 $Y2=0.34
r49 16 25 2.69937 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=20.502 $Y=0.425
+ $X2=20.502 $Y2=0.34
r50 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=20.502 $Y=0.425
+ $X2=20.502 $Y2=0.715
r51 14 17 7.55824 $w=1.7e-07 $l=1.898e-07 $layer=LI1_cond $X=20.35 $Y=0.8
+ $X2=20.502 $Y2=0.715
r52 14 15 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=20.35 $Y=0.8
+ $X2=19.795 $Y2=0.8
r53 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=19.63 $Y=0.715
+ $X2=19.795 $Y2=0.8
r54 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=19.63 $Y=0.715
+ $X2=19.63 $Y2=0.38
r55 3 22 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=21.275
+ $Y=0.345 $X2=21.41 $Y2=0.605
r56 2 25 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=20.335
+ $Y=0.235 $X2=20.495 $Y2=0.42
r57 1 12 91 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_NDIFF $count=2 $X=19.455
+ $Y=0.235 $X2=19.63 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUXB8TO1_2%A_4709_69# 1 2 3 12 14 15 16 18 19 22
c46 16 0 1.81988e-19 $X=24.577 $Y=0.425
r47 20 22 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=25.45 $Y=0.715
+ $X2=25.45 $Y2=0.38
r48 18 20 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=25.285 $Y=0.8
+ $X2=25.45 $Y2=0.715
r49 18 19 36.2086 $w=1.68e-07 $l=5.55e-07 $layer=LI1_cond $X=25.285 $Y=0.8
+ $X2=24.73 $Y2=0.8
r50 17 19 7.55824 $w=1.7e-07 $l=1.90825e-07 $layer=LI1_cond $X=24.577 $Y=0.715
+ $X2=24.73 $Y2=0.8
r51 16 25 2.71076 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=24.577 $Y=0.425
+ $X2=24.577 $Y2=0.34
r52 16 17 10.9577 $w=3.03e-07 $l=2.9e-07 $layer=LI1_cond $X=24.577 $Y=0.425
+ $X2=24.577 $Y2=0.715
r53 14 25 4.84748 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=24.425 $Y=0.34
+ $X2=24.577 $Y2=0.34
r54 14 15 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=24.425 $Y=0.34
+ $X2=23.755 $Y2=0.34
r55 10 15 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=23.67 $Y=0.425
+ $X2=23.755 $Y2=0.34
r56 10 12 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=23.67 $Y=0.425
+ $X2=23.67 $Y2=0.605
r57 3 22 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=25.315
+ $Y=0.235 $X2=25.45 $Y2=0.38
r58 2 25 91 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=2 $X=24.375
+ $Y=0.345 $X2=24.585 $Y2=0.42
r59 1 12 182 $w=1.7e-07 $l=3.16386e-07 $layer=licon1_NDIFF $count=1 $X=23.545
+ $Y=0.345 $X2=23.67 $Y2=0.605
.ends

