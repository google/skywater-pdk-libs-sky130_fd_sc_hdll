* File: sky130_fd_sc_hdll__muxb8to1_1.pxi.spice
* Created: Thu Aug 27 19:12:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[0] N_D[0]_c_272_n N_D[0]_M1040_g
+ N_D[0]_c_273_n N_D[0]_M1015_g N_D[0]_c_274_n N_D[0]_c_275_n D[0]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_184_265# N_A_184_265#_M1029_s
+ N_A_184_265#_M1023_s N_A_184_265#_M1019_g N_A_184_265#_c_300_n
+ N_A_184_265#_c_301_n N_A_184_265#_c_305_n N_A_184_265#_c_302_n
+ N_A_184_265#_c_303_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_184_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[0] N_S[0]_c_356_n N_S[0]_M1044_g
+ N_S[0]_c_357_n N_S[0]_c_358_n N_S[0]_c_359_n N_S[0]_M1023_g N_S[0]_c_360_n
+ N_S[0]_M1029_g S[0] N_S[0]_c_361_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[0]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[1] N_S[1]_c_403_n N_S[1]_M1020_g
+ N_S[1]_c_404_n N_S[1]_M1028_g N_S[1]_c_405_n N_S[1]_c_406_n N_S[1]_M1014_g
+ S[1] N_S[1]_c_407_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_533_47# N_A_533_47#_M1028_d
+ N_A_533_47#_M1020_d N_A_533_47#_M1009_g N_A_533_47#_c_452_n
+ N_A_533_47#_c_447_n N_A_533_47#_c_448_n N_A_533_47#_c_449_n
+ N_A_533_47#_c_450_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_533_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[1] N_D[1]_c_502_n N_D[1]_M1035_g
+ N_D[1]_c_503_n N_D[1]_M1032_g N_D[1]_c_504_n N_D[1]_c_505_n D[1]
+ N_D[1]_c_534_p PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[1]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[2] N_D[2]_c_539_n N_D[2]_M1001_g
+ N_D[2]_c_540_n N_D[2]_M1021_g N_D[2]_c_541_n N_D[2]_c_542_n D[2]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1012_265# N_A_1012_265#_M1042_s
+ N_A_1012_265#_M1025_s N_A_1012_265#_M1022_g N_A_1012_265#_c_576_n
+ N_A_1012_265#_c_577_n N_A_1012_265#_c_581_n N_A_1012_265#_c_578_n
+ N_A_1012_265#_c_579_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1012_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[2] N_S[2]_c_632_n N_S[2]_M1010_g
+ N_S[2]_c_633_n N_S[2]_c_634_n N_S[2]_c_635_n N_S[2]_M1025_g N_S[2]_c_636_n
+ N_S[2]_M1042_g S[2] N_S[2]_c_637_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[2]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[3] N_S[3]_c_679_n N_S[3]_M1005_g
+ N_S[3]_c_680_n N_S[3]_M1027_g N_S[3]_c_681_n N_S[3]_c_682_n N_S[3]_M1008_g
+ S[3] N_S[3]_c_683_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1361_47# N_A_1361_47#_M1027_d
+ N_A_1361_47#_M1005_d N_A_1361_47#_M1013_g N_A_1361_47#_c_728_n
+ N_A_1361_47#_c_723_n N_A_1361_47#_c_724_n N_A_1361_47#_c_725_n
+ N_A_1361_47#_c_726_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1361_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[3] N_D[3]_c_778_n N_D[3]_M1016_g
+ N_D[3]_c_779_n N_D[3]_M1039_g N_D[3]_c_780_n N_D[3]_c_781_n D[3]
+ N_D[3]_c_810_p PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[3]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[4] N_D[4]_c_815_n N_D[4]_M1000_g
+ N_D[4]_c_816_n N_D[4]_M1003_g N_D[4]_c_817_n N_D[4]_c_818_n D[4]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1840_265# N_A_1840_265#_M1046_s
+ N_A_1840_265#_M1038_s N_A_1840_265#_M1007_g N_A_1840_265#_c_852_n
+ N_A_1840_265#_c_853_n N_A_1840_265#_c_857_n N_A_1840_265#_c_854_n
+ N_A_1840_265#_c_855_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_1840_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[4] N_S[4]_c_908_n N_S[4]_M1018_g
+ N_S[4]_c_909_n N_S[4]_c_910_n N_S[4]_c_911_n N_S[4]_M1038_g N_S[4]_c_912_n
+ N_S[4]_M1046_g S[4] N_S[4]_c_913_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[4]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[5] N_S[5]_c_955_n N_S[5]_M1024_g
+ N_S[5]_c_956_n N_S[5]_M1037_g N_S[5]_c_957_n N_S[5]_c_958_n N_S[5]_M1012_g
+ S[5] N_S[5]_c_959_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2189_47# N_A_2189_47#_M1037_d
+ N_A_2189_47#_M1024_d N_A_2189_47#_M1030_g N_A_2189_47#_c_1004_n
+ N_A_2189_47#_c_999_n N_A_2189_47#_c_1000_n N_A_2189_47#_c_1001_n
+ N_A_2189_47#_c_1002_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2189_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[5] N_D[5]_c_1054_n N_D[5]_M1036_g
+ N_D[5]_c_1055_n N_D[5]_M1041_g N_D[5]_c_1056_n N_D[5]_c_1057_n D[5]
+ N_D[5]_c_1086_p PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[5]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[6] N_D[6]_c_1091_n N_D[6]_M1002_g
+ N_D[6]_c_1092_n N_D[6]_M1017_g N_D[6]_c_1093_n N_D[6]_c_1094_n D[6]
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2668_265# N_A_2668_265#_M1004_s
+ N_A_2668_265#_M1034_s N_A_2668_265#_M1026_g N_A_2668_265#_c_1128_n
+ N_A_2668_265#_c_1129_n N_A_2668_265#_c_1133_n N_A_2668_265#_c_1130_n
+ N_A_2668_265#_c_1131_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_2668_265#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[6] N_S[6]_c_1184_n N_S[6]_M1033_g
+ N_S[6]_c_1185_n N_S[6]_c_1186_n N_S[6]_c_1187_n N_S[6]_M1034_g N_S[6]_c_1188_n
+ N_S[6]_M1004_g S[6] N_S[6]_c_1189_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[6]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[7] N_S[7]_c_1231_n N_S[7]_M1011_g
+ N_S[7]_c_1232_n N_S[7]_M1047_g N_S[7]_c_1233_n N_S[7]_c_1234_n N_S[7]_M1031_g
+ S[7] N_S[7]_c_1235_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%S[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_3017_47# N_A_3017_47#_M1047_d
+ N_A_3017_47#_M1011_d N_A_3017_47#_M1045_g N_A_3017_47#_c_1280_n
+ N_A_3017_47#_c_1275_n N_A_3017_47#_c_1276_n N_A_3017_47#_c_1277_n
+ N_A_3017_47#_c_1278_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%A_3017_47#
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[7] N_D[7]_c_1330_n N_D[7]_M1006_g
+ N_D[7]_c_1331_n N_D[7]_M1043_g N_D[7]_c_1332_n N_D[7]_c_1333_n D[7]
+ N_D[7]_c_1353_p PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%D[7]
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VPWR N_VPWR_M1015_s N_VPWR_M1023_d
+ N_VPWR_M1035_d N_VPWR_M1025_d N_VPWR_M1016_d N_VPWR_M1038_d N_VPWR_M1036_d
+ N_VPWR_M1034_d N_VPWR_M1006_d N_VPWR_c_1359_n N_VPWR_c_1360_n N_VPWR_c_1361_n
+ N_VPWR_c_1362_n N_VPWR_c_1363_n N_VPWR_c_1364_n N_VPWR_c_1365_n
+ N_VPWR_c_1366_n N_VPWR_c_1367_n N_VPWR_c_1368_n N_VPWR_c_1369_n
+ N_VPWR_c_1370_n N_VPWR_c_1371_n N_VPWR_c_1372_n N_VPWR_c_1373_n
+ N_VPWR_c_1374_n N_VPWR_c_1375_n N_VPWR_c_1376_n N_VPWR_c_1377_n VPWR VPWR VPWR
+ VPWR VPWR N_VPWR_c_1379_n N_VPWR_c_1380_n N_VPWR_c_1381_n N_VPWR_c_1382_n
+ N_VPWR_c_1383_n N_VPWR_c_1384_n N_VPWR_c_1385_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VPWR
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%Z N_Z_M1044_d N_Z_M1014_s N_Z_M1010_d
+ N_Z_M1008_s N_Z_M1018_d N_Z_M1012_s N_Z_M1033_d N_Z_M1031_s N_Z_M1019_d
+ N_Z_M1009_s N_Z_M1022_d N_Z_M1013_s N_Z_M1007_d N_Z_M1030_s N_Z_M1026_d
+ N_Z_M1045_s N_Z_c_1624_n N_Z_c_1625_n N_Z_c_1626_n N_Z_c_1649_n N_Z_c_1650_n
+ N_Z_c_1627_n N_Z_c_1628_n N_Z_c_1629_n N_Z_c_1630_n N_Z_c_1631_n N_Z_c_1653_n
+ N_Z_c_1654_n N_Z_c_1632_n N_Z_c_1633_n N_Z_c_1634_n N_Z_c_1635_n N_Z_c_1636_n
+ N_Z_c_1657_n N_Z_c_1658_n N_Z_c_1637_n N_Z_c_1638_n N_Z_c_1639_n N_Z_c_1640_n
+ N_Z_c_1641_n N_Z_c_1661_n N_Z_c_1662_n N_Z_c_1642_n N_Z_c_1643_n N_Z_c_1644_n
+ N_Z_c_1645_n N_Z_c_1646_n N_Z_c_1647_n N_Z_c_1664_n N_Z_c_1696_n N_Z_c_1743_n
+ N_Z_c_1730_n N_Z_c_1665_n N_Z_c_1769_n N_Z_c_1816_n N_Z_c_1803_n N_Z_c_1666_n
+ N_Z_c_1842_n N_Z_c_1889_n N_Z_c_1876_n N_Z_c_1667_n N_Z_c_1915_n Z Z Z Z Z Z Z
+ Z N_Z_c_1668_n N_Z_c_1669_n N_Z_c_1670_n N_Z_c_1671_n N_Z_c_1672_n
+ N_Z_c_1673_n N_Z_c_1674_n N_Z_c_1675_n PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%Z
x_PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VGND N_VGND_M1040_s N_VGND_M1029_d
+ N_VGND_M1032_d N_VGND_M1042_d N_VGND_M1039_d N_VGND_M1046_d N_VGND_M1041_d
+ N_VGND_M1004_d N_VGND_M1043_d N_VGND_c_2109_n N_VGND_c_2110_n N_VGND_c_2111_n
+ N_VGND_c_2112_n N_VGND_c_2113_n N_VGND_c_2114_n N_VGND_c_2115_n
+ N_VGND_c_2116_n N_VGND_c_2117_n N_VGND_c_2118_n N_VGND_c_2119_n
+ N_VGND_c_2120_n N_VGND_c_2121_n N_VGND_c_2122_n N_VGND_c_2123_n
+ N_VGND_c_2124_n N_VGND_c_2125_n N_VGND_c_2126_n N_VGND_c_2127_n VGND VGND VGND
+ VGND VGND N_VGND_c_2129_n N_VGND_c_2130_n N_VGND_c_2131_n N_VGND_c_2132_n
+ N_VGND_c_2133_n N_VGND_c_2134_n N_VGND_c_2135_n
+ PM_SKY130_FD_SC_HDLL__MUXB8TO1_1%VGND
cc_1 VNB N_D[0]_c_272_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_D[0]_c_273_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_D[0]_c_274_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_4 VNB N_D[0]_c_275_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_5 VNB N_A_184_265#_c_300_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_6 VNB N_A_184_265#_c_301_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_184_265#_c_302_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_184_265#_c_303_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_S[0]_c_356_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_S[0]_c_357_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_S[0]_c_358_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_S[0]_c_359_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_13 VNB N_S[0]_c_360_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_14 VNB N_S[0]_c_361_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_15 VNB N_S[1]_c_403_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_16 VNB N_S[1]_c_404_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_S[1]_c_405_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_18 VNB N_S[1]_c_406_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_19 VNB N_S[1]_c_407_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_20 VNB N_A_533_47#_c_447_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_533_47#_c_448_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_533_47#_c_449_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_533_47#_c_450_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_D[1]_c_502_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_25 VNB N_D[1]_c_503_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_26 VNB N_D[1]_c_504_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_27 VNB N_D[1]_c_505_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_D[2]_c_539_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_29 VNB N_D[2]_c_540_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_30 VNB N_D[2]_c_541_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_31 VNB N_D[2]_c_542_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_32 VNB N_A_1012_265#_c_576_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_33 VNB N_A_1012_265#_c_577_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_1012_265#_c_578_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_1012_265#_c_579_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_S[2]_c_632_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_37 VNB N_S[2]_c_633_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_38 VNB N_S[2]_c_634_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_39 VNB N_S[2]_c_635_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_40 VNB N_S[2]_c_636_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_41 VNB N_S[2]_c_637_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_42 VNB N_S[3]_c_679_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_43 VNB N_S[3]_c_680_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_44 VNB N_S[3]_c_681_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_45 VNB N_S[3]_c_682_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_46 VNB N_S[3]_c_683_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_47 VNB N_A_1361_47#_c_723_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_1361_47#_c_724_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_1361_47#_c_725_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_1361_47#_c_726_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_D[3]_c_778_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_52 VNB N_D[3]_c_779_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_53 VNB N_D[3]_c_780_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_54 VNB N_D[3]_c_781_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_D[4]_c_815_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_56 VNB N_D[4]_c_816_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_57 VNB N_D[4]_c_817_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_58 VNB N_D[4]_c_818_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_59 VNB N_A_1840_265#_c_852_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_60 VNB N_A_1840_265#_c_853_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_A_1840_265#_c_854_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_A_1840_265#_c_855_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_S[4]_c_908_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_64 VNB N_S[4]_c_909_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_65 VNB N_S[4]_c_910_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_66 VNB N_S[4]_c_911_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_67 VNB N_S[4]_c_912_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_68 VNB N_S[4]_c_913_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_69 VNB N_S[5]_c_955_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_70 VNB N_S[5]_c_956_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_71 VNB N_S[5]_c_957_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_72 VNB N_S[5]_c_958_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_73 VNB N_S[5]_c_959_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_74 VNB N_A_2189_47#_c_999_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_A_2189_47#_c_1000_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_A_2189_47#_c_1001_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_A_2189_47#_c_1002_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_D[5]_c_1054_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_79 VNB N_D[5]_c_1055_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_80 VNB N_D[5]_c_1056_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_81 VNB N_D[5]_c_1057_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_D[6]_c_1091_n 0.0174886f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_83 VNB N_D[6]_c_1092_n 0.0251359f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_84 VNB N_D[6]_c_1093_n 0.00253531f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_85 VNB N_D[6]_c_1094_n 0.00430529f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.19
cc_86 VNB N_A_2668_265#_c_1128_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_87 VNB N_A_2668_265#_c_1129_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_A_2668_265#_c_1130_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_A_2668_265#_c_1131_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_S[6]_c_1184_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_91 VNB N_S[6]_c_1185_n 0.0502713f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_92 VNB N_S[6]_c_1186_n 0.00937382f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_93 VNB N_S[6]_c_1187_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_94 VNB N_S[6]_c_1188_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_95 VNB N_S[6]_c_1189_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_96 VNB N_S[7]_c_1231_n 0.0331443f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_97 VNB N_S[7]_c_1232_n 0.0188277f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_98 VNB N_S[7]_c_1233_n 0.0596452f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=0.625
cc_99 VNB N_S[7]_c_1234_n 0.0178443f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.19
cc_100 VNB N_S[7]_c_1235_n 0.00873659f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.16
cc_101 VNB N_A_3017_47#_c_1275_n 0.00489787f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_A_3017_47#_c_1276_n 0.00322081f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_A_3017_47#_c_1277_n 0.0120668f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_A_3017_47#_c_1278_n 0.0089001f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_D[7]_c_1330_n 0.0309471f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_106 VNB N_D[7]_c_1331_n 0.0226847f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_107 VNB N_D[7]_c_1332_n 0.00249376f $X=-0.19 $Y=-0.24 $X2=0.645 $Y2=1.055
cc_108 VNB N_D[7]_c_1333_n 0.012124f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB VPWR 0.706209f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_Z_c_1624_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_Z_c_1625_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_Z_c_1626_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_Z_c_1627_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_Z_c_1628_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_Z_c_1629_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_Z_c_1630_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VNB N_Z_c_1631_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_118 VNB N_Z_c_1632_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_119 VNB N_Z_c_1633_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_120 VNB N_Z_c_1634_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_121 VNB N_Z_c_1635_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_122 VNB N_Z_c_1636_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_123 VNB N_Z_c_1637_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_124 VNB N_Z_c_1638_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_125 VNB N_Z_c_1639_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_126 VNB N_Z_c_1640_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_127 VNB N_Z_c_1641_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_128 VNB N_Z_c_1642_n 0.00516268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_129 VNB N_Z_c_1643_n 0.00523842f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_130 VNB N_Z_c_1644_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_131 VNB N_Z_c_1645_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_132 VNB N_Z_c_1646_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_133 VNB N_Z_c_1647_n 0.00277891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_134 VNB N_VGND_c_2109_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_135 VNB N_VGND_c_2110_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_136 VNB N_VGND_c_2111_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_137 VNB N_VGND_c_2112_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_138 VNB N_VGND_c_2113_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_139 VNB N_VGND_c_2114_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_140 VNB N_VGND_c_2115_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_141 VNB N_VGND_c_2116_n 0.00902444f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_142 VNB N_VGND_c_2117_n 0.00561737f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_143 VNB N_VGND_c_2118_n 0.0113488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_144 VNB N_VGND_c_2119_n 0.0320435f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_145 VNB N_VGND_c_2120_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_146 VNB N_VGND_c_2121_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_147 VNB N_VGND_c_2122_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_148 VNB N_VGND_c_2123_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_149 VNB N_VGND_c_2124_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_150 VNB N_VGND_c_2125_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_151 VNB N_VGND_c_2126_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_152 VNB N_VGND_c_2127_n 0.00634747f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_153 VNB VGND 0.799771f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_154 VNB N_VGND_c_2129_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_155 VNB N_VGND_c_2130_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_156 VNB N_VGND_c_2131_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_157 VNB N_VGND_c_2132_n 0.0485067f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_158 VNB N_VGND_c_2133_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_159 VNB N_VGND_c_2134_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_160 VNB N_VGND_c_2135_n 0.00615512f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_161 VPB N_D[0]_c_273_n 0.0335483f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_162 VPB N_D[0]_c_275_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_163 VPB N_A_184_265#_M1019_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_164 VPB N_A_184_265#_c_305_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.425
cc_165 VPB N_A_184_265#_c_302_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_A_184_265#_c_303_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_S[0]_c_359_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_168 VPB N_S[1]_c_403_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_169 VPB N_A_533_47#_M1009_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_170 VPB N_A_533_47#_c_452_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_171 VPB N_A_533_47#_c_448_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_A_533_47#_c_449_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_D[1]_c_502_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_174 VPB N_D[1]_c_505_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_D[2]_c_540_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_176 VPB N_D[2]_c_542_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_177 VPB N_A_1012_265#_M1022_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_178 VPB N_A_1012_265#_c_581_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_179 VPB N_A_1012_265#_c_578_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_A_1012_265#_c_579_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_S[2]_c_635_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_182 VPB N_S[3]_c_679_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_183 VPB N_A_1361_47#_M1013_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_184 VPB N_A_1361_47#_c_728_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_185 VPB N_A_1361_47#_c_724_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_A_1361_47#_c_725_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_D[3]_c_778_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_188 VPB N_D[3]_c_781_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_D[4]_c_816_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_190 VPB N_D[4]_c_818_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_191 VPB N_A_1840_265#_M1007_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_192 VPB N_A_1840_265#_c_857_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_193 VPB N_A_1840_265#_c_854_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_A_1840_265#_c_855_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_S[4]_c_911_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_196 VPB N_S[5]_c_955_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_197 VPB N_A_2189_47#_M1030_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_198 VPB N_A_2189_47#_c_1004_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_199 VPB N_A_2189_47#_c_1000_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_A_2189_47#_c_1001_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_D[5]_c_1054_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_202 VPB N_D[5]_c_1057_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_D[6]_c_1092_n 0.0267097f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_204 VPB N_D[6]_c_1094_n 0.00206353f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_205 VPB N_A_2668_265#_M1026_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_206 VPB N_A_2668_265#_c_1133_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.605
+ $Y2=0.425
cc_207 VPB N_A_2668_265#_c_1130_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_A_2668_265#_c_1131_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_S[6]_c_1187_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_210 VPB N_S[7]_c_1231_n 0.0280248f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_211 VPB N_A_3017_47#_M1045_g 0.0269712f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.19
cc_212 VPB N_A_3017_47#_c_1280_n 0.0075635f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.19
cc_213 VPB N_A_3017_47#_c_1276_n 0.0108568f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_A_3017_47#_c_1277_n 0.0306622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_D[7]_c_1330_n 0.0335483f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_216 VPB N_D[7]_c_1333_n 0.00458905f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_VPWR_c_1359_n 0.0103693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_VPWR_c_1360_n 0.0425009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_VPWR_c_1361_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB N_VPWR_c_1362_n 4.89801e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB N_VPWR_c_1363_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 VPB N_VPWR_c_1364_n 4.89801e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_223 VPB N_VPWR_c_1365_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_224 VPB N_VPWR_c_1366_n 4.89801e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_225 VPB N_VPWR_c_1367_n 0.0150686f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_226 VPB N_VPWR_c_1368_n 0.0103693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_227 VPB N_VPWR_c_1369_n 0.0425009f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_228 VPB N_VPWR_c_1370_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_229 VPB N_VPWR_c_1371_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_230 VPB N_VPWR_c_1372_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_231 VPB N_VPWR_c_1373_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_232 VPB N_VPWR_c_1374_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_233 VPB N_VPWR_c_1375_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_234 VPB N_VPWR_c_1376_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_235 VPB N_VPWR_c_1377_n 0.00632158f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_236 VPB VPWR 0.0724189f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_237 VPB N_VPWR_c_1379_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_238 VPB N_VPWR_c_1380_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_239 VPB N_VPWR_c_1381_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_240 VPB N_VPWR_c_1382_n 0.0461673f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_241 VPB N_VPWR_c_1383_n 0.0051677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_242 VPB N_VPWR_c_1384_n 0.0051677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_243 VPB N_VPWR_c_1385_n 0.0051677f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_244 VPB N_Z_c_1624_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_245 VPB N_Z_c_1649_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_246 VPB N_Z_c_1650_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_247 VPB N_Z_c_1628_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_248 VPB N_Z_c_1629_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_249 VPB N_Z_c_1653_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_250 VPB N_Z_c_1654_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_251 VPB N_Z_c_1633_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_252 VPB N_Z_c_1634_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_253 VPB N_Z_c_1657_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_254 VPB N_Z_c_1658_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_255 VPB N_Z_c_1638_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_256 VPB N_Z_c_1639_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_257 VPB N_Z_c_1661_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_258 VPB N_Z_c_1662_n 0.00457032f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_259 VPB N_Z_c_1643_n 0.00365513f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_260 VPB N_Z_c_1664_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_261 VPB N_Z_c_1665_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_262 VPB N_Z_c_1666_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_263 VPB N_Z_c_1667_n 0.00809084f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_264 VPB N_Z_c_1668_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_265 VPB N_Z_c_1669_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_266 VPB N_Z_c_1670_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_267 VPB N_Z_c_1671_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_268 VPB N_Z_c_1672_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_269 VPB N_Z_c_1673_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_270 VPB N_Z_c_1674_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_271 VPB N_Z_c_1675_n 0.00133145f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_272 N_D[0]_c_273_n N_A_184_265#_M1019_g 0.0381613f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_273 N_D[0]_c_273_n N_A_184_265#_c_303_n 0.00712672f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_274 N_D[0]_c_272_n N_S[0]_c_356_n 0.0286599f $X=0.47 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_275 N_D[0]_c_274_n N_S[0]_c_356_n 0.00289497f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_276 N_D[0]_c_273_n N_VPWR_c_1360_n 0.0245615f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_277 N_D[0]_c_275_n N_VPWR_c_1360_n 0.00471543f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_278 N_D[0]_c_273_n N_VPWR_c_1370_n 0.00622633f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_279 N_D[0]_c_273_n VPWR 0.0106352f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_280 N_D[0]_c_273_n N_Z_c_1624_n 0.00605747f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_281 N_D[0]_c_274_n N_Z_c_1624_n 0.00376465f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_282 N_D[0]_c_275_n N_Z_c_1624_n 0.0216525f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_283 N_D[0]_c_274_n N_Z_c_1625_n 0.0128881f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_284 N_D[0]_c_274_n N_Z_c_1626_n 0.00686805f $X=0.645 $Y=1.055 $X2=0 $Y2=0
cc_285 N_D[0]_c_273_n N_Z_c_1649_n 0.00145364f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_286 N_D[0]_c_272_n N_VGND_c_2110_n 0.00487865f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_287 N_D[0]_c_275_n N_VGND_c_2110_n 0.00222881f $X=0.645 $Y=1.19 $X2=0 $Y2=0
cc_288 N_D[0]_c_272_n N_VGND_c_2120_n 0.00585385f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_289 D[0] N_VGND_c_2120_n 0.00842546f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_290 N_D[0]_c_272_n VGND 0.011617f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_291 D[0] VGND 0.00942277f $X=0.605 $Y=0.425 $X2=0 $Y2=0
cc_292 N_D[0]_c_274_n A_109_47# 0.00426617f $X=0.645 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_293 D[0] A_109_47# 0.00894235f $X=0.605 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_294 N_A_184_265#_c_300_n N_S[0]_c_357_n 0.00827389f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_295 N_A_184_265#_c_301_n N_S[0]_c_357_n 0.0164662f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_296 N_A_184_265#_c_302_n N_S[0]_c_357_n 0.00928634f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_297 N_A_184_265#_c_303_n N_S[0]_c_357_n 0.0184911f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_298 N_A_184_265#_c_303_n N_S[0]_c_358_n 0.00820745f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_299 N_A_184_265#_c_301_n N_S[0]_c_359_n 0.0012443f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_300 N_A_184_265#_c_305_n N_S[0]_c_359_n 0.00903826f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_301 N_A_184_265#_c_302_n N_S[0]_c_359_n 0.00767015f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_302 N_A_184_265#_c_303_n N_S[0]_c_359_n 0.00659591f $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_303 N_A_184_265#_c_301_n N_S[0]_c_360_n 0.00219336f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_304 N_A_184_265#_c_300_n N_S[0]_c_361_n 0.00603567f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_305 N_A_184_265#_c_301_n N_S[0]_c_361_n 0.0178233f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_306 N_A_184_265#_c_302_n N_S[0]_c_361_n 0.0214702f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_307 N_A_184_265#_c_303_n N_S[0]_c_361_n 2.59957e-19 $X=1.02 $Y=1.34 $X2=0
+ $Y2=0
cc_308 N_A_184_265#_M1019_g N_VPWR_c_1360_n 0.00298082f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_309 N_A_184_265#_c_305_n N_VPWR_c_1361_n 0.0292866f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_310 N_A_184_265#_c_302_n N_VPWR_c_1361_n 0.00688579f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_311 N_A_184_265#_M1019_g N_VPWR_c_1370_n 0.00522699f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_312 N_A_184_265#_c_305_n N_VPWR_c_1370_n 0.0210596f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_313 N_A_184_265#_M1023_s VPWR 0.00179197f $X=1.65 $Y=1.485 $X2=0 $Y2=0
cc_314 N_A_184_265#_M1019_g VPWR 0.00828927f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_315 N_A_184_265#_c_305_n VPWR 0.00594162f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_316 N_A_184_265#_M1019_g N_Z_c_1624_n 0.00862328f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_317 N_A_184_265#_c_301_n N_Z_c_1624_n 0.00719188f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_318 N_A_184_265#_c_305_n N_Z_c_1624_n 0.00378484f $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_319 N_A_184_265#_c_302_n N_Z_c_1624_n 0.0304368f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_320 N_A_184_265#_c_303_n N_Z_c_1624_n 0.00814206f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_321 N_A_184_265#_c_301_n N_Z_c_1625_n 0.0124144f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_322 N_A_184_265#_c_302_n N_Z_c_1625_n 0.00398133f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_323 N_A_184_265#_c_303_n N_Z_c_1625_n 0.00349316f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_324 N_A_184_265#_c_300_n N_Z_c_1626_n 0.0259454f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_325 N_A_184_265#_c_301_n N_Z_c_1626_n 0.00611965f $X=1.545 $Y=1.175 $X2=0
+ $Y2=0
cc_326 N_A_184_265#_M1019_g N_Z_c_1649_n 0.00988241f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_327 N_A_184_265#_c_305_n N_Z_c_1649_n 0.0369227f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_328 N_A_184_265#_c_305_n N_Z_c_1664_n 0.0291787f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_329 N_A_184_265#_c_302_n N_Z_c_1664_n 0.0126642f $X=1.775 $Y=1.63 $X2=0 $Y2=0
cc_330 N_A_184_265#_M1019_g N_Z_c_1696_n 0.00289142f $X=1.02 $Y=2.075 $X2=0
+ $Y2=0
cc_331 N_A_184_265#_c_305_n N_Z_c_1696_n 6.03258e-19 $X=1.775 $Y=2.31 $X2=0
+ $Y2=0
cc_332 N_A_184_265#_c_302_n N_Z_c_1696_n 4.25753e-19 $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_333 N_A_184_265#_M1019_g N_Z_c_1668_n 0.0105217f $X=1.02 $Y=2.075 $X2=0 $Y2=0
cc_334 N_A_184_265#_c_305_n N_Z_c_1668_n 0.0139746f $X=1.775 $Y=2.31 $X2=0 $Y2=0
cc_335 N_A_184_265#_c_302_n N_Z_c_1668_n 0.00749676f $X=1.775 $Y=1.63 $X2=0
+ $Y2=0
cc_336 N_A_184_265#_c_303_n N_Z_c_1668_n 0.00449162f $X=1.02 $Y=1.34 $X2=0 $Y2=0
cc_337 N_A_184_265#_c_300_n N_VGND_c_2120_n 0.015238f $X=1.545 $Y=0.755 $X2=0
+ $Y2=0
cc_338 N_A_184_265#_M1029_s VGND 0.00358139f $X=1.65 $Y=0.235 $X2=0 $Y2=0
cc_339 N_A_184_265#_c_300_n VGND 0.0150148f $X=1.545 $Y=0.755 $X2=0 $Y2=0
cc_340 N_S[0]_c_359_n N_S[1]_c_403_n 0.0578733f $X=2.01 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_341 N_S[0]_c_361_n N_S[1]_c_403_n 0.00112057f $X=1.975 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_342 N_S[0]_c_360_n N_S[1]_c_404_n 0.0091402f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_343 N_S[0]_c_359_n N_S[1]_c_407_n 0.00112057f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_344 N_S[0]_c_361_n N_S[1]_c_407_n 0.0277403f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_345 N_S[0]_c_359_n N_VPWR_c_1361_n 0.00965725f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_346 N_S[0]_c_361_n N_VPWR_c_1361_n 0.00587376f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_347 N_S[0]_c_359_n N_VPWR_c_1370_n 0.00673617f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_348 N_S[0]_c_359_n VPWR 0.00871384f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_349 N_S[0]_c_358_n N_Z_c_1624_n 7.46972e-19 $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_350 N_S[0]_c_357_n N_Z_c_1625_n 0.00806549f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_351 N_S[0]_c_358_n N_Z_c_1625_n 0.00605736f $X=1.02 $Y=0.905 $X2=0 $Y2=0
cc_352 N_S[0]_c_356_n N_Z_c_1626_n 0.00316445f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_353 N_S[0]_c_357_n N_Z_c_1626_n 0.00501353f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_354 N_S[0]_c_359_n N_Z_c_1664_n 0.0062071f $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_355 N_S[0]_c_361_n N_Z_c_1664_n 0.00659242f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_356 N_S[0]_c_360_n N_VGND_c_2111_n 0.00570474f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_357 N_S[0]_c_361_n N_VGND_c_2111_n 0.00391126f $X=1.975 $Y=1.03 $X2=0 $Y2=0
cc_358 N_S[0]_c_356_n N_VGND_c_2120_n 0.00585385f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_359 N_S[0]_c_360_n N_VGND_c_2120_n 0.00585385f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_360 N_S[0]_c_356_n VGND 0.00880034f $X=0.945 $Y=0.83 $X2=0 $Y2=0
cc_361 N_S[0]_c_357_n VGND 0.00349917f $X=1.84 $Y=0.905 $X2=0 $Y2=0
cc_362 N_S[0]_c_359_n VGND 6.15795e-19 $X=2.01 $Y=1.41 $X2=0 $Y2=0
cc_363 N_S[0]_c_360_n VGND 0.0124506f $X=2.01 $Y=0.83 $X2=0 $Y2=0
cc_364 N_S[1]_c_403_n N_A_533_47#_c_452_n 0.00903826f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_365 N_S[1]_c_403_n N_A_533_47#_c_447_n 0.0012443f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_366 N_S[1]_c_404_n N_A_533_47#_c_447_n 0.00219336f $X=2.59 $Y=0.83 $X2=0
+ $Y2=0
cc_367 N_S[1]_c_405_n N_A_533_47#_c_447_n 0.0164662f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_368 N_S[1]_c_407_n N_A_533_47#_c_447_n 0.0178233f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_369 N_S[1]_c_403_n N_A_533_47#_c_448_n 0.00767015f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_370 N_S[1]_c_405_n N_A_533_47#_c_448_n 0.00928634f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_371 N_S[1]_c_407_n N_A_533_47#_c_448_n 0.0214702f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_372 N_S[1]_c_403_n N_A_533_47#_c_449_n 0.00659591f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_373 N_S[1]_c_405_n N_A_533_47#_c_449_n 0.0266986f $X=3.58 $Y=0.905 $X2=0
+ $Y2=0
cc_374 N_S[1]_c_407_n N_A_533_47#_c_449_n 2.59957e-19 $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_375 N_S[1]_c_403_n N_A_533_47#_c_450_n 0.00827389f $X=2.59 $Y=1.41 $X2=0
+ $Y2=0
cc_376 N_S[1]_c_407_n N_A_533_47#_c_450_n 0.00603567f $X=2.625 $Y=1.03 $X2=0
+ $Y2=0
cc_377 N_S[1]_c_406_n N_D[1]_c_503_n 0.0286599f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_378 N_S[1]_c_406_n N_D[1]_c_504_n 0.00289497f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_379 N_S[1]_c_403_n N_VPWR_c_1361_n 0.00965725f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_380 N_S[1]_c_407_n N_VPWR_c_1361_n 0.00587376f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_381 N_S[1]_c_403_n VPWR 0.00871384f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_382 N_S[1]_c_403_n N_VPWR_c_1379_n 0.00673617f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_383 N_S[1]_c_405_n N_Z_c_1627_n 0.00501353f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_384 N_S[1]_c_406_n N_Z_c_1627_n 0.00316445f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_385 N_S[1]_c_405_n N_Z_c_1628_n 7.46972e-19 $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_386 N_S[1]_c_405_n N_Z_c_1644_n 0.0141229f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_387 N_S[1]_c_403_n N_Z_c_1664_n 0.0062071f $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_388 N_S[1]_c_407_n N_Z_c_1664_n 0.00659242f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_389 N_S[1]_c_404_n N_VGND_c_2111_n 0.00570474f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_390 N_S[1]_c_407_n N_VGND_c_2111_n 0.00391126f $X=2.625 $Y=1.03 $X2=0 $Y2=0
cc_391 N_S[1]_c_403_n VGND 6.15795e-19 $X=2.59 $Y=1.41 $X2=0 $Y2=0
cc_392 N_S[1]_c_404_n VGND 0.0124506f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_393 N_S[1]_c_405_n VGND 0.00349917f $X=3.58 $Y=0.905 $X2=0 $Y2=0
cc_394 N_S[1]_c_406_n VGND 0.00880034f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_395 N_S[1]_c_404_n N_VGND_c_2129_n 0.00585385f $X=2.59 $Y=0.83 $X2=0 $Y2=0
cc_396 N_S[1]_c_406_n N_VGND_c_2129_n 0.00585385f $X=3.655 $Y=0.83 $X2=0 $Y2=0
cc_397 N_A_533_47#_M1009_g N_D[1]_c_502_n 0.0388862f $X=3.58 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_398 N_A_533_47#_c_449_n N_D[1]_c_502_n 0.00712672f $X=3.275 $Y=1.34 $X2=-0.19
+ $Y2=-0.24
cc_399 N_A_533_47#_c_452_n N_VPWR_c_1361_n 0.0292866f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_400 N_A_533_47#_c_448_n N_VPWR_c_1361_n 0.00688579f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_401 N_A_533_47#_M1009_g N_VPWR_c_1362_n 0.0030953f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_402 N_A_533_47#_M1020_d VPWR 0.00179197f $X=2.68 $Y=1.485 $X2=0 $Y2=0
cc_403 N_A_533_47#_M1009_g VPWR 0.00809563f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_404 N_A_533_47#_c_452_n VPWR 0.00594162f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_405 N_A_533_47#_M1009_g N_VPWR_c_1379_n 0.00522699f $X=3.58 $Y=2.075 $X2=0
+ $Y2=0
cc_406 N_A_533_47#_c_452_n N_VPWR_c_1379_n 0.0210596f $X=2.825 $Y=2.31 $X2=0
+ $Y2=0
cc_407 N_A_533_47#_M1009_g N_Z_c_1650_n 0.00988241f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_408 N_A_533_47#_c_452_n N_Z_c_1650_n 0.0369227f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_409 N_A_533_47#_c_447_n N_Z_c_1627_n 0.00611965f $X=3.055 $Y=1.175 $X2=0
+ $Y2=0
cc_410 N_A_533_47#_c_450_n N_Z_c_1627_n 0.0259454f $X=2.825 $Y=0.495 $X2=0 $Y2=0
cc_411 N_A_533_47#_M1009_g N_Z_c_1628_n 0.00862328f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_412 N_A_533_47#_c_452_n N_Z_c_1628_n 0.00378484f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_413 N_A_533_47#_c_447_n N_Z_c_1628_n 0.00719188f $X=3.055 $Y=1.175 $X2=0
+ $Y2=0
cc_414 N_A_533_47#_c_448_n N_Z_c_1628_n 0.0304368f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_415 N_A_533_47#_c_449_n N_Z_c_1628_n 0.00814206f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_416 N_A_533_47#_c_447_n N_Z_c_1644_n 0.0124144f $X=3.055 $Y=1.175 $X2=0 $Y2=0
cc_417 N_A_533_47#_c_448_n N_Z_c_1644_n 0.00398133f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_418 N_A_533_47#_c_449_n N_Z_c_1644_n 0.00349316f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_419 N_A_533_47#_c_452_n N_Z_c_1664_n 0.0291787f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_420 N_A_533_47#_c_448_n N_Z_c_1664_n 0.0126642f $X=3.055 $Y=1.405 $X2=0 $Y2=0
cc_421 N_A_533_47#_M1009_g N_Z_c_1730_n 0.00289142f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_422 N_A_533_47#_c_452_n N_Z_c_1730_n 6.03258e-19 $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_423 N_A_533_47#_c_448_n N_Z_c_1730_n 4.25753e-19 $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_424 N_A_533_47#_M1009_g N_Z_c_1669_n 0.0105217f $X=3.58 $Y=2.075 $X2=0 $Y2=0
cc_425 N_A_533_47#_c_452_n N_Z_c_1669_n 0.0139746f $X=2.825 $Y=2.31 $X2=0 $Y2=0
cc_426 N_A_533_47#_c_448_n N_Z_c_1669_n 0.00749676f $X=3.055 $Y=1.405 $X2=0
+ $Y2=0
cc_427 N_A_533_47#_c_449_n N_Z_c_1669_n 0.00449162f $X=3.275 $Y=1.34 $X2=0 $Y2=0
cc_428 N_A_533_47#_M1028_d VGND 0.00358139f $X=2.665 $Y=0.235 $X2=0 $Y2=0
cc_429 N_A_533_47#_c_450_n VGND 0.0150148f $X=2.825 $Y=0.495 $X2=0 $Y2=0
cc_430 N_A_533_47#_c_450_n N_VGND_c_2129_n 0.015238f $X=2.825 $Y=0.495 $X2=0
+ $Y2=0
cc_431 N_D[1]_c_503_n N_D[2]_c_539_n 0.00915308f $X=4.13 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_432 N_D[1]_c_502_n N_D[2]_c_540_n 0.0270908f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_433 N_D[1]_c_505_n N_D[2]_c_540_n 9.4377e-19 $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_434 N_D[1]_c_504_n N_D[2]_c_541_n 0.00442615f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_435 N_D[1]_c_502_n N_D[2]_c_542_n 9.4377e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_436 N_D[1]_c_505_n N_D[2]_c_542_n 0.0199139f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_437 N_D[1]_c_502_n N_VPWR_c_1362_n 0.0231278f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_438 N_D[1]_c_505_n N_VPWR_c_1362_n 0.0044581f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_439 N_D[1]_c_502_n VPWR 0.00594051f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_440 N_D[1]_c_502_n N_VPWR_c_1379_n 0.00622633f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_441 N_D[1]_c_502_n N_Z_c_1650_n 0.00145364f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_442 N_D[1]_c_504_n N_Z_c_1627_n 0.00686805f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_443 N_D[1]_c_502_n N_Z_c_1628_n 0.00605747f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_444 N_D[1]_c_504_n N_Z_c_1628_n 0.00376465f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_445 N_D[1]_c_505_n N_Z_c_1628_n 0.0216525f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_446 N_D[1]_c_504_n N_Z_c_1644_n 0.0128881f $X=3.955 $Y=1.055 $X2=0 $Y2=0
cc_447 N_D[1]_c_502_n N_Z_c_1743_n 0.00719456f $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_448 N_D[1]_c_505_n N_Z_c_1743_n 0.00989895f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_449 N_D[1]_c_502_n N_Z_c_1669_n 8.42164e-19 $X=4.105 $Y=1.41 $X2=0 $Y2=0
cc_450 N_D[1]_c_503_n N_VGND_c_2112_n 0.00322791f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_451 N_D[1]_c_505_n N_VGND_c_2112_n 0.00222881f $X=4.1 $Y=1.16 $X2=0 $Y2=0
cc_452 N_D[1]_c_503_n VGND 0.0108306f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_453 N_D[1]_c_534_p VGND 0.00942277f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_454 N_D[1]_c_503_n N_VGND_c_2129_n 0.00585385f $X=4.13 $Y=0.995 $X2=0 $Y2=0
cc_455 N_D[1]_c_534_p N_VGND_c_2129_n 0.00842546f $X=3.955 $Y=0.51 $X2=0 $Y2=0
cc_456 N_D[1]_c_504_n A_746_47# 0.00426617f $X=3.955 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_457 N_D[1]_c_534_p A_746_47# 0.00894235f $X=3.955 $Y=0.51 $X2=-0.19 $Y2=-0.24
cc_458 N_D[2]_c_540_n N_A_1012_265#_M1022_g 0.0388862f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_459 N_D[2]_c_540_n N_A_1012_265#_c_579_n 0.00712672f $X=4.635 $Y=1.41 $X2=0
+ $Y2=0
cc_460 N_D[2]_c_539_n N_S[2]_c_632_n 0.0286599f $X=4.61 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_461 N_D[2]_c_541_n N_S[2]_c_632_n 0.00289497f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_462 N_D[2]_c_540_n N_VPWR_c_1362_n 0.0231278f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_463 N_D[2]_c_542_n N_VPWR_c_1362_n 0.0044581f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_464 N_D[2]_c_540_n N_VPWR_c_1372_n 0.00622633f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_465 N_D[2]_c_540_n VPWR 0.00594051f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_466 N_D[2]_c_540_n N_Z_c_1629_n 0.00605747f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_467 N_D[2]_c_541_n N_Z_c_1629_n 0.00376465f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_468 N_D[2]_c_542_n N_Z_c_1629_n 0.0216525f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_469 N_D[2]_c_541_n N_Z_c_1630_n 0.0128881f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_470 N_D[2]_c_541_n N_Z_c_1631_n 0.00686805f $X=4.785 $Y=1.055 $X2=0 $Y2=0
cc_471 N_D[2]_c_540_n N_Z_c_1653_n 0.00145364f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_472 N_D[2]_c_540_n N_Z_c_1743_n 0.00719456f $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_473 N_D[2]_c_542_n N_Z_c_1743_n 0.00989895f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_474 N_D[2]_c_540_n N_Z_c_1670_n 8.42164e-19 $X=4.635 $Y=1.41 $X2=0 $Y2=0
cc_475 N_D[2]_c_539_n N_VGND_c_2112_n 0.00322791f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_476 N_D[2]_c_542_n N_VGND_c_2112_n 0.00222881f $X=4.785 $Y=1.19 $X2=0 $Y2=0
cc_477 N_D[2]_c_539_n N_VGND_c_2122_n 0.00585385f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_478 D[2] N_VGND_c_2122_n 0.00842546f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_479 N_D[2]_c_539_n VGND 0.0108306f $X=4.61 $Y=0.995 $X2=0 $Y2=0
cc_480 D[2] VGND 0.00942277f $X=4.745 $Y=0.425 $X2=0 $Y2=0
cc_481 N_D[2]_c_541_n A_937_47# 0.00426617f $X=4.785 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_482 D[2] A_937_47# 0.00894235f $X=4.745 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_483 N_A_1012_265#_c_576_n N_S[2]_c_633_n 0.00827389f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_484 N_A_1012_265#_c_577_n N_S[2]_c_633_n 0.0164662f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_485 N_A_1012_265#_c_578_n N_S[2]_c_633_n 0.00928634f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_486 N_A_1012_265#_c_579_n N_S[2]_c_633_n 0.0184911f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_487 N_A_1012_265#_c_579_n N_S[2]_c_634_n 0.00820745f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_488 N_A_1012_265#_c_577_n N_S[2]_c_635_n 0.0012443f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_489 N_A_1012_265#_c_581_n N_S[2]_c_635_n 0.00903826f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_490 N_A_1012_265#_c_578_n N_S[2]_c_635_n 0.00767015f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_491 N_A_1012_265#_c_579_n N_S[2]_c_635_n 0.00659591f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_492 N_A_1012_265#_c_577_n N_S[2]_c_636_n 0.00219336f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_493 N_A_1012_265#_c_576_n N_S[2]_c_637_n 0.00603567f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_494 N_A_1012_265#_c_577_n N_S[2]_c_637_n 0.0178233f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_495 N_A_1012_265#_c_578_n N_S[2]_c_637_n 0.0214702f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_496 N_A_1012_265#_c_579_n N_S[2]_c_637_n 2.59957e-19 $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_497 N_A_1012_265#_M1022_g N_VPWR_c_1362_n 0.0030953f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_498 N_A_1012_265#_c_581_n N_VPWR_c_1363_n 0.0292866f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_499 N_A_1012_265#_c_578_n N_VPWR_c_1363_n 0.00688579f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_500 N_A_1012_265#_M1022_g N_VPWR_c_1372_n 0.00522699f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_501 N_A_1012_265#_c_581_n N_VPWR_c_1372_n 0.0210596f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_502 N_A_1012_265#_M1025_s VPWR 0.00179197f $X=5.79 $Y=1.485 $X2=0 $Y2=0
cc_503 N_A_1012_265#_M1022_g VPWR 0.00809563f $X=5.16 $Y=2.075 $X2=0 $Y2=0
cc_504 N_A_1012_265#_c_581_n VPWR 0.00594162f $X=5.915 $Y=2.31 $X2=0 $Y2=0
cc_505 N_A_1012_265#_M1022_g N_Z_c_1629_n 0.00862328f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_506 N_A_1012_265#_c_577_n N_Z_c_1629_n 0.00719188f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_507 N_A_1012_265#_c_581_n N_Z_c_1629_n 0.00378484f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_508 N_A_1012_265#_c_578_n N_Z_c_1629_n 0.0304368f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_509 N_A_1012_265#_c_579_n N_Z_c_1629_n 0.00814206f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_510 N_A_1012_265#_c_577_n N_Z_c_1630_n 0.0124144f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_511 N_A_1012_265#_c_578_n N_Z_c_1630_n 0.00398133f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_512 N_A_1012_265#_c_579_n N_Z_c_1630_n 0.00349316f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_513 N_A_1012_265#_c_576_n N_Z_c_1631_n 0.0259454f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_514 N_A_1012_265#_c_577_n N_Z_c_1631_n 0.00611965f $X=5.685 $Y=1.175 $X2=0
+ $Y2=0
cc_515 N_A_1012_265#_M1022_g N_Z_c_1653_n 0.00988241f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_516 N_A_1012_265#_c_581_n N_Z_c_1653_n 0.0369227f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_517 N_A_1012_265#_c_581_n N_Z_c_1665_n 0.0291787f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_518 N_A_1012_265#_c_578_n N_Z_c_1665_n 0.0126642f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_519 N_A_1012_265#_M1022_g N_Z_c_1769_n 0.00289142f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_520 N_A_1012_265#_c_581_n N_Z_c_1769_n 6.03258e-19 $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_521 N_A_1012_265#_c_578_n N_Z_c_1769_n 4.25753e-19 $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_522 N_A_1012_265#_M1022_g N_Z_c_1670_n 0.0105217f $X=5.16 $Y=2.075 $X2=0
+ $Y2=0
cc_523 N_A_1012_265#_c_581_n N_Z_c_1670_n 0.0139746f $X=5.915 $Y=2.31 $X2=0
+ $Y2=0
cc_524 N_A_1012_265#_c_578_n N_Z_c_1670_n 0.00749676f $X=5.915 $Y=1.63 $X2=0
+ $Y2=0
cc_525 N_A_1012_265#_c_579_n N_Z_c_1670_n 0.00449162f $X=5.16 $Y=1.34 $X2=0
+ $Y2=0
cc_526 N_A_1012_265#_c_576_n N_VGND_c_2122_n 0.015238f $X=5.685 $Y=0.755 $X2=0
+ $Y2=0
cc_527 N_A_1012_265#_M1042_s VGND 0.00358139f $X=5.79 $Y=0.235 $X2=0 $Y2=0
cc_528 N_A_1012_265#_c_576_n VGND 0.0150148f $X=5.685 $Y=0.755 $X2=0 $Y2=0
cc_529 N_S[2]_c_635_n N_S[3]_c_679_n 0.0578733f $X=6.15 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_530 N_S[2]_c_637_n N_S[3]_c_679_n 0.00112057f $X=6.115 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_531 N_S[2]_c_636_n N_S[3]_c_680_n 0.0091402f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_532 N_S[2]_c_635_n N_S[3]_c_683_n 0.00112057f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_533 N_S[2]_c_637_n N_S[3]_c_683_n 0.0277403f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_534 N_S[2]_c_635_n N_VPWR_c_1363_n 0.00965725f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_535 N_S[2]_c_637_n N_VPWR_c_1363_n 0.00587376f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_536 N_S[2]_c_635_n N_VPWR_c_1372_n 0.00673617f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_537 N_S[2]_c_635_n VPWR 0.00871384f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_538 N_S[2]_c_634_n N_Z_c_1629_n 7.46972e-19 $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_539 N_S[2]_c_633_n N_Z_c_1630_n 0.00806549f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_540 N_S[2]_c_634_n N_Z_c_1630_n 0.00605736f $X=5.16 $Y=0.905 $X2=0 $Y2=0
cc_541 N_S[2]_c_632_n N_Z_c_1631_n 0.00316445f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_542 N_S[2]_c_633_n N_Z_c_1631_n 0.00501353f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_543 N_S[2]_c_635_n N_Z_c_1665_n 0.0062071f $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_544 N_S[2]_c_637_n N_Z_c_1665_n 0.00659242f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_545 N_S[2]_c_636_n N_VGND_c_2113_n 0.00570474f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_546 N_S[2]_c_637_n N_VGND_c_2113_n 0.00391126f $X=6.115 $Y=1.03 $X2=0 $Y2=0
cc_547 N_S[2]_c_632_n N_VGND_c_2122_n 0.00585385f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_548 N_S[2]_c_636_n N_VGND_c_2122_n 0.00585385f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_549 N_S[2]_c_632_n VGND 0.00880034f $X=5.085 $Y=0.83 $X2=0 $Y2=0
cc_550 N_S[2]_c_633_n VGND 0.00349917f $X=5.98 $Y=0.905 $X2=0 $Y2=0
cc_551 N_S[2]_c_635_n VGND 6.15795e-19 $X=6.15 $Y=1.41 $X2=0 $Y2=0
cc_552 N_S[2]_c_636_n VGND 0.0124506f $X=6.15 $Y=0.83 $X2=0 $Y2=0
cc_553 N_S[3]_c_679_n N_A_1361_47#_c_728_n 0.00903826f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_554 N_S[3]_c_679_n N_A_1361_47#_c_723_n 0.0012443f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_555 N_S[3]_c_680_n N_A_1361_47#_c_723_n 0.00219336f $X=6.73 $Y=0.83 $X2=0
+ $Y2=0
cc_556 N_S[3]_c_681_n N_A_1361_47#_c_723_n 0.0164662f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_557 N_S[3]_c_683_n N_A_1361_47#_c_723_n 0.0178233f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_558 N_S[3]_c_679_n N_A_1361_47#_c_724_n 0.00767015f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_559 N_S[3]_c_681_n N_A_1361_47#_c_724_n 0.00928634f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_560 N_S[3]_c_683_n N_A_1361_47#_c_724_n 0.0214702f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_561 N_S[3]_c_679_n N_A_1361_47#_c_725_n 0.00659591f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_562 N_S[3]_c_681_n N_A_1361_47#_c_725_n 0.0266986f $X=7.72 $Y=0.905 $X2=0
+ $Y2=0
cc_563 N_S[3]_c_683_n N_A_1361_47#_c_725_n 2.59957e-19 $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_564 N_S[3]_c_679_n N_A_1361_47#_c_726_n 0.00827389f $X=6.73 $Y=1.41 $X2=0
+ $Y2=0
cc_565 N_S[3]_c_683_n N_A_1361_47#_c_726_n 0.00603567f $X=6.765 $Y=1.03 $X2=0
+ $Y2=0
cc_566 N_S[3]_c_682_n N_D[3]_c_779_n 0.0286599f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_567 N_S[3]_c_682_n N_D[3]_c_780_n 0.00289497f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_568 N_S[3]_c_679_n N_VPWR_c_1363_n 0.00965725f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_569 N_S[3]_c_683_n N_VPWR_c_1363_n 0.00587376f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_570 N_S[3]_c_679_n VPWR 0.00871384f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_571 N_S[3]_c_679_n N_VPWR_c_1380_n 0.00673617f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_572 N_S[3]_c_681_n N_Z_c_1632_n 0.00501353f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_573 N_S[3]_c_682_n N_Z_c_1632_n 0.00316445f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_574 N_S[3]_c_681_n N_Z_c_1633_n 7.46972e-19 $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_575 N_S[3]_c_681_n N_Z_c_1645_n 0.0141229f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_576 N_S[3]_c_679_n N_Z_c_1665_n 0.0062071f $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_577 N_S[3]_c_683_n N_Z_c_1665_n 0.00659242f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_578 N_S[3]_c_680_n N_VGND_c_2113_n 0.00570474f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_579 N_S[3]_c_683_n N_VGND_c_2113_n 0.00391126f $X=6.765 $Y=1.03 $X2=0 $Y2=0
cc_580 N_S[3]_c_679_n VGND 6.15795e-19 $X=6.73 $Y=1.41 $X2=0 $Y2=0
cc_581 N_S[3]_c_680_n VGND 0.0124506f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_582 N_S[3]_c_681_n VGND 0.00349917f $X=7.72 $Y=0.905 $X2=0 $Y2=0
cc_583 N_S[3]_c_682_n VGND 0.00880034f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_584 N_S[3]_c_680_n N_VGND_c_2130_n 0.00585385f $X=6.73 $Y=0.83 $X2=0 $Y2=0
cc_585 N_S[3]_c_682_n N_VGND_c_2130_n 0.00585385f $X=7.795 $Y=0.83 $X2=0 $Y2=0
cc_586 N_A_1361_47#_M1013_g N_D[3]_c_778_n 0.0388862f $X=7.72 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_587 N_A_1361_47#_c_725_n N_D[3]_c_778_n 0.00712672f $X=7.415 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_588 N_A_1361_47#_c_728_n N_VPWR_c_1363_n 0.0292866f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_589 N_A_1361_47#_c_724_n N_VPWR_c_1363_n 0.00688579f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_590 N_A_1361_47#_M1013_g N_VPWR_c_1364_n 0.0030953f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_591 N_A_1361_47#_M1005_d VPWR 0.00179197f $X=6.82 $Y=1.485 $X2=0 $Y2=0
cc_592 N_A_1361_47#_M1013_g VPWR 0.00809563f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_593 N_A_1361_47#_c_728_n VPWR 0.00594162f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_594 N_A_1361_47#_M1013_g N_VPWR_c_1380_n 0.00522699f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_595 N_A_1361_47#_c_728_n N_VPWR_c_1380_n 0.0210596f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_596 N_A_1361_47#_M1013_g N_Z_c_1654_n 0.00988241f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_597 N_A_1361_47#_c_728_n N_Z_c_1654_n 0.0369227f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_598 N_A_1361_47#_c_723_n N_Z_c_1632_n 0.00611965f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_599 N_A_1361_47#_c_726_n N_Z_c_1632_n 0.0259454f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_600 N_A_1361_47#_M1013_g N_Z_c_1633_n 0.00862328f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_601 N_A_1361_47#_c_728_n N_Z_c_1633_n 0.00378484f $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_602 N_A_1361_47#_c_723_n N_Z_c_1633_n 0.00719188f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_603 N_A_1361_47#_c_724_n N_Z_c_1633_n 0.0304368f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_604 N_A_1361_47#_c_725_n N_Z_c_1633_n 0.00814206f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_605 N_A_1361_47#_c_723_n N_Z_c_1645_n 0.0124144f $X=7.195 $Y=1.175 $X2=0
+ $Y2=0
cc_606 N_A_1361_47#_c_724_n N_Z_c_1645_n 0.00398133f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_607 N_A_1361_47#_c_725_n N_Z_c_1645_n 0.00349316f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_608 N_A_1361_47#_c_728_n N_Z_c_1665_n 0.0291787f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_609 N_A_1361_47#_c_724_n N_Z_c_1665_n 0.0126642f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_610 N_A_1361_47#_M1013_g N_Z_c_1803_n 0.00289142f $X=7.72 $Y=2.075 $X2=0
+ $Y2=0
cc_611 N_A_1361_47#_c_728_n N_Z_c_1803_n 6.03258e-19 $X=6.965 $Y=2.31 $X2=0
+ $Y2=0
cc_612 N_A_1361_47#_c_724_n N_Z_c_1803_n 4.25753e-19 $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_613 N_A_1361_47#_M1013_g N_Z_c_1671_n 0.0105217f $X=7.72 $Y=2.075 $X2=0 $Y2=0
cc_614 N_A_1361_47#_c_728_n N_Z_c_1671_n 0.0139746f $X=6.965 $Y=2.31 $X2=0 $Y2=0
cc_615 N_A_1361_47#_c_724_n N_Z_c_1671_n 0.00749676f $X=7.195 $Y=1.405 $X2=0
+ $Y2=0
cc_616 N_A_1361_47#_c_725_n N_Z_c_1671_n 0.00449162f $X=7.415 $Y=1.34 $X2=0
+ $Y2=0
cc_617 N_A_1361_47#_M1027_d VGND 0.00358139f $X=6.805 $Y=0.235 $X2=0 $Y2=0
cc_618 N_A_1361_47#_c_726_n VGND 0.0150148f $X=6.965 $Y=0.495 $X2=0 $Y2=0
cc_619 N_A_1361_47#_c_726_n N_VGND_c_2130_n 0.015238f $X=6.965 $Y=0.495 $X2=0
+ $Y2=0
cc_620 N_D[3]_c_779_n N_D[4]_c_815_n 0.00915308f $X=8.27 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_621 N_D[3]_c_778_n N_D[4]_c_816_n 0.0270908f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_622 N_D[3]_c_781_n N_D[4]_c_816_n 9.4377e-19 $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_623 N_D[3]_c_780_n N_D[4]_c_817_n 0.00442615f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_624 N_D[3]_c_778_n N_D[4]_c_818_n 9.4377e-19 $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_625 N_D[3]_c_781_n N_D[4]_c_818_n 0.0199139f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_626 N_D[3]_c_778_n N_VPWR_c_1364_n 0.0231278f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_627 N_D[3]_c_781_n N_VPWR_c_1364_n 0.0044581f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_628 N_D[3]_c_778_n VPWR 0.00594051f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_629 N_D[3]_c_778_n N_VPWR_c_1380_n 0.00622633f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_630 N_D[3]_c_778_n N_Z_c_1654_n 0.00145364f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_631 N_D[3]_c_780_n N_Z_c_1632_n 0.00686805f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_632 N_D[3]_c_778_n N_Z_c_1633_n 0.00605747f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_633 N_D[3]_c_780_n N_Z_c_1633_n 0.00376465f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_634 N_D[3]_c_781_n N_Z_c_1633_n 0.0216525f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_635 N_D[3]_c_780_n N_Z_c_1645_n 0.0128881f $X=8.095 $Y=1.055 $X2=0 $Y2=0
cc_636 N_D[3]_c_778_n N_Z_c_1816_n 0.00719456f $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_637 N_D[3]_c_781_n N_Z_c_1816_n 0.00989895f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_638 N_D[3]_c_778_n N_Z_c_1671_n 8.42164e-19 $X=8.245 $Y=1.41 $X2=0 $Y2=0
cc_639 N_D[3]_c_779_n N_VGND_c_2114_n 0.00322791f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_640 N_D[3]_c_781_n N_VGND_c_2114_n 0.00222881f $X=8.24 $Y=1.16 $X2=0 $Y2=0
cc_641 N_D[3]_c_779_n VGND 0.0108306f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_642 N_D[3]_c_810_p VGND 0.00942277f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_643 N_D[3]_c_779_n N_VGND_c_2130_n 0.00585385f $X=8.27 $Y=0.995 $X2=0 $Y2=0
cc_644 N_D[3]_c_810_p N_VGND_c_2130_n 0.00842546f $X=8.095 $Y=0.51 $X2=0 $Y2=0
cc_645 N_D[3]_c_780_n A_1574_47# 0.00426617f $X=8.095 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_646 N_D[3]_c_810_p A_1574_47# 0.00894235f $X=8.095 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_647 N_D[4]_c_816_n N_A_1840_265#_M1007_g 0.0388862f $X=8.775 $Y=1.41 $X2=0
+ $Y2=0
cc_648 N_D[4]_c_816_n N_A_1840_265#_c_855_n 0.00712672f $X=8.775 $Y=1.41 $X2=0
+ $Y2=0
cc_649 N_D[4]_c_815_n N_S[4]_c_908_n 0.0286599f $X=8.75 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_650 N_D[4]_c_817_n N_S[4]_c_908_n 0.00289497f $X=8.925 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_651 N_D[4]_c_816_n N_VPWR_c_1364_n 0.0231278f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_652 N_D[4]_c_818_n N_VPWR_c_1364_n 0.0044581f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_653 N_D[4]_c_816_n N_VPWR_c_1374_n 0.00622633f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_654 N_D[4]_c_816_n VPWR 0.00594051f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_655 N_D[4]_c_816_n N_Z_c_1634_n 0.00605747f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_656 N_D[4]_c_817_n N_Z_c_1634_n 0.00376465f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_657 N_D[4]_c_818_n N_Z_c_1634_n 0.0216525f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_658 N_D[4]_c_817_n N_Z_c_1635_n 0.0128881f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_659 N_D[4]_c_817_n N_Z_c_1636_n 0.00686805f $X=8.925 $Y=1.055 $X2=0 $Y2=0
cc_660 N_D[4]_c_816_n N_Z_c_1657_n 0.00145364f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_661 N_D[4]_c_816_n N_Z_c_1816_n 0.00719456f $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_662 N_D[4]_c_818_n N_Z_c_1816_n 0.00989895f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_663 N_D[4]_c_816_n N_Z_c_1672_n 8.42164e-19 $X=8.775 $Y=1.41 $X2=0 $Y2=0
cc_664 N_D[4]_c_815_n N_VGND_c_2114_n 0.00322791f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_665 N_D[4]_c_818_n N_VGND_c_2114_n 0.00222881f $X=8.925 $Y=1.19 $X2=0 $Y2=0
cc_666 N_D[4]_c_815_n N_VGND_c_2124_n 0.00585385f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_667 D[4] N_VGND_c_2124_n 0.00842546f $X=8.885 $Y=0.425 $X2=0 $Y2=0
cc_668 N_D[4]_c_815_n VGND 0.0108306f $X=8.75 $Y=0.995 $X2=0 $Y2=0
cc_669 D[4] VGND 0.00942277f $X=8.885 $Y=0.425 $X2=0 $Y2=0
cc_670 N_D[4]_c_817_n A_1765_47# 0.00426617f $X=8.925 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_671 D[4] A_1765_47# 0.00894235f $X=8.885 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_672 N_A_1840_265#_c_852_n N_S[4]_c_909_n 0.00827389f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_673 N_A_1840_265#_c_853_n N_S[4]_c_909_n 0.0164662f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_674 N_A_1840_265#_c_854_n N_S[4]_c_909_n 0.00928634f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_675 N_A_1840_265#_c_855_n N_S[4]_c_909_n 0.0184911f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_676 N_A_1840_265#_c_855_n N_S[4]_c_910_n 0.00820745f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_677 N_A_1840_265#_c_853_n N_S[4]_c_911_n 0.0012443f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_678 N_A_1840_265#_c_857_n N_S[4]_c_911_n 0.00903826f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_679 N_A_1840_265#_c_854_n N_S[4]_c_911_n 0.00767015f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_680 N_A_1840_265#_c_855_n N_S[4]_c_911_n 0.00659591f $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_681 N_A_1840_265#_c_853_n N_S[4]_c_912_n 0.00219336f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_682 N_A_1840_265#_c_852_n N_S[4]_c_913_n 0.00603567f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_683 N_A_1840_265#_c_853_n N_S[4]_c_913_n 0.0178233f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_684 N_A_1840_265#_c_854_n N_S[4]_c_913_n 0.0214702f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_685 N_A_1840_265#_c_855_n N_S[4]_c_913_n 2.59957e-19 $X=9.3 $Y=1.34 $X2=0
+ $Y2=0
cc_686 N_A_1840_265#_M1007_g N_VPWR_c_1364_n 0.0030953f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_687 N_A_1840_265#_c_857_n N_VPWR_c_1365_n 0.0292866f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_688 N_A_1840_265#_c_854_n N_VPWR_c_1365_n 0.00688579f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_689 N_A_1840_265#_M1007_g N_VPWR_c_1374_n 0.00522699f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_690 N_A_1840_265#_c_857_n N_VPWR_c_1374_n 0.0210596f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_691 N_A_1840_265#_M1038_s VPWR 0.00179197f $X=9.93 $Y=1.485 $X2=0 $Y2=0
cc_692 N_A_1840_265#_M1007_g VPWR 0.00809563f $X=9.3 $Y=2.075 $X2=0 $Y2=0
cc_693 N_A_1840_265#_c_857_n VPWR 0.00594162f $X=10.055 $Y=2.31 $X2=0 $Y2=0
cc_694 N_A_1840_265#_M1007_g N_Z_c_1634_n 0.00862328f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_695 N_A_1840_265#_c_853_n N_Z_c_1634_n 0.00719188f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_696 N_A_1840_265#_c_857_n N_Z_c_1634_n 0.00378484f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_697 N_A_1840_265#_c_854_n N_Z_c_1634_n 0.0304368f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_698 N_A_1840_265#_c_855_n N_Z_c_1634_n 0.00814206f $X=9.3 $Y=1.34 $X2=0 $Y2=0
cc_699 N_A_1840_265#_c_853_n N_Z_c_1635_n 0.0124144f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_700 N_A_1840_265#_c_854_n N_Z_c_1635_n 0.00398133f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_701 N_A_1840_265#_c_855_n N_Z_c_1635_n 0.00349316f $X=9.3 $Y=1.34 $X2=0 $Y2=0
cc_702 N_A_1840_265#_c_852_n N_Z_c_1636_n 0.0259454f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_703 N_A_1840_265#_c_853_n N_Z_c_1636_n 0.00611965f $X=9.825 $Y=1.175 $X2=0
+ $Y2=0
cc_704 N_A_1840_265#_M1007_g N_Z_c_1657_n 0.00988241f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_705 N_A_1840_265#_c_857_n N_Z_c_1657_n 0.0369227f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_706 N_A_1840_265#_c_857_n N_Z_c_1666_n 0.0291787f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_707 N_A_1840_265#_c_854_n N_Z_c_1666_n 0.0126642f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_708 N_A_1840_265#_M1007_g N_Z_c_1842_n 0.00289142f $X=9.3 $Y=2.075 $X2=0
+ $Y2=0
cc_709 N_A_1840_265#_c_857_n N_Z_c_1842_n 6.03258e-19 $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_710 N_A_1840_265#_c_854_n N_Z_c_1842_n 4.25753e-19 $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_711 N_A_1840_265#_M1007_g N_Z_c_1672_n 0.0105217f $X=9.3 $Y=2.075 $X2=0 $Y2=0
cc_712 N_A_1840_265#_c_857_n N_Z_c_1672_n 0.0139746f $X=10.055 $Y=2.31 $X2=0
+ $Y2=0
cc_713 N_A_1840_265#_c_854_n N_Z_c_1672_n 0.00749676f $X=10.055 $Y=1.63 $X2=0
+ $Y2=0
cc_714 N_A_1840_265#_c_855_n N_Z_c_1672_n 0.00449162f $X=9.3 $Y=1.34 $X2=0 $Y2=0
cc_715 N_A_1840_265#_c_852_n N_VGND_c_2124_n 0.015238f $X=9.825 $Y=0.755 $X2=0
+ $Y2=0
cc_716 N_A_1840_265#_M1046_s VGND 0.00358139f $X=9.93 $Y=0.235 $X2=0 $Y2=0
cc_717 N_A_1840_265#_c_852_n VGND 0.0150148f $X=9.825 $Y=0.755 $X2=0 $Y2=0
cc_718 N_S[4]_c_911_n N_S[5]_c_955_n 0.0578733f $X=10.29 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_719 N_S[4]_c_913_n N_S[5]_c_955_n 0.00112057f $X=10.255 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_720 N_S[4]_c_912_n N_S[5]_c_956_n 0.0091402f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_721 N_S[4]_c_911_n N_S[5]_c_959_n 0.00112057f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_722 N_S[4]_c_913_n N_S[5]_c_959_n 0.0277403f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_723 N_S[4]_c_911_n N_VPWR_c_1365_n 0.00965725f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_724 N_S[4]_c_913_n N_VPWR_c_1365_n 0.00587376f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_725 N_S[4]_c_911_n N_VPWR_c_1374_n 0.00673617f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_726 N_S[4]_c_911_n VPWR 0.00871384f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_727 N_S[4]_c_910_n N_Z_c_1634_n 7.46972e-19 $X=9.3 $Y=0.905 $X2=0 $Y2=0
cc_728 N_S[4]_c_909_n N_Z_c_1635_n 0.00806549f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_729 N_S[4]_c_910_n N_Z_c_1635_n 0.00605736f $X=9.3 $Y=0.905 $X2=0 $Y2=0
cc_730 N_S[4]_c_908_n N_Z_c_1636_n 0.00316445f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_731 N_S[4]_c_909_n N_Z_c_1636_n 0.00501353f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_732 N_S[4]_c_911_n N_Z_c_1666_n 0.0062071f $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_733 N_S[4]_c_913_n N_Z_c_1666_n 0.00659242f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_734 N_S[4]_c_912_n N_VGND_c_2115_n 0.00570474f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_735 N_S[4]_c_913_n N_VGND_c_2115_n 0.00391126f $X=10.255 $Y=1.03 $X2=0 $Y2=0
cc_736 N_S[4]_c_908_n N_VGND_c_2124_n 0.00585385f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_737 N_S[4]_c_912_n N_VGND_c_2124_n 0.00585385f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_738 N_S[4]_c_908_n VGND 0.00880034f $X=9.225 $Y=0.83 $X2=0 $Y2=0
cc_739 N_S[4]_c_909_n VGND 0.00349917f $X=10.12 $Y=0.905 $X2=0 $Y2=0
cc_740 N_S[4]_c_911_n VGND 6.15795e-19 $X=10.29 $Y=1.41 $X2=0 $Y2=0
cc_741 N_S[4]_c_912_n VGND 0.0124506f $X=10.29 $Y=0.83 $X2=0 $Y2=0
cc_742 N_S[5]_c_955_n N_A_2189_47#_c_1004_n 0.00903826f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_743 N_S[5]_c_955_n N_A_2189_47#_c_999_n 0.0012443f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_744 N_S[5]_c_956_n N_A_2189_47#_c_999_n 0.00219336f $X=10.87 $Y=0.83 $X2=0
+ $Y2=0
cc_745 N_S[5]_c_957_n N_A_2189_47#_c_999_n 0.0164662f $X=11.86 $Y=0.905 $X2=0
+ $Y2=0
cc_746 N_S[5]_c_959_n N_A_2189_47#_c_999_n 0.0178233f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_747 N_S[5]_c_955_n N_A_2189_47#_c_1000_n 0.00767015f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_748 N_S[5]_c_957_n N_A_2189_47#_c_1000_n 0.00928634f $X=11.86 $Y=0.905 $X2=0
+ $Y2=0
cc_749 N_S[5]_c_959_n N_A_2189_47#_c_1000_n 0.0214702f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_750 N_S[5]_c_955_n N_A_2189_47#_c_1001_n 0.00659591f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_751 N_S[5]_c_957_n N_A_2189_47#_c_1001_n 0.0266986f $X=11.86 $Y=0.905 $X2=0
+ $Y2=0
cc_752 N_S[5]_c_959_n N_A_2189_47#_c_1001_n 2.59957e-19 $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_753 N_S[5]_c_955_n N_A_2189_47#_c_1002_n 0.00827389f $X=10.87 $Y=1.41 $X2=0
+ $Y2=0
cc_754 N_S[5]_c_959_n N_A_2189_47#_c_1002_n 0.00603567f $X=10.905 $Y=1.03 $X2=0
+ $Y2=0
cc_755 N_S[5]_c_958_n N_D[5]_c_1055_n 0.0286599f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_756 N_S[5]_c_958_n N_D[5]_c_1056_n 0.00289497f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_757 N_S[5]_c_955_n N_VPWR_c_1365_n 0.00965725f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_758 N_S[5]_c_959_n N_VPWR_c_1365_n 0.00587376f $X=10.905 $Y=1.03 $X2=0 $Y2=0
cc_759 N_S[5]_c_955_n VPWR 0.00871384f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_760 N_S[5]_c_955_n N_VPWR_c_1381_n 0.00673617f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_761 N_S[5]_c_957_n N_Z_c_1637_n 0.00501353f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_762 N_S[5]_c_958_n N_Z_c_1637_n 0.00316445f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_763 N_S[5]_c_957_n N_Z_c_1638_n 7.46972e-19 $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_764 N_S[5]_c_957_n N_Z_c_1646_n 0.0141229f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_765 N_S[5]_c_955_n N_Z_c_1666_n 0.0062071f $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_766 N_S[5]_c_959_n N_Z_c_1666_n 0.00659242f $X=10.905 $Y=1.03 $X2=0 $Y2=0
cc_767 N_S[5]_c_956_n N_VGND_c_2115_n 0.00570474f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_768 N_S[5]_c_959_n N_VGND_c_2115_n 0.00391126f $X=10.905 $Y=1.03 $X2=0 $Y2=0
cc_769 N_S[5]_c_955_n VGND 6.15795e-19 $X=10.87 $Y=1.41 $X2=0 $Y2=0
cc_770 N_S[5]_c_956_n VGND 0.0124506f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_771 N_S[5]_c_957_n VGND 0.00349917f $X=11.86 $Y=0.905 $X2=0 $Y2=0
cc_772 N_S[5]_c_958_n VGND 0.00880034f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_773 N_S[5]_c_956_n N_VGND_c_2131_n 0.00585385f $X=10.87 $Y=0.83 $X2=0 $Y2=0
cc_774 N_S[5]_c_958_n N_VGND_c_2131_n 0.00585385f $X=11.935 $Y=0.83 $X2=0 $Y2=0
cc_775 N_A_2189_47#_M1030_g N_D[5]_c_1054_n 0.0388862f $X=11.86 $Y=2.075
+ $X2=-0.19 $Y2=-0.24
cc_776 N_A_2189_47#_c_1001_n N_D[5]_c_1054_n 0.00712672f $X=11.555 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_777 N_A_2189_47#_c_1004_n N_VPWR_c_1365_n 0.0292866f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_778 N_A_2189_47#_c_1000_n N_VPWR_c_1365_n 0.00688579f $X=11.335 $Y=1.405
+ $X2=0 $Y2=0
cc_779 N_A_2189_47#_M1030_g N_VPWR_c_1366_n 0.0030953f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_780 N_A_2189_47#_M1024_d VPWR 0.00179197f $X=10.96 $Y=1.485 $X2=0 $Y2=0
cc_781 N_A_2189_47#_M1030_g VPWR 0.00809563f $X=11.86 $Y=2.075 $X2=0 $Y2=0
cc_782 N_A_2189_47#_c_1004_n VPWR 0.00594162f $X=11.105 $Y=2.31 $X2=0 $Y2=0
cc_783 N_A_2189_47#_M1030_g N_VPWR_c_1381_n 0.00522699f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_784 N_A_2189_47#_c_1004_n N_VPWR_c_1381_n 0.0210596f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_785 N_A_2189_47#_M1030_g N_Z_c_1658_n 0.00988241f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_786 N_A_2189_47#_c_1004_n N_Z_c_1658_n 0.0369227f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_787 N_A_2189_47#_c_999_n N_Z_c_1637_n 0.00611965f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_788 N_A_2189_47#_c_1002_n N_Z_c_1637_n 0.0259454f $X=11.105 $Y=0.495 $X2=0
+ $Y2=0
cc_789 N_A_2189_47#_M1030_g N_Z_c_1638_n 0.00862328f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_790 N_A_2189_47#_c_1004_n N_Z_c_1638_n 0.00378484f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_791 N_A_2189_47#_c_999_n N_Z_c_1638_n 0.00719188f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_792 N_A_2189_47#_c_1000_n N_Z_c_1638_n 0.0304368f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_793 N_A_2189_47#_c_1001_n N_Z_c_1638_n 0.00814206f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_794 N_A_2189_47#_c_999_n N_Z_c_1646_n 0.0124144f $X=11.335 $Y=1.175 $X2=0
+ $Y2=0
cc_795 N_A_2189_47#_c_1000_n N_Z_c_1646_n 0.00398133f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_796 N_A_2189_47#_c_1001_n N_Z_c_1646_n 0.00349316f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_797 N_A_2189_47#_c_1004_n N_Z_c_1666_n 0.0291787f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_798 N_A_2189_47#_c_1000_n N_Z_c_1666_n 0.0126642f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_799 N_A_2189_47#_M1030_g N_Z_c_1876_n 0.00289142f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_800 N_A_2189_47#_c_1004_n N_Z_c_1876_n 6.03258e-19 $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_801 N_A_2189_47#_c_1000_n N_Z_c_1876_n 4.25753e-19 $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_802 N_A_2189_47#_M1030_g N_Z_c_1673_n 0.0105217f $X=11.86 $Y=2.075 $X2=0
+ $Y2=0
cc_803 N_A_2189_47#_c_1004_n N_Z_c_1673_n 0.0139746f $X=11.105 $Y=2.31 $X2=0
+ $Y2=0
cc_804 N_A_2189_47#_c_1000_n N_Z_c_1673_n 0.00749676f $X=11.335 $Y=1.405 $X2=0
+ $Y2=0
cc_805 N_A_2189_47#_c_1001_n N_Z_c_1673_n 0.00449162f $X=11.555 $Y=1.34 $X2=0
+ $Y2=0
cc_806 N_A_2189_47#_M1037_d VGND 0.00358139f $X=10.945 $Y=0.235 $X2=0 $Y2=0
cc_807 N_A_2189_47#_c_1002_n VGND 0.0150148f $X=11.105 $Y=0.495 $X2=0 $Y2=0
cc_808 N_A_2189_47#_c_1002_n N_VGND_c_2131_n 0.015238f $X=11.105 $Y=0.495 $X2=0
+ $Y2=0
cc_809 N_D[5]_c_1055_n N_D[6]_c_1091_n 0.00915308f $X=12.41 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_810 N_D[5]_c_1054_n N_D[6]_c_1092_n 0.0270908f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_811 N_D[5]_c_1057_n N_D[6]_c_1092_n 9.4377e-19 $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_812 N_D[5]_c_1056_n N_D[6]_c_1093_n 0.00442615f $X=12.235 $Y=1.055 $X2=0
+ $Y2=0
cc_813 N_D[5]_c_1054_n N_D[6]_c_1094_n 9.4377e-19 $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_814 N_D[5]_c_1057_n N_D[6]_c_1094_n 0.0199139f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_815 N_D[5]_c_1054_n N_VPWR_c_1366_n 0.0231278f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_816 N_D[5]_c_1057_n N_VPWR_c_1366_n 0.0044581f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_817 N_D[5]_c_1054_n VPWR 0.00594051f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_818 N_D[5]_c_1054_n N_VPWR_c_1381_n 0.00622633f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_819 N_D[5]_c_1054_n N_Z_c_1658_n 0.00145364f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_820 N_D[5]_c_1056_n N_Z_c_1637_n 0.00686805f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_821 N_D[5]_c_1054_n N_Z_c_1638_n 0.00605747f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_822 N_D[5]_c_1056_n N_Z_c_1638_n 0.00376465f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_823 N_D[5]_c_1057_n N_Z_c_1638_n 0.0216525f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_824 N_D[5]_c_1056_n N_Z_c_1646_n 0.0128881f $X=12.235 $Y=1.055 $X2=0 $Y2=0
cc_825 N_D[5]_c_1054_n N_Z_c_1889_n 0.00719456f $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_826 N_D[5]_c_1057_n N_Z_c_1889_n 0.00989895f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_827 N_D[5]_c_1054_n N_Z_c_1673_n 8.42164e-19 $X=12.385 $Y=1.41 $X2=0 $Y2=0
cc_828 N_D[5]_c_1055_n N_VGND_c_2116_n 0.00322791f $X=12.41 $Y=0.995 $X2=0 $Y2=0
cc_829 N_D[5]_c_1057_n N_VGND_c_2116_n 0.00222881f $X=12.38 $Y=1.16 $X2=0 $Y2=0
cc_830 N_D[5]_c_1055_n VGND 0.0108306f $X=12.41 $Y=0.995 $X2=0 $Y2=0
cc_831 N_D[5]_c_1086_p VGND 0.00942277f $X=12.235 $Y=0.51 $X2=0 $Y2=0
cc_832 N_D[5]_c_1055_n N_VGND_c_2131_n 0.00585385f $X=12.41 $Y=0.995 $X2=0 $Y2=0
cc_833 N_D[5]_c_1086_p N_VGND_c_2131_n 0.00842546f $X=12.235 $Y=0.51 $X2=0 $Y2=0
cc_834 N_D[5]_c_1056_n A_2402_47# 0.00426617f $X=12.235 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_835 N_D[5]_c_1086_p A_2402_47# 0.00894235f $X=12.235 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_836 N_D[6]_c_1092_n N_A_2668_265#_M1026_g 0.0388862f $X=12.915 $Y=1.41 $X2=0
+ $Y2=0
cc_837 N_D[6]_c_1092_n N_A_2668_265#_c_1131_n 0.00712672f $X=12.915 $Y=1.41
+ $X2=0 $Y2=0
cc_838 N_D[6]_c_1091_n N_S[6]_c_1184_n 0.0286599f $X=12.89 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_839 N_D[6]_c_1093_n N_S[6]_c_1184_n 0.00289497f $X=13.065 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_840 N_D[6]_c_1092_n N_VPWR_c_1366_n 0.0231278f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_841 N_D[6]_c_1094_n N_VPWR_c_1366_n 0.0044581f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_842 N_D[6]_c_1092_n N_VPWR_c_1376_n 0.00622633f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_843 N_D[6]_c_1092_n VPWR 0.00594051f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_844 N_D[6]_c_1092_n N_Z_c_1639_n 0.00605747f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_845 N_D[6]_c_1093_n N_Z_c_1639_n 0.00376465f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_846 N_D[6]_c_1094_n N_Z_c_1639_n 0.0216525f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_847 N_D[6]_c_1093_n N_Z_c_1640_n 0.0128881f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_848 N_D[6]_c_1093_n N_Z_c_1641_n 0.00686805f $X=13.065 $Y=1.055 $X2=0 $Y2=0
cc_849 N_D[6]_c_1092_n N_Z_c_1661_n 0.00145364f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_850 N_D[6]_c_1092_n N_Z_c_1889_n 0.00719456f $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_851 N_D[6]_c_1094_n N_Z_c_1889_n 0.00989895f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_852 N_D[6]_c_1092_n N_Z_c_1674_n 8.42164e-19 $X=12.915 $Y=1.41 $X2=0 $Y2=0
cc_853 N_D[6]_c_1091_n N_VGND_c_2116_n 0.00322791f $X=12.89 $Y=0.995 $X2=0 $Y2=0
cc_854 N_D[6]_c_1094_n N_VGND_c_2116_n 0.00222881f $X=13.065 $Y=1.19 $X2=0 $Y2=0
cc_855 N_D[6]_c_1091_n N_VGND_c_2126_n 0.00585385f $X=12.89 $Y=0.995 $X2=0 $Y2=0
cc_856 D[6] N_VGND_c_2126_n 0.00842546f $X=13.025 $Y=0.425 $X2=0 $Y2=0
cc_857 N_D[6]_c_1091_n VGND 0.0108306f $X=12.89 $Y=0.995 $X2=0 $Y2=0
cc_858 D[6] VGND 0.00942277f $X=13.025 $Y=0.425 $X2=0 $Y2=0
cc_859 N_D[6]_c_1093_n A_2593_47# 0.00426617f $X=13.065 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_860 D[6] A_2593_47# 0.00894235f $X=13.025 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_861 N_A_2668_265#_c_1128_n N_S[6]_c_1185_n 0.00827389f $X=13.965 $Y=0.755
+ $X2=0 $Y2=0
cc_862 N_A_2668_265#_c_1129_n N_S[6]_c_1185_n 0.0164662f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_863 N_A_2668_265#_c_1130_n N_S[6]_c_1185_n 0.00928634f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_864 N_A_2668_265#_c_1131_n N_S[6]_c_1185_n 0.0184911f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_865 N_A_2668_265#_c_1131_n N_S[6]_c_1186_n 0.00820745f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_866 N_A_2668_265#_c_1129_n N_S[6]_c_1187_n 0.0012443f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_867 N_A_2668_265#_c_1133_n N_S[6]_c_1187_n 0.00903826f $X=14.195 $Y=2.31
+ $X2=0 $Y2=0
cc_868 N_A_2668_265#_c_1130_n N_S[6]_c_1187_n 0.00767015f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_869 N_A_2668_265#_c_1131_n N_S[6]_c_1187_n 0.00659591f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_870 N_A_2668_265#_c_1129_n N_S[6]_c_1188_n 0.00219336f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_871 N_A_2668_265#_c_1128_n N_S[6]_c_1189_n 0.00603567f $X=13.965 $Y=0.755
+ $X2=0 $Y2=0
cc_872 N_A_2668_265#_c_1129_n N_S[6]_c_1189_n 0.0178233f $X=13.965 $Y=1.175
+ $X2=0 $Y2=0
cc_873 N_A_2668_265#_c_1130_n N_S[6]_c_1189_n 0.0214702f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_874 N_A_2668_265#_c_1131_n N_S[6]_c_1189_n 2.59957e-19 $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_875 N_A_2668_265#_M1026_g N_VPWR_c_1366_n 0.0030953f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_876 N_A_2668_265#_c_1133_n N_VPWR_c_1367_n 0.0292866f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_877 N_A_2668_265#_c_1130_n N_VPWR_c_1367_n 0.00688579f $X=14.195 $Y=1.63
+ $X2=0 $Y2=0
cc_878 N_A_2668_265#_M1026_g N_VPWR_c_1376_n 0.00522699f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_879 N_A_2668_265#_c_1133_n N_VPWR_c_1376_n 0.0210596f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_880 N_A_2668_265#_M1034_s VPWR 0.00179197f $X=14.07 $Y=1.485 $X2=0 $Y2=0
cc_881 N_A_2668_265#_M1026_g VPWR 0.00809563f $X=13.44 $Y=2.075 $X2=0 $Y2=0
cc_882 N_A_2668_265#_c_1133_n VPWR 0.00594162f $X=14.195 $Y=2.31 $X2=0 $Y2=0
cc_883 N_A_2668_265#_M1026_g N_Z_c_1639_n 0.00862328f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_884 N_A_2668_265#_c_1129_n N_Z_c_1639_n 0.00719188f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_885 N_A_2668_265#_c_1133_n N_Z_c_1639_n 0.00378484f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_886 N_A_2668_265#_c_1130_n N_Z_c_1639_n 0.0304368f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_887 N_A_2668_265#_c_1131_n N_Z_c_1639_n 0.00814206f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_888 N_A_2668_265#_c_1129_n N_Z_c_1640_n 0.0124144f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_889 N_A_2668_265#_c_1130_n N_Z_c_1640_n 0.00398133f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_890 N_A_2668_265#_c_1131_n N_Z_c_1640_n 0.00349316f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_891 N_A_2668_265#_c_1128_n N_Z_c_1641_n 0.0259454f $X=13.965 $Y=0.755 $X2=0
+ $Y2=0
cc_892 N_A_2668_265#_c_1129_n N_Z_c_1641_n 0.00611965f $X=13.965 $Y=1.175 $X2=0
+ $Y2=0
cc_893 N_A_2668_265#_M1026_g N_Z_c_1661_n 0.00988241f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_894 N_A_2668_265#_c_1133_n N_Z_c_1661_n 0.0369227f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_895 N_A_2668_265#_c_1133_n N_Z_c_1667_n 0.0291787f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_896 N_A_2668_265#_c_1130_n N_Z_c_1667_n 0.0126642f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_897 N_A_2668_265#_M1026_g N_Z_c_1915_n 0.00289142f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_898 N_A_2668_265#_c_1133_n N_Z_c_1915_n 6.03258e-19 $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_899 N_A_2668_265#_c_1130_n N_Z_c_1915_n 4.25753e-19 $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_900 N_A_2668_265#_M1026_g N_Z_c_1674_n 0.0105217f $X=13.44 $Y=2.075 $X2=0
+ $Y2=0
cc_901 N_A_2668_265#_c_1133_n N_Z_c_1674_n 0.0139746f $X=14.195 $Y=2.31 $X2=0
+ $Y2=0
cc_902 N_A_2668_265#_c_1130_n N_Z_c_1674_n 0.00749676f $X=14.195 $Y=1.63 $X2=0
+ $Y2=0
cc_903 N_A_2668_265#_c_1131_n N_Z_c_1674_n 0.00449162f $X=13.44 $Y=1.34 $X2=0
+ $Y2=0
cc_904 N_A_2668_265#_c_1128_n N_VGND_c_2126_n 0.015238f $X=13.965 $Y=0.755 $X2=0
+ $Y2=0
cc_905 N_A_2668_265#_M1004_s VGND 0.00358139f $X=14.07 $Y=0.235 $X2=0 $Y2=0
cc_906 N_A_2668_265#_c_1128_n VGND 0.0150148f $X=13.965 $Y=0.755 $X2=0 $Y2=0
cc_907 N_S[6]_c_1187_n N_S[7]_c_1231_n 0.0578733f $X=14.43 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_908 N_S[6]_c_1189_n N_S[7]_c_1231_n 0.00112057f $X=14.395 $Y=1.03 $X2=-0.19
+ $Y2=-0.24
cc_909 N_S[6]_c_1188_n N_S[7]_c_1232_n 0.0091402f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_910 N_S[6]_c_1187_n N_S[7]_c_1235_n 0.00112057f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_911 N_S[6]_c_1189_n N_S[7]_c_1235_n 0.0277403f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_912 N_S[6]_c_1187_n N_VPWR_c_1367_n 0.00965725f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_913 N_S[6]_c_1189_n N_VPWR_c_1367_n 0.00587376f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_914 N_S[6]_c_1187_n N_VPWR_c_1376_n 0.00673617f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_915 N_S[6]_c_1187_n VPWR 0.00871384f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_916 N_S[6]_c_1186_n N_Z_c_1639_n 7.46972e-19 $X=13.44 $Y=0.905 $X2=0 $Y2=0
cc_917 N_S[6]_c_1185_n N_Z_c_1640_n 0.00806549f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_918 N_S[6]_c_1186_n N_Z_c_1640_n 0.00605736f $X=13.44 $Y=0.905 $X2=0 $Y2=0
cc_919 N_S[6]_c_1184_n N_Z_c_1641_n 0.00316445f $X=13.365 $Y=0.83 $X2=0 $Y2=0
cc_920 N_S[6]_c_1185_n N_Z_c_1641_n 0.00501353f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_921 N_S[6]_c_1187_n N_Z_c_1667_n 0.0062071f $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_922 N_S[6]_c_1189_n N_Z_c_1667_n 0.00659242f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_923 N_S[6]_c_1188_n N_VGND_c_2117_n 0.00570474f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_924 N_S[6]_c_1189_n N_VGND_c_2117_n 0.00391126f $X=14.395 $Y=1.03 $X2=0 $Y2=0
cc_925 N_S[6]_c_1184_n N_VGND_c_2126_n 0.00585385f $X=13.365 $Y=0.83 $X2=0 $Y2=0
cc_926 N_S[6]_c_1188_n N_VGND_c_2126_n 0.00585385f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_927 N_S[6]_c_1184_n VGND 0.00880034f $X=13.365 $Y=0.83 $X2=0 $Y2=0
cc_928 N_S[6]_c_1185_n VGND 0.00349917f $X=14.26 $Y=0.905 $X2=0 $Y2=0
cc_929 N_S[6]_c_1187_n VGND 6.15795e-19 $X=14.43 $Y=1.41 $X2=0 $Y2=0
cc_930 N_S[6]_c_1188_n VGND 0.0124506f $X=14.43 $Y=0.83 $X2=0 $Y2=0
cc_931 N_S[7]_c_1231_n N_A_3017_47#_c_1280_n 0.00903826f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_932 N_S[7]_c_1231_n N_A_3017_47#_c_1275_n 0.0012443f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_933 N_S[7]_c_1232_n N_A_3017_47#_c_1275_n 0.00219336f $X=15.01 $Y=0.83 $X2=0
+ $Y2=0
cc_934 N_S[7]_c_1233_n N_A_3017_47#_c_1275_n 0.0164662f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_935 N_S[7]_c_1235_n N_A_3017_47#_c_1275_n 0.0178233f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_936 N_S[7]_c_1231_n N_A_3017_47#_c_1276_n 0.00767015f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_937 N_S[7]_c_1233_n N_A_3017_47#_c_1276_n 0.00928634f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_938 N_S[7]_c_1235_n N_A_3017_47#_c_1276_n 0.0214702f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_939 N_S[7]_c_1231_n N_A_3017_47#_c_1277_n 0.00659591f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_940 N_S[7]_c_1233_n N_A_3017_47#_c_1277_n 0.0266986f $X=16 $Y=0.905 $X2=0
+ $Y2=0
cc_941 N_S[7]_c_1235_n N_A_3017_47#_c_1277_n 2.59957e-19 $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_942 N_S[7]_c_1231_n N_A_3017_47#_c_1278_n 0.00827389f $X=15.01 $Y=1.41 $X2=0
+ $Y2=0
cc_943 N_S[7]_c_1235_n N_A_3017_47#_c_1278_n 0.00603567f $X=15.045 $Y=1.03 $X2=0
+ $Y2=0
cc_944 N_S[7]_c_1234_n N_D[7]_c_1331_n 0.0286599f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_945 N_S[7]_c_1234_n N_D[7]_c_1332_n 0.00289497f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_946 N_S[7]_c_1231_n N_VPWR_c_1367_n 0.00965725f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_947 N_S[7]_c_1235_n N_VPWR_c_1367_n 0.00587376f $X=15.045 $Y=1.03 $X2=0 $Y2=0
cc_948 N_S[7]_c_1231_n VPWR 0.00871384f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_949 N_S[7]_c_1231_n N_VPWR_c_1382_n 0.00673617f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_950 N_S[7]_c_1233_n N_Z_c_1642_n 0.00501353f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_951 N_S[7]_c_1234_n N_Z_c_1642_n 0.00316445f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_952 N_S[7]_c_1233_n N_Z_c_1643_n 7.46972e-19 $X=16 $Y=0.905 $X2=0 $Y2=0
cc_953 N_S[7]_c_1233_n N_Z_c_1647_n 0.0141229f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_954 N_S[7]_c_1231_n N_Z_c_1667_n 0.0062071f $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_955 N_S[7]_c_1235_n N_Z_c_1667_n 0.00659242f $X=15.045 $Y=1.03 $X2=0 $Y2=0
cc_956 N_S[7]_c_1232_n N_VGND_c_2117_n 0.00570474f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_957 N_S[7]_c_1235_n N_VGND_c_2117_n 0.00391126f $X=15.045 $Y=1.03 $X2=0 $Y2=0
cc_958 N_S[7]_c_1231_n VGND 6.15795e-19 $X=15.01 $Y=1.41 $X2=0 $Y2=0
cc_959 N_S[7]_c_1232_n VGND 0.0124506f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_960 N_S[7]_c_1233_n VGND 0.00349917f $X=16 $Y=0.905 $X2=0 $Y2=0
cc_961 N_S[7]_c_1234_n VGND 0.00880034f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_962 N_S[7]_c_1232_n N_VGND_c_2132_n 0.00585385f $X=15.01 $Y=0.83 $X2=0 $Y2=0
cc_963 N_S[7]_c_1234_n N_VGND_c_2132_n 0.00585385f $X=16.075 $Y=0.83 $X2=0 $Y2=0
cc_964 N_A_3017_47#_M1045_g N_D[7]_c_1330_n 0.0381613f $X=16 $Y=2.075 $X2=-0.19
+ $Y2=-0.24
cc_965 N_A_3017_47#_c_1277_n N_D[7]_c_1330_n 0.00712672f $X=15.695 $Y=1.34
+ $X2=-0.19 $Y2=-0.24
cc_966 N_A_3017_47#_c_1280_n N_VPWR_c_1367_n 0.0292866f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_967 N_A_3017_47#_c_1276_n N_VPWR_c_1367_n 0.00688579f $X=15.475 $Y=1.405
+ $X2=0 $Y2=0
cc_968 N_A_3017_47#_M1045_g N_VPWR_c_1369_n 0.00298082f $X=16 $Y=2.075 $X2=0
+ $Y2=0
cc_969 N_A_3017_47#_M1011_d VPWR 0.00179197f $X=15.1 $Y=1.485 $X2=0 $Y2=0
cc_970 N_A_3017_47#_M1045_g VPWR 0.00828927f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_971 N_A_3017_47#_c_1280_n VPWR 0.00594162f $X=15.245 $Y=2.31 $X2=0 $Y2=0
cc_972 N_A_3017_47#_M1045_g N_VPWR_c_1382_n 0.00522699f $X=16 $Y=2.075 $X2=0
+ $Y2=0
cc_973 N_A_3017_47#_c_1280_n N_VPWR_c_1382_n 0.0210596f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_974 N_A_3017_47#_M1045_g N_Z_c_1662_n 0.00988241f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_975 N_A_3017_47#_c_1280_n N_Z_c_1662_n 0.0369227f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_976 N_A_3017_47#_c_1275_n N_Z_c_1642_n 0.00611965f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_977 N_A_3017_47#_c_1278_n N_Z_c_1642_n 0.0259454f $X=15.245 $Y=0.495 $X2=0
+ $Y2=0
cc_978 N_A_3017_47#_M1045_g N_Z_c_1643_n 0.00862328f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_979 N_A_3017_47#_c_1280_n N_Z_c_1643_n 0.00378484f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_980 N_A_3017_47#_c_1275_n N_Z_c_1643_n 0.00719188f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_981 N_A_3017_47#_c_1276_n N_Z_c_1643_n 0.0304368f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_982 N_A_3017_47#_c_1277_n N_Z_c_1643_n 0.00814206f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_983 N_A_3017_47#_c_1275_n N_Z_c_1647_n 0.0124144f $X=15.475 $Y=1.175 $X2=0
+ $Y2=0
cc_984 N_A_3017_47#_c_1276_n N_Z_c_1647_n 0.00398133f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_985 N_A_3017_47#_c_1277_n N_Z_c_1647_n 0.00349316f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_986 N_A_3017_47#_c_1280_n N_Z_c_1667_n 0.0291787f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_987 N_A_3017_47#_c_1276_n N_Z_c_1667_n 0.0126642f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_988 N_A_3017_47#_M1045_g Z 0.00289142f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_989 N_A_3017_47#_c_1280_n Z 6.03258e-19 $X=15.245 $Y=2.31 $X2=0 $Y2=0
cc_990 N_A_3017_47#_c_1276_n Z 4.25753e-19 $X=15.475 $Y=1.405 $X2=0 $Y2=0
cc_991 N_A_3017_47#_M1045_g N_Z_c_1675_n 0.0105217f $X=16 $Y=2.075 $X2=0 $Y2=0
cc_992 N_A_3017_47#_c_1280_n N_Z_c_1675_n 0.0139746f $X=15.245 $Y=2.31 $X2=0
+ $Y2=0
cc_993 N_A_3017_47#_c_1276_n N_Z_c_1675_n 0.00749676f $X=15.475 $Y=1.405 $X2=0
+ $Y2=0
cc_994 N_A_3017_47#_c_1277_n N_Z_c_1675_n 0.00449162f $X=15.695 $Y=1.34 $X2=0
+ $Y2=0
cc_995 N_A_3017_47#_M1047_d VGND 0.00358139f $X=15.085 $Y=0.235 $X2=0 $Y2=0
cc_996 N_A_3017_47#_c_1278_n VGND 0.0150148f $X=15.245 $Y=0.495 $X2=0 $Y2=0
cc_997 N_A_3017_47#_c_1278_n N_VGND_c_2132_n 0.015238f $X=15.245 $Y=0.495 $X2=0
+ $Y2=0
cc_998 N_D[7]_c_1330_n N_VPWR_c_1369_n 0.0245615f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_999 N_D[7]_c_1333_n N_VPWR_c_1369_n 0.00471543f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_1000 N_D[7]_c_1330_n VPWR 0.0106352f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_1001 N_D[7]_c_1330_n N_VPWR_c_1382_n 0.00622633f $X=16.525 $Y=1.41 $X2=0
+ $Y2=0
cc_1002 N_D[7]_c_1330_n N_Z_c_1662_n 0.00145364f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_1003 N_D[7]_c_1332_n N_Z_c_1642_n 0.00686805f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_1004 N_D[7]_c_1330_n N_Z_c_1643_n 0.00605747f $X=16.525 $Y=1.41 $X2=0 $Y2=0
cc_1005 N_D[7]_c_1332_n N_Z_c_1643_n 0.00376465f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_1006 N_D[7]_c_1333_n N_Z_c_1643_n 0.0216525f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_1007 N_D[7]_c_1332_n N_Z_c_1647_n 0.0128881f $X=16.375 $Y=1.055 $X2=0 $Y2=0
cc_1008 N_D[7]_c_1331_n N_VGND_c_2119_n 0.00487865f $X=16.55 $Y=0.995 $X2=0
+ $Y2=0
cc_1009 N_D[7]_c_1333_n N_VGND_c_2119_n 0.00222881f $X=16.52 $Y=1.16 $X2=0 $Y2=0
cc_1010 N_D[7]_c_1331_n VGND 0.011617f $X=16.55 $Y=0.995 $X2=0 $Y2=0
cc_1011 N_D[7]_c_1353_p VGND 0.00942277f $X=16.375 $Y=0.51 $X2=0 $Y2=0
cc_1012 N_D[7]_c_1331_n N_VGND_c_2132_n 0.00585385f $X=16.55 $Y=0.995 $X2=0
+ $Y2=0
cc_1013 N_D[7]_c_1353_p N_VGND_c_2132_n 0.00842546f $X=16.375 $Y=0.51 $X2=0
+ $Y2=0
cc_1014 N_D[7]_c_1332_n A_3230_47# 0.00426617f $X=16.375 $Y=1.055 $X2=-0.19
+ $Y2=-0.24
cc_1015 N_D[7]_c_1353_p A_3230_47# 0.00894235f $X=16.375 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_1016 VPWR A_117_297# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1017 VPWR N_Z_M1019_d 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1018 VPWR N_Z_M1009_s 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1019 VPWR N_Z_M1022_d 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1020 VPWR N_Z_M1013_s 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1021 VPWR N_Z_M1007_d 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1022 VPWR N_Z_M1030_s 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1023 VPWR N_Z_M1026_d 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1024 VPWR N_Z_M1045_s 0.00174926f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1025 N_VPWR_c_1360_n N_Z_c_1624_n 0.00734981f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_1026 N_VPWR_c_1360_n N_Z_c_1649_n 0.0115091f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_1027 N_VPWR_c_1370_n N_Z_c_1649_n 0.0210727f $X=2.135 $Y=2.72 $X2=0 $Y2=0
cc_1028 VPWR N_Z_c_1649_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1029 N_VPWR_c_1362_n N_Z_c_1650_n 0.0116583f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1030 VPWR N_Z_c_1650_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1031 N_VPWR_c_1379_n N_Z_c_1650_n 0.0210727f $X=4.175 $Y=2.72 $X2=0 $Y2=0
cc_1032 N_VPWR_c_1362_n N_Z_c_1628_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1033 N_VPWR_c_1362_n N_Z_c_1629_n 0.0074594f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1034 N_VPWR_c_1362_n N_Z_c_1653_n 0.0116583f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1035 N_VPWR_c_1372_n N_Z_c_1653_n 0.0210727f $X=6.275 $Y=2.72 $X2=0 $Y2=0
cc_1036 VPWR N_Z_c_1653_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1037 N_VPWR_c_1364_n N_Z_c_1654_n 0.0116583f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1038 VPWR N_Z_c_1654_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1039 N_VPWR_c_1380_n N_Z_c_1654_n 0.0210727f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_1040 N_VPWR_c_1364_n N_Z_c_1633_n 0.0074594f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1041 N_VPWR_c_1364_n N_Z_c_1634_n 0.0074594f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1042 N_VPWR_c_1364_n N_Z_c_1657_n 0.0116583f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1043 N_VPWR_c_1374_n N_Z_c_1657_n 0.0210727f $X=10.415 $Y=2.72 $X2=0 $Y2=0
cc_1044 VPWR N_Z_c_1657_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1045 N_VPWR_c_1366_n N_Z_c_1658_n 0.0116583f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1046 VPWR N_Z_c_1658_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1047 N_VPWR_c_1381_n N_Z_c_1658_n 0.0210727f $X=12.455 $Y=2.72 $X2=0 $Y2=0
cc_1048 N_VPWR_c_1366_n N_Z_c_1638_n 0.0074594f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1049 N_VPWR_c_1366_n N_Z_c_1639_n 0.0074594f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1050 N_VPWR_c_1366_n N_Z_c_1661_n 0.0116583f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1051 N_VPWR_c_1376_n N_Z_c_1661_n 0.0210727f $X=14.555 $Y=2.72 $X2=0 $Y2=0
cc_1052 VPWR N_Z_c_1661_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1053 N_VPWR_c_1369_n N_Z_c_1662_n 0.0115091f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_1054 VPWR N_Z_c_1662_n 0.00577491f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1055 N_VPWR_c_1382_n N_Z_c_1662_n 0.0210727f $X=16.595 $Y=2.72 $X2=0 $Y2=0
cc_1056 N_VPWR_c_1369_n N_Z_c_1643_n 0.00734981f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_1057 N_VPWR_M1023_d N_Z_c_1664_n 0.001769f $X=2.1 $Y=1.485 $X2=0 $Y2=0
cc_1058 N_VPWR_c_1361_n N_Z_c_1664_n 0.0291114f $X=2.3 $Y=1.63 $X2=0 $Y2=0
cc_1059 VPWR N_Z_c_1664_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1060 N_VPWR_c_1360_n N_Z_c_1696_n 0.00119119f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_1061 VPWR N_Z_c_1696_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1062 N_VPWR_c_1362_n N_Z_c_1743_n 0.0355595f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1063 VPWR N_Z_c_1743_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1064 N_VPWR_c_1362_n N_Z_c_1730_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1065 VPWR N_Z_c_1730_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1066 N_VPWR_M1025_d N_Z_c_1665_n 0.001769f $X=6.24 $Y=1.485 $X2=0 $Y2=0
cc_1067 N_VPWR_c_1363_n N_Z_c_1665_n 0.0291114f $X=6.44 $Y=1.63 $X2=0 $Y2=0
cc_1068 VPWR N_Z_c_1665_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1069 N_VPWR_c_1362_n N_Z_c_1769_n 4.83404e-19 $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1070 VPWR N_Z_c_1769_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1071 N_VPWR_c_1364_n N_Z_c_1816_n 0.0355595f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1072 VPWR N_Z_c_1816_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1073 N_VPWR_c_1364_n N_Z_c_1803_n 4.83404e-19 $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1074 VPWR N_Z_c_1803_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1075 N_VPWR_M1038_d N_Z_c_1666_n 0.001769f $X=10.38 $Y=1.485 $X2=0 $Y2=0
cc_1076 N_VPWR_c_1365_n N_Z_c_1666_n 0.0291114f $X=10.58 $Y=1.63 $X2=0 $Y2=0
cc_1077 VPWR N_Z_c_1666_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1078 N_VPWR_c_1364_n N_Z_c_1842_n 4.83404e-19 $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1079 VPWR N_Z_c_1842_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1080 N_VPWR_c_1366_n N_Z_c_1889_n 0.0355595f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1081 VPWR N_Z_c_1889_n 0.0739714f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1082 N_VPWR_c_1366_n N_Z_c_1876_n 4.83404e-19 $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1083 VPWR N_Z_c_1876_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1084 N_VPWR_M1034_d N_Z_c_1667_n 0.001769f $X=14.52 $Y=1.485 $X2=0 $Y2=0
cc_1085 N_VPWR_c_1367_n N_Z_c_1667_n 0.0291114f $X=14.72 $Y=1.63 $X2=0 $Y2=0
cc_1086 VPWR N_Z_c_1667_n 0.094685f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1087 N_VPWR_c_1366_n N_Z_c_1915_n 4.83404e-19 $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1088 VPWR N_Z_c_1915_n 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1089 N_VPWR_c_1369_n Z 0.00119119f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_1090 VPWR Z 0.0144722f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1091 N_VPWR_c_1370_n N_Z_c_1668_n 0.00233997f $X=2.135 $Y=2.72 $X2=0 $Y2=0
cc_1092 VPWR N_Z_c_1668_n 0.00317613f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1093 N_VPWR_c_1362_n N_Z_c_1669_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1094 VPWR N_Z_c_1669_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1095 N_VPWR_c_1379_n N_Z_c_1669_n 0.00233997f $X=4.175 $Y=2.72 $X2=0 $Y2=0
cc_1096 N_VPWR_c_1362_n N_Z_c_1670_n 0.00305596f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1097 N_VPWR_c_1372_n N_Z_c_1670_n 0.00233997f $X=6.275 $Y=2.72 $X2=0 $Y2=0
cc_1098 VPWR N_Z_c_1670_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1099 N_VPWR_c_1364_n N_Z_c_1671_n 0.00305596f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1100 VPWR N_Z_c_1671_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1101 N_VPWR_c_1380_n N_Z_c_1671_n 0.00233997f $X=8.315 $Y=2.72 $X2=0 $Y2=0
cc_1102 N_VPWR_c_1364_n N_Z_c_1672_n 0.00305596f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1103 N_VPWR_c_1374_n N_Z_c_1672_n 0.00233997f $X=10.415 $Y=2.72 $X2=0 $Y2=0
cc_1104 VPWR N_Z_c_1672_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1105 N_VPWR_c_1366_n N_Z_c_1673_n 0.00305596f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1106 VPWR N_Z_c_1673_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1107 N_VPWR_c_1381_n N_Z_c_1673_n 0.00233997f $X=12.455 $Y=2.72 $X2=0 $Y2=0
cc_1108 N_VPWR_c_1366_n N_Z_c_1674_n 0.00305596f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1109 N_VPWR_c_1376_n N_Z_c_1674_n 0.00233997f $X=14.555 $Y=2.72 $X2=0 $Y2=0
cc_1110 VPWR N_Z_c_1674_n 0.00180522f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1111 VPWR N_Z_c_1675_n 0.00317613f $X=16.705 $Y=2.635 $X2=0 $Y2=0
cc_1112 N_VPWR_c_1382_n N_Z_c_1675_n 0.00233997f $X=16.595 $Y=2.72 $X2=0 $Y2=0
cc_1113 VPWR A_734_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1114 VPWR A_945_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1115 VPWR A_1562_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1116 VPWR A_1773_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1117 VPWR A_2390_333# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1118 VPWR A_2601_297# 0.00481681f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1119 VPWR A_3218_333# 0.0138589f $X=16.705 $Y=2.635 $X2=-0.19 $Y2=-0.24
cc_1120 N_VPWR_c_1360_n N_VGND_c_2110_n 0.00704239f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_1121 N_VPWR_c_1362_n N_VGND_c_2112_n 0.00723368f $X=4.37 $Y=1.66 $X2=0 $Y2=0
cc_1122 N_VPWR_c_1364_n N_VGND_c_2114_n 0.00723368f $X=8.51 $Y=1.66 $X2=0 $Y2=0
cc_1123 N_VPWR_c_1366_n N_VGND_c_2116_n 0.00723368f $X=12.65 $Y=1.66 $X2=0 $Y2=0
cc_1124 N_VPWR_c_1369_n N_VGND_c_2119_n 0.00704239f $X=16.76 $Y=1.66 $X2=0 $Y2=0
cc_1125 N_Z_c_1743_n A_734_333# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_1126 N_Z_c_1743_n A_945_297# 0.0127078f $X=5.145 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_1127 N_Z_c_1816_n A_1562_333# 0.0127078f $X=9.285 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_1128 N_Z_c_1816_n A_1773_297# 0.0127078f $X=9.285 $Y=1.87 $X2=-0.19 $Y2=-0.24
cc_1129 N_Z_c_1889_n A_2390_333# 0.0127078f $X=13.425 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_1130 N_Z_c_1889_n A_2601_297# 0.0127078f $X=13.425 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_1131 N_Z_c_1626_n N_VGND_c_2120_n 0.0106022f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_1132 N_Z_c_1631_n N_VGND_c_2122_n 0.0106022f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_1133 N_Z_c_1636_n N_VGND_c_2124_n 0.0106022f $X=9.435 $Y=0.495 $X2=0 $Y2=0
cc_1134 N_Z_c_1641_n N_VGND_c_2126_n 0.0106022f $X=13.575 $Y=0.495 $X2=0 $Y2=0
cc_1135 N_Z_M1044_d VGND 0.00232956f $X=1.02 $Y=0.235 $X2=0 $Y2=0
cc_1136 N_Z_M1014_s VGND 0.00232956f $X=3.32 $Y=0.235 $X2=0 $Y2=0
cc_1137 N_Z_M1010_d VGND 0.00232956f $X=5.16 $Y=0.235 $X2=0 $Y2=0
cc_1138 N_Z_M1008_s VGND 0.00232956f $X=7.46 $Y=0.235 $X2=0 $Y2=0
cc_1139 N_Z_M1018_d VGND 0.00232956f $X=9.3 $Y=0.235 $X2=0 $Y2=0
cc_1140 N_Z_M1012_s VGND 0.00232956f $X=11.6 $Y=0.235 $X2=0 $Y2=0
cc_1141 N_Z_M1033_d VGND 0.00232956f $X=13.44 $Y=0.235 $X2=0 $Y2=0
cc_1142 N_Z_M1031_s VGND 0.00232956f $X=15.74 $Y=0.235 $X2=0 $Y2=0
cc_1143 N_Z_c_1625_n VGND 0.00409585f $X=1.167 $Y=0.835 $X2=0 $Y2=0
cc_1144 N_Z_c_1626_n VGND 0.00891193f $X=1.155 $Y=0.495 $X2=0 $Y2=0
cc_1145 N_Z_c_1627_n VGND 0.00891193f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_1146 N_Z_c_1630_n VGND 0.00409585f $X=5.307 $Y=0.835 $X2=0 $Y2=0
cc_1147 N_Z_c_1631_n VGND 0.00891193f $X=5.295 $Y=0.495 $X2=0 $Y2=0
cc_1148 N_Z_c_1632_n VGND 0.00891193f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_1149 N_Z_c_1635_n VGND 0.00409585f $X=9.447 $Y=0.835 $X2=0 $Y2=0
cc_1150 N_Z_c_1636_n VGND 0.00891193f $X=9.435 $Y=0.495 $X2=0 $Y2=0
cc_1151 N_Z_c_1637_n VGND 0.00891193f $X=11.725 $Y=0.495 $X2=0 $Y2=0
cc_1152 N_Z_c_1640_n VGND 0.00409585f $X=13.587 $Y=0.835 $X2=0 $Y2=0
cc_1153 N_Z_c_1641_n VGND 0.00891193f $X=13.575 $Y=0.495 $X2=0 $Y2=0
cc_1154 N_Z_c_1642_n VGND 0.00891193f $X=15.865 $Y=0.495 $X2=0 $Y2=0
cc_1155 N_Z_c_1644_n VGND 0.00409585f $X=3.615 $Y=0.92 $X2=0 $Y2=0
cc_1156 N_Z_c_1645_n VGND 0.00409585f $X=7.755 $Y=0.92 $X2=0 $Y2=0
cc_1157 N_Z_c_1646_n VGND 0.00409585f $X=11.895 $Y=0.92 $X2=0 $Y2=0
cc_1158 N_Z_c_1647_n VGND 0.00409585f $X=16.035 $Y=0.92 $X2=0 $Y2=0
cc_1159 N_Z_c_1627_n N_VGND_c_2129_n 0.0106022f $X=3.445 $Y=0.495 $X2=0 $Y2=0
cc_1160 N_Z_c_1632_n N_VGND_c_2130_n 0.0106022f $X=7.585 $Y=0.495 $X2=0 $Y2=0
cc_1161 N_Z_c_1637_n N_VGND_c_2131_n 0.0106022f $X=11.725 $Y=0.495 $X2=0 $Y2=0
cc_1162 N_Z_c_1642_n N_VGND_c_2132_n 0.0106022f $X=15.865 $Y=0.495 $X2=0 $Y2=0
cc_1163 VGND A_109_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1164 VGND A_746_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1165 VGND A_937_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1166 VGND A_1574_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1167 VGND A_1765_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1168 VGND A_2402_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1169 VGND A_2593_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
cc_1170 VGND A_3230_47# 0.00453173f $X=16.705 $Y=-0.085 $X2=-0.19 $Y2=-0.24
