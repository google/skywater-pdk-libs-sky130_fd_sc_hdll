# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o21ba_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o21ba_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  6.440000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.540000 1.075000 6.355000 1.275000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.180000 1.075000 5.320000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.425000 1.075000 0.935000 1.285000 ;
        RECT 0.605000 1.285000 0.935000 1.705000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.155000 0.255000 1.485000 0.725000 ;
        RECT 1.155000 0.725000 2.375000 0.910000 ;
        RECT 1.155000 0.910000 1.705000 1.445000 ;
        RECT 1.155000 1.445000 2.425000 1.705000 ;
        RECT 2.045000 0.255000 2.375000 0.725000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 6.440000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.630000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 6.440000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 6.440000 0.085000 ;
      RECT 0.000000  2.635000 6.440000 2.805000 ;
      RECT 0.085000  0.265000 0.545000 0.855000 ;
      RECT 0.085000  0.855000 0.255000 1.455000 ;
      RECT 0.085000  1.455000 0.435000 1.875000 ;
      RECT 0.085000  1.875000 2.815000 2.045000 ;
      RECT 0.085000  2.045000 0.435000 2.465000 ;
      RECT 0.635000  2.215000 1.015000 2.635000 ;
      RECT 0.765000  0.085000 0.935000 0.905000 ;
      RECT 1.575000  2.215000 1.955000 2.635000 ;
      RECT 1.705000  0.085000 1.875000 0.555000 ;
      RECT 1.875000  1.080000 2.815000 1.250000 ;
      RECT 2.515000  2.215000 2.895000 2.635000 ;
      RECT 2.565000  0.085000 2.895000 0.475000 ;
      RECT 2.645000  0.645000 3.935000 0.895000 ;
      RECT 2.645000  0.895000 2.815000 1.080000 ;
      RECT 2.645000  1.445000 3.205000 1.615000 ;
      RECT 2.645000  1.615000 2.815000 1.875000 ;
      RECT 2.985000  1.075000 3.435000 1.245000 ;
      RECT 2.985000  1.245000 3.205000 1.445000 ;
      RECT 3.105000  0.255000 4.405000 0.475000 ;
      RECT 3.115000  1.795000 4.830000 1.965000 ;
      RECT 3.115000  1.965000 3.285000 2.465000 ;
      RECT 3.550000  2.135000 3.800000 2.635000 ;
      RECT 3.745000  0.895000 3.935000 1.795000 ;
      RECT 4.035000  2.135000 4.325000 2.295000 ;
      RECT 4.035000  2.295000 5.265000 2.465000 ;
      RECT 4.155000  0.475000 4.405000 0.725000 ;
      RECT 4.155000  0.725000 6.310000 0.905000 ;
      RECT 4.585000  1.445000 4.830000 1.795000 ;
      RECT 4.585000  1.965000 4.830000 2.125000 ;
      RECT 4.625000  0.085000 4.795000 0.555000 ;
      RECT 4.965000  0.255000 5.345000 0.725000 ;
      RECT 5.095000  1.455000 6.310000 1.665000 ;
      RECT 5.095000  1.665000 5.265000 2.295000 ;
      RECT 5.435000  1.835000 5.815000 2.635000 ;
      RECT 5.565000  0.085000 5.735000 0.555000 ;
      RECT 5.905000  0.265000 6.310000 0.725000 ;
      RECT 6.035000  1.665000 6.310000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21ba_4
END LIBRARY
