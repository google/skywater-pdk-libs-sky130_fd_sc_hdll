* File: sky130_fd_sc_hdll__o21ai_2.pex.spice
* Created: Thu Aug 27 19:19:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%A1 1 3 4 6 7 9 10 12 13 16 21 22
c70 21 0 1.57685e-19 $X=0.225 $Y=1.19
c71 10 0 1.33462e-19 $X=2.085 $Y=0.995
r72 21 22 8.20134 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=0.285 $Y=1.16
+ $X2=0.285 $Y2=1.445
r73 21 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.285
+ $Y=1.16 $X2=0.285 $Y2=1.16
r74 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.015
+ $Y=1.16 $X2=2.015 $Y2=1.16
r75 14 22 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.45 $Y=1.53
+ $X2=0.285 $Y2=1.53
r76 13 16 8.12016 $w=5.43e-07 $l=3.7e-07 $layer=LI1_cond $X=2.022 $Y=1.53
+ $X2=2.022 $Y2=1.16
r77 13 14 84.8128 $w=1.68e-07 $l=1.3e-06 $layer=LI1_cond $X=1.75 $Y=1.53
+ $X2=0.45 $Y2=1.53
r78 10 17 38.7084 $w=3.43e-07 $l=1.86145e-07 $layer=POLY_cond $X=2.085 $Y=0.995
+ $X2=2.04 $Y2=1.16
r79 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.085 $Y=0.995
+ $X2=2.085 $Y2=0.56
r80 7 17 45.964 $w=3.43e-07 $l=2.59808e-07 $layer=POLY_cond $X=2.02 $Y=1.41
+ $X2=2.04 $Y2=1.16
r81 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.02 $Y=1.41 $X2=2.02
+ $Y2=1.985
r82 4 27 44.0391 $w=4.22e-07 $l=2.72029e-07 $layer=POLY_cond $X=0.535 $Y=0.96
+ $X2=0.365 $Y2=1.16
r83 4 6 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=0.535 $Y=0.96 $X2=0.535
+ $Y2=0.56
r84 1 27 44.7429 $w=4.22e-07 $l=3.14245e-07 $layer=POLY_cond $X=0.51 $Y=1.41
+ $X2=0.365 $Y2=1.16
r85 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.51 $Y=1.41 $X2=0.51
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%A2 1 3 4 6 7 9 10 12 13 19 20 23
c51 1 0 1.57685e-19 $X=0.99 $Y=1.41
r52 20 21 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=1.47 $Y=1.202
+ $X2=1.495 $Y2=1.202
r53 18 20 15.424 $w=3.75e-07 $l=1.2e-07 $layer=POLY_cond $X=1.35 $Y=1.202
+ $X2=1.47 $Y2=1.202
r54 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.35
+ $Y=1.16 $X2=1.35 $Y2=1.16
r55 16 18 43.0587 $w=3.75e-07 $l=3.35e-07 $layer=POLY_cond $X=1.015 $Y=1.202
+ $X2=1.35 $Y2=1.202
r56 15 16 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.015 $Y2=1.202
r57 13 19 5.82273 $w=1.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.245 $Y=1.175
+ $X2=1.35 $Y2=1.175
r58 13 23 5.54545 $w=1.98e-07 $l=1e-07 $layer=LI1_cond $X=1.245 $Y=1.175
+ $X2=1.145 $Y2=1.175
r59 10 21 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.202
r60 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r61 7 20 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.47 $Y=1.41
+ $X2=1.47 $Y2=1.202
r62 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.47 $Y=1.41 $X2=1.47
+ $Y2=1.985
r63 4 16 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=1.202
r64 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.015 $Y=0.995
+ $X2=1.015 $Y2=0.56
r65 1 15 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.99 $Y=1.41
+ $X2=0.99 $Y2=1.202
r66 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.99 $Y=1.41 $X2=0.99
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%B1 1 3 5 6 8 9 11 13 14 16 17 19 20 21 25
+ 31 34
c55 5 0 8.49032e-20 $X=2.54 $Y=1.31
r56 21 34 2.38436 $w=2.88e-07 $l=6e-08 $layer=LI1_cond $X=3.425 $Y=1.16
+ $X2=3.425 $Y2=1.22
r57 21 31 11.127 $w=2.88e-07 $l=2.8e-07 $layer=LI1_cond $X=3.425 $Y=1.16
+ $X2=3.425 $Y2=0.88
r58 21 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.365
+ $Y=1.16 $X2=3.365 $Y2=1.16
r59 20 31 1.19218 $w=2.88e-07 $l=3e-08 $layer=LI1_cond $X=3.425 $Y=0.85
+ $X2=3.425 $Y2=0.88
r60 18 25 42.841 $w=3.3e-07 $l=2.45e-07 $layer=POLY_cond $X=3.12 $Y=1.16
+ $X2=3.365 $Y2=1.16
r61 18 19 6.791 $w=3.3e-07 $l=2.82843e-07 $layer=POLY_cond $X=3.12 $Y=1.16
+ $X2=2.92 $Y2=0.96
r62 14 19 18.3167 $w=1.8e-07 $l=4.97494e-07 $layer=POLY_cond $X=3.02 $Y=1.41
+ $X2=2.92 $Y2=0.96
r63 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.02 $Y=1.41
+ $X2=3.02 $Y2=1.985
r64 11 19 18.3167 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.995 $Y=0.96
+ $X2=2.92 $Y2=0.96
r65 11 13 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.995 $Y=0.96
+ $X2=2.995 $Y2=0.56
r66 10 17 3.07963 $w=2.05e-07 $l=1e-07 $layer=POLY_cond $X=2.64 $Y=1.062
+ $X2=2.54 $Y2=1.062
r67 9 19 6.791 $w=2.05e-07 $l=1.02e-07 $layer=POLY_cond $X=2.92 $Y=1.062
+ $X2=2.92 $Y2=0.96
r68 9 10 90.5772 $w=2.05e-07 $l=2.8e-07 $layer=POLY_cond $X=2.92 $Y=1.062
+ $X2=2.64 $Y2=1.062
r69 6 8 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.54 $Y=1.41 $X2=2.54
+ $Y2=1.985
r70 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.54 $Y=1.31 $X2=2.54
+ $Y2=1.41
r71 4 17 23.2339 $w=1.75e-07 $l=1.03e-07 $layer=POLY_cond $X=2.54 $Y=1.165
+ $X2=2.54 $Y2=1.062
r72 4 5 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=2.54 $Y=1.165 $X2=2.54
+ $Y2=1.31
r73 1 17 23.2339 $w=1.75e-07 $l=1.13816e-07 $layer=POLY_cond $X=2.515 $Y=0.96
+ $X2=2.54 $Y2=1.062
r74 1 3 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.515 $Y=0.96 $X2=2.515
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%VPWR 1 2 3 10 12 16 18 20 22 24 29 38 42
r54 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r55 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r56 33 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r57 33 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r59 30 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.44 $Y=2.72 $X2=2.25
+ $Y2=2.72
r60 30 32 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=2.44 $Y=2.72
+ $X2=2.99 $Y2=2.72
r61 29 41 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=3.28 $Y=2.72 $X2=3.48
+ $Y2=2.72
r62 29 32 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=3.28 $Y=2.72
+ $X2=2.99 $Y2=2.72
r63 28 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.07 $Y2=2.72
r64 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r65 25 35 4.75569 $w=1.7e-07 $l=2.18e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.217 $Y2=2.72
r66 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.435 $Y=2.72
+ $X2=0.69 $Y2=2.72
r67 24 38 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.06 $Y=2.72 $X2=2.25
+ $Y2=2.72
r68 24 27 89.3797 $w=1.68e-07 $l=1.37e-06 $layer=LI1_cond $X=2.06 $Y=2.72
+ $X2=0.69 $Y2=2.72
r69 22 28 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.225 $Y=2.72
+ $X2=0.69 $Y2=2.72
r70 22 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 18 41 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.48 $Y2=2.72
r72 18 20 41.4879 $w=2.48e-07 $l=9e-07 $layer=LI1_cond $X=3.405 $Y=2.635
+ $X2=3.405 $Y2=1.735
r73 14 38 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.25 $Y=2.635
+ $X2=2.25 $Y2=2.72
r74 14 16 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.25 $Y=2.635
+ $X2=2.25 $Y2=2.34
r75 10 35 3.01048 $w=3.3e-07 $l=1.08305e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.217 $Y2=2.72
r76 10 12 23.9219 $w=3.28e-07 $l=6.85e-07 $layer=LI1_cond $X=0.27 $Y=2.635
+ $X2=0.27 $Y2=1.95
r77 3 20 300 $w=1.7e-07 $l=3.58852e-07 $layer=licon1_PDIFF $count=2 $X=3.11
+ $Y=1.485 $X2=3.365 $Y2=1.735
r78 2 16 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=2.11
+ $Y=1.485 $X2=2.275 $Y2=2.34
r79 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.145
+ $Y=1.485 $X2=0.27 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%A_120_297# 1 2 9 11 12 14
r21 11 14 1.386 $w=1.7e-07 $l=1.28938e-07 $layer=LI1_cond $X=1.675 $Y=2.38
+ $X2=1.77 $Y2=2.3
r22 11 12 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=1.675 $Y=2.38
+ $X2=0.875 $Y2=2.38
r23 7 12 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.765 $Y=2.295
+ $X2=0.875 $Y2=2.38
r24 7 9 18.0724 $w=2.18e-07 $l=3.45e-07 $layer=LI1_cond $X=0.765 $Y=2.295
+ $X2=0.765 $Y2=1.95
r25 2 14 600 $w=1.7e-07 $l=9.09519e-07 $layer=licon1_PDIFF $count=1 $X=1.56
+ $Y=1.485 $X2=1.76 $Y2=2.3
r26 1 9 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=0.6
+ $Y=1.485 $X2=0.75 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%Y 1 2 3 10 13 14 15 16 23 26 30 34 44 45
c45 34 0 1.33462e-19 $X=2.78 $Y=0.76
r46 44 45 7.1142 $w=3.38e-07 $l=1.35e-07 $layer=LI1_cond $X=1.26 $Y=1.955
+ $X2=1.395 $Y2=1.955
r47 34 37 24.1596 $w=4.13e-07 $l=8.7e-07 $layer=LI1_cond $X=2.902 $Y=0.76
+ $X2=2.902 $Y2=1.63
r48 26 45 21.5657 $w=1.78e-07 $l=3.5e-07 $layer=LI1_cond $X=1.745 $Y=1.875
+ $X2=1.395 $Y2=1.875
r49 16 23 4.46552 $w=1.8e-07 $l=2.07e-07 $layer=LI1_cond $X=2.902 $Y=1.875
+ $X2=2.695 $Y2=1.875
r50 16 37 4.18249 $w=5.78e-07 $l=1.55e-07 $layer=LI1_cond $X=2.902 $Y=1.785
+ $X2=2.902 $Y2=1.63
r51 16 23 0.184848 $w=1.78e-07 $l=3e-09 $layer=LI1_cond $X=2.692 $Y=1.875
+ $X2=2.695 $Y2=1.875
r52 16 30 25.0778 $w=1.78e-07 $l=4.07e-07 $layer=LI1_cond $X=2.692 $Y=1.875
+ $X2=2.285 $Y2=1.875
r53 15 30 1.23232 $w=1.78e-07 $l=2e-08 $layer=LI1_cond $X=2.265 $Y=1.875
+ $X2=2.285 $Y2=1.875
r54 14 15 31.4242 $w=1.78e-07 $l=5.1e-07 $layer=LI1_cond $X=1.755 $Y=1.875
+ $X2=2.265 $Y2=1.875
r55 14 26 0.616162 $w=1.78e-07 $l=1e-08 $layer=LI1_cond $X=1.755 $Y=1.875
+ $X2=1.745 $Y2=1.875
r56 13 44 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=1.245 $Y=1.955
+ $X2=1.26 $Y2=1.955
r57 13 40 0.508431 $w=3.38e-07 $l=1.5e-08 $layer=LI1_cond $X=1.245 $Y=1.955
+ $X2=1.23 $Y2=1.955
r58 10 16 2.46455 $w=4.15e-07 $l=9e-08 $layer=LI1_cond $X=2.902 $Y=1.965
+ $X2=2.902 $Y2=1.875
r59 10 12 3.6747 $w=4.15e-07 $l=1.25e-07 $layer=LI1_cond $X=2.902 $Y=1.965
+ $X2=2.902 $Y2=2.09
r60 3 37 600 $w=1.7e-07 $l=2.10357e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.78 $Y2=1.63
r61 3 12 600 $w=1.7e-07 $l=6.75851e-07 $layer=licon1_PDIFF $count=1 $X=2.63
+ $Y=1.485 $X2=2.78 $Y2=2.09
r62 2 40 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=1.08
+ $Y=1.485 $X2=1.23 $Y2=1.96
r63 1 34 182 $w=1.7e-07 $l=6.12679e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.235 $X2=2.78 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%A_29_47# 1 2 3 4 15 17 18 21 23 25 26 27
+ 29 32
r69 32 35 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.405 $Y=0.34
+ $X2=3.405 $Y2=0.43
r70 28 31 5.12568 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.465 $Y=0.34
+ $X2=2.3 $Y2=0.34
r71 27 32 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.28 $Y=0.34
+ $X2=3.405 $Y2=0.34
r72 27 28 53.1711 $w=1.68e-07 $l=8.15e-07 $layer=LI1_cond $X=3.28 $Y=0.34
+ $X2=2.465 $Y2=0.34
r73 25 31 2.6405 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.3 $Y=0.425 $X2=2.3
+ $Y2=0.34
r74 25 26 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=2.3 $Y=0.425 $X2=2.3
+ $Y2=0.715
r75 24 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.395 $Y=0.8
+ $X2=1.205 $Y2=0.8
r76 23 26 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.135 $Y=0.8
+ $X2=2.3 $Y2=0.715
r77 23 24 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=2.135 $Y=0.8
+ $X2=1.395 $Y2=0.8
r78 19 29 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.205 $Y=0.715
+ $X2=1.205 $Y2=0.8
r79 19 21 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.205 $Y=0.715
+ $X2=1.205 $Y2=0.4
r80 17 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.015 $Y=0.8
+ $X2=1.205 $Y2=0.8
r81 17 18 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=1.015 $Y=0.8
+ $X2=0.435 $Y2=0.8
r82 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.27 $Y=0.715
+ $X2=0.435 $Y2=0.8
r83 13 15 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=0.27 $Y=0.715
+ $X2=0.27 $Y2=0.4
r84 4 35 182 $w=1.7e-07 $l=3.80197e-07 $layer=licon1_NDIFF $count=1 $X=3.07
+ $Y=0.235 $X2=3.365 $Y2=0.43
r85 3 31 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=2.16
+ $Y=0.235 $X2=2.3 $Y2=0.4
r86 2 21 91 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=2 $X=1.09
+ $Y=0.235 $X2=1.23 $Y2=0.4
r87 1 15 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.145
+ $Y=0.235 $X2=0.27 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21AI_2%VGND 1 2 11 15 18 19 20 30 31 34
r52 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r53 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 28 31 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r55 27 30 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.07 $Y=0 $X2=3.45
+ $Y2=0
r56 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r57 25 28 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r58 25 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=0.69
+ $Y2=0
r59 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r60 22 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.835 $Y=0 $X2=0.75
+ $Y2=0
r61 22 24 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=0.835 $Y=0 $X2=1.61
+ $Y2=0
r62 20 35 0.132312 $w=4.8e-07 $l=4.65e-07 $layer=MET1_cond $X=0.225 $Y=0
+ $X2=0.69 $Y2=0
r63 18 24 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.61
+ $Y2=0
r64 18 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.675 $Y=0 $X2=1.76
+ $Y2=0
r65 17 27 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.845 $Y=0 $X2=2.07
+ $Y2=0
r66 17 19 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.845 $Y=0 $X2=1.76
+ $Y2=0
r67 13 19 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0
r68 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.76 $Y=0.085
+ $X2=1.76 $Y2=0.38
r69 9 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=0.085 $X2=0.75
+ $Y2=0
r70 9 11 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.75 $Y=0.085
+ $X2=0.75 $Y2=0.38
r71 2 15 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.57
+ $Y=0.235 $X2=1.76 $Y2=0.38
r72 1 11 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=0.61
+ $Y=0.235 $X2=0.75 $Y2=0.38
.ends

