* File: sky130_fd_sc_hdll__o22a_4.pex.spice
* Created: Thu Aug 27 19:21:14 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A_96_21# 1 2 3 4 13 15 16 18 19 21 22 24 25
+ 27 28 30 31 33 34 36 37 46 48 50 51 52 53 57 59 61 62 63 68 81
c146 57 0 1.91072e-19 $X=4.155 $Y=0.73
r147 81 82 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r148 78 79 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.495 $Y=1.202
+ $X2=1.52 $Y2=1.202
r149 77 78 57.6586 $w=3.72e-07 $l=4.45e-07 $layer=POLY_cond $X=1.05 $Y=1.202
+ $X2=1.495 $Y2=1.202
r150 76 77 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=1.025 $Y=1.202
+ $X2=1.05 $Y2=1.202
r151 73 74 3.23925 $w=3.72e-07 $l=2.5e-08 $layer=POLY_cond $X=0.555 $Y=1.202
+ $X2=0.58 $Y2=1.202
r152 68 71 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=5.645 $Y=1.87
+ $X2=5.645 $Y2=1.96
r153 63 66 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=3.685 $Y=1.87
+ $X2=3.685 $Y2=1.96
r154 60 63 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.81 $Y=1.87
+ $X2=3.685 $Y2=1.87
r155 59 68 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.52 $Y=1.87
+ $X2=5.645 $Y2=1.87
r156 59 60 111.561 $w=1.68e-07 $l=1.71e-06 $layer=LI1_cond $X=5.52 $Y=1.87
+ $X2=3.81 $Y2=1.87
r157 55 57 41.6652 $w=2.58e-07 $l=9.4e-07 $layer=LI1_cond $X=3.215 $Y=0.775
+ $X2=4.155 $Y2=0.775
r158 53 62 7.14225 $w=2.58e-07 $l=1.3e-07 $layer=LI1_cond $X=2.745 $Y=0.775
+ $X2=2.615 $Y2=0.775
r159 53 55 20.8326 $w=2.58e-07 $l=4.7e-07 $layer=LI1_cond $X=2.745 $Y=0.775
+ $X2=3.215 $Y2=0.775
r160 51 63 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.56 $Y=1.87
+ $X2=3.685 $Y2=1.87
r161 51 52 73.7219 $w=1.68e-07 $l=1.13e-06 $layer=LI1_cond $X=3.56 $Y=1.87
+ $X2=2.43 $Y2=1.87
r162 50 62 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.43 $Y=0.82
+ $X2=2.615 $Y2=0.82
r163 48 61 3.53812 $w=3.1e-07 $l=1.09545e-07 $layer=LI1_cond $X=2.285 $Y=1.075
+ $X2=2.265 $Y2=1.175
r164 47 50 7.43784 $w=1.7e-07 $l=1.8262e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.43 $Y2=0.82
r165 47 48 6.7557 $w=2.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.285 $Y=0.905
+ $X2=2.285 $Y2=1.075
r166 46 52 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=2.265 $Y=1.785
+ $X2=2.43 $Y2=1.87
r167 45 61 3.53812 $w=3.1e-07 $l=1e-07 $layer=LI1_cond $X=2.265 $Y=1.275
+ $X2=2.265 $Y2=1.175
r168 45 46 17.8105 $w=3.28e-07 $l=5.1e-07 $layer=LI1_cond $X=2.265 $Y=1.275
+ $X2=2.265 $Y2=1.785
r169 44 81 14.9005 $w=3.72e-07 $l=1.15e-07 $layer=POLY_cond $X=1.875 $Y=1.202
+ $X2=1.99 $Y2=1.202
r170 44 79 45.9973 $w=3.72e-07 $l=3.55e-07 $layer=POLY_cond $X=1.875 $Y=1.202
+ $X2=1.52 $Y2=1.202
r171 43 44 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.875
+ $Y=1.16 $X2=1.875 $Y2=1.16
r172 40 76 41.4624 $w=3.72e-07 $l=3.2e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=1.025 $Y2=1.202
r173 40 74 16.1962 $w=3.72e-07 $l=1.25e-07 $layer=POLY_cond $X=0.705 $Y=1.202
+ $X2=0.58 $Y2=1.202
r174 39 43 64.8818 $w=1.98e-07 $l=1.17e-06 $layer=LI1_cond $X=0.705 $Y=1.175
+ $X2=1.875 $Y2=1.175
r175 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.705
+ $Y=1.16 $X2=0.705 $Y2=1.16
r176 37 61 2.95888 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.1 $Y=1.175
+ $X2=2.265 $Y2=1.175
r177 37 43 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=2.1 $Y=1.175
+ $X2=1.875 $Y2=1.175
r178 34 82 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.202
r179 34 36 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r180 31 81 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.202
r181 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.985
r182 28 79 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.202
r183 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.52 $Y=1.41
+ $X2=1.52 $Y2=1.985
r184 25 78 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=1.202
r185 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.495 $Y=0.995
+ $X2=1.495 $Y2=0.56
r186 22 77 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.05 $Y2=1.202
r187 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.05 $Y=1.41
+ $X2=1.05 $Y2=1.985
r188 19 76 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=1.202
r189 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.025 $Y=0.995
+ $X2=1.025 $Y2=0.56
r190 16 74 19.7411 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.58 $Y2=1.202
r191 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.58 $Y=1.41
+ $X2=0.58 $Y2=1.985
r192 13 73 24.0971 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=1.202
r193 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.555 $Y=0.995
+ $X2=0.555 $Y2=0.56
r194 4 71 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=5.5
+ $Y=1.485 $X2=5.645 $Y2=1.96
r195 3 66 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=3.54
+ $Y=1.485 $X2=3.685 $Y2=1.96
r196 2 57 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=4.02
+ $Y=0.235 $X2=4.155 $Y2=0.73
r197 1 55 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.08
+ $Y=0.235 $X2=3.215 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%B1 1 3 4 6 7 9 10 12 13 17 20 29 31
c77 10 0 1.91072e-19 $X=4.415 $Y=0.995
r78 24 31 11.0969 $w=5.38e-07 $l=2.25e-07 $layer=LI1_cond $X=2.955 $Y=1.345
+ $X2=3.18 $Y2=1.345
r79 24 29 2.9902 $w=5.38e-07 $l=1.35e-07 $layer=LI1_cond $X=2.955 $Y=1.345
+ $X2=2.82 $Y2=1.345
r80 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.955
+ $Y=1.16 $X2=2.955 $Y2=1.16
r81 20 29 1.55047 $w=5.38e-07 $l=7e-08 $layer=LI1_cond $X=2.75 $Y=1.345 $X2=2.82
+ $Y2=1.345
r82 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.365
+ $Y=1.16 $X2=4.365 $Y2=1.16
r83 15 17 9.66018 $w=3.38e-07 $l=2.85e-07 $layer=LI1_cond $X=4.37 $Y=1.445
+ $X2=4.37 $Y2=1.16
r84 13 15 7.85115 $w=1.7e-07 $l=2.08207e-07 $layer=LI1_cond $X=4.2 $Y=1.53
+ $X2=4.37 $Y2=1.445
r85 13 31 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=4.2 $Y=1.53
+ $X2=3.18 $Y2=1.53
r86 10 18 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.39 $Y2=1.16
r87 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.415 $Y=0.995
+ $X2=4.415 $Y2=0.56
r88 7 18 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.39 $Y=1.41
+ $X2=4.39 $Y2=1.16
r89 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.39 $Y=1.41 $X2=4.39
+ $Y2=1.985
r90 4 23 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=2.98 $Y2=1.16
r91 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=0.56
r92 1 23 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.98 $Y=1.41
+ $X2=2.98 $Y2=1.16
r93 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.98 $Y=1.41 $X2=2.98
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%B2 1 3 4 6 7 9 10 12 13 20 24
r43 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.92 $Y=1.202
+ $X2=3.945 $Y2=1.202
r44 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.685 $Y=1.202
+ $X2=3.92 $Y2=1.202
r45 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.685
+ $Y=1.16 $X2=3.685 $Y2=1.16
r46 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=3.45 $Y=1.202
+ $X2=3.685 $Y2=1.202
r47 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.425 $Y=1.202
+ $X2=3.45 $Y2=1.202
r48 13 24 4.71364 $w=1.98e-07 $l=8.5e-08 $layer=LI1_cond $X=3.77 $Y=1.175
+ $X2=3.685 $Y2=1.175
r49 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.945 $Y=0.995
+ $X2=3.945 $Y2=0.56
r51 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.92 $Y=1.41
+ $X2=3.92 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.92 $Y=1.41 $X2=3.92
+ $Y2=1.985
r53 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.45 $Y=1.41
+ $X2=3.45 $Y2=1.202
r54 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.45 $Y=1.41 $X2=3.45
+ $Y2=1.985
r55 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=1.202
r56 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.425 $Y=0.995
+ $X2=3.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A1 1 3 4 6 7 9 10 12 13 16 21 22 32
c75 7 0 3.17292e-19 $X=6.35 $Y=1.41
c76 4 0 2.98731e-20 $X=4.965 $Y=0.995
r77 30 32 2.44 $w=2e-07 $l=4e-08 $layer=LI1_cond $X=6.285 $Y=1.175 $X2=6.325
+ $Y2=1.175
r78 28 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.325
+ $Y=1.16 $X2=6.325 $Y2=1.16
r79 22 30 3.49408 $w=2e-07 $l=1.05e-07 $layer=LI1_cond $X=6.18 $Y=1.175
+ $X2=6.285 $Y2=1.175
r80 22 32 1.342 $w=2e-07 $l=2.2e-08 $layer=LI1_cond $X=6.347 $Y=1.175 $X2=6.325
+ $Y2=1.175
r81 21 22 8.07595 $w=2.53e-07 $l=1.7e-07 $layer=LI1_cond $X=6.18 $Y=1.445
+ $X2=6.18 $Y2=1.275
r82 16 19 10.1525 $w=4.18e-07 $l=3.7e-07 $layer=LI1_cond $X=4.92 $Y=1.16
+ $X2=4.92 $Y2=1.53
r83 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.915
+ $Y=1.16 $X2=4.915 $Y2=1.16
r84 14 19 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=5.13 $Y=1.53 $X2=4.92
+ $Y2=1.53
r85 13 21 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=6.075 $Y=1.53
+ $X2=6.18 $Y2=1.445
r86 13 14 61.6524 $w=1.68e-07 $l=9.45e-07 $layer=LI1_cond $X=6.075 $Y=1.53
+ $X2=5.13 $Y2=1.53
r87 10 28 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.35 $Y2=1.16
r88 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.375 $Y=0.995
+ $X2=6.375 $Y2=0.56
r89 7 28 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=6.35 $Y=1.41
+ $X2=6.35 $Y2=1.16
r90 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.35 $Y=1.41 $X2=6.35
+ $Y2=1.985
r91 4 17 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.94 $Y2=1.16
r92 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.965 $Y=0.995
+ $X2=4.965 $Y2=0.56
r93 1 17 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=4.94 $Y=1.41
+ $X2=4.94 $Y2=1.16
r94 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.94 $Y=1.41 $X2=4.94
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A2 1 3 4 6 7 9 10 12 13 20 23
c46 13 0 1.74489e-19 $X=5.725 $Y=1.105
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.88 $Y=1.202
+ $X2=5.905 $Y2=1.202
r48 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=5.645 $Y=1.202
+ $X2=5.88 $Y2=1.202
r49 18 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.645
+ $Y=1.16 $X2=5.645 $Y2=1.16
r50 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=5.41 $Y=1.202
+ $X2=5.645 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=5.385 $Y=1.202
+ $X2=5.41 $Y2=1.202
r52 13 23 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=5.81 $Y=1.175
+ $X2=5.575 $Y2=1.175
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.905 $Y=0.995
+ $X2=5.905 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.905 $Y=0.995
+ $X2=5.905 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.88 $Y=1.41
+ $X2=5.88 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.88 $Y=1.41 $X2=5.88
+ $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.41 $Y=1.41
+ $X2=5.41 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.41 $Y=1.41 $X2=5.41
+ $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.385 $Y=0.995
+ $X2=5.385 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.385 $Y=0.995
+ $X2=5.385 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%VPWR 1 2 3 4 5 16 18 22 26 28 30 35 36 38
+ 39 40 57 70 73 76
r90 75 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r91 72 73 9.97279 $w=6.78e-07 $l=1.25e-07 $layer=LI1_cond $X=2.745 $Y=2.465
+ $X2=2.87 $Y2=2.465
r92 68 72 3.78172 $w=6.78e-07 $l=2.15e-07 $layer=LI1_cond $X=2.53 $Y=2.465
+ $X2=2.745 $Y2=2.465
r93 68 70 15.3376 $w=6.78e-07 $l=4.3e-07 $layer=LI1_cond $X=2.53 $Y=2.465
+ $X2=2.1 $Y2=2.465
r94 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r95 63 76 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r96 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r97 60 63 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r98 59 62 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=6.21 $Y2=2.72
r99 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r100 57 75 3.60244 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.702 $Y2=2.72
r101 57 62 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.505 $Y=2.72
+ $X2=6.21 $Y2=2.72
r102 56 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r103 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r104 53 56 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r105 53 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r106 52 55 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=4.37 $Y2=2.72
r107 52 73 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.87 $Y2=2.72
r108 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r109 49 69 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r110 48 70 1.95722 $w=1.68e-07 $l=3e-08 $layer=LI1_cond $X=2.07 $Y=2.72 $X2=2.1
+ $Y2=2.72
r111 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 45 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r114 42 65 3.90382 $w=1.7e-07 $l=2.35e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=0.235 $Y2=2.72
r115 42 44 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.47 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 40 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r117 40 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r118 39 59 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.665 $Y=2.72
+ $X2=4.83 $Y2=2.72
r119 38 55 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=4.5 $Y=2.72
+ $X2=4.37 $Y2=2.72
r120 38 39 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.5 $Y=2.72
+ $X2=4.665 $Y2=2.72
r121 35 44 0.652406 $w=1.68e-07 $l=1e-08 $layer=LI1_cond $X=1.16 $Y=2.72
+ $X2=1.15 $Y2=2.72
r122 35 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.16 $Y=2.72
+ $X2=1.285 $Y2=2.72
r123 34 48 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=2.07 $Y2=2.72
r124 34 36 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.41 $Y=2.72
+ $X2=1.285 $Y2=2.72
r125 30 33 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.607 $Y=1.62
+ $X2=6.607 $Y2=2.3
r126 28 75 3.29157 $w=2.05e-07 $l=1.30767e-07 $layer=LI1_cond $X=6.607 $Y=2.635
+ $X2=6.702 $Y2=2.72
r127 28 33 18.1242 $w=2.03e-07 $l=3.35e-07 $layer=LI1_cond $X=6.607 $Y=2.635
+ $X2=6.607 $Y2=2.3
r128 24 39 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.665 $Y=2.635
+ $X2=4.665 $Y2=2.72
r129 24 26 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=4.665 $Y=2.635
+ $X2=4.665 $Y2=2.3
r130 20 36 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=2.72
r131 20 22 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=1.285 $Y=2.635
+ $X2=1.285 $Y2=1.99
r132 16 65 3.23934 $w=2.5e-07 $l=1.46458e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.235 $Y2=2.72
r133 16 18 29.733 $w=2.48e-07 $l=6.45e-07 $layer=LI1_cond $X=0.345 $Y=2.635
+ $X2=0.345 $Y2=1.99
r134 5 33 400 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.485 $X2=6.59 $Y2=2.3
r135 5 30 400 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=6.44
+ $Y=1.485 $X2=6.59 $Y2=1.62
r136 4 26 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.48
+ $Y=1.485 $X2=4.625 $Y2=2.3
r137 3 72 300 $w=1.7e-07 $l=1.09827e-06 $layer=licon1_PDIFF $count=2 $X=2.08
+ $Y=1.485 $X2=2.745 $Y2=2.3
r138 2 22 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=1.14
+ $Y=1.485 $X2=1.285 $Y2=1.99
r139 1 18 300 $w=1.7e-07 $l=5.72931e-07 $layer=licon1_PDIFF $count=2 $X=0.2
+ $Y=1.485 $X2=0.345 $Y2=1.99
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%X 1 2 3 4 13 14 15 16 19 23 27 29 33 37 43
+ 44 45
r73 42 45 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=0.227 $Y=1.445
+ $X2=0.227 $Y2=1.19
r74 41 45 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=0.227 $Y=0.905
+ $X2=0.227 $Y2=1.19
r75 37 39 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=1.755 $Y=1.62
+ $X2=1.755 $Y2=2.3
r76 35 37 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=1.755 $Y=1.615
+ $X2=1.755 $Y2=1.62
r77 31 33 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.73 $Y=0.725
+ $X2=1.73 $Y2=0.39
r78 30 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.98 $Y=0.815
+ $X2=0.79 $Y2=0.815
r79 29 31 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=1.54 $Y=0.815
+ $X2=1.73 $Y2=0.725
r80 29 30 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.54 $Y=0.815
+ $X2=0.98 $Y2=0.815
r81 28 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.94 $Y=1.53
+ $X2=0.815 $Y2=1.53
r82 27 35 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.63 $Y=1.53
+ $X2=1.755 $Y2=1.615
r83 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.63 $Y=1.53 $X2=0.94
+ $Y2=1.53
r84 23 25 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=0.815 $Y=1.62
+ $X2=0.815 $Y2=2.3
r85 21 44 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=1.615
+ $X2=0.815 $Y2=1.53
r86 21 23 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.815 $Y=1.615
+ $X2=0.815 $Y2=1.62
r87 17 43 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=0.79 $Y=0.725 $X2=0.79
+ $Y2=0.815
r88 17 19 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.79 $Y=0.725
+ $X2=0.79 $Y2=0.39
r89 16 42 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=0.37 $Y=1.53
+ $X2=0.227 $Y2=1.445
r90 15 44 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.69 $Y=1.53
+ $X2=0.815 $Y2=1.53
r91 15 16 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.69 $Y=1.53 $X2=0.37
+ $Y2=1.53
r92 14 41 7.27854 $w=1.8e-07 $l=1.82535e-07 $layer=LI1_cond $X=0.37 $Y=0.815
+ $X2=0.227 $Y2=0.905
r93 13 43 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=0.6 $Y=0.815 $X2=0.79
+ $Y2=0.815
r94 13 14 14.1717 $w=1.78e-07 $l=2.3e-07 $layer=LI1_cond $X=0.6 $Y=0.815
+ $X2=0.37 $Y2=0.815
r95 4 39 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=2.3
r96 4 37 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.61
+ $Y=1.485 $X2=1.755 $Y2=1.62
r97 3 25 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.485 $X2=0.815 $Y2=2.3
r98 3 23 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.67
+ $Y=1.485 $X2=0.815 $Y2=1.62
r99 2 33 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.57
+ $Y=0.235 $X2=1.755 $Y2=0.39
r100 1 19 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.63
+ $Y=0.235 $X2=0.815 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A_614_297# 1 2 7 10 15
r21 15 17 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.155 $Y=2.3 $X2=4.155
+ $Y2=2.38
r22 10 12 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=3.215 $Y=2.3 $X2=3.215
+ $Y2=2.38
r23 8 12 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.34 $Y=2.38
+ $X2=3.215 $Y2=2.38
r24 7 17 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.03 $Y=2.38
+ $X2=4.155 $Y2=2.38
r25 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.03 $Y=2.38 $X2=3.34
+ $Y2=2.38
r26 2 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.01
+ $Y=1.485 $X2=4.155 $Y2=2.3
r27 1 10 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.07
+ $Y=1.485 $X2=3.215 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A_1006_297# 1 2 7 11 14
c17 11 0 1.42804e-19 $X=6.115 $Y=1.96
r18 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=5.175 $Y=2.3 $X2=5.175
+ $Y2=2.38
r19 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=6.115 $Y=2.295
+ $X2=6.115 $Y2=1.96
r20 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.3 $Y=2.38 $X2=5.175
+ $Y2=2.38
r21 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=5.99 $Y=2.38
+ $X2=6.115 $Y2=2.295
r22 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=5.99 $Y=2.38 $X2=5.3
+ $Y2=2.38
r23 2 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=5.97
+ $Y=1.485 $X2=6.115 $Y2=1.96
r24 1 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.03
+ $Y=1.485 $X2=5.175 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 43 44 46 47 48 50 67 68
r102 71 74 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=0.23 $Y=0
+ $X2=0.345 $Y2=0
r103 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r104 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r105 64 65 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r106 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r107 61 62 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r108 59 62 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r109 58 61 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=4.83
+ $Y2=0
r110 58 59 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r111 56 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r112 55 56 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r113 53 56 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r114 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r115 50 74 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=0.43 $Y=0 $X2=0.345
+ $Y2=0
r116 50 52 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=0.43 $Y=0 $X2=1.15
+ $Y2=0
r117 48 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r118 48 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r119 46 64 18.2674 $w=1.68e-07 $l=2.8e-07 $layer=LI1_cond $X=6.03 $Y=0 $X2=5.75
+ $Y2=0
r120 46 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.03 $Y=0 $X2=6.115
+ $Y2=0
r121 45 67 30.6631 $w=1.68e-07 $l=4.7e-07 $layer=LI1_cond $X=6.2 $Y=0 $X2=6.67
+ $Y2=0
r122 45 47 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.2 $Y=0 $X2=6.115
+ $Y2=0
r123 43 61 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=5.09 $Y=0 $X2=4.83
+ $Y2=0
r124 43 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.09 $Y=0 $X2=5.175
+ $Y2=0
r125 42 64 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.75
+ $Y2=0
r126 42 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.26 $Y=0 $X2=5.175
+ $Y2=0
r127 40 55 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.07
+ $Y2=0
r128 40 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0 $X2=2.225
+ $Y2=0
r129 39 58 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.53
+ $Y2=0
r130 39 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.225
+ $Y2=0
r131 37 52 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.15
+ $Y2=0
r132 37 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0 $X2=1.285
+ $Y2=0
r133 36 55 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.37 $Y=0 $X2=2.07
+ $Y2=0
r134 36 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.37 $Y=0 $X2=1.285
+ $Y2=0
r135 32 47 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.115 $Y=0.085
+ $X2=6.115 $Y2=0
r136 32 34 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=6.115 $Y=0.085
+ $X2=6.115 $Y2=0.39
r137 28 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.175 $Y=0.085
+ $X2=5.175 $Y2=0
r138 28 30 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.175 $Y=0.085
+ $X2=5.175 $Y2=0.39
r139 24 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0
r140 24 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.225 $Y=0.085
+ $X2=2.225 $Y2=0.39
r141 20 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0
r142 20 22 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.285 $Y=0.085
+ $X2=1.285 $Y2=0.39
r143 16 74 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0
r144 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.345 $Y=0.085
+ $X2=0.345 $Y2=0.39
r145 5 34 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.98
+ $Y=0.235 $X2=6.115 $Y2=0.39
r146 4 30 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=5.04
+ $Y=0.235 $X2=5.175 $Y2=0.39
r147 3 26 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.225 $Y2=0.39
r148 2 22 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=1.1
+ $Y=0.235 $X2=1.285 $Y2=0.39
r149 1 18 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=0.2
+ $Y=0.235 $X2=0.345 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O22A_4%A_524_47# 1 2 3 4 5 16 22 26 27 30 32 36 40
c69 40 0 2.98731e-20 $X=5.62 $Y=0.815
r70 34 36 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.56 $Y=0.725
+ $X2=6.56 $Y2=0.39
r71 33 40 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=5.81 $Y=0.815
+ $X2=5.62 $Y2=0.815
r72 32 34 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=6.37 $Y=0.815
+ $X2=6.56 $Y2=0.725
r73 32 33 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=6.37 $Y=0.815
+ $X2=5.81 $Y2=0.815
r74 28 40 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=5.62 $Y=0.725 $X2=5.62
+ $Y2=0.815
r75 28 30 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.62 $Y=0.725
+ $X2=5.62 $Y2=0.39
r76 26 40 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=5.43 $Y=0.82
+ $X2=5.62 $Y2=0.815
r77 26 27 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.43 $Y=0.82
+ $X2=4.87 $Y2=0.82
r78 23 27 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=4.705 $Y=0.735
+ $X2=4.87 $Y2=0.82
r79 23 25 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=4.705 $Y=0.735
+ $X2=4.705 $Y2=0.73
r80 22 39 2.87089 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=4.705 $Y=0.475
+ $X2=4.705 $Y2=0.365
r81 22 25 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=4.705 $Y=0.475
+ $X2=4.705 $Y2=0.73
r82 18 21 49.2407 $w=2.18e-07 $l=9.4e-07 $layer=LI1_cond $X=2.745 $Y=0.365
+ $X2=3.685 $Y2=0.365
r83 16 39 4.30634 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=4.54 $Y=0.365
+ $X2=4.705 $Y2=0.365
r84 16 21 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=4.54 $Y=0.365
+ $X2=3.685 $Y2=0.365
r85 5 36 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=6.45
+ $Y=0.235 $X2=6.585 $Y2=0.39
r86 4 30 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.46
+ $Y=0.235 $X2=5.645 $Y2=0.39
r87 3 39 182 $w=1.7e-07 $l=2.45561e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.235 $X2=4.67 $Y2=0.39
r88 3 25 182 $w=1.7e-07 $l=5.78035e-07 $layer=licon1_NDIFF $count=1 $X=4.49
+ $Y=0.235 $X2=4.67 $Y2=0.73
r89 2 21 182 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=1 $X=3.5
+ $Y=0.235 $X2=3.685 $Y2=0.39
r90 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.62
+ $Y=0.235 $X2=2.745 $Y2=0.39
.ends

