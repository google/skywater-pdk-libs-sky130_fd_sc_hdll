* File: sky130_fd_sc_hdll__and2_8.pex.spice
* Created: Thu Aug 27 18:57:24 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2_8%B 1 3 4 6 7 9 10 12 13 14 15 16 18 19 24 28
c81 18 0 1.22108e-19 $X=1.795 $Y=1.465
c82 15 0 1.48863e-19 $X=1.705 $Y=1.55
c83 10 0 1.60887e-19 $X=1.905 $Y=1.41
c84 7 0 7.31881e-20 $X=1.82 $Y=0.995
r85 24 27 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.835 $Y=1.16
+ $X2=1.835 $Y2=1.325
r86 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.88
+ $Y=1.16 $X2=1.88 $Y2=1.16
r87 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.49
+ $Y=1.16 $X2=0.49 $Y2=1.16
r88 19 28 7.15912 $w=3.28e-07 $l=2.05e-07 $layer=LI1_cond $X=0.435 $Y=1.16
+ $X2=0.23 $Y2=1.16
r89 19 21 2.68691 $w=3.3e-07 $l=9e-08 $layer=LI1_cond $X=0.435 $Y=1.16 $X2=0.525
+ $Y2=1.16
r90 18 27 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=1.795 $Y=1.465
+ $X2=1.795 $Y2=1.325
r91 15 18 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.705 $Y=1.55
+ $X2=1.795 $Y2=1.465
r92 15 16 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.705 $Y=1.55
+ $X2=0.615 $Y2=1.55
r93 14 16 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=0.525 $Y=1.465
+ $X2=0.615 $Y2=1.55
r94 13 21 4.92601 $w=1.8e-07 $l=1.65e-07 $layer=LI1_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.16
r95 13 14 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=0.525 $Y=1.325
+ $X2=0.525 $Y2=1.465
r96 10 25 49.2447 $w=2.79e-07 $l=2.54951e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.895 $Y2=1.16
r97 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r98 7 25 38.7444 $w=2.79e-07 $l=1.98997e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.895 $Y2=1.16
r99 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.56
r100 4 22 38.5416 $w=3.03e-07 $l=2.05122e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.49 $Y2=1.16
r101 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.58 $Y=0.995
+ $X2=0.58 $Y2=0.56
r102 1 22 47.6478 $w=3.03e-07 $l=2.52488e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.49 $Y2=1.16
r103 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_8%A 1 3 4 6 7 9 10 12 13 19 20
r48 20 21 5.70789 $w=3.8e-07 $l=4.5e-08 $layer=POLY_cond $X=1.39 $Y=1.202
+ $X2=1.435 $Y2=1.202
r49 18 20 2.53684 $w=3.8e-07 $l=2e-08 $layer=POLY_cond $X=1.37 $Y=1.202 $X2=1.39
+ $Y2=1.202
r50 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.37
+ $Y=1.16 $X2=1.37 $Y2=1.16
r51 16 18 50.7368 $w=3.8e-07 $l=4e-07 $layer=POLY_cond $X=0.97 $Y=1.202 $X2=1.37
+ $Y2=1.202
r52 15 16 0.634211 $w=3.8e-07 $l=5e-09 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.97 $Y2=1.202
r53 13 19 8.45125 $w=2.98e-07 $l=2.2e-07 $layer=LI1_cond $X=1.15 $Y=1.145
+ $X2=1.37 $Y2=1.145
r54 10 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r55 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r56 7 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.39 $Y=0.995
+ $X2=1.39 $Y2=1.202
r57 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.39 $Y=0.995 $X2=1.39
+ $Y2=0.56
r58 4 16 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.97 $Y=0.995
+ $X2=0.97 $Y2=1.202
r59 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.97 $Y=0.995 $X2=0.97
+ $Y2=0.56
r60 1 15 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r61 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_8%A_117_297# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 36 37 39 40 42 43 45 46 48 49 51 52 54 55 57 60 64 66
+ 67 70 73 75 81 85 87 88 105
c196 105 0 7.45138e-20 $X=5.64 $Y=1.202
c197 87 0 1.60887e-19 $X=1.67 $Y=1.96
c198 10 0 1.96457e-19 $X=2.375 $Y=1.41
r199 105 106 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.202
+ $X2=5.665 $Y2=1.202
r200 104 105 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=5.22 $Y=1.202
+ $X2=5.64 $Y2=1.202
r201 103 104 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=5.195 $Y=1.202
+ $X2=5.22 $Y2=1.202
r202 100 101 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.202
+ $X2=4.725 $Y2=1.202
r203 99 100 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=4.28 $Y=1.202
+ $X2=4.7 $Y2=1.202
r204 98 99 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=4.255 $Y=1.202
+ $X2=4.28 $Y2=1.202
r205 97 98 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=3.785 $Y=1.202
+ $X2=4.255 $Y2=1.202
r206 96 97 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.202
+ $X2=3.785 $Y2=1.202
r207 95 96 55.0109 $w=3.68e-07 $l=4.2e-07 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.76 $Y2=1.202
r208 94 95 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=3.315 $Y=1.202
+ $X2=3.34 $Y2=1.202
r209 93 94 61.5598 $w=3.68e-07 $l=4.7e-07 $layer=POLY_cond $X=2.845 $Y=1.202
+ $X2=3.315 $Y2=1.202
r210 92 93 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.82 $Y=1.202
+ $X2=2.845 $Y2=1.202
r211 89 90 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.202
+ $X2=2.4 $Y2=1.202
r212 82 103 4.58424 $w=3.68e-07 $l=3.5e-08 $layer=POLY_cond $X=5.16 $Y=1.202
+ $X2=5.195 $Y2=1.202
r213 82 101 56.9755 $w=3.68e-07 $l=4.35e-07 $layer=POLY_cond $X=5.16 $Y=1.202
+ $X2=4.725 $Y2=1.202
r214 81 82 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=5.16
+ $Y=1.16 $X2=5.16 $Y2=1.16
r215 79 92 49.7717 $w=3.68e-07 $l=3.8e-07 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.82 $Y2=1.202
r216 79 90 5.23913 $w=3.68e-07 $l=4e-08 $layer=POLY_cond $X=2.44 $Y=1.202
+ $X2=2.4 $Y2=1.202
r217 78 81 143.654 $w=2.08e-07 $l=2.72e-06 $layer=LI1_cond $X=2.44 $Y=1.16
+ $X2=5.16 $Y2=1.16
r218 78 79 32.2844 $w=1.7e-07 $l=7.65e-07 $layer=licon1_POLY $count=4 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r219 76 88 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.305 $Y=1.16
+ $X2=2.22 $Y2=1.16
r220 76 78 7.12987 $w=2.08e-07 $l=1.35e-07 $layer=LI1_cond $X=2.305 $Y=1.16
+ $X2=2.44 $Y2=1.16
r221 74 88 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.22 $Y=1.265
+ $X2=2.22 $Y2=1.16
r222 74 75 35.2299 $w=1.68e-07 $l=5.4e-07 $layer=LI1_cond $X=2.22 $Y=1.265
+ $X2=2.22 $Y2=1.805
r223 73 88 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.22 $Y=1.055
+ $X2=2.22 $Y2=1.16
r224 72 73 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=2.22 $Y=0.825
+ $X2=2.22 $Y2=1.055
r225 71 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.805 $Y=1.89
+ $X2=1.67 $Y2=1.89
r226 70 75 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=2.22 $Y2=1.805
r227 70 71 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.135 $Y=1.89
+ $X2=1.805 $Y2=1.89
r228 66 72 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=2.22 $Y2=0.825
r229 66 67 51.5401 $w=1.68e-07 $l=7.9e-07 $layer=LI1_cond $X=2.135 $Y=0.74
+ $X2=1.345 $Y2=0.74
r230 62 67 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.345 $Y2=0.74
r231 62 64 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.18 $Y=0.655
+ $X2=1.18 $Y2=0.38
r232 61 85 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.865 $Y=1.89
+ $X2=0.715 $Y2=1.89
r233 60 87 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=1.535 $Y=1.89
+ $X2=1.67 $Y2=1.89
r234 60 61 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.535 $Y=1.89
+ $X2=0.865 $Y2=1.89
r235 55 106 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.202
r236 55 57 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r237 52 105 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.64 $Y=0.995
+ $X2=5.64 $Y2=1.202
r238 52 54 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.64 $Y=0.995
+ $X2=5.64 $Y2=0.56
r239 49 104 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=1.202
r240 49 51 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.22 $Y=0.995
+ $X2=5.22 $Y2=0.56
r241 46 103 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.202
r242 46 48 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r243 43 101 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.202
r244 43 45 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r245 40 100 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=1.202
r246 40 42 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.7 $Y=0.995
+ $X2=4.7 $Y2=0.56
r247 37 99 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=1.202
r248 37 39 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.28 $Y=0.995
+ $X2=4.28 $Y2=0.56
r249 34 98 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.202
r250 34 36 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r251 31 97 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.202
r252 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r253 28 96 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=1.202
r254 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.76 $Y=0.995
+ $X2=3.76 $Y2=0.56
r255 25 95 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=1.202
r256 25 27 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.34 $Y=0.995
+ $X2=3.34 $Y2=0.56
r257 22 94 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.202
r258 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r259 19 93 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.202
r260 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r261 16 92 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=1.202
r262 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.82 $Y=0.995
+ $X2=2.82 $Y2=0.56
r263 13 90 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=1.202
r264 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.4 $Y=0.995
+ $X2=2.4 $Y2=0.56
r265 10 89 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.202
r266 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r267 3 87 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r268 2 85 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.96
r269 1 64 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.045
+ $Y=0.235 $X2=1.18 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_8%VPWR 1 2 3 4 5 6 7 22 24 28 32 34 38 40 44
+ 46 50 52 56 58 60 65 72 73 79 82 85 88 91 94
r108 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r109 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r110 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r111 89 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r112 88 89 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 86 89 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r114 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r115 83 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r116 82 83 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r117 79 80 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 73 95 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r119 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r120 70 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=5.9 $Y2=2.72
r121 70 72 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.065 $Y=2.72
+ $X2=6.21 $Y2=2.72
r122 69 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r123 69 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r124 68 69 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r125 66 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.2 $Y2=2.72
r126 66 68 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=1.365 $Y=2.72
+ $X2=1.61 $Y2=2.72
r127 65 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=2.14 $Y2=2.72
r128 65 68 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.975 $Y=2.72
+ $X2=1.61 $Y2=2.72
r129 64 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r130 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r131 61 76 4.49698 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.197 $Y2=2.72
r132 61 63 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=2.72
+ $X2=0.69 $Y2=2.72
r133 60 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=1.2 $Y2=2.72
r134 60 63 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=1.035 $Y=2.72
+ $X2=0.69 $Y2=2.72
r135 58 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 58 76 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r137 54 94 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635 $X2=5.9
+ $Y2=2.72
r138 54 56 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=1.89
r139 53 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=2.72
+ $X2=4.96 $Y2=2.72
r140 52 94 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.9 $Y2=2.72
r141 52 53 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=2.72
+ $X2=5.125 $Y2=2.72
r142 48 91 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r143 48 50 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=1.89
r144 47 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=2.72
+ $X2=4.02 $Y2=2.72
r145 46 91 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.96 $Y2=2.72
r146 46 47 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=2.72
+ $X2=4.185 $Y2=2.72
r147 42 88 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r148 42 44 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=1.89
r149 41 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=2.72
+ $X2=3.08 $Y2=2.72
r150 40 88 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=4.02 $Y2=2.72
r151 40 41 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=2.72
+ $X2=3.245 $Y2=2.72
r152 36 85 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r153 36 38 26.0173 $w=3.28e-07 $l=7.45e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=1.89
r154 35 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.305 $Y=2.72
+ $X2=2.14 $Y2=2.72
r155 34 85 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.08 $Y2=2.72
r156 34 35 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.305 $Y2=2.72
r157 30 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r158 30 32 13.6198 $w=3.28e-07 $l=3.9e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.245
r159 26 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635 $X2=1.2
+ $Y2=2.72
r160 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.34
r161 22 76 3.0207 $w=3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.197 $Y2=2.72
r162 22 24 24.3934 $w=2.98e-07 $l=6.35e-07 $layer=LI1_cond $X=0.245 $Y=2.635
+ $X2=0.245 $Y2=2
r163 7 56 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=1.89
r164 6 50 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=1.89
r165 5 44 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=1.89
r166 4 38 300 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=1.89
r167 3 32 600 $w=1.7e-07 $l=8.29337e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.245
r168 2 28 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r169 1 24 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_8%X 1 2 3 4 5 6 7 8 27 31 35 36 37 38 41 45
+ 49 51 55 59 63 65 69 73 77 78 79 80 82 84 85
c114 36 0 7.31881e-20 $X=2.745 $Y=0.8
r115 83 85 6.99698 $w=4.18e-07 $l=2.55e-07 $layer=LI1_cond $X=5.705 $Y=1.445
+ $X2=5.705 $Y2=1.19
r116 83 84 2.7724 $w=3.45e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.705 $Y=1.445
+ $X2=5.605 $Y2=1.53
r117 81 85 8.36893 $w=4.18e-07 $l=3.05e-07 $layer=LI1_cond $X=5.705 $Y=0.885
+ $X2=5.705 $Y2=1.19
r118 81 82 2.7724 $w=3.45e-07 $l=1.36015e-07 $layer=LI1_cond $X=5.705 $Y=0.885
+ $X2=5.605 $Y2=0.8
r119 73 75 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=5.43 $Y=1.62
+ $X2=5.43 $Y2=2.3
r120 71 84 2.7724 $w=3.45e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.43 $Y=1.615
+ $X2=5.605 $Y2=1.53
r121 71 73 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=5.43 $Y=1.615
+ $X2=5.43 $Y2=1.62
r122 67 82 2.7724 $w=3.45e-07 $l=2.13307e-07 $layer=LI1_cond $X=5.43 $Y=0.715
+ $X2=5.605 $Y2=0.8
r123 67 69 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=5.43 $Y=0.715
+ $X2=5.43 $Y2=0.42
r124 66 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=1.53
+ $X2=4.49 $Y2=1.53
r125 65 84 3.97867 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=5.295 $Y=1.53
+ $X2=5.605 $Y2=1.53
r126 65 66 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=1.53
+ $X2=4.625 $Y2=1.53
r127 64 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.625 $Y=0.8
+ $X2=4.49 $Y2=0.8
r128 63 82 3.97867 $w=1.7e-07 $l=3.1e-07 $layer=LI1_cond $X=5.295 $Y=0.8
+ $X2=5.605 $Y2=0.8
r129 63 64 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=5.295 $Y=0.8
+ $X2=4.625 $Y2=0.8
r130 59 61 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=4.49 $Y=1.62
+ $X2=4.49 $Y2=2.3
r131 57 80 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.53
r132 57 59 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=4.49 $Y=1.615
+ $X2=4.49 $Y2=1.62
r133 53 79 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.49 $Y2=0.8
r134 53 55 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.49 $Y=0.715
+ $X2=4.49 $Y2=0.42
r135 52 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=1.53
+ $X2=3.55 $Y2=1.53
r136 51 80 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=1.53
+ $X2=4.49 $Y2=1.53
r137 51 52 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=1.53
+ $X2=3.685 $Y2=1.53
r138 50 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.685 $Y=0.8
+ $X2=3.55 $Y2=0.8
r139 49 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=4.355 $Y=0.8
+ $X2=4.49 $Y2=0.8
r140 49 50 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.355 $Y=0.8
+ $X2=3.685 $Y2=0.8
r141 45 47 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=3.55 $Y=1.62
+ $X2=3.55 $Y2=2.3
r142 43 78 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.53
r143 43 45 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=3.55 $Y=1.615
+ $X2=3.55 $Y2=1.62
r144 39 77 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.8
r145 39 41 12.5915 $w=2.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.55 $Y=0.715
+ $X2=3.55 $Y2=0.42
r146 37 78 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=3.55 $Y2=1.53
r147 37 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=1.53
+ $X2=2.745 $Y2=1.53
r148 35 77 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=3.415 $Y=0.8
+ $X2=3.55 $Y2=0.8
r149 35 36 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=3.415 $Y=0.8
+ $X2=2.745 $Y2=0.8
r150 31 33 29.0245 $w=2.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.61 $Y=1.62
+ $X2=2.61 $Y2=2.3
r151 29 38 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.745 $Y2=1.53
r152 29 31 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=2.61 $Y=1.615
+ $X2=2.61 $Y2=1.62
r153 25 36 7.28469 $w=1.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.745 $Y2=0.8
r154 25 27 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=2.61 $Y=0.715
+ $X2=2.61 $Y2=0.56
r155 8 75 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.3
r156 8 73 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.62
r157 7 61 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.3
r158 7 59 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.62
r159 6 47 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.3
r160 6 45 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.62
r161 5 33 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.3
r162 5 31 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.62
r163 4 69 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=5.295
+ $Y=0.235 $X2=5.43 $Y2=0.42
r164 3 55 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=4.355
+ $Y=0.235 $X2=4.49 $Y2=0.42
r165 2 41 91 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=2 $X=3.415
+ $Y=0.235 $X2=3.55 $Y2=0.42
r166 1 27 182 $w=1.7e-07 $l=3.86652e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2_8%VGND 1 2 3 4 5 6 19 21 25 27 31 33 37 39 43
+ 45 49 51 53 63 64 70 73 76 79 82
r98 82 83 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r99 80 83 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r100 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r101 77 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r102 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r103 74 77 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.91
+ $Y2=0
r104 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r105 71 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r106 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r107 64 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=5.75
+ $Y2=0
r108 63 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r109 61 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=6.065 $Y=0 $X2=5.9
+ $Y2=0
r110 61 63 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=6.065 $Y=0
+ $X2=6.21 $Y2=0
r111 60 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.07
+ $Y2=0
r112 59 60 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r113 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r114 56 59 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r115 56 57 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r116 54 67 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r117 54 56 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r118 53 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=2.105
+ $Y2=0
r119 53 59 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=1.94 $Y=0 $X2=1.61
+ $Y2=0
r120 51 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r121 51 67 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r122 47 82 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.085 $X2=5.9
+ $Y2=0
r123 47 49 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0.44
r124 46 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.125 $Y=0 $X2=4.96
+ $Y2=0
r125 45 82 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.735 $Y=0 $X2=5.9
+ $Y2=0
r126 45 46 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=5.735 $Y=0
+ $X2=5.125 $Y2=0
r127 41 79 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r128 41 43 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.44
r129 40 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.185 $Y=0 $X2=4.02
+ $Y2=0
r130 39 79 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.795 $Y=0 $X2=4.96
+ $Y2=0
r131 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=4.795 $Y=0
+ $X2=4.185 $Y2=0
r132 35 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r133 35 37 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.44
r134 34 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.245 $Y=0 $X2=3.08
+ $Y2=0
r135 33 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.855 $Y=0 $X2=4.02
+ $Y2=0
r136 33 34 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.855 $Y=0
+ $X2=3.245 $Y2=0
r137 29 73 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r138 29 31 12.3975 $w=3.28e-07 $l=3.55e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.44
r139 28 70 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.27 $Y=0 $X2=2.105
+ $Y2=0
r140 27 73 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.08
+ $Y2=0
r141 27 28 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=2.915 $Y=0
+ $X2=2.27 $Y2=0
r142 23 70 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0
r143 23 25 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.105 $Y=0.085
+ $X2=2.105 $Y2=0.36
r144 19 67 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r145 19 21 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r146 6 49 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.44
r147 5 43 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.44
r148 4 37 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.44
r149 3 31 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=2.895
+ $Y=0.235 $X2=3.08 $Y2=0.44
r150 2 25 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.105 $Y2=0.36
r151 1 21 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

