* File: sky130_fd_sc_hdll__clkbuf_16.pex.spice
* Created: Thu Aug 27 19:01:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_16%A 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 44
r64 43 44 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=1.94 $Y=1.155
+ $X2=1.965 $Y2=1.155
r65 42 43 47.733 $w=5.1e-07 $l=4.55e-07 $layer=POLY_cond $X=1.485 $Y=1.155
+ $X2=1.94 $Y2=1.155
r66 41 42 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=1.46 $Y=1.155
+ $X2=1.485 $Y2=1.155
r67 40 41 47.733 $w=5.1e-07 $l=4.55e-07 $layer=POLY_cond $X=1.005 $Y=1.155
+ $X2=1.46 $Y2=1.155
r68 39 40 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=0.98 $Y=1.155
+ $X2=1.005 $Y2=1.155
r69 38 39 47.733 $w=5.1e-07 $l=4.55e-07 $layer=POLY_cond $X=0.525 $Y=1.155
+ $X2=0.98 $Y2=1.155
r70 37 38 2.62269 $w=5.1e-07 $l=2.5e-08 $layer=POLY_cond $X=0.5 $Y=1.155
+ $X2=0.525 $Y2=1.155
r71 34 37 24.1288 $w=5.1e-07 $l=2.3e-07 $layer=POLY_cond $X=0.27 $Y=1.155
+ $X2=0.5 $Y2=1.155
r72 30 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.27
+ $Y=1.16 $X2=0.27 $Y2=1.16
r73 29 30 11.3415 $w=3.13e-07 $l=3.1e-07 $layer=LI1_cond $X=0.242 $Y=0.85
+ $X2=0.242 $Y2=1.16
r74 25 44 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.965 $Y=0.9
+ $X2=1.965 $Y2=1.155
r75 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.965 $Y=0.9
+ $X2=1.965 $Y2=0.445
r76 22 43 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.155
r77 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.94 $Y=1.41
+ $X2=1.94 $Y2=1.985
r78 18 42 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.485 $Y=0.9
+ $X2=1.485 $Y2=1.155
r79 18 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.485 $Y=0.9
+ $X2=1.485 $Y2=0.445
r80 15 41 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.155
r81 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.46 $Y=1.41
+ $X2=1.46 $Y2=1.985
r82 11 40 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=1.005 $Y=0.9
+ $X2=1.005 $Y2=1.155
r83 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.005 $Y=0.9
+ $X2=1.005 $Y2=0.445
r84 8 39 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.155
r85 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.98 $Y=1.41
+ $X2=0.98 $Y2=1.985
r86 4 38 31.9091 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=0.525 $Y=0.9
+ $X2=0.525 $Y2=1.155
r87 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.525 $Y=0.9
+ $X2=0.525 $Y2=0.445
r88 1 37 27.3507 $w=1.8e-07 $l=2.55e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.155
r89 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41 $X2=0.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_16%A_118_297# 1 2 3 4 15 17 19 22 24 26 29
+ 31 33 36 38 40 43 45 47 50 52 54 57 59 61 64 66 68 71 73 75 78 80 82 85 87 89
+ 92 94 96 99 101 103 106 108 110 113 115 117 118 120 123 127 131 133 137 141
+ 148 151 152 185
r277 185 186 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=9.615 $Y=1.18
+ $X2=9.64 $Y2=1.18
r278 184 185 56.292 $w=4.11e-07 $l=4.8e-07 $layer=POLY_cond $X=9.135 $Y=1.18
+ $X2=9.615 $Y2=1.18
r279 183 184 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=9.11 $Y=1.18
+ $X2=9.135 $Y2=1.18
r280 182 183 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=8.655 $Y=1.18
+ $X2=9.11 $Y2=1.18
r281 181 182 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=8.63 $Y=1.18
+ $X2=8.655 $Y2=1.18
r282 178 179 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=8.15 $Y=1.18
+ $X2=8.175 $Y2=1.18
r283 177 178 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=7.695 $Y=1.18
+ $X2=8.15 $Y2=1.18
r284 176 177 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=7.67 $Y=1.18
+ $X2=7.695 $Y2=1.18
r285 175 176 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=7.215 $Y=1.18
+ $X2=7.67 $Y2=1.18
r286 174 175 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=7.19 $Y=1.18
+ $X2=7.215 $Y2=1.18
r287 173 174 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=6.735 $Y=1.18
+ $X2=7.19 $Y2=1.18
r288 172 173 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=6.71 $Y=1.18
+ $X2=6.735 $Y2=1.18
r289 171 172 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=6.255 $Y=1.18
+ $X2=6.71 $Y2=1.18
r290 170 171 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=6.23 $Y=1.18
+ $X2=6.255 $Y2=1.18
r291 169 170 52.7737 $w=4.11e-07 $l=4.5e-07 $layer=POLY_cond $X=5.78 $Y=1.18
+ $X2=6.23 $Y2=1.18
r292 168 169 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=5.755 $Y=1.18
+ $X2=5.78 $Y2=1.18
r293 167 168 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=5.3 $Y=1.18
+ $X2=5.755 $Y2=1.18
r294 166 167 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=5.275 $Y=1.18
+ $X2=5.3 $Y2=1.18
r295 165 166 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=4.82 $Y=1.18
+ $X2=5.275 $Y2=1.18
r296 164 165 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=4.795 $Y=1.18
+ $X2=4.82 $Y2=1.18
r297 163 164 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=4.34 $Y=1.18
+ $X2=4.795 $Y2=1.18
r298 162 163 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=4.315 $Y=1.18
+ $X2=4.34 $Y2=1.18
r299 161 162 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=3.86 $Y=1.18
+ $X2=4.315 $Y2=1.18
r300 160 161 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.18
+ $X2=3.86 $Y2=1.18
r301 159 160 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=3.38 $Y=1.18
+ $X2=3.835 $Y2=1.18
r302 158 159 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=3.355 $Y=1.18
+ $X2=3.38 $Y2=1.18
r303 157 158 53.3601 $w=4.11e-07 $l=4.55e-07 $layer=POLY_cond $X=2.9 $Y=1.18
+ $X2=3.355 $Y2=1.18
r304 156 157 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=2.875 $Y=1.18
+ $X2=2.9 $Y2=1.18
r305 153 154 2.93187 $w=4.11e-07 $l=2.5e-08 $layer=POLY_cond $X=2.395 $Y=1.18
+ $X2=2.42 $Y2=1.18
r306 149 181 38.1144 $w=4.11e-07 $l=3.25e-07 $layer=POLY_cond $X=8.305 $Y=1.18
+ $X2=8.63 $Y2=1.18
r307 149 179 15.2457 $w=4.11e-07 $l=1.3e-07 $layer=POLY_cond $X=8.305 $Y=1.18
+ $X2=8.175 $Y2=1.18
r308 148 149 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=8.305
+ $Y=1.16 $X2=8.305 $Y2=1.16
r309 146 156 25.8005 $w=4.11e-07 $l=2.2e-07 $layer=POLY_cond $X=2.655 $Y=1.18
+ $X2=2.875 $Y2=1.18
r310 146 154 27.5596 $w=4.11e-07 $l=2.35e-07 $layer=POLY_cond $X=2.655 $Y=1.18
+ $X2=2.42 $Y2=1.18
r311 145 148 260.452 $w=2.48e-07 $l=5.65e-06 $layer=LI1_cond $X=2.655 $Y=1.2
+ $X2=8.305 $Y2=1.2
r312 145 146 18.16 $w=1.7e-07 $l=1.36e-06 $layer=licon1_POLY $count=8 $X=2.655
+ $Y=1.16 $X2=2.655 $Y2=1.16
r313 143 152 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.83 $Y=1.2 $X2=1.705
+ $Y2=1.2
r314 143 145 38.0306 $w=2.48e-07 $l=8.25e-07 $layer=LI1_cond $X=1.83 $Y=1.2
+ $X2=2.655 $Y2=1.2
r315 139 152 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=1.325
+ $X2=1.705 $Y2=1.2
r316 139 141 27.4281 $w=2.48e-07 $l=5.95e-07 $layer=LI1_cond $X=1.705 $Y=1.325
+ $X2=1.705 $Y2=1.92
r317 135 152 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.705 $Y=1.075
+ $X2=1.705 $Y2=1.2
r318 135 137 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=1.705 $Y=1.075
+ $X2=1.705 $Y2=0.445
r319 134 151 1.3064 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=0.87 $Y=1.2
+ $X2=0.745 $Y2=1.2
r320 133 152 6.1 $w=2.5e-07 $l=1.25e-07 $layer=LI1_cond $X=1.58 $Y=1.2 $X2=1.705
+ $Y2=1.2
r321 133 134 32.7294 $w=2.48e-07 $l=7.1e-07 $layer=LI1_cond $X=1.58 $Y=1.2
+ $X2=0.87 $Y2=1.2
r322 129 151 5.20938 $w=2.47e-07 $l=1.26491e-07 $layer=LI1_cond $X=0.742
+ $Y=1.325 $X2=0.745 $Y2=1.2
r323 129 131 29.8694 $w=2.43e-07 $l=6.35e-07 $layer=LI1_cond $X=0.742 $Y=1.325
+ $X2=0.742 $Y2=1.96
r324 125 151 5.20938 $w=2.47e-07 $l=1.25e-07 $layer=LI1_cond $X=0.745 $Y=1.075
+ $X2=0.745 $Y2=1.2
r325 125 127 29.0416 $w=2.48e-07 $l=6.3e-07 $layer=LI1_cond $X=0.745 $Y=1.075
+ $X2=0.745 $Y2=0.445
r326 121 186 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=9.64 $Y=0.95
+ $X2=9.64 $Y2=1.18
r327 121 123 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.64 $Y=0.95
+ $X2=9.64 $Y2=0.445
r328 118 185 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=9.615 $Y=1.41
+ $X2=9.615 $Y2=1.18
r329 118 120 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.615 $Y=1.41
+ $X2=9.615 $Y2=1.985
r330 115 184 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=9.135 $Y=1.41
+ $X2=9.135 $Y2=1.18
r331 115 117 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.135 $Y=1.41
+ $X2=9.135 $Y2=1.985
r332 111 183 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=9.11 $Y=0.95
+ $X2=9.11 $Y2=1.18
r333 111 113 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=9.11 $Y=0.95
+ $X2=9.11 $Y2=0.445
r334 108 182 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=8.655 $Y=1.41
+ $X2=8.655 $Y2=1.18
r335 108 110 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.655 $Y=1.41
+ $X2=8.655 $Y2=1.985
r336 104 181 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=8.63 $Y=0.95
+ $X2=8.63 $Y2=1.18
r337 104 106 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.63 $Y=0.95
+ $X2=8.63 $Y2=0.445
r338 101 179 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=8.175 $Y=1.41
+ $X2=8.175 $Y2=1.18
r339 101 103 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.175 $Y=1.41
+ $X2=8.175 $Y2=1.985
r340 97 178 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=8.15 $Y=0.95
+ $X2=8.15 $Y2=1.18
r341 97 99 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=8.15 $Y=0.95
+ $X2=8.15 $Y2=0.445
r342 94 177 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=7.695 $Y=1.41
+ $X2=7.695 $Y2=1.18
r343 94 96 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.695 $Y=1.41
+ $X2=7.695 $Y2=1.985
r344 90 176 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.67 $Y=0.95
+ $X2=7.67 $Y2=1.18
r345 90 92 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.67 $Y=0.95
+ $X2=7.67 $Y2=0.445
r346 87 175 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=7.215 $Y=1.41
+ $X2=7.215 $Y2=1.18
r347 87 89 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.215 $Y=1.41
+ $X2=7.215 $Y2=1.985
r348 83 174 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=7.19 $Y=0.95
+ $X2=7.19 $Y2=1.18
r349 83 85 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=7.19 $Y=0.95
+ $X2=7.19 $Y2=0.445
r350 80 173 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=6.735 $Y=1.41
+ $X2=6.735 $Y2=1.18
r351 80 82 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.735 $Y=1.41
+ $X2=6.735 $Y2=1.985
r352 76 172 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.71 $Y=0.95
+ $X2=6.71 $Y2=1.18
r353 76 78 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.71 $Y=0.95
+ $X2=6.71 $Y2=0.445
r354 73 171 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=6.255 $Y=1.41
+ $X2=6.255 $Y2=1.18
r355 73 75 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.255 $Y=1.41
+ $X2=6.255 $Y2=1.985
r356 69 170 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=6.23 $Y=0.95
+ $X2=6.23 $Y2=1.18
r357 69 71 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=6.23 $Y=0.95
+ $X2=6.23 $Y2=0.445
r358 66 169 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.78 $Y=1.41
+ $X2=5.78 $Y2=1.18
r359 66 68 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.78 $Y=1.41
+ $X2=5.78 $Y2=1.985
r360 62 168 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.755 $Y=0.95
+ $X2=5.755 $Y2=1.18
r361 62 64 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.755 $Y=0.95
+ $X2=5.755 $Y2=0.445
r362 59 167 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=5.3 $Y=1.41
+ $X2=5.3 $Y2=1.18
r363 59 61 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.3 $Y=1.41
+ $X2=5.3 $Y2=1.985
r364 55 166 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=5.275 $Y=0.95
+ $X2=5.275 $Y2=1.18
r365 55 57 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=5.275 $Y=0.95
+ $X2=5.275 $Y2=0.445
r366 52 165 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.18
r367 52 54 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.985
r368 48 164 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.795 $Y=0.95
+ $X2=4.795 $Y2=1.18
r369 48 50 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.795 $Y=0.95
+ $X2=4.795 $Y2=0.445
r370 45 163 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.18
r371 45 47 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.34 $Y=1.41
+ $X2=4.34 $Y2=1.985
r372 41 162 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=4.315 $Y=0.95
+ $X2=4.315 $Y2=1.18
r373 41 43 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=4.315 $Y=0.95
+ $X2=4.315 $Y2=0.445
r374 38 161 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.18
r375 38 40 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.86 $Y=1.41
+ $X2=3.86 $Y2=1.985
r376 34 160 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.835 $Y=0.95
+ $X2=3.835 $Y2=1.18
r377 34 36 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.835 $Y=0.95
+ $X2=3.835 $Y2=0.445
r378 31 159 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.18
r379 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.38 $Y=1.41
+ $X2=3.38 $Y2=1.985
r380 27 158 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=3.355 $Y=0.95
+ $X2=3.355 $Y2=1.18
r381 27 29 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=3.355 $Y=0.95
+ $X2=3.355 $Y2=0.445
r382 24 157 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.9 $Y=1.41
+ $X2=2.9 $Y2=1.18
r383 24 26 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.9 $Y=1.41
+ $X2=2.9 $Y2=1.985
r384 20 156 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.875 $Y=0.95
+ $X2=2.875 $Y2=1.18
r385 20 22 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.875 $Y=0.95
+ $X2=2.875 $Y2=0.445
r386 17 154 22.1098 $w=1.8e-07 $l=2.3e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.18
r387 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.42 $Y2=1.985
r388 13 153 26.5265 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=2.395 $Y=0.95
+ $X2=2.395 $Y2=1.18
r389 13 15 258.947 $w=1.5e-07 $l=5.05e-07 $layer=POLY_cond $X=2.395 $Y=0.95
+ $X2=2.395 $Y2=0.445
r390 4 141 300 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=2 $X=1.55
+ $Y=1.485 $X2=1.7 $Y2=1.92
r391 3 131 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=1.96
r392 2 137 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.7 $Y2=0.445
r393 1 127 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=0.6
+ $Y=0.235 $X2=0.74 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 34 36 38 42
+ 44 48 52 56 60 64 68 72 76 78 80 83 84 86 87 89 90 92 93 95 96 98 99 101 102
+ 103 127 135 138 142
r146 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r147 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r148 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r149 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r150 130 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=9.89 $Y2=2.72
r151 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r152 127 141 4.22234 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=9.755 $Y=2.72
+ $X2=9.937 $Y2=2.72
r153 127 129 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=9.755 $Y=2.72
+ $X2=9.43 $Y2=2.72
r154 126 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r155 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r156 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r157 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r158 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r159 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r160 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r161 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r162 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r163 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r164 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r165 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r166 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r167 108 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r168 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r169 105 138 7.16073 $w=1.72e-07 $l=1.3e-07 $layer=LI1_cond $X=2.31 $Y=2.717
+ $X2=2.18 $Y2=2.717
r170 105 107 43.0961 $w=1.73e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=2.717
+ $X2=2.99 $Y2=2.717
r171 103 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r172 103 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r173 101 125 16.4779 $w=1.73e-07 $l=2.6e-07 $layer=LI1_cond $X=8.77 $Y=2.717
+ $X2=8.51 $Y2=2.717
r174 101 102 7.05609 $w=1.72e-07 $l=1.27e-07 $layer=LI1_cond $X=8.77 $Y=2.717
+ $X2=8.897 $Y2=2.717
r175 100 129 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.025 $Y=2.72
+ $X2=9.43 $Y2=2.72
r176 100 102 7.05609 $w=1.72e-07 $l=1.29491e-07 $layer=LI1_cond $X=9.025 $Y=2.72
+ $X2=8.897 $Y2=2.717
r177 98 122 13.9429 $w=1.73e-07 $l=2.2e-07 $layer=LI1_cond $X=7.81 $Y=2.717
+ $X2=7.59 $Y2=2.717
r178 98 99 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=7.81 $Y=2.717
+ $X2=7.932 $Y2=2.717
r179 97 125 28.8364 $w=1.73e-07 $l=4.55e-07 $layer=LI1_cond $X=8.055 $Y=2.717
+ $X2=8.51 $Y2=2.717
r180 97 99 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=8.055 $Y=2.717
+ $X2=7.932 $Y2=2.717
r181 95 119 11.4078 $w=1.73e-07 $l=1.8e-07 $layer=LI1_cond $X=6.85 $Y=2.717
+ $X2=6.67 $Y2=2.717
r182 95 96 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=6.85 $Y=2.717
+ $X2=6.972 $Y2=2.717
r183 94 122 31.3714 $w=1.73e-07 $l=4.95e-07 $layer=LI1_cond $X=7.095 $Y=2.717
+ $X2=7.59 $Y2=2.717
r184 94 96 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=7.095 $Y=2.717
+ $X2=6.972 $Y2=2.717
r185 92 116 8.87273 $w=1.73e-07 $l=1.4e-07 $layer=LI1_cond $X=5.89 $Y=2.717
+ $X2=5.75 $Y2=2.717
r186 92 93 6.76825 $w=1.75e-07 $l=1.22e-07 $layer=LI1_cond $X=5.89 $Y=2.717
+ $X2=6.012 $Y2=2.717
r187 91 119 33.9065 $w=1.73e-07 $l=5.35e-07 $layer=LI1_cond $X=6.135 $Y=2.717
+ $X2=6.67 $Y2=2.717
r188 91 93 6.76825 $w=1.75e-07 $l=1.23e-07 $layer=LI1_cond $X=6.135 $Y=2.717
+ $X2=6.012 $Y2=2.717
r189 89 113 6.33766 $w=1.73e-07 $l=1e-07 $layer=LI1_cond $X=4.93 $Y=2.717
+ $X2=4.83 $Y2=2.717
r190 89 90 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.93 $Y=2.717
+ $X2=5.06 $Y2=2.717
r191 88 116 35.4909 $w=1.73e-07 $l=5.6e-07 $layer=LI1_cond $X=5.19 $Y=2.717
+ $X2=5.75 $Y2=2.717
r192 88 90 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=5.19 $Y=2.717
+ $X2=5.06 $Y2=2.717
r193 86 110 3.8026 $w=1.73e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=2.717
+ $X2=3.91 $Y2=2.717
r194 86 87 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=3.97 $Y=2.717
+ $X2=4.1 $Y2=2.717
r195 85 113 38.026 $w=1.73e-07 $l=6e-07 $layer=LI1_cond $X=4.23 $Y=2.717
+ $X2=4.83 $Y2=2.717
r196 85 87 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=4.23 $Y=2.717
+ $X2=4.1 $Y2=2.717
r197 83 107 1.26753 $w=1.73e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=2.717
+ $X2=2.99 $Y2=2.717
r198 83 84 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=3.01 $Y=2.717
+ $X2=3.14 $Y2=2.717
r199 82 110 40.561 $w=1.73e-07 $l=6.4e-07 $layer=LI1_cond $X=3.27 $Y=2.717
+ $X2=3.91 $Y2=2.717
r200 82 84 7.08309 $w=1.75e-07 $l=1.3e-07 $layer=LI1_cond $X=3.27 $Y=2.717
+ $X2=3.14 $Y2=2.717
r201 78 141 3.06235 $w=2.7e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.89 $Y=2.635
+ $X2=9.937 $Y2=2.72
r202 78 80 17.7135 $w=2.68e-07 $l=4.15e-07 $layer=LI1_cond $X=9.89 $Y=2.635
+ $X2=9.89 $Y2=2.22
r203 74 102 0.0190999 $w=2.55e-07 $l=8.7e-08 $layer=LI1_cond $X=8.897 $Y=2.63
+ $X2=8.897 $Y2=2.717
r204 74 76 18.5295 $w=2.53e-07 $l=4.1e-07 $layer=LI1_cond $X=8.897 $Y=2.63
+ $X2=8.897 $Y2=2.22
r205 70 99 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=7.932 $Y=2.63
+ $X2=7.932 $Y2=2.717
r206 70 72 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=7.932 $Y=2.63
+ $X2=7.932 $Y2=2.22
r207 66 96 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=6.972 $Y=2.63
+ $X2=6.972 $Y2=2.717
r208 66 68 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=6.972 $Y=2.63
+ $X2=6.972 $Y2=2.22
r209 62 93 0.164012 $w=2.45e-07 $l=8.7e-08 $layer=LI1_cond $X=6.012 $Y=2.63
+ $X2=6.012 $Y2=2.717
r210 62 64 19.2858 $w=2.43e-07 $l=4.1e-07 $layer=LI1_cond $X=6.012 $Y=2.63
+ $X2=6.012 $Y2=2.22
r211 58 90 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=5.06 $Y=2.63
+ $X2=5.06 $Y2=2.717
r212 58 60 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=5.06 $Y=2.63
+ $X2=5.06 $Y2=2.22
r213 54 87 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=4.1 $Y=2.63
+ $X2=4.1 $Y2=2.717
r214 54 56 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=4.1 $Y=2.63 $X2=4.1
+ $Y2=2.22
r215 50 84 0.0359085 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=3.14 $Y=2.63
+ $X2=3.14 $Y2=2.717
r216 50 52 18.1731 $w=2.58e-07 $l=4.1e-07 $layer=LI1_cond $X=3.14 $Y=2.63
+ $X2=3.14 $Y2=2.22
r217 46 138 0.0838798 $w=2.6e-07 $l=8.7e-08 $layer=LI1_cond $X=2.18 $Y=2.63
+ $X2=2.18 $Y2=2.717
r218 46 48 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=2.18 $Y=2.63
+ $X2=2.18 $Y2=2
r219 45 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=2.72
+ $X2=1.22 $Y2=2.72
r220 44 138 7.16073 $w=1.72e-07 $l=1.31491e-07 $layer=LI1_cond $X=2.05 $Y=2.72
+ $X2=2.18 $Y2=2.717
r221 44 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.05 $Y=2.72 $X2=1.35
+ $Y2=2.72
r222 40 135 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r223 40 42 28.1462 $w=2.58e-07 $l=6.35e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2
r224 39 132 4.45907 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=2.72
+ $X2=0.195 $Y2=2.72
r225 38 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=2.72
+ $X2=1.22 $Y2=2.72
r226 38 39 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=2.72 $X2=0.39
+ $Y2=2.72
r227 34 132 3.01845 $w=2.95e-07 $l=1.05924e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.195 $Y2=2.72
r228 34 36 24.8068 $w=2.93e-07 $l=6.35e-07 $layer=LI1_cond $X=0.242 $Y=2.635
+ $X2=0.242 $Y2=2
r229 11 80 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=9.705
+ $Y=1.485 $X2=9.855 $Y2=2.22
r230 10 76 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=8.745
+ $Y=1.485 $X2=8.895 $Y2=2.22
r231 9 72 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=7.785
+ $Y=1.485 $X2=7.935 $Y2=2.22
r232 8 68 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=6.825
+ $Y=1.485 $X2=6.975 $Y2=2.22
r233 7 64 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=5.87
+ $Y=1.485 $X2=6.02 $Y2=2.22
r234 6 60 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.485 $X2=5.06 $Y2=2.22
r235 5 56 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=3.95
+ $Y=1.485 $X2=4.1 $Y2=2.22
r236 4 52 600 $w=1.7e-07 $l=8.0652e-07 $layer=licon1_PDIFF $count=1 $X=2.99
+ $Y=1.485 $X2=3.14 $Y2=2.22
r237 3 48 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=2.03
+ $Y=1.485 $X2=2.18 $Y2=2
r238 2 42 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=1.07
+ $Y=1.485 $X2=1.22 $Y2=2
r239 1 36 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16
+ 51 55 56 57 61 65 67 71 75 77 81 85 87 91 95 97 101 105 107 111 113 119 124
+ 125 127 128 130 131 133 134 136 137 139 140 141 144 157 161 163
c220 144 0 7.59816e-20 $X=9.375 $Y=1.445
r221 161 163 1.02191 $w=7.76e-07 $l=6.5e-08 $layer=LI1_cond $X=9.375 $Y=1.235
+ $X2=9.44 $Y2=1.235
r222 157 161 6.21005 $w=7.76e-07 $l=3.95e-07 $layer=LI1_cond $X=8.98 $Y=1.235
+ $X2=9.375 $Y2=1.235
r223 144 163 0.314433 $w=7.76e-07 $l=2e-08 $layer=LI1_cond $X=9.46 $Y=1.235
+ $X2=9.44 $Y2=1.235
r224 141 157 0.471649 $w=7.76e-07 $l=3e-08 $layer=LI1_cond $X=8.95 $Y=1.235
+ $X2=8.98 $Y2=1.235
r225 117 161 7.24882 $w=2.6e-07 $l=5e-07 $layer=LI1_cond $X=9.375 $Y=0.735
+ $X2=9.375 $Y2=1.235
r226 117 119 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=9.375 $Y=0.735
+ $X2=9.375 $Y2=0.445
r227 116 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.535 $Y=0.82
+ $X2=8.405 $Y2=0.82
r228 113 141 8.5683 $w=7.76e-07 $l=7.54669e-07 $layer=LI1_cond $X=8.405 $Y=1.735
+ $X2=8.95 $Y2=1.235
r229 109 140 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.405 $Y=0.735
+ $X2=8.405 $Y2=0.82
r230 109 111 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=8.405 $Y=0.735
+ $X2=8.405 $Y2=0.445
r231 108 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=7.575 $Y=1.615
+ $X2=7.445 $Y2=1.615
r232 107 113 14.4985 $w=7.76e-07 $l=1.07798e-06 $layer=LI1_cond $X=8.76 $Y=0.82
+ $X2=8.405 $Y2=1.735
r233 107 116 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=8.76 $Y=0.82
+ $X2=8.535 $Y2=0.82
r234 107 108 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=8.275 $Y=1.615
+ $X2=7.575 $Y2=1.615
r235 106 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.575 $Y=0.82
+ $X2=7.445 $Y2=0.82
r236 105 140 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=8.405 $Y2=0.82
r237 105 106 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=8.275 $Y=0.82
+ $X2=7.575 $Y2=0.82
r238 99 137 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=7.445 $Y=0.735
+ $X2=7.445 $Y2=0.82
r239 99 101 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=7.445 $Y=0.735
+ $X2=7.445 $Y2=0.445
r240 98 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.615 $Y=1.615
+ $X2=6.485 $Y2=1.615
r241 97 139 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=7.315 $Y=1.615
+ $X2=7.445 $Y2=1.615
r242 97 98 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=7.315 $Y=1.615
+ $X2=6.615 $Y2=1.615
r243 96 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.615 $Y=0.82
+ $X2=6.485 $Y2=0.82
r244 95 137 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=7.315 $Y=0.82
+ $X2=7.445 $Y2=0.82
r245 95 96 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=7.315 $Y=0.82
+ $X2=6.615 $Y2=0.82
r246 89 134 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=6.485 $Y=0.735
+ $X2=6.485 $Y2=0.82
r247 89 91 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=6.485 $Y=0.735
+ $X2=6.485 $Y2=0.445
r248 88 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.67 $Y=1.615
+ $X2=5.54 $Y2=1.615
r249 87 136 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=6.355 $Y=1.615
+ $X2=6.485 $Y2=1.615
r250 87 88 32.8926 $w=2.38e-07 $l=6.85e-07 $layer=LI1_cond $X=6.355 $Y=1.615
+ $X2=5.67 $Y2=1.615
r251 86 131 8.5188 $w=1.7e-07 $l=1.63e-07 $layer=LI1_cond $X=5.67 $Y=0.82
+ $X2=5.507 $Y2=0.82
r252 85 134 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=6.355 $Y=0.82
+ $X2=6.485 $Y2=0.82
r253 85 86 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=6.355 $Y=0.82
+ $X2=5.67 $Y2=0.82
r254 79 131 0.848899 $w=3.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.507 $Y=0.735
+ $X2=5.507 $Y2=0.82
r255 79 81 10.2833 $w=3.23e-07 $l=2.9e-07 $layer=LI1_cond $X=5.507 $Y=0.735
+ $X2=5.507 $Y2=0.445
r256 78 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.71 $Y=1.615
+ $X2=4.58 $Y2=1.615
r257 77 133 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=5.41 $Y=1.615
+ $X2=5.54 $Y2=1.615
r258 77 78 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=5.41 $Y=1.615
+ $X2=4.71 $Y2=1.615
r259 76 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.71 $Y=0.82
+ $X2=4.58 $Y2=0.82
r260 75 131 8.5188 $w=1.7e-07 $l=1.62e-07 $layer=LI1_cond $X=5.345 $Y=0.82
+ $X2=5.507 $Y2=0.82
r261 75 76 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.345 $Y=0.82
+ $X2=4.71 $Y2=0.82
r262 69 128 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.58 $Y=0.735
+ $X2=4.58 $Y2=0.82
r263 69 71 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=4.58 $Y=0.735
+ $X2=4.58 $Y2=0.445
r264 68 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.75 $Y=1.615
+ $X2=3.62 $Y2=1.615
r265 67 130 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=4.45 $Y=1.615
+ $X2=4.58 $Y2=1.615
r266 67 68 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=4.45 $Y=1.615
+ $X2=3.75 $Y2=1.615
r267 66 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.75 $Y=0.82
+ $X2=3.62 $Y2=0.82
r268 65 128 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.45 $Y=0.82
+ $X2=4.58 $Y2=0.82
r269 65 66 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.45 $Y=0.82 $X2=3.75
+ $Y2=0.82
r270 59 125 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.82
r271 59 61 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=3.62 $Y=0.735
+ $X2=3.62 $Y2=0.445
r272 58 124 3.55196 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=2.79 $Y=1.615
+ $X2=2.66 $Y2=1.615
r273 57 127 5.51899 $w=2.4e-07 $l=1.3e-07 $layer=LI1_cond $X=3.49 $Y=1.615
+ $X2=3.62 $Y2=1.615
r274 57 58 33.6129 $w=2.38e-07 $l=7e-07 $layer=LI1_cond $X=3.49 $Y=1.615
+ $X2=2.79 $Y2=1.615
r275 55 125 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.49 $Y=0.82
+ $X2=3.62 $Y2=0.82
r276 55 56 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=3.49 $Y=0.82 $X2=2.79
+ $Y2=0.82
r277 49 56 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=2.66 $Y=0.735
+ $X2=2.79 $Y2=0.82
r278 49 51 12.8542 $w=2.58e-07 $l=2.9e-07 $layer=LI1_cond $X=2.66 $Y=0.735
+ $X2=2.66 $Y2=0.445
r279 16 161 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=9.225
+ $Y=1.485 $X2=9.375 $Y2=1.69
r280 15 113 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=8.265
+ $Y=1.485 $X2=8.415 $Y2=1.69
r281 14 139 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=7.305
+ $Y=1.485 $X2=7.455 $Y2=1.69
r282 13 136 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=6.345
+ $Y=1.485 $X2=6.495 $Y2=1.69
r283 12 133 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=5.39
+ $Y=1.485 $X2=5.54 $Y2=1.69
r284 11 130 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=4.43
+ $Y=1.485 $X2=4.58 $Y2=1.69
r285 10 127 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=3.47
+ $Y=1.485 $X2=3.62 $Y2=1.69
r286 9 124 300 $w=1.7e-07 $l=2.69768e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=1.485 $X2=2.66 $Y2=1.69
r287 8 119 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=9.185
+ $Y=0.235 $X2=9.375 $Y2=0.445
r288 7 111 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=8.225
+ $Y=0.235 $X2=8.415 $Y2=0.445
r289 6 101 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=7.265
+ $Y=0.235 $X2=7.455 $Y2=0.445
r290 5 91 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=6.305
+ $Y=0.235 $X2=6.495 $Y2=0.445
r291 4 81 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=5.35
+ $Y=0.235 $X2=5.54 $Y2=0.445
r292 3 71 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=4.39
+ $Y=0.235 $X2=4.58 $Y2=0.445
r293 2 61 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=3.43
+ $Y=0.235 $X2=3.62 $Y2=0.445
r294 1 51 182 $w=1.7e-07 $l=2.89828e-07 $layer=licon1_NDIFF $count=1 $X=2.47
+ $Y=0.235 $X2=2.66 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__CLKBUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 34 36 38 42
+ 44 48 52 56 60 64 68 72 76 78 80 83 84 86 87 89 90 92 93 95 96 98 99 101 102
+ 103 127 135 138 142
c160 101 0 7.59816e-20 $X=8.765 $Y=0
r161 141 142 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.89 $Y=0
+ $X2=9.89 $Y2=0
r162 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r163 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r164 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r165 130 142 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=9.89 $Y2=0
r166 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r167 127 141 4.50146 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=9.725 $Y=0
+ $X2=9.922 $Y2=0
r168 127 129 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.725 $Y=0
+ $X2=9.43 $Y2=0
r169 126 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r170 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r171 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r172 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r173 120 123 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r174 119 120 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r175 117 120 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r176 116 117 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r177 114 117 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r178 113 114 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r179 111 114 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r180 110 111 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r181 108 111 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r182 108 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r183 107 108 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r184 105 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.31 $Y=0 $X2=2.18
+ $Y2=0
r185 105 107 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=2.31 $Y=0
+ $X2=2.99 $Y2=0
r186 103 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r187 103 132 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r188 101 125 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.51 $Y2=0
r189 101 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=8.765 $Y=0
+ $X2=8.895 $Y2=0
r190 100 129 26.4225 $w=1.68e-07 $l=4.05e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=9.43 $Y2=0
r191 100 102 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=9.025 $Y=0
+ $X2=8.895 $Y2=0
r192 98 122 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=7.805 $Y=0
+ $X2=7.59 $Y2=0
r193 98 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.805 $Y=0 $X2=7.93
+ $Y2=0
r194 97 125 29.6845 $w=1.68e-07 $l=4.55e-07 $layer=LI1_cond $X=8.055 $Y=0
+ $X2=8.51 $Y2=0
r195 97 99 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.055 $Y=0 $X2=7.93
+ $Y2=0
r196 95 119 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.845 $Y=0
+ $X2=6.67 $Y2=0
r197 95 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=6.845 $Y=0 $X2=6.97
+ $Y2=0
r198 94 122 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=7.095 $Y=0
+ $X2=7.59 $Y2=0
r199 94 96 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=7.095 $Y=0 $X2=6.97
+ $Y2=0
r200 92 116 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=5.75
+ $Y2=0
r201 92 93 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=5.89 $Y=0 $X2=6.012
+ $Y2=0
r202 91 119 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.135 $Y=0
+ $X2=6.67 $Y2=0
r203 91 93 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=6.135 $Y=0
+ $X2=6.012 $Y2=0
r204 89 113 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=4.83
+ $Y2=0
r205 89 90 6.92067 $w=1.7e-07 $l=1.22e-07 $layer=LI1_cond $X=4.93 $Y=0 $X2=5.052
+ $Y2=0
r206 88 116 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.75 $Y2=0
r207 88 90 6.92067 $w=1.7e-07 $l=1.23e-07 $layer=LI1_cond $X=5.175 $Y=0
+ $X2=5.052 $Y2=0
r208 86 110 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.97 $Y=0 $X2=3.91
+ $Y2=0
r209 86 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.97 $Y=0 $X2=4.1
+ $Y2=0
r210 85 113 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.83
+ $Y2=0
r211 85 87 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.23 $Y=0 $X2=4.1
+ $Y2=0
r212 83 107 1.30481 $w=1.68e-07 $l=2e-08 $layer=LI1_cond $X=3.01 $Y=0 $X2=2.99
+ $Y2=0
r213 83 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.01 $Y=0 $X2=3.14
+ $Y2=0
r214 82 110 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.91
+ $Y2=0
r215 82 84 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=3.27 $Y=0 $X2=3.14
+ $Y2=0
r216 78 141 3.01621 $w=3e-07 $l=1.05924e-07 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.922 $Y2=0
r217 78 80 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=9.875 $Y=0.085
+ $X2=9.875 $Y2=0.4
r218 74 102 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=8.895 $Y=0.085
+ $X2=8.895 $Y2=0
r219 74 76 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=8.895 $Y=0.085
+ $X2=8.895 $Y2=0.4
r220 70 99 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0
r221 70 72 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=7.93 $Y=0.085
+ $X2=7.93 $Y2=0.4
r222 66 96 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=6.97 $Y=0.085
+ $X2=6.97 $Y2=0
r223 66 68 14.5208 $w=2.48e-07 $l=3.15e-07 $layer=LI1_cond $X=6.97 $Y=0.085
+ $X2=6.97 $Y2=0.4
r224 62 93 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=6.012 $Y=0.085
+ $X2=6.012 $Y2=0
r225 62 64 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=6.012 $Y=0.085
+ $X2=6.012 $Y2=0.4
r226 58 90 0.066131 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=5.052 $Y=0.085
+ $X2=5.052 $Y2=0
r227 58 60 14.8171 $w=2.43e-07 $l=3.15e-07 $layer=LI1_cond $X=5.052 $Y=0.085
+ $X2=5.052 $Y2=0.4
r228 54 87 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.1 $Y=0.085
+ $X2=4.1 $Y2=0
r229 54 56 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=4.1 $Y=0.085
+ $X2=4.1 $Y2=0.4
r230 50 84 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0
r231 50 52 13.9623 $w=2.58e-07 $l=3.15e-07 $layer=LI1_cond $X=3.14 $Y=0.085
+ $X2=3.14 $Y2=0.4
r232 46 138 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r233 46 48 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.445
r234 45 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.35 $Y=0 $X2=1.22
+ $Y2=0
r235 44 138 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=2.18
+ $Y2=0
r236 44 45 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=2.05 $Y=0 $X2=1.35
+ $Y2=0
r237 40 135 0.132371 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r238 40 42 15.9569 $w=2.58e-07 $l=3.6e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.445
r239 39 132 4.57719 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=0.39 $Y=0
+ $X2=0.195 $Y2=0
r240 38 135 7.24004 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=1.22
+ $Y2=0
r241 38 39 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.09 $Y=0 $X2=0.39
+ $Y2=0
r242 34 132 2.98104 $w=3.05e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.195 $Y2=0
r243 34 36 11.1466 $w=3.03e-07 $l=2.95e-07 $layer=LI1_cond $X=0.237 $Y=0.085
+ $X2=0.237 $Y2=0.38
r244 11 80 182 $w=1.7e-07 $l=2.24332e-07 $layer=licon1_NDIFF $count=1 $X=9.715
+ $Y=0.235 $X2=9.855 $Y2=0.4
r245 10 76 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=8.705
+ $Y=0.235 $X2=8.895 $Y2=0.4
r246 9 72 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.935 $Y2=0.4
r247 8 68 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=6.785
+ $Y=0.235 $X2=6.975 $Y2=0.4
r248 7 64 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=5.83
+ $Y=0.235 $X2=6.02 $Y2=0.4
r249 6 60 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=5.06 $Y2=0.4
r250 5 56 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=3.91
+ $Y=0.235 $X2=4.1 $Y2=0.4
r251 4 52 182 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=1 $X=2.95
+ $Y=0.235 $X2=3.14 $Y2=0.4
r252 3 48 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=2.04
+ $Y=0.235 $X2=2.18 $Y2=0.445
r253 2 42 182 $w=1.7e-07 $l=2.71109e-07 $layer=licon1_NDIFF $count=1 $X=1.08
+ $Y=0.235 $X2=1.22 $Y2=0.445
r254 1 36 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

