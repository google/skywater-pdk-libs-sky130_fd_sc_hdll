* File: sky130_fd_sc_hdll__inputiso1p_1.pxi.spice
* Created: Thu Aug 27 19:08:50 2020
* 
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A N_A_c_36_n N_A_M1004_g N_A_M1000_g A A
+ PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%SLEEP N_SLEEP_M1003_g N_SLEEP_c_60_n
+ N_SLEEP_M1001_g SLEEP SLEEP PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%SLEEP
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A_44_297# N_A_44_297#_M1000_d
+ N_A_44_297#_M1004_s N_A_44_297#_c_89_n N_A_44_297#_M1002_g N_A_44_297#_c_90_n
+ N_A_44_297#_M1005_g N_A_44_297#_c_91_n N_A_44_297#_c_109_n N_A_44_297#_c_95_n
+ N_A_44_297#_c_92_n N_A_44_297#_c_102_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%A_44_297#
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VPWR N_VPWR_M1001_d N_VPWR_c_138_n
+ N_VPWR_c_139_n N_VPWR_c_140_n VPWR N_VPWR_c_141_n N_VPWR_c_137_n
+ PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VPWR
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%X N_X_M1002_d N_X_M1005_d N_X_c_157_n X X
+ PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%X
x_PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VGND N_VGND_M1000_s N_VGND_M1003_d
+ N_VGND_c_175_n N_VGND_c_176_n N_VGND_c_177_n N_VGND_c_178_n N_VGND_c_179_n
+ VGND N_VGND_c_180_n N_VGND_c_181_n PM_SKY130_FD_SC_HDLL__INPUTISO1P_1%VGND
cc_1 VNB N_A_c_36_n 0.0408906f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.41
cc_2 VNB N_A_M1000_g 0.0331738f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.445
cc_3 VNB A 0.0261632f $X=-0.19 $Y=-0.24 $X2=0.085 $Y2=0.765
cc_4 VNB N_SLEEP_M1003_g 0.0293131f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.695
cc_5 VNB N_SLEEP_c_60_n 0.0244764f $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=0.445
cc_6 VNB SLEEP 0.00535294f $X=-0.19 $Y=-0.24 $X2=0.085 $Y2=0.765
cc_7 VNB N_A_44_297#_c_89_n 0.0206197f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_44_297#_c_90_n 0.0245003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_44_297#_c_91_n 0.00425168f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_10 VNB N_A_44_297#_c_92_n 0.00161632f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_VPWR_c_137_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_X_c_157_n 0.0285407f $X=-0.19 $Y=-0.24 $X2=0.085 $Y2=1.105
cc_13 VNB X 0.0262965f $X=-0.19 $Y=-0.24 $X2=0.435 $Y2=1.16
cc_14 VNB N_VGND_c_175_n 0.0124942f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_176_n 0.0185131f $X=-0.19 $Y=-0.24 $X2=0.085 $Y2=1.105
cc_16 VNB N_VGND_c_177_n 0.00498362f $X=-0.19 $Y=-0.24 $X2=0.355 $Y2=1.16
cc_17 VNB N_VGND_c_178_n 0.0220497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_179_n 0.00410958f $X=-0.19 $Y=-0.24 $X2=0.262 $Y2=1.16
cc_19 VNB N_VGND_c_180_n 0.0245139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_181_n 0.144549f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VPB N_A_c_36_n 0.0411351f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.41
cc_22 VPB A 0.00599725f $X=-0.19 $Y=1.305 $X2=0.085 $Y2=0.765
cc_23 VPB N_SLEEP_c_60_n 0.0290484f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.445
cc_24 VPB SLEEP 0.00166667f $X=-0.19 $Y=1.305 $X2=0.085 $Y2=0.765
cc_25 VPB N_A_44_297#_c_90_n 0.032781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_44_297#_c_91_n 0.00166053f $X=-0.19 $Y=1.305 $X2=0.355 $Y2=1.16
cc_27 VPB N_A_44_297#_c_95_n 0.0176291f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_28 VPB N_A_44_297#_c_92_n 0.0015314f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_138_n 0.0216266f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=0.445
cc_30 VPB N_VPWR_c_139_n 0.0398524f $X=-0.19 $Y=1.305 $X2=0.085 $Y2=1.105
cc_31 VPB N_VPWR_c_140_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_141_n 0.0221444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_137_n 0.0808613f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB X 0.0251137f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_35 VPB X 0.0276962f $X=-0.19 $Y=1.305 $X2=0.262 $Y2=1.19
cc_36 N_A_M1000_g N_SLEEP_M1003_g 0.020427f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_37 N_A_c_36_n N_SLEEP_c_60_n 0.0479471f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_38 N_A_M1000_g SLEEP 5.08993e-19 $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_39 N_A_c_36_n N_A_44_297#_c_91_n 0.0181419f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_40 N_A_M1000_g N_A_44_297#_c_91_n 0.0134287f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_41 A N_A_44_297#_c_91_n 0.0419086f $X=0.085 $Y=0.765 $X2=0 $Y2=0
cc_42 N_A_c_36_n N_A_44_297#_c_95_n 0.0235594f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_43 A N_A_44_297#_c_95_n 0.0236956f $X=0.085 $Y=0.765 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_A_44_297#_c_102_n 0.00521178f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_45 N_A_c_36_n N_VPWR_c_139_n 0.00393512f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_46 N_A_c_36_n N_VPWR_c_137_n 0.00500987f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_47 A N_VGND_c_175_n 0.00162397f $X=0.085 $Y=0.765 $X2=0 $Y2=0
cc_48 N_A_c_36_n N_VGND_c_176_n 0.00111494f $X=0.58 $Y=1.41 $X2=0 $Y2=0
cc_49 N_A_M1000_g N_VGND_c_176_n 0.00561241f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_50 A N_VGND_c_176_n 0.0209296f $X=0.085 $Y=0.765 $X2=0 $Y2=0
cc_51 N_A_M1000_g N_VGND_c_178_n 0.00481596f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_52 N_A_M1000_g N_VGND_c_181_n 0.00923392f $X=0.605 $Y=0.445 $X2=0 $Y2=0
cc_53 A N_VGND_c_181_n 0.00421253f $X=0.085 $Y=0.765 $X2=0 $Y2=0
cc_54 N_SLEEP_M1003_g N_A_44_297#_c_89_n 0.0190472f $X=1.025 $Y=0.445 $X2=0
+ $Y2=0
cc_55 SLEEP N_A_44_297#_c_89_n 0.00523523f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_56 N_SLEEP_c_60_n N_A_44_297#_c_90_n 0.038401f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_57 N_SLEEP_M1003_g N_A_44_297#_c_91_n 0.00941806f $X=1.025 $Y=0.445 $X2=0
+ $Y2=0
cc_58 N_SLEEP_c_60_n N_A_44_297#_c_91_n 0.0019407f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_59 SLEEP N_A_44_297#_c_91_n 0.0427403f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_60 N_SLEEP_c_60_n N_A_44_297#_c_109_n 0.0190232f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_61 SLEEP N_A_44_297#_c_109_n 0.0219959f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_62 N_SLEEP_c_60_n N_A_44_297#_c_95_n 8.48903e-19 $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_63 N_SLEEP_c_60_n N_A_44_297#_c_92_n 0.00131322f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_64 SLEEP N_A_44_297#_c_92_n 0.0204828f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_65 N_SLEEP_c_60_n N_VPWR_c_138_n 0.0040866f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_66 N_SLEEP_c_60_n N_VPWR_c_139_n 0.00393512f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_67 N_SLEEP_c_60_n N_VPWR_c_137_n 0.00500987f $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_68 SLEEP X 0.00413293f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_69 SLEEP N_VGND_M1003_d 0.00251175f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_70 N_SLEEP_M1003_g N_VGND_c_177_n 0.00614826f $X=1.025 $Y=0.445 $X2=0 $Y2=0
cc_71 N_SLEEP_c_60_n N_VGND_c_177_n 2.29546e-19 $X=1.05 $Y=1.41 $X2=0 $Y2=0
cc_72 SLEEP N_VGND_c_177_n 0.0080166f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_73 N_SLEEP_M1003_g N_VGND_c_178_n 0.00585385f $X=1.025 $Y=0.445 $X2=0 $Y2=0
cc_74 N_SLEEP_M1003_g N_VGND_c_181_n 0.00801125f $X=1.025 $Y=0.445 $X2=0 $Y2=0
cc_75 SLEEP N_VGND_c_181_n 0.00864001f $X=1.055 $Y=0.765 $X2=0 $Y2=0
cc_76 N_A_44_297#_c_109_n A_134_297# 0.0054944f $X=1.535 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_44_297#_c_95_n A_134_297# 0.00460127f $X=0.83 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_44_297#_c_109_n N_VPWR_M1001_d 0.0083705f $X=1.535 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_44_297#_c_90_n N_VPWR_c_138_n 0.0164735f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_44_297#_c_109_n N_VPWR_c_138_n 0.0210126f $X=1.535 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_44_297#_c_90_n N_VPWR_c_141_n 0.00622633f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_44_297#_c_90_n N_VPWR_c_137_n 0.0115811f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_44_297#_c_90_n N_X_c_157_n 0.00242142f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_44_297#_c_92_n N_X_c_157_n 0.00213172f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_44_297#_c_89_n X 0.0025624f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_86 N_A_44_297#_c_90_n X 0.0144663f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_44_297#_c_92_n X 0.0342014f $X=1.62 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_44_297#_c_90_n X 0.0144362f $X=1.585 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_44_297#_c_102_n N_VGND_c_176_n 0.0239215f $X=0.815 $Y=0.43 $X2=0 $Y2=0
cc_90 N_A_44_297#_c_89_n N_VGND_c_177_n 0.00291856f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A_44_297#_c_102_n N_VGND_c_178_n 0.0179341f $X=0.815 $Y=0.43 $X2=0 $Y2=0
cc_92 N_A_44_297#_c_89_n N_VGND_c_180_n 0.00585385f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_44_297#_M1000_d N_VGND_c_181_n 0.00250238f $X=0.68 $Y=0.235 $X2=0
+ $Y2=0
cc_94 N_A_44_297#_c_89_n N_VGND_c_181_n 0.0120719f $X=1.56 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_44_297#_c_102_n N_VGND_c_181_n 0.0121054f $X=0.815 $Y=0.43 $X2=0 $Y2=0
cc_96 N_VPWR_c_137_n N_X_M1005_d 0.00753152f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_97 N_VPWR_c_138_n X 0.0334613f $X=1.35 $Y=1.92 $X2=0 $Y2=0
cc_98 N_VPWR_c_141_n X 0.029522f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_99 N_VPWR_c_137_n X 0.0160882f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_100 N_X_c_157_n N_VGND_c_180_n 0.03773f $X=1.88 $Y=0.39 $X2=0 $Y2=0
cc_101 N_X_M1002_d N_VGND_c_181_n 0.00407918f $X=1.635 $Y=0.235 $X2=0 $Y2=0
cc_102 N_X_c_157_n N_VGND_c_181_n 0.0210632f $X=1.88 $Y=0.39 $X2=0 $Y2=0
