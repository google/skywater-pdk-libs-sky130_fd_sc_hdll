* File: sky130_fd_sc_hdll__nor4b_1.pxi.spice
* Created: Thu Aug 27 19:17:28 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%A_91_199# N_A_91_199#_M1008_d
+ N_A_91_199#_M1002_d N_A_91_199#_c_53_n N_A_91_199#_M1001_g N_A_91_199#_c_54_n
+ N_A_91_199#_M1006_g N_A_91_199#_c_55_n N_A_91_199#_c_60_n N_A_91_199#_c_85_p
+ N_A_91_199#_c_56_n N_A_91_199#_c_57_n PM_SKY130_FD_SC_HDLL__NOR4B_1%A_91_199#
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%C N_C_c_111_n N_C_M1000_g N_C_c_112_n
+ N_C_M1004_g C C PM_SKY130_FD_SC_HDLL__NOR4B_1%C
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%B N_B_c_139_n N_B_M1009_g N_B_c_140_n
+ N_B_M1003_g B B PM_SKY130_FD_SC_HDLL__NOR4B_1%B
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%A N_A_c_167_n N_A_M1007_g N_A_c_168_n
+ N_A_M1005_g A A PM_SKY130_FD_SC_HDLL__NOR4B_1%A
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%D_N N_D_N_M1008_g N_D_N_c_198_n N_D_N_c_199_n
+ N_D_N_M1002_g D_N N_D_N_c_196_n N_D_N_c_197_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_1%D_N
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_M1001_s
+ N_Y_c_226_n N_Y_c_227_n N_Y_c_253_p N_Y_c_239_n N_Y_c_260_p N_Y_c_242_n Y
+ PM_SKY130_FD_SC_HDLL__NOR4B_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%VPWR N_VPWR_M1005_d N_VPWR_c_278_n VPWR
+ N_VPWR_c_279_n N_VPWR_c_280_n N_VPWR_c_277_n N_VPWR_c_282_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4B_1%VGND N_VGND_M1006_s N_VGND_M1004_d
+ N_VGND_M1007_d N_VGND_c_309_n N_VGND_c_310_n N_VGND_c_311_n N_VGND_c_312_n
+ N_VGND_c_313_n N_VGND_c_314_n N_VGND_c_315_n VGND N_VGND_c_316_n
+ N_VGND_c_317_n N_VGND_c_318_n N_VGND_c_319_n
+ PM_SKY130_FD_SC_HDLL__NOR4B_1%VGND
cc_1 VNB N_A_91_199#_c_53_n 0.0325448f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_2 VNB N_A_91_199#_c_54_n 0.0203255f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.995
cc_3 VNB N_A_91_199#_c_55_n 0.0016809f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_4 VNB N_A_91_199#_c_56_n 0.0233369f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=1.795
cc_5 VNB N_A_91_199#_c_57_n 0.0195983f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.66
cc_6 VNB N_C_c_111_n 0.0229469f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.465
cc_7 VNB N_C_c_112_n 0.0178891f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB C 0.00309854f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_9 VNB N_B_c_139_n 0.0209862f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.465
cc_10 VNB N_B_c_140_n 0.0174501f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB B 0.00532903f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.41
cc_12 VNB N_A_c_167_n 0.0192807f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=0.465
cc_13 VNB N_A_c_168_n 0.0252199f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB A 0.00420726f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_15 VNB D_N 0.00623652f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.985
cc_16 VNB N_D_N_c_196_n 0.0314533f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_17 VNB N_D_N_c_197_n 0.0219832f $X=-0.19 $Y=-0.24 $X2=0.635 $Y2=1.16
cc_18 VNB N_Y_c_226_n 0.00144477f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.995
cc_19 VNB N_Y_c_227_n 0.0120961f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_20 VNB Y 0.0257734f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.655
cc_21 VNB N_VPWR_c_277_n 0.155873f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=1.9
cc_22 VNB N_VGND_c_309_n 0.0144276f $X=-0.19 $Y=-0.24 $X2=0.78 $Y2=0.56
cc_23 VNB N_VGND_c_310_n 0.00443151f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_24 VNB N_VGND_c_311_n 0.00362637f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=1.9
cc_25 VNB N_VGND_c_312_n 0.0122893f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=1.795
cc_26 VNB N_VGND_c_313_n 0.00631534f $X=-0.19 $Y=-0.24 $X2=3.175 $Y2=0.655
cc_27 VNB N_VGND_c_314_n 0.0167009f $X=-0.19 $Y=-0.24 $X2=3.48 $Y2=0.655
cc_28 VNB N_VGND_c_315_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0.655 $Y2=1.16
cc_29 VNB N_VGND_c_316_n 0.0150439f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_317_n 0.0297181f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_318_n 0.218721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_319_n 0.00818228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VPB N_A_91_199#_c_53_n 0.0351565f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_34 VPB N_A_91_199#_c_55_n 0.00150521f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_35 VPB N_A_91_199#_c_60_n 0.017699f $X=-0.19 $Y=1.305 $X2=3.395 $Y2=1.9
cc_36 VPB N_A_91_199#_c_56_n 0.0239135f $X=-0.19 $Y=1.305 $X2=3.48 $Y2=1.795
cc_37 VPB N_C_c_111_n 0.0265666f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=0.465
cc_38 VPB C 0.00109619f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_39 VPB N_B_c_139_n 0.025448f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=0.465
cc_40 VPB B 0.00236344f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.41
cc_41 VPB N_A_c_168_n 0.0297228f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB A 0.00130397f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_43 VPB N_D_N_c_198_n 0.012551f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_D_N_c_199_n 0.0308124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_45 VPB D_N 0.00723933f $X=-0.19 $Y=1.305 $X2=0.755 $Y2=1.985
cc_46 VPB N_D_N_c_196_n 0.00487631f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.56
cc_47 VPB Y 0.0464602f $X=-0.19 $Y=1.305 $X2=3.175 $Y2=0.655
cc_48 VPB N_VPWR_c_278_n 0.00590885f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_VPWR_c_279_n 0.066956f $X=-0.19 $Y=1.305 $X2=0.78 $Y2=0.995
cc_50 VPB N_VPWR_c_280_n 0.0298965f $X=-0.19 $Y=1.305 $X2=3.175 $Y2=1.9
cc_51 VPB N_VPWR_c_277_n 0.0548418f $X=-0.19 $Y=1.305 $X2=3.175 $Y2=1.9
cc_52 VPB N_VPWR_c_282_n 0.00727973f $X=-0.19 $Y=1.305 $X2=3.175 $Y2=0.655
cc_53 N_A_91_199#_c_53_n N_C_c_111_n 0.0800421f $X=0.755 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_91_199#_c_55_n N_C_c_111_n 0.00145018f $X=0.62 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A_91_199#_c_60_n N_C_c_111_n 0.0181666f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_56 N_A_91_199#_c_54_n N_C_c_112_n 0.0206964f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A_91_199#_c_53_n C 0.00459353f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_91_199#_c_55_n C 0.0438802f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_59 N_A_91_199#_c_60_n C 0.0221118f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_60 N_A_91_199#_c_60_n N_B_c_139_n 0.0163381f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_61 N_A_91_199#_c_60_n B 0.0260965f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_62 N_A_91_199#_c_60_n N_A_c_168_n 0.0185467f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_63 N_A_91_199#_c_60_n A 0.0323235f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_64 N_A_91_199#_c_56_n N_D_N_c_198_n 0.00127516f $X=3.48 $Y=1.795 $X2=0 $Y2=0
cc_65 N_A_91_199#_c_60_n N_D_N_c_199_n 0.0135648f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_66 N_A_91_199#_c_56_n N_D_N_c_199_n 0.00387776f $X=3.48 $Y=1.795 $X2=0 $Y2=0
cc_67 N_A_91_199#_c_60_n D_N 0.0277253f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_68 N_A_91_199#_c_56_n D_N 0.0499816f $X=3.48 $Y=1.795 $X2=0 $Y2=0
cc_69 N_A_91_199#_c_57_n D_N 0.0115587f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_70 N_A_91_199#_c_60_n N_D_N_c_196_n 3.7104e-19 $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_71 N_A_91_199#_c_56_n N_D_N_c_196_n 0.00192392f $X=3.48 $Y=1.795 $X2=0 $Y2=0
cc_72 N_A_91_199#_c_57_n N_D_N_c_196_n 0.0014913f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_73 N_A_91_199#_c_56_n N_D_N_c_197_n 0.00411682f $X=3.48 $Y=1.795 $X2=0 $Y2=0
cc_74 N_A_91_199#_c_57_n N_D_N_c_197_n 0.00336376f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_75 N_A_91_199#_c_55_n N_Y_M1001_s 0.00339944f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_91_199#_c_85_p N_Y_M1001_s 0.00402256f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_77 N_A_91_199#_c_53_n N_Y_c_226_n 0.00380065f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_91_199#_c_54_n N_Y_c_226_n 0.016961f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_91_199#_c_55_n N_Y_c_226_n 0.014961f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_91_199#_c_53_n Y 0.0258784f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_91_199#_c_54_n Y 0.00497439f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_91_199#_c_55_n Y 0.0587008f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_91_199#_c_85_p Y 0.0168523f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_84 N_A_91_199#_c_60_n A_169_297# 0.00621636f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_85 N_A_91_199#_c_60_n A_263_297# 0.00968698f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_91_199#_c_60_n A_369_297# 0.00931379f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_91_199#_c_60_n N_VPWR_M1005_d 0.0156566f $X=3.395 $Y=1.9 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_91_199#_c_60_n N_VPWR_c_278_n 0.0250066f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_89 N_A_91_199#_c_53_n N_VPWR_c_279_n 0.00523711f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_91_199#_c_60_n N_VPWR_c_279_n 0.0204801f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_91 N_A_91_199#_c_85_p N_VPWR_c_279_n 0.0030042f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_92 N_A_91_199#_c_60_n N_VPWR_c_280_n 0.0123248f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_93 N_A_91_199#_c_53_n N_VPWR_c_277_n 0.00822286f $X=0.755 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_91_199#_c_60_n N_VPWR_c_277_n 0.0639154f $X=3.395 $Y=1.9 $X2=0 $Y2=0
cc_95 N_A_91_199#_c_85_p N_VPWR_c_277_n 0.00581552f $X=0.745 $Y=1.9 $X2=0 $Y2=0
cc_96 N_A_91_199#_c_54_n N_VGND_c_309_n 0.00341589f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_91_199#_c_57_n N_VGND_c_311_n 0.0199887f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_98 N_A_91_199#_c_54_n N_VGND_c_314_n 0.00428022f $X=0.78 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_91_199#_c_57_n N_VGND_c_317_n 0.0116646f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_100 N_A_91_199#_c_54_n N_VGND_c_318_n 0.00698263f $X=0.78 $Y=0.995 $X2=0
+ $Y2=0
cc_101 N_A_91_199#_c_57_n N_VGND_c_318_n 0.0147176f $X=3.175 $Y=0.66 $X2=0 $Y2=0
cc_102 N_C_c_111_n N_B_c_139_n 0.0697151f $X=1.225 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_103 C N_B_c_139_n 5.48905e-19 $X=1.095 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_104 N_C_c_112_n N_B_c_140_n 0.0225663f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_105 N_C_c_111_n B 0.00450333f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_106 C B 0.0465599f $X=1.095 $Y=1.105 $X2=0 $Y2=0
cc_107 N_C_c_111_n N_Y_c_239_n 0.00287627f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_108 N_C_c_112_n N_Y_c_239_n 0.0133461f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_109 C N_Y_c_239_n 0.0116012f $X=1.095 $Y=1.105 $X2=0 $Y2=0
cc_110 N_C_c_111_n N_Y_c_242_n 9.23565e-19 $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_111 C N_Y_c_242_n 0.0149833f $X=1.095 $Y=1.105 $X2=0 $Y2=0
cc_112 C A_169_297# 0.00282179f $X=1.095 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_113 N_C_c_111_n N_VPWR_c_279_n 0.00523784f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_114 N_C_c_111_n N_VPWR_c_277_n 0.00727071f $X=1.225 $Y=1.41 $X2=0 $Y2=0
cc_115 N_C_c_112_n N_VGND_c_310_n 0.0018911f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_116 N_C_c_112_n N_VGND_c_314_n 0.00427293f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_117 N_C_c_112_n N_VGND_c_318_n 0.00605079f $X=1.25 $Y=0.995 $X2=0 $Y2=0
cc_118 N_B_c_140_n N_A_c_167_n 0.0241813f $X=1.78 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_119 N_B_c_139_n N_A_c_168_n 0.0798081f $X=1.755 $Y=1.41 $X2=0 $Y2=0
cc_120 B N_A_c_168_n 0.00416163f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_121 N_B_c_139_n A 6.7133e-19 $X=1.755 $Y=1.41 $X2=0 $Y2=0
cc_122 B A 0.0399166f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_123 N_B_c_139_n N_Y_c_239_n 0.00332807f $X=1.755 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_c_140_n N_Y_c_239_n 0.0115708f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_125 B N_Y_c_239_n 0.0320021f $X=1.625 $Y=1.105 $X2=0 $Y2=0
cc_126 B A_263_297# 0.00266339f $X=1.625 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_127 B A_369_297# 0.00166074f $X=1.625 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_128 N_B_c_139_n N_VPWR_c_279_n 0.00523784f $X=1.755 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B_c_139_n N_VPWR_c_277_n 0.00727071f $X=1.755 $Y=1.41 $X2=0 $Y2=0
cc_130 N_B_c_140_n N_VGND_c_310_n 0.00299011f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B_c_140_n N_VGND_c_311_n 8.85533e-19 $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_132 N_B_c_140_n N_VGND_c_316_n 0.00428022f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_140_n N_VGND_c_318_n 0.00611511f $X=1.78 $Y=0.995 $X2=0 $Y2=0
cc_134 N_A_c_168_n N_D_N_c_198_n 0.00496577f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_135 N_A_c_168_n N_D_N_c_199_n 0.0147764f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A_c_168_n D_N 0.00138594f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_137 A D_N 0.0539856f $X=2.51 $Y=1.19 $X2=0 $Y2=0
cc_138 N_A_c_168_n N_D_N_c_196_n 0.0093861f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_139 A N_D_N_c_196_n 0.00247252f $X=2.51 $Y=1.19 $X2=0 $Y2=0
cc_140 N_A_c_167_n N_D_N_c_197_n 0.011174f $X=2.2 $Y=0.995 $X2=0 $Y2=0
cc_141 A N_VPWR_M1005_d 0.0052813f $X=2.51 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_142 N_A_c_168_n N_VPWR_c_278_n 0.0107179f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_168_n N_VPWR_c_279_n 0.00523784f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_168_n N_VPWR_c_277_n 0.00821171f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_167_n N_VGND_c_311_n 0.0232412f $X=2.2 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_168_n N_VGND_c_311_n 0.00395521f $X=2.225 $Y=1.41 $X2=0 $Y2=0
cc_147 A N_VGND_c_311_n 0.0336371f $X=2.51 $Y=1.19 $X2=0 $Y2=0
cc_148 N_A_c_167_n N_VGND_c_316_n 0.0046653f $X=2.2 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A_c_167_n N_VGND_c_318_n 0.00799591f $X=2.2 $Y=0.995 $X2=0 $Y2=0
cc_150 N_D_N_c_199_n N_VPWR_c_278_n 0.00124992f $X=2.94 $Y=1.605 $X2=0 $Y2=0
cc_151 N_D_N_c_199_n N_VPWR_c_280_n 0.00393205f $X=2.94 $Y=1.605 $X2=0 $Y2=0
cc_152 N_D_N_c_199_n N_VPWR_c_277_n 0.00561636f $X=2.94 $Y=1.605 $X2=0 $Y2=0
cc_153 N_D_N_c_197_n N_VGND_c_311_n 0.00759411f $X=2.997 $Y=0.995 $X2=0 $Y2=0
cc_154 N_D_N_c_197_n N_VGND_c_317_n 0.00510437f $X=2.997 $Y=0.995 $X2=0 $Y2=0
cc_155 N_D_N_c_197_n N_VGND_c_318_n 0.00512902f $X=2.997 $Y=0.995 $X2=0 $Y2=0
cc_156 Y N_VPWR_c_279_n 0.0166143f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_157 N_Y_M1001_s N_VPWR_c_277_n 0.0112757f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_158 Y N_VPWR_c_277_n 0.00986501f $X=0.145 $Y=1.785 $X2=0 $Y2=0
cc_159 N_Y_c_226_n N_VGND_M1006_s 0.00904954f $X=0.905 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_160 N_Y_c_239_n N_VGND_M1004_d 0.00806359f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_161 N_Y_c_226_n N_VGND_c_309_n 0.021906f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_162 N_Y_c_253_p N_VGND_c_310_n 0.0121114f $X=0.99 $Y=0.495 $X2=0 $Y2=0
cc_163 N_Y_c_239_n N_VGND_c_310_n 0.0204201f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_164 N_Y_c_227_n N_VGND_c_312_n 0.00506771f $X=0.345 $Y=0.74 $X2=0 $Y2=0
cc_165 N_Y_c_226_n N_VGND_c_314_n 0.0029785f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_166 N_Y_c_253_p N_VGND_c_314_n 0.0104406f $X=0.99 $Y=0.495 $X2=0 $Y2=0
cc_167 N_Y_c_239_n N_VGND_c_314_n 0.00306813f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_168 N_Y_c_239_n N_VGND_c_316_n 0.0029785f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_169 N_Y_c_260_p N_VGND_c_316_n 0.00906533f $X=1.99 $Y=0.495 $X2=0 $Y2=0
cc_170 N_Y_M1006_d N_VGND_c_318_n 0.00304673f $X=0.855 $Y=0.235 $X2=0 $Y2=0
cc_171 N_Y_M1003_d N_VGND_c_318_n 0.00403782f $X=1.855 $Y=0.235 $X2=0 $Y2=0
cc_172 N_Y_c_226_n N_VGND_c_318_n 0.00706381f $X=0.905 $Y=0.74 $X2=0 $Y2=0
cc_173 N_Y_c_227_n N_VGND_c_318_n 0.00770874f $X=0.345 $Y=0.74 $X2=0 $Y2=0
cc_174 N_Y_c_253_p N_VGND_c_318_n 0.00739742f $X=0.99 $Y=0.495 $X2=0 $Y2=0
cc_175 N_Y_c_239_n N_VGND_c_318_n 0.012146f $X=1.875 $Y=0.74 $X2=0 $Y2=0
cc_176 N_Y_c_260_p N_VGND_c_318_n 0.00735151f $X=1.99 $Y=0.495 $X2=0 $Y2=0
cc_177 A_169_297# N_VPWR_c_277_n 0.0037272f $X=0.845 $Y=1.485 $X2=3.175 $Y2=1.9
cc_178 A_263_297# N_VPWR_c_277_n 0.00449835f $X=1.315 $Y=1.485 $X2=3.175 $Y2=1.9
cc_179 A_369_297# N_VPWR_c_277_n 0.0037272f $X=1.845 $Y=1.485 $X2=3.175 $Y2=1.9
