* File: sky130_fd_sc_hdll__o21bai_4.spice
* Created: Wed Sep  2 08:44:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o21bai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o21bai_4  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1009 N_A_33_297#_M1009_d N_B1_N_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.2145 PD=1.82 PS=1.96 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.3 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1006 N_A_245_47#_M1006_d N_A_33_297#_M1006_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1013 N_A_245_47#_M1013_d N_A_33_297#_M1013_g N_Y_M1006_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1019 N_A_245_47#_M1013_d N_A_33_297#_M1019_g N_Y_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1024 N_A_245_47#_M1024_d N_A_33_297#_M1024_g N_Y_M1019_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.6 SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1004 N_A_245_47#_M1024_d N_A2_M1004_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.104 PD=0.92 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1010 N_A_245_47#_M1010_d N_A2_M1010_g N_VGND_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1017 N_A_245_47#_M1010_d N_A2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1018 N_A_245_47#_M1018_d N_A2_M1018_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A1_M1005_g N_A_245_47#_M1018_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.9
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1005_d N_A1_M1007_g N_A_245_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.4
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1020 N_VGND_M1020_d N_A1_M1020_g N_A_245_47#_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75004.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1020_d N_A1_M1023_g N_A_245_47#_M1023_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.169 PD=1.02 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_B1_N_M1008_g N_A_33_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_A_33_297#_M1001_g N_VPWR_M1008_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1001_d N_A_33_297#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1014 N_Y_M1014_d N_A_33_297#_M1014_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1021 N_Y_M1014_d N_A_33_297#_M1021_g N_VPWR_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1002 N_Y_M1002_d N_A2_M1002_g N_A_621_297#_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1012 N_Y_M1002_d N_A2_M1012_g N_A_621_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90003 A=0.18 P=2.36 MULT=1
MM1016 N_Y_M1016_d N_A2_M1016_g N_A_621_297#_M1012_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1025 N_Y_M1016_d N_A2_M1025_g N_A_621_297#_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1000 N_A_621_297#_M1025_s N_A1_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_621_297#_M1003_d N_A1_M1003_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1015 N_A_621_297#_M1003_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1022 N_A_621_297#_M1022_d N_A1_M1022_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.145 PD=2.58 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX26_noxref VNB VPB NWDIODE A=12.4227 P=18.69
pX27_noxref noxref_12 B1_N B1_N PROBETYPE=1
pX28_noxref noxref_13 A2 A2 PROBETYPE=1
pX29_noxref noxref_14 A1 A1 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o21bai_4.pxi.spice"
*
.ends
*
*
