* File: sky130_fd_sc_hdll__xor3_1.pex.spice
* Created: Thu Aug 27 19:30:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_116_21# 1 2 7 9 10 12 16 18 19 20 21 23
+ 25 27 28 30 33 34
c102 19 0 1.62085e-19 $X=1 $Y=0.78
r103 33 34 13.3132 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=2.725 $Y=0.355
+ $X2=2.49 $Y2=0.355
r104 28 30 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=1.57 $Y=2.32
+ $X2=2.73 $Y2=2.32
r105 27 34 67.8503 $w=1.68e-07 $l=1.04e-06 $layer=LI1_cond $X=1.45 $Y=0.34
+ $X2=2.49 $Y2=0.34
r106 25 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.46 $Y=2.235
+ $X2=1.57 $Y2=2.32
r107 24 25 9.95292 $w=2.18e-07 $l=1.9e-07 $layer=LI1_cond $X=1.46 $Y=2.045
+ $X2=1.46 $Y2=2.235
r108 22 27 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.45 $Y2=0.34
r109 22 23 14.1436 $w=2.18e-07 $l=2.7e-07 $layer=LI1_cond $X=1.34 $Y=0.425
+ $X2=1.34 $Y2=0.695
r110 20 24 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.35 $Y=1.96
+ $X2=1.46 $Y2=2.045
r111 20 21 22.8342 $w=1.68e-07 $l=3.5e-07 $layer=LI1_cond $X=1.35 $Y=1.96 $X2=1
+ $Y2=1.96
r112 18 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.23 $Y=0.78
+ $X2=1.34 $Y2=0.695
r113 18 19 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.23 $Y=0.78 $X2=1
+ $Y2=0.78
r114 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.885
+ $Y=1.16 $X2=0.885 $Y2=1.16
r115 14 21 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.9 $Y=1.875
+ $X2=1 $Y2=1.96
r116 14 16 39.65 $w=1.98e-07 $l=7.15e-07 $layer=LI1_cond $X=0.9 $Y=1.875 $X2=0.9
+ $Y2=1.16
r117 13 19 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=0.9 $Y=0.865
+ $X2=1 $Y2=0.78
r118 13 16 16.3591 $w=1.98e-07 $l=2.95e-07 $layer=LI1_cond $X=0.9 $Y=0.865
+ $X2=0.9 $Y2=1.16
r119 10 17 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=0.68 $Y=1.41
+ $X2=0.8 $Y2=1.16
r120 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.68 $Y=1.41
+ $X2=0.68 $Y2=1.985
r121 7 17 39.3952 $w=3.9e-07 $l=2.26164e-07 $layer=POLY_cond $X=0.655 $Y=0.995
+ $X2=0.8 $Y2=1.16
r122 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.655 $Y=0.995
+ $X2=0.655 $Y2=0.56
r123 2 30 600 $w=1.7e-07 $l=7.84267e-07 $layer=licon1_PDIFF $count=1 $X=2.54
+ $Y=1.625 $X2=2.73 $Y2=2.32
r124 1 33 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.59
+ $Y=0.245 $X2=2.725 $Y2=0.37
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%C 1 3 7 8 10 12 13 15 16 18 22 24
r64 18 22 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=2.105 $Y=1.16
+ $X2=2.41 $Y2=1.16
r65 18 24 1.22229 $w=3.28e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=1.16
+ $X2=2.07 $Y2=1.16
r66 13 15 134.96 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=2.515 $Y=0.985
+ $X2=2.515 $Y2=0.565
r67 10 12 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=2.45 $Y=1.55
+ $X2=2.45 $Y2=2.045
r68 9 16 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.43 $Y=1.16
+ $X2=1.33 $Y2=1.202
r69 8 10 85.013 $w=2.27e-07 $l=4.00849e-07 $layer=POLY_cond $X=2.472 $Y=1.16
+ $X2=2.45 $Y2=1.55
r70 8 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=2.41 $Y=1.16
+ $X2=2.41 $Y2=1.16
r71 8 13 42.7097 $w=2.27e-07 $l=1.9532e-07 $layer=POLY_cond $X=2.472 $Y=1.16
+ $X2=2.515 $Y2=0.985
r72 8 9 160.872 $w=3.3e-07 $l=9.2e-07 $layer=POLY_cond $X=2.35 $Y=1.16 $X2=1.43
+ $Y2=1.16
r73 4 16 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.33 $Y=1.41
+ $X2=1.33 $Y2=1.202
r74 4 7 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.33 $Y=1.41 $X2=1.33
+ $Y2=1.805
r75 1 16 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.305 $Y=0.995
+ $X2=1.33 $Y2=1.202
r76 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.305 $Y=0.995
+ $X2=1.305 $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_276_93# 1 2 7 9 10 12 13 18 20 23 24 28
r75 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.005
+ $Y=1.16 $X2=3.005 $Y2=1.16
r76 25 28 3.66686 $w=3.28e-07 $l=1.05e-07 $layer=LI1_cond $X=2.9 $Y=1.16
+ $X2=3.005 $Y2=1.16
r77 22 25 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.9 $Y=1.325 $X2=2.9
+ $Y2=1.16
r78 22 23 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=2.9 $Y=1.325 $X2=2.9
+ $Y2=1.535
r79 21 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.79 $Y=1.62
+ $X2=1.705 $Y2=1.62
r80 20 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.815 $Y=1.62
+ $X2=2.9 $Y2=1.535
r81 20 21 66.8717 $w=1.68e-07 $l=1.025e-06 $layer=LI1_cond $X=2.815 $Y=1.62
+ $X2=1.79 $Y2=1.62
r82 16 24 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.705 $Y=1.535
+ $X2=1.705 $Y2=1.62
r83 16 18 50.5615 $w=1.68e-07 $l=7.75e-07 $layer=LI1_cond $X=1.705 $Y=1.535
+ $X2=1.705 $Y2=0.76
r84 13 24 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=1.62
+ $X2=1.705 $Y2=1.62
r85 13 15 3.94706 $w=1.7e-07 $l=5.5e-08 $layer=LI1_cond $X=1.62 $Y=1.62
+ $X2=1.565 $Y2=1.62
r86 10 29 38.8824 $w=2.71e-07 $l=2.03101e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.03 $Y2=1.16
r87 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=3.115 $Y=0.995
+ $X2=3.115 $Y2=0.565
r88 7 29 74.8096 $w=2.71e-07 $l=3.9e-07 $layer=POLY_cond $X=3.03 $Y=1.55
+ $X2=3.03 $Y2=1.16
r89 7 9 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=3.03 $Y=1.55 $X2=3.03
+ $Y2=2.045
r90 2 15 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.42
+ $Y=1.485 $X2=1.565 $Y2=1.62
r91 1 18 182 $w=1.7e-07 $l=4.48888e-07 $layer=licon1_NDIFF $count=1 $X=1.38
+ $Y=0.465 $X2=1.705 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_875_297# 1 2 7 9 12 15 16 18 21 22 23 27
+ 35 37 38 39 40 47 49 50 55 57 60
c181 55 0 1.24749e-19 $X=7.7 $Y=1.11
r182 55 58 37.8858 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.722 $Y=1.11
+ $X2=7.722 $Y2=1.275
r183 55 57 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=7.722 $Y=1.11
+ $X2=7.722 $Y2=0.945
r184 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.7
+ $Y=1.11 $X2=7.7 $Y2=1.11
r185 50 56 11.8358 $w=2.68e-07 $l=2.6e-07 $layer=LI1_cond $X=7.63 $Y=0.85
+ $X2=7.63 $Y2=1.11
r186 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.58 $Y=0.85
+ $X2=7.58 $Y2=0.85
r187 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=0.85 $X2=6.1
+ $Y2=0.85
r188 42 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.62 $Y=0.85
+ $X2=4.62 $Y2=0.85
r189 40 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=6.245 $Y=0.85
+ $X2=6.1 $Y2=0.85
r190 39 49 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.435 $Y=0.85
+ $X2=7.58 $Y2=0.85
r191 39 40 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=7.435 $Y=0.85
+ $X2=6.245 $Y2=0.85
r192 38 42 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.765 $Y=0.85
+ $X2=4.62 $Y2=0.85
r193 37 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=0.85
+ $X2=6.1 $Y2=0.85
r194 37 38 1.47277 $w=1.4e-07 $l=1.19e-06 $layer=MET1_cond $X=5.955 $Y=0.85
+ $X2=4.765 $Y2=0.85
r195 35 47 7.77229 $w=2.13e-07 $l=1.45e-07 $layer=LI1_cond $X=6.077 $Y=0.995
+ $X2=6.077 $Y2=0.85
r196 31 35 6.36987 $w=2.73e-07 $l=1.52e-07 $layer=LI1_cond $X=5.925 $Y=1.132
+ $X2=6.077 $Y2=1.132
r197 31 32 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.925
+ $Y=1.16 $X2=5.925 $Y2=1.16
r198 28 60 28.8111 $w=2.88e-07 $l=7.25e-07 $layer=LI1_cond $X=4.675 $Y=1.445
+ $X2=4.675 $Y2=0.72
r199 27 28 0.275955 $w=2.9e-07 $l=1.35e-07 $layer=LI1_cond $X=4.675 $Y=1.58
+ $X2=4.675 $Y2=1.445
r200 25 27 6.61588 $w=2.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.52 $Y=1.58
+ $X2=4.675 $Y2=1.58
r201 22 32 46.3382 $w=3.3e-07 $l=2.65e-07 $layer=POLY_cond $X=6.19 $Y=1.16
+ $X2=5.925 $Y2=1.16
r202 22 23 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=6.19 $Y=1.16
+ $X2=6.29 $Y2=1.202
r203 21 57 131.747 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=7.805 $Y=0.535
+ $X2=7.805 $Y2=0.945
r204 16 18 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=7.78 $Y=1.57
+ $X2=7.78 $Y2=2.065
r205 15 16 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.78 $Y=1.47 $X2=7.78
+ $Y2=1.57
r206 15 58 64.6575 $w=2e-07 $l=1.95e-07 $layer=POLY_cond $X=7.78 $Y=1.47
+ $X2=7.78 $Y2=1.275
r207 10 23 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=6.315 $Y=0.995
+ $X2=6.29 $Y2=1.202
r208 10 12 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=6.315 $Y=0.995
+ $X2=6.315 $Y2=0.455
r209 7 23 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.202
r210 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=6.29 $Y=1.41
+ $X2=6.29 $Y2=1.805
r211 2 25 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.375
+ $Y=1.485 $X2=4.52 $Y2=1.63
r212 1 60 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=4.6
+ $Y=0.235 $X2=4.735 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%B 1 3 6 8 9 13 16 18 19 22 24 25 28 31 33
+ 35 36 40 42 45
c137 42 0 1.94872e-19 $X=7.495 $Y=1.5
r138 38 42 11.3186 $w=2.78e-07 $l=2.75e-07 $layer=LI1_cond $X=7.305 $Y=1.585
+ $X2=7.58 $Y2=1.585
r139 38 40 3.05577 $w=2.8e-07 $l=1.1e-07 $layer=LI1_cond $X=7.305 $Y=1.585
+ $X2=7.195 $Y2=1.585
r140 36 46 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.16
+ $X2=7.195 $Y2=1.325
r141 36 45 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.195 $Y=1.16
+ $X2=7.195 $Y2=0.995
r142 35 36 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.17
+ $Y=1.16 $X2=7.17 $Y2=1.16
r143 33 40 3.88917 $w=2.2e-07 $l=1.4e-07 $layer=LI1_cond $X=7.195 $Y=1.445
+ $X2=7.195 $Y2=1.585
r144 33 35 14.9294 $w=2.18e-07 $l=2.85e-07 $layer=LI1_cond $X=7.195 $Y=1.445
+ $X2=7.195 $Y2=1.16
r145 31 32 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=5.48 $Y=1.16 $X2=5.48
+ $Y2=1.085
r146 26 28 174.919 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=7.215 $Y=2.415
+ $X2=7.215 $Y2=1.965
r147 25 28 153.54 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=7.215 $Y=1.57
+ $X2=7.215 $Y2=1.965
r148 24 25 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.215 $Y=1.47 $X2=7.215
+ $Y2=1.57
r149 24 46 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=7.215 $Y=1.47
+ $X2=7.215 $Y2=1.325
r150 22 45 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=7.11 $Y=0.565
+ $X2=7.11 $Y2=0.995
r151 18 26 27.2212 $w=1.5e-07 $l=1.67705e-07 $layer=POLY_cond $X=7.115 $Y=2.54
+ $X2=7.215 $Y2=2.415
r152 18 19 787.096 $w=1.5e-07 $l=1.535e-06 $layer=POLY_cond $X=7.115 $Y=2.54
+ $X2=5.58 $Y2=2.54
r153 16 32 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=5.505 $Y=0.565
+ $X2=5.505 $Y2=1.085
r154 11 19 27.2212 $w=1.5e-07 $l=1.36015e-07 $layer=POLY_cond $X=5.48 $Y=2.455
+ $X2=5.58 $Y2=2.54
r155 11 13 213.79 $w=1.8e-07 $l=5.5e-07 $layer=POLY_cond $X=5.48 $Y=2.455
+ $X2=5.48 $Y2=1.905
r156 10 31 83.702 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=5.48 $Y=1.41 $X2=5.48
+ $Y2=1.16
r157 10 13 192.411 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=5.48 $Y=1.41
+ $X2=5.48 $Y2=1.905
r158 8 31 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=5.38 $Y=1.16 $X2=5.48
+ $Y2=1.16
r159 8 9 399.957 $w=1.5e-07 $l=7.8e-07 $layer=POLY_cond $X=5.38 $Y=1.16 $X2=4.6
+ $Y2=1.16
r160 4 9 21.6409 $w=2.34e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.525 $Y=1.085
+ $X2=4.6 $Y2=1.16
r161 4 6 269.202 $w=1.5e-07 $l=5.25e-07 $layer=POLY_cond $X=4.525 $Y=1.085
+ $X2=4.525 $Y2=0.56
r162 1 4 49.4359 $w=2.34e-07 $l=3.38349e-07 $layer=POLY_cond $X=4.285 $Y=1.322
+ $X2=4.525 $Y2=1.085
r163 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.285 $Y=1.41
+ $X2=4.285 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A 1 3 4 6 7 15
c37 1 0 1.94872e-19 $X=8.335 $Y=1.41
r38 11 15 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=8.23 $Y=1.2
+ $X2=8.505 $Y2=1.2
r39 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.23
+ $Y=1.16 $X2=8.23 $Y2=1.16
r40 7 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=8.51 $Y=1.2 $X2=8.505
+ $Y2=1.2
r41 4 10 38.532 $w=3.11e-07 $l=2.07123e-07 $layer=POLY_cond $X=8.36 $Y=0.995
+ $X2=8.265 $Y2=1.16
r42 4 6 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.36 $Y=0.995 $X2=8.36
+ $Y2=0.555
r43 1 10 47.2262 $w=3.11e-07 $l=2.82843e-07 $layer=POLY_cond $X=8.335 $Y=1.41
+ $X2=8.265 $Y2=1.16
r44 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.335 $Y=1.41
+ $X2=8.335 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_991_365# 1 2 3 4 13 15 16 18 21 23 27 28
+ 29 30 36 37 40 43 44
c129 30 0 1.4108e-19 $X=9.03 $Y=1.495
c130 27 0 1.2773e-19 $X=8.945 $Y=0.82
r131 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.09 $Y=0.51
+ $X2=8.09 $Y2=0.51
r132 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.13 $Y=0.51
+ $X2=5.13 $Y2=0.51
r133 37 39 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.275 $Y=0.51
+ $X2=5.13 $Y2=0.51
r134 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=7.945 $Y=0.51
+ $X2=8.09 $Y2=0.51
r135 36 37 3.30445 $w=1.4e-07 $l=2.67e-06 $layer=MET1_cond $X=7.945 $Y=0.51
+ $X2=5.275 $Y2=0.51
r136 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.09
+ $Y=1.16 $X2=9.09 $Y2=1.16
r137 32 34 17.9567 $w=2.31e-07 $l=3.4e-07 $layer=LI1_cond $X=9.085 $Y=0.82
+ $X2=9.085 $Y2=1.16
r138 31 44 8.94137 $w=2.88e-07 $l=2.25e-07 $layer=LI1_cond $X=8.12 $Y=0.735
+ $X2=8.12 $Y2=0.51
r139 29 34 9.58904 $w=2.31e-07 $l=1.90526e-07 $layer=LI1_cond $X=9.03 $Y=1.325
+ $X2=9.085 $Y2=1.16
r140 29 30 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=9.03 $Y=1.325
+ $X2=9.03 $Y2=1.495
r141 28 31 14.5133 $w=1.17e-07 $l=1.8262e-07 $layer=LI1_cond $X=8.265 $Y=0.82
+ $X2=8.12 $Y2=0.735
r142 27 32 2.5345 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=8.945 $Y=0.82
+ $X2=9.085 $Y2=0.82
r143 27 28 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=8.945 $Y=0.82
+ $X2=8.265 $Y2=0.82
r144 23 30 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=8.945 $Y=1.6
+ $X2=9.03 $Y2=1.495
r145 23 25 44.6277 $w=2.08e-07 $l=8.45e-07 $layer=LI1_cond $X=8.945 $Y=1.6
+ $X2=8.1 $Y2=1.6
r146 19 40 3.61456 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.08 $Y=0.595
+ $X2=5.08 $Y2=0.43
r147 19 21 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=5.08 $Y=0.595
+ $X2=5.08 $Y2=1.94
r148 16 35 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=9.14 $Y=0.995
+ $X2=9.115 $Y2=1.16
r149 16 18 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=9.14 $Y=0.995
+ $X2=9.14 $Y2=0.555
r150 13 35 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=9.115 $Y=1.41
+ $X2=9.115 $Y2=1.16
r151 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.115 $Y=1.41
+ $X2=9.115 $Y2=1.985
r152 4 25 600 $w=1.7e-07 $l=2.42178e-07 $layer=licon1_PDIFF $count=1 $X=7.87
+ $Y=1.645 $X2=8.1 $Y2=1.62
r153 3 21 600 $w=1.7e-07 $l=1.73205e-07 $layer=licon1_PDIFF $count=1 $X=4.955
+ $Y=1.825 $X2=5.08 $Y2=1.94
r154 2 44 182 $w=1.7e-07 $l=4.8775e-07 $layer=licon1_NDIFF $count=1 $X=7.88
+ $Y=0.235 $X2=8.1 $Y2=0.625
r155 1 40 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=5.12
+ $Y=0.245 $X2=5.245 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%X 1 2 10 15 16 17
r24 17 22 9.79645 $w=5.23e-07 $l=4.3e-07 $layer=LI1_cond $X=0.347 $Y=1.87
+ $X2=0.347 $Y2=2.3
r25 15 16 5.99972 $w=5.23e-07 $l=1.8e-07 $layer=LI1_cond $X=0.347 $Y=1.62
+ $X2=0.347 $Y2=1.44
r26 13 17 3.82745 $w=5.23e-07 $l=1.68e-07 $layer=LI1_cond $X=0.347 $Y=1.702
+ $X2=0.347 $Y2=1.87
r27 13 15 1.86816 $w=5.23e-07 $l=8.2e-08 $layer=LI1_cond $X=0.347 $Y=1.702
+ $X2=0.347 $Y2=1.62
r28 12 16 18.8415 $w=3.13e-07 $l=5.15e-07 $layer=LI1_cond $X=0.242 $Y=0.925
+ $X2=0.242 $Y2=1.44
r29 10 12 10.3285 $w=5.03e-07 $l=3.65e-07 $layer=LI1_cond $X=0.337 $Y=0.56
+ $X2=0.337 $Y2=0.925
r30 2 22 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=2.3
r31 2 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.3
+ $Y=1.485 $X2=0.445 $Y2=1.62
r32 1 10 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.3
+ $Y=0.235 $X2=0.425 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%VPWR 1 2 3 12 14 18 20 22 37 38 41 44 48 52
c97 3 0 1.4108e-19 $X=8.425 $Y=1.485
r98 50 52 7.78613 $w=5.28e-07 $l=8e-08 $layer=LI1_cond $X=8.97 $Y=2.54 $X2=9.05
+ $Y2=2.54
r99 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r100 47 50 5.52904 $w=5.28e-07 $l=2.45e-07 $layer=LI1_cond $X=8.725 $Y=2.54
+ $X2=8.97 $Y2=2.54
r101 47 48 14.3307 $w=5.28e-07 $l=3.7e-07 $layer=LI1_cond $X=8.725 $Y=2.54
+ $X2=8.355 $Y2=2.54
r102 44 45 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r103 42 45 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r104 41 42 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r105 38 51 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=8.97 $Y2=2.72
r106 37 52 24.7914 $w=1.68e-07 $l=3.8e-07 $layer=LI1_cond $X=9.43 $Y=2.72
+ $X2=9.05 $Y2=2.72
r107 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r108 34 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=2.72
+ $X2=8.97 $Y2=2.72
r109 33 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=8.05 $Y=2.72
+ $X2=8.355 $Y2=2.72
r110 33 34 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=8.05 $Y=2.72
+ $X2=8.05 $Y2=2.72
r111 31 34 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r112 31 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r113 30 33 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=8.05 $Y2=2.72
r114 30 31 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 28 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=4.05 $Y2=2.72
r116 28 30 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=4.215 $Y=2.72
+ $X2=4.37 $Y2=2.72
r117 25 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 24 25 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r119 22 41 8.70163 $w=1.7e-07 $l=1.67e-07 $layer=LI1_cond $X=0.83 $Y=2.72
+ $X2=0.997 $Y2=2.72
r120 22 24 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=0.83 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 20 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.05 $Y=2.635
+ $X2=4.05 $Y2=2.72
r123 16 18 11.0006 $w=3.28e-07 $l=3.15e-07 $layer=LI1_cond $X=4.05 $Y=2.635
+ $X2=4.05 $Y2=2.32
r124 15 41 8.70163 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=1.165 $Y=2.72
+ $X2=0.997 $Y2=2.72
r125 14 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=4.05 $Y2=2.72
r126 14 15 177.455 $w=1.68e-07 $l=2.72e-06 $layer=LI1_cond $X=3.885 $Y=2.72
+ $X2=1.165 $Y2=2.72
r127 10 41 0.942324 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=0.997 $Y=2.635
+ $X2=0.997 $Y2=2.72
r128 10 12 11.5244 $w=3.33e-07 $l=3.35e-07 $layer=LI1_cond $X=0.997 $Y=2.635
+ $X2=0.997 $Y2=2.3
r129 3 47 600 $w=1.7e-07 $l=1.01396e-06 $layer=licon1_PDIFF $count=1 $X=8.425
+ $Y=1.485 $X2=8.725 $Y2=2.36
r130 2 18 600 $w=1.7e-07 $l=8.95321e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.05 $Y2=2.32
r131 1 12 600 $w=1.7e-07 $l=9.22862e-07 $layer=licon1_PDIFF $count=1 $X=0.77
+ $Y=1.485 $X2=1 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_406_325# 1 2 3 4 13 18 21 23 25 27 30 32
+ 33 35 37 38 39 45 49
c147 35 0 1.24749e-19 $X=7.38 $Y=0.38
r148 48 49 11.956 $w=2.5e-07 $l=2.45e-07 $layer=LI1_cond $X=3.29 $Y=1.535
+ $X2=3.535 $Y2=1.535
r149 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.1 $Y=1.53 $X2=6.1
+ $Y2=1.53
r150 42 49 5.612 $w=2.5e-07 $l=1.15e-07 $layer=LI1_cond $X=3.65 $Y=1.535
+ $X2=3.535 $Y2=1.535
r151 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.65 $Y=1.53
+ $X2=3.65 $Y2=1.53
r152 39 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.795 $Y=1.53
+ $X2=3.65 $Y2=1.53
r153 38 45 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.955 $Y=1.53
+ $X2=6.1 $Y2=1.53
r154 38 39 2.67326 $w=1.4e-07 $l=2.16e-06 $layer=MET1_cond $X=5.955 $Y=1.53
+ $X2=3.795 $Y2=1.53
r155 33 37 11.5258 $w=2.08e-07 $l=2.1e-07 $layer=LI1_cond $X=7.295 $Y=0.36
+ $X2=7.085 $Y2=0.36
r156 33 35 4.48918 $w=2.08e-07 $l=8.5e-08 $layer=LI1_cond $X=7.295 $Y=0.36
+ $X2=7.38 $Y2=0.36
r157 32 37 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=6.575 $Y=0.34
+ $X2=7.085 $Y2=0.34
r158 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.49 $Y=0.425
+ $X2=6.575 $Y2=0.34
r159 29 30 66.5455 $w=1.68e-07 $l=1.02e-06 $layer=LI1_cond $X=6.49 $Y=0.425
+ $X2=6.49 $Y2=1.445
r160 28 46 6.03523 $w=1.7e-07 $l=2.08e-07 $layer=LI1_cond $X=6.16 $Y=1.53
+ $X2=5.952 $Y2=1.53
r161 27 30 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.405 $Y=1.53
+ $X2=6.49 $Y2=1.445
r162 27 28 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=6.405 $Y=1.53
+ $X2=6.16 $Y2=1.53
r163 23 46 2.46632 $w=4.15e-07 $l=8.5e-08 $layer=LI1_cond $X=5.952 $Y=1.615
+ $X2=5.952 $Y2=1.53
r164 23 25 0.138849 $w=4.13e-07 $l=5e-09 $layer=LI1_cond $X=5.952 $Y=1.615
+ $X2=5.952 $Y2=1.62
r165 19 49 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.535 $Y=1.375
+ $X2=3.535 $Y2=1.535
r166 19 21 40.123 $w=1.68e-07 $l=6.15e-07 $layer=LI1_cond $X=3.535 $Y=1.375
+ $X2=3.535 $Y2=0.76
r167 17 48 2.99516 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=3.29 $Y=1.695
+ $X2=3.29 $Y2=1.535
r168 17 18 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.29 $Y=1.695
+ $X2=3.29 $Y2=1.895
r169 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.205 $Y=1.98
+ $X2=3.29 $Y2=1.895
r170 13 15 64.5882 $w=1.68e-07 $l=9.9e-07 $layer=LI1_cond $X=3.205 $Y=1.98
+ $X2=2.215 $Y2=1.98
r171 4 25 300 $w=1.7e-07 $l=4.12007e-07 $layer=licon1_PDIFF $count=2 $X=5.57
+ $Y=1.485 $X2=5.92 $Y2=1.62
r172 3 15 600 $w=1.7e-07 $l=4.37836e-07 $layer=licon1_PDIFF $count=1 $X=2.03
+ $Y=1.625 $X2=2.215 $Y2=1.98
r173 2 35 182 $w=1.7e-07 $l=2.53673e-07 $layer=licon1_NDIFF $count=1 $X=7.185
+ $Y=0.245 $X2=7.38 $Y2=0.38
r174 1 21 182 $w=1.7e-07 $l=6.65507e-07 $layer=licon1_NDIFF $count=1 $X=3.19
+ $Y=0.245 $X2=3.535 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_424_49# 1 2 3 4 13 18 19 20 22 23 24 26
+ 28 29 32 33 34 36 39 43 48 52 54 55 57
r187 55 56 17.995 $w=2e-07 $l=2.95e-07 $layer=LI1_cond $X=5.42 $Y=0.772
+ $X2=5.715 $Y2=0.772
r188 50 52 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.875 $Y=1.12
+ $X2=3.99 $Y2=1.12
r189 46 48 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=3.515 $Y=2.32
+ $X2=3.63 $Y2=2.32
r190 41 56 1.68994 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=5.715 $Y=0.655
+ $X2=5.715 $Y2=0.772
r191 41 43 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=5.715 $Y=0.655
+ $X2=5.715 $Y2=0.545
r192 37 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.505 $Y=2.36
+ $X2=5.42 $Y2=2.36
r193 37 39 132.439 $w=1.68e-07 $l=2.03e-06 $layer=LI1_cond $X=5.505 $Y=2.36
+ $X2=7.535 $Y2=2.36
r194 36 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.42 $Y=2.275
+ $X2=5.42 $Y2=2.36
r195 35 55 1.68994 $w=1.7e-07 $l=1.18e-07 $layer=LI1_cond $X=5.42 $Y=0.89
+ $X2=5.42 $Y2=0.772
r196 35 36 90.3583 $w=1.68e-07 $l=1.385e-06 $layer=LI1_cond $X=5.42 $Y=0.89
+ $X2=5.42 $Y2=2.275
r197 33 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.335 $Y=2.36
+ $X2=5.42 $Y2=2.36
r198 33 34 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=5.335 $Y=2.36
+ $X2=4.82 $Y2=2.36
r199 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.735 $Y=2.275
+ $X2=4.82 $Y2=2.36
r200 31 32 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=4.735 $Y=2.065
+ $X2=4.735 $Y2=2.275
r201 30 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=1.98
+ $X2=3.99 $Y2=1.98
r202 29 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=4.65 $Y=1.98
+ $X2=4.735 $Y2=2.065
r203 29 30 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=4.65 $Y=1.98
+ $X2=4.075 $Y2=1.98
r204 28 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.895
+ $X2=3.99 $Y2=1.98
r205 27 52 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.99 $Y=1.205
+ $X2=3.99 $Y2=1.12
r206 27 28 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.99 $Y=1.205
+ $X2=3.99 $Y2=1.895
r207 26 50 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.875 $Y=1.035
+ $X2=3.875 $Y2=1.12
r208 25 26 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.875 $Y=0.425
+ $X2=3.875 $Y2=1.035
r209 23 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.905 $Y=1.98
+ $X2=3.99 $Y2=1.98
r210 23 24 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=3.905 $Y=1.98
+ $X2=3.715 $Y2=1.98
r211 22 48 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.63 $Y=2.235
+ $X2=3.63 $Y2=2.32
r212 21 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.63 $Y=2.065
+ $X2=3.715 $Y2=1.98
r213 21 22 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.63 $Y=2.065
+ $X2=3.63 $Y2=2.235
r214 19 25 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.79 $Y=0.34
+ $X2=3.875 $Y2=0.425
r215 19 20 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=3.79 $Y=0.34
+ $X2=3.28 $Y2=0.34
r216 17 20 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.17 $Y=0.425
+ $X2=3.28 $Y2=0.34
r217 17 18 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=3.17 $Y=0.425
+ $X2=3.17 $Y2=0.655
r218 13 18 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.06 $Y=0.74
+ $X2=3.17 $Y2=0.655
r219 13 15 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=3.06 $Y=0.74
+ $X2=2.255 $Y2=0.74
r220 4 39 600 $w=1.7e-07 $l=8.21995e-07 $layer=licon1_PDIFF $count=1 $X=7.305
+ $Y=1.645 $X2=7.535 $Y2=2.36
r221 3 46 600 $w=1.7e-07 $l=8.70373e-07 $layer=licon1_PDIFF $count=1 $X=3.12
+ $Y=1.625 $X2=3.515 $Y2=2.32
r222 2 43 182 $w=1.7e-07 $l=3.61248e-07 $layer=licon1_NDIFF $count=1 $X=5.58
+ $Y=0.245 $X2=5.715 $Y2=0.545
r223 1 15 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.12
+ $Y=0.245 $X2=2.255 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%A_1276_297# 1 2 3 4 15 18 23 26 29 31 36
r66 34 36 4.53993 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=9.35 $Y=0.42
+ $X2=9.48 $Y2=0.42
r67 28 29 17.0922 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=9.355 $Y=1.99
+ $X2=9.03 $Y2=1.99
r68 26 31 2.50919 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=9.48 $Y=1.875
+ $X2=9.48 $Y2=1.99
r69 25 36 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=9.48 $Y=0.585
+ $X2=9.48 $Y2=0.42
r70 25 26 84.1604 $w=1.68e-07 $l=1.29e-06 $layer=LI1_cond $X=9.48 $Y=0.585
+ $X2=9.48 $Y2=1.875
r71 21 31 3.15669 $w=2.28e-07 $l=6.3e-08 $layer=LI1_cond $X=9.417 $Y=1.99
+ $X2=9.48 $Y2=1.99
r72 21 28 3.10659 $w=2.28e-07 $l=6.2e-08 $layer=LI1_cond $X=9.417 $Y=1.99
+ $X2=9.355 $Y2=1.99
r73 21 23 7.61784 $w=2.93e-07 $l=1.95e-07 $layer=LI1_cond $X=9.417 $Y=2.105
+ $X2=9.417 $Y2=2.3
r74 20 29 133.743 $w=1.68e-07 $l=2.05e-06 $layer=LI1_cond $X=6.98 $Y=2.02
+ $X2=9.03 $Y2=2.02
r75 18 20 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.915 $Y=2.02
+ $X2=6.98 $Y2=2.02
r76 13 18 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.83 $Y=1.935
+ $X2=6.915 $Y2=2.02
r77 13 15 76.6578 $w=1.68e-07 $l=1.175e-06 $layer=LI1_cond $X=6.83 $Y=1.935
+ $X2=6.83 $Y2=0.76
r78 4 28 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=9.205
+ $Y=1.485 $X2=9.355 $Y2=1.96
r79 4 23 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=9.205
+ $Y=1.485 $X2=9.355 $Y2=2.3
r80 3 20 600 $w=1.7e-07 $l=8.25227e-07 $layer=licon1_PDIFF $count=1 $X=6.38
+ $Y=1.485 $X2=6.98 $Y2=2.02
r81 2 34 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=9.215
+ $Y=0.235 $X2=9.35 $Y2=0.42
r82 1 15 182 $w=1.7e-07 $l=7.01302e-07 $layer=licon1_NDIFF $count=1 $X=6.39
+ $Y=0.245 $X2=6.83 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__XOR3_1%VGND 1 2 3 12 16 20 23 24 26 27 28 40 46 47
+ 50
c105 46 0 1.2773e-19 $X=9.43 $Y=0
c106 23 0 1.62085e-19 $X=0.81 $Y=0
r107 50 51 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r108 47 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0 $X2=8.51
+ $Y2=0
r109 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r110 44 50 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.935 $Y=0 $X2=8.71
+ $Y2=0
r111 44 46 32.2941 $w=1.68e-07 $l=4.95e-07 $layer=LI1_cond $X=8.935 $Y=0
+ $X2=9.43 $Y2=0
r112 43 51 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=4.37 $Y=0 $X2=8.51
+ $Y2=0
r113 42 43 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r114 40 50 10.5822 $w=1.7e-07 $l=2.25e-07 $layer=LI1_cond $X=8.485 $Y=0 $X2=8.71
+ $Y2=0
r115 40 42 268.465 $w=1.68e-07 $l=4.115e-06 $layer=LI1_cond $X=8.485 $Y=0
+ $X2=4.37 $Y2=0
r116 39 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r117 38 39 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r118 36 39 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=3.91 $Y2=0
r119 35 38 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=3.91
+ $Y2=0
r120 35 36 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r121 32 36 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r122 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r123 28 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r124 26 38 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=4.13 $Y=0 $X2=3.91
+ $Y2=0
r125 26 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.13 $Y=0 $X2=4.215
+ $Y2=0
r126 25 42 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.37
+ $Y2=0
r127 25 27 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.3 $Y=0 $X2=4.215
+ $Y2=0
r128 23 31 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.69
+ $Y2=0
r129 23 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.81 $Y=0 $X2=0.935
+ $Y2=0
r130 22 35 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=1.06 $Y=0 $X2=1.15
+ $Y2=0
r131 22 24 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.06 $Y=0 $X2=0.935
+ $Y2=0
r132 18 50 1.79621 $w=4.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.71 $Y=0.085
+ $X2=8.71 $Y2=0
r133 18 20 8.37255 $w=4.48e-07 $l=3.15e-07 $layer=LI1_cond $X=8.71 $Y=0.085
+ $X2=8.71 $Y2=0.4
r134 14 27 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r135 14 16 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.36
r136 10 24 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0
r137 10 12 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=0.935 $Y=0.085
+ $X2=0.935 $Y2=0.36
r138 3 20 182 $w=1.7e-07 $l=3.52987e-07 $layer=licon1_NDIFF $count=1 $X=8.435
+ $Y=0.235 $X2=8.715 $Y2=0.4
r139 2 16 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=4.05
+ $Y=0.235 $X2=4.215 $Y2=0.36
r140 1 12 182 $w=1.7e-07 $l=3.01081e-07 $layer=licon1_NDIFF $count=1 $X=0.73
+ $Y=0.235 $X2=0.975 $Y2=0.36
.ends

