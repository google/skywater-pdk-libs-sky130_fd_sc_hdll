* File: sky130_fd_sc_hdll__nor2b_4.pxi.spice
* Created: Thu Aug 27 19:16:04 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%A N_A_c_80_n N_A_M1003_g N_A_c_86_n N_A_M1002_g
+ N_A_c_81_n N_A_M1008_g N_A_c_87_n N_A_M1004_g N_A_c_82_n N_A_M1009_g
+ N_A_c_88_n N_A_M1007_g N_A_c_89_n N_A_M1013_g N_A_c_83_n N_A_M1016_g A
+ N_A_c_84_n N_A_c_85_n A PM_SKY130_FD_SC_HDLL__NOR2B_4%A
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%A_459_21# N_A_459_21#_M1012_s
+ N_A_459_21#_M1011_s N_A_459_21#_c_158_n N_A_459_21#_M1001_g
+ N_A_459_21#_c_165_n N_A_459_21#_M1000_g N_A_459_21#_c_159_n
+ N_A_459_21#_M1005_g N_A_459_21#_c_166_n N_A_459_21#_M1010_g
+ N_A_459_21#_c_160_n N_A_459_21#_M1006_g N_A_459_21#_c_167_n
+ N_A_459_21#_M1015_g N_A_459_21#_c_161_n N_A_459_21#_M1014_g
+ N_A_459_21#_c_168_n N_A_459_21#_M1017_g N_A_459_21#_c_196_p
+ N_A_459_21#_c_162_n N_A_459_21#_c_163_n N_A_459_21#_c_170_n
+ N_A_459_21#_c_179_p N_A_459_21#_c_164_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_4%A_459_21#
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%B_N N_B_N_c_263_n N_B_N_M1012_g N_B_N_c_266_n
+ N_B_N_M1011_g B_N N_B_N_c_265_n B_N PM_SKY130_FD_SC_HDLL__NOR2B_4%B_N
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%A_27_297# N_A_27_297#_M1002_s
+ N_A_27_297#_M1004_s N_A_27_297#_M1013_s N_A_27_297#_M1010_s
+ N_A_27_297#_M1017_s N_A_27_297#_c_288_n N_A_27_297#_c_289_n
+ N_A_27_297#_c_290_n N_A_27_297#_c_335_p N_A_27_297#_c_291_n
+ N_A_27_297#_c_292_n N_A_27_297#_c_308_n N_A_27_297#_c_316_n
+ N_A_27_297#_c_318_n N_A_27_297#_c_293_n N_A_27_297#_c_294_n
+ N_A_27_297#_c_295_n N_A_27_297#_c_327_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%VPWR N_VPWR_M1002_d N_VPWR_M1007_d
+ N_VPWR_M1011_d N_VPWR_c_377_n N_VPWR_c_378_n N_VPWR_c_379_n N_VPWR_c_380_n
+ VPWR N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n N_VPWR_c_384_n
+ N_VPWR_c_385_n N_VPWR_c_376_n PM_SKY130_FD_SC_HDLL__NOR2B_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%Y N_Y_M1003_s N_Y_M1009_s N_Y_M1001_s
+ N_Y_M1006_s N_Y_M1000_d N_Y_M1015_d N_Y_c_458_n N_Y_c_447_n N_Y_c_448_n
+ N_Y_c_469_n N_Y_c_449_n N_Y_c_473_n N_Y_c_450_n N_Y_c_511_n N_Y_c_451_n
+ N_Y_c_493_n N_Y_c_455_n N_Y_c_515_n N_Y_c_452_n N_Y_c_453_n N_Y_c_456_n
+ N_Y_c_457_n Y Y PM_SKY130_FD_SC_HDLL__NOR2B_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR2B_4%VGND N_VGND_M1003_d N_VGND_M1008_d
+ N_VGND_M1016_d N_VGND_M1005_d N_VGND_M1014_d N_VGND_M1012_d N_VGND_c_561_n
+ N_VGND_c_562_n N_VGND_c_563_n N_VGND_c_564_n N_VGND_c_565_n N_VGND_c_566_n
+ N_VGND_c_567_n N_VGND_c_568_n N_VGND_c_569_n N_VGND_c_570_n N_VGND_c_571_n
+ N_VGND_c_572_n N_VGND_c_573_n N_VGND_c_574_n N_VGND_c_575_n VGND
+ N_VGND_c_576_n N_VGND_c_577_n N_VGND_c_578_n
+ PM_SKY130_FD_SC_HDLL__NOR2B_4%VGND
cc_1 VNB N_A_c_80_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_81_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_82_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_c_83_n 0.0169164f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_A_c_84_n 0.0105081f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_6 VNB N_A_c_85_n 0.081832f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_A_459_21#_c_158_n 0.0164599f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_8 VNB N_A_459_21#_c_159_n 0.0163741f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_9 VNB N_A_459_21#_c_160_n 0.016732f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_10 VNB N_A_459_21#_c_161_n 0.0202448f $X=-0.19 $Y=-0.24 $X2=0.66 $Y2=1.105
cc_11 VNB N_A_459_21#_c_162_n 0.0468993f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.16
cc_12 VNB N_A_459_21#_c_163_n 0.0083181f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_13 VNB N_A_459_21#_c_164_n 0.0722105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_B_N_c_263_n 0.0254042f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_15 VNB B_N 0.0152983f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_16 VNB N_B_N_c_265_n 0.0415667f $X=-0.19 $Y=-0.24 $X2=0.985 $Y2=1.41
cc_17 VNB N_VPWR_c_376_n 0.231782f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_447_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_19 VNB N_Y_c_448_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_20 VNB N_Y_c_449_n 0.0042799f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.202
cc_21 VNB N_Y_c_450_n 8.90776e-19 $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.202
cc_22 VNB N_Y_c_451_n 0.0054182f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_23 VNB N_Y_c_452_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_Y_c_453_n 0.00375367f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_561_n 0.0102948f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.41
cc_26 VNB N_VGND_c_562_n 0.0354575f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.985
cc_27 VNB N_VGND_c_563_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.56
cc_28 VNB N_VGND_c_564_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_29 VNB N_VGND_c_565_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_30 VNB N_VGND_c_566_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_31 VNB N_VGND_c_567_n 0.00611401f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_32 VNB N_VGND_c_568_n 0.0159132f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.175
cc_33 VNB N_VGND_c_569_n 0.0336329f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.175
cc_34 VNB N_VGND_c_570_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=1.77 $Y2=1.175
cc_35 VNB N_VGND_c_571_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_572_n 0.019174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_573_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_574_n 0.0200006f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_575_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_576_n 0.023488f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_577_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_578_n 0.291384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VPB N_A_c_86_n 0.0198936f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_44 VPB N_A_c_87_n 0.0158033f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_45 VPB N_A_c_88_n 0.015524f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_46 VPB N_A_c_89_n 0.0160204f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_47 VPB N_A_c_85_n 0.0483884f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_48 VPB N_A_459_21#_c_165_n 0.0161571f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_49 VPB N_A_459_21#_c_166_n 0.0155647f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_50 VPB N_A_459_21#_c_167_n 0.015551f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.995
cc_51 VPB N_A_459_21#_c_168_n 0.0195715f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_52 VPB N_A_459_21#_c_162_n 0.0217619f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.16
cc_53 VPB N_A_459_21#_c_170_n 0.012489f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.175
cc_54 VPB N_A_459_21#_c_164_n 0.0496374f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_B_N_c_266_n 0.0244499f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_56 VPB B_N 0.00364731f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=0.995
cc_57 VPB N_B_N_c_265_n 0.0197674f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_58 VPB N_A_27_297#_c_288_n 0.0133505f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_59 VPB N_A_27_297#_c_289_n 0.0309889f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_60 VPB N_A_27_297#_c_290_n 0.00262139f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_61 VPB N_A_27_297#_c_291_n 0.00210179f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_297#_c_292_n 0.00441003f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_63 VPB N_A_27_297#_c_293_n 0.00179369f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=1.202
cc_64 VPB N_A_27_297#_c_294_n 0.0066054f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_65 VPB N_A_27_297#_c_295_n 0.00104475f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.175
cc_66 VPB N_VPWR_c_377_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_67 VPB N_VPWR_c_378_n 0.00229677f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_68 VPB N_VPWR_c_379_n 0.014431f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_69 VPB N_VPWR_c_380_n 0.0516989f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_70 VPB N_VPWR_c_381_n 0.0155059f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_382_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_72 VPB N_VPWR_c_383_n 0.0760872f $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_73 VPB N_VPWR_c_384_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0.745 $Y2=1.175
cc_74 VPB N_VPWR_c_385_n 0.00426137f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_376_n 0.0537008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_Y_c_450_n 8.36437e-19 $X=-0.19 $Y=1.305 $X2=1.77 $Y2=1.202
cc_77 VPB N_Y_c_455_n 0.00184951f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_Y_c_456_n 6.23625e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_Y_c_457_n 0.002236f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 N_A_c_83_n N_A_459_21#_c_158_n 0.0243795f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_c_89_n N_A_459_21#_c_165_n 0.00965936f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_84_n N_A_459_21#_c_164_n 8.57065e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A_c_85_n N_A_459_21#_c_164_n 0.0243795f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_84 N_A_c_84_n N_A_27_297#_c_288_n 4.10066e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_85 N_A_c_86_n N_A_27_297#_c_290_n 0.0151455f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_c_87_n N_A_27_297#_c_290_n 0.0164876f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_c_84_n N_A_27_297#_c_290_n 0.0530179f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_88 N_A_c_85_n N_A_27_297#_c_290_n 0.00953178f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_89 N_A_c_88_n N_A_27_297#_c_291_n 0.01491f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_c_89_n N_A_27_297#_c_291_n 0.0111858f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_91 N_A_c_84_n N_A_27_297#_c_291_n 0.0439319f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_c_85_n N_A_27_297#_c_291_n 0.00905881f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_c_89_n N_A_27_297#_c_292_n 0.00359583f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_c_84_n N_A_27_297#_c_292_n 3.67829e-19 $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_95 N_A_c_85_n N_A_27_297#_c_292_n 3.8543e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_96 N_A_c_88_n N_A_27_297#_c_308_n 4.84481e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_c_89_n N_A_27_297#_c_308_n 0.0132763f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_c_84_n N_A_27_297#_c_295_n 0.0132791f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_99 N_A_c_85_n N_A_27_297#_c_295_n 0.00435155f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_100 N_A_c_86_n N_VPWR_c_377_n 0.0171285f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_87_n N_VPWR_c_377_n 0.0117009f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_c_88_n N_VPWR_c_377_n 6.2189e-19 $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_c_87_n N_VPWR_c_378_n 6.52114e-19 $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_c_88_n N_VPWR_c_378_n 0.014932f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_c_89_n N_VPWR_c_378_n 0.00519421f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_c_86_n N_VPWR_c_381_n 0.00427505f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_c_87_n N_VPWR_c_382_n 0.00622633f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_c_88_n N_VPWR_c_382_n 0.00427505f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_109 N_A_c_89_n N_VPWR_c_383_n 0.00596194f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_86_n N_VPWR_c_376_n 0.00825932f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_c_87_n N_VPWR_c_376_n 0.0104011f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_c_88_n N_VPWR_c_376_n 0.00732977f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_c_89_n N_VPWR_c_376_n 0.0099828f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_c_80_n N_Y_c_458_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A_c_81_n N_Y_c_458_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A_c_82_n N_Y_c_458_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A_c_81_n N_Y_c_447_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A_c_82_n N_Y_c_447_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_119 N_A_c_84_n N_Y_c_447_n 0.0397461f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A_c_85_n N_Y_c_447_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_121 N_A_c_80_n N_Y_c_448_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_122 N_A_c_81_n N_Y_c_448_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_c_84_n N_Y_c_448_n 0.0306016f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_85_n N_Y_c_448_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_c_81_n N_Y_c_469_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_126 N_A_c_82_n N_Y_c_469_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A_c_83_n N_Y_c_449_n 0.01152f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_c_84_n N_Y_c_449_n 0.00658691f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_129 N_A_c_83_n N_Y_c_473_n 5.32212e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_130 N_A_c_84_n N_Y_c_450_n 0.0055903f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_85_n N_Y_c_450_n 0.0012283f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_c_82_n N_Y_c_452_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_133 N_A_c_84_n N_Y_c_452_n 0.0307352f $X=1.77 $Y=1.16 $X2=0 $Y2=0
cc_134 N_A_c_85_n N_Y_c_452_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_135 N_A_c_80_n N_VGND_c_562_n 0.00497314f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A_c_80_n N_VGND_c_563_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A_c_81_n N_VGND_c_563_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_c_81_n N_VGND_c_564_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_139 N_A_c_82_n N_VGND_c_564_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_c_83_n N_VGND_c_565_n 0.00268723f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A_c_82_n N_VGND_c_570_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A_c_83_n N_VGND_c_570_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A_c_80_n N_VGND_c_578_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_c_81_n N_VGND_c_578_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_145 N_A_c_82_n N_VGND_c_578_n 0.00608558f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_c_83_n N_VGND_c_578_n 0.00615622f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_147 N_A_459_21#_c_163_n N_B_N_c_263_n 0.0143944f $X=4.59 $Y=0.39 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_459_21#_c_170_n N_B_N_c_266_n 0.0173173f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_149 N_A_459_21#_c_170_n B_N 0.00576373f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_150 N_A_459_21#_c_179_p B_N 0.013979f $X=4.575 $Y=1.16 $X2=0 $Y2=0
cc_151 N_A_459_21#_c_162_n N_B_N_c_265_n 0.0215718f $X=4.38 $Y=1.16 $X2=0 $Y2=0
cc_152 N_A_459_21#_c_163_n N_B_N_c_265_n 0.00450679f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_153 N_A_459_21#_c_170_n N_B_N_c_265_n 0.0080525f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_154 N_A_459_21#_c_179_p N_B_N_c_265_n 0.00447418f $X=4.575 $Y=1.16 $X2=0
+ $Y2=0
cc_155 N_A_459_21#_c_165_n N_A_27_297#_c_292_n 0.00336534f $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_156 N_A_459_21#_c_164_n N_A_27_297#_c_292_n 3.8543e-19 $X=3.905 $Y=1.16 $X2=0
+ $Y2=0
cc_157 N_A_459_21#_c_165_n N_A_27_297#_c_308_n 0.00892871f $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_158 N_A_459_21#_c_166_n N_A_27_297#_c_308_n 5.45102e-19 $X=2.865 $Y=1.41
+ $X2=0 $Y2=0
cc_159 N_A_459_21#_c_165_n N_A_27_297#_c_316_n 0.0129846f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_160 N_A_459_21#_c_166_n N_A_27_297#_c_316_n 0.0080971f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_161 N_A_459_21#_c_167_n N_A_27_297#_c_318_n 0.010646f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A_459_21#_c_168_n N_A_27_297#_c_318_n 0.00955151f $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_163 N_A_459_21#_c_168_n N_A_27_297#_c_293_n 0.00169565f $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_164 N_A_459_21#_c_170_n N_A_27_297#_c_293_n 0.0151324f $X=4.59 $Y=1.66 $X2=0
+ $Y2=0
cc_165 N_A_459_21#_c_167_n N_A_27_297#_c_294_n 5.76911e-19 $X=3.335 $Y=1.41
+ $X2=0 $Y2=0
cc_166 N_A_459_21#_c_168_n N_A_27_297#_c_294_n 0.0127777f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_167 N_A_459_21#_c_196_p N_A_27_297#_c_294_n 0.0171609f $X=4.395 $Y=1.16 $X2=0
+ $Y2=0
cc_168 N_A_459_21#_c_162_n N_A_27_297#_c_294_n 0.00720567f $X=4.38 $Y=1.16 $X2=0
+ $Y2=0
cc_169 N_A_459_21#_c_170_n N_A_27_297#_c_294_n 0.0611923f $X=4.59 $Y=1.66 $X2=0
+ $Y2=0
cc_170 N_A_459_21#_c_165_n N_A_27_297#_c_327_n 6.08324e-19 $X=2.395 $Y=1.41
+ $X2=0 $Y2=0
cc_171 N_A_459_21#_c_166_n N_A_27_297#_c_327_n 0.00957505f $X=2.865 $Y=1.41
+ $X2=0 $Y2=0
cc_172 N_A_459_21#_c_167_n N_A_27_297#_c_327_n 0.00657656f $X=3.335 $Y=1.41
+ $X2=0 $Y2=0
cc_173 N_A_459_21#_c_168_n N_A_27_297#_c_327_n 5.59969e-19 $X=3.805 $Y=1.41
+ $X2=0 $Y2=0
cc_174 N_A_459_21#_c_170_n N_VPWR_c_380_n 0.0631564f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_175 N_A_459_21#_c_165_n N_VPWR_c_383_n 0.00429425f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_459_21#_c_166_n N_VPWR_c_383_n 0.00430873f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_177 N_A_459_21#_c_167_n N_VPWR_c_383_n 0.00430943f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A_459_21#_c_168_n N_VPWR_c_383_n 0.00429355f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_459_21#_c_170_n N_VPWR_c_383_n 0.0231967f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_180 N_A_459_21#_M1011_s N_VPWR_c_376_n 0.00225715f $X=4.455 $Y=1.485 $X2=0
+ $Y2=0
cc_181 N_A_459_21#_c_165_n N_VPWR_c_376_n 0.00609019f $X=2.395 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_459_21#_c_166_n N_VPWR_c_376_n 0.00605584f $X=2.865 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_459_21#_c_167_n N_VPWR_c_376_n 0.0060559f $X=3.335 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_459_21#_c_168_n N_VPWR_c_376_n 0.00734727f $X=3.805 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_459_21#_c_170_n N_VPWR_c_376_n 0.0136279f $X=4.59 $Y=1.66 $X2=0 $Y2=0
cc_186 N_A_459_21#_c_158_n N_Y_c_449_n 0.0117455f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_459_21#_c_158_n N_Y_c_473_n 0.00644736f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_459_21#_c_159_n N_Y_c_473_n 0.00686626f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A_459_21#_c_160_n N_Y_c_473_n 5.45498e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_190 N_A_459_21#_c_158_n N_Y_c_450_n 0.00232392f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_459_21#_c_159_n N_Y_c_450_n 0.00309297f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_192 N_A_459_21#_c_160_n N_Y_c_450_n 4.96717e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_459_21#_c_196_p N_Y_c_450_n 0.012261f $X=4.395 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A_459_21#_c_164_n N_Y_c_450_n 0.0410234f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_195 N_A_459_21#_c_159_n N_Y_c_451_n 0.0049614f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_459_21#_c_160_n N_Y_c_451_n 0.0101838f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_459_21#_c_161_n N_Y_c_451_n 0.00289584f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_198 N_A_459_21#_c_196_p N_Y_c_451_n 0.0506253f $X=4.395 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A_459_21#_c_164_n N_Y_c_451_n 0.00728851f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A_459_21#_c_159_n N_Y_c_493_n 5.24597e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_459_21#_c_160_n N_Y_c_493_n 0.00651696f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_459_21#_c_161_n N_Y_c_493_n 0.00600712f $X=3.78 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A_459_21#_c_168_n N_Y_c_455_n 0.00532752f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_459_21#_c_196_p N_Y_c_455_n 0.0137657f $X=4.395 $Y=1.16 $X2=0 $Y2=0
cc_205 N_A_459_21#_c_164_n N_Y_c_455_n 0.0045351f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A_459_21#_c_158_n N_Y_c_453_n 0.00224457f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_207 N_A_459_21#_c_159_n N_Y_c_453_n 0.00412844f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_208 N_A_459_21#_c_164_n N_Y_c_453_n 4.78733e-19 $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_209 N_A_459_21#_c_165_n N_Y_c_456_n 0.00280211f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_459_21#_c_166_n N_Y_c_456_n 0.00645246f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A_459_21#_c_166_n N_Y_c_457_n 0.00957657f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A_459_21#_c_167_n N_Y_c_457_n 0.0172194f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_213 N_A_459_21#_c_196_p N_Y_c_457_n 0.0309323f $X=4.395 $Y=1.16 $X2=0 $Y2=0
cc_214 N_A_459_21#_c_164_n N_Y_c_457_n 0.010263f $X=3.905 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_459_21#_c_158_n N_VGND_c_565_n 0.00268723f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_216 N_A_459_21#_c_159_n N_VGND_c_566_n 0.00379224f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_217 N_A_459_21#_c_160_n N_VGND_c_566_n 0.00276126f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_218 N_A_459_21#_c_161_n N_VGND_c_567_n 0.00678411f $X=3.78 $Y=0.995 $X2=0
+ $Y2=0
cc_219 N_A_459_21#_c_196_p N_VGND_c_567_n 0.0135533f $X=4.395 $Y=1.16 $X2=0
+ $Y2=0
cc_220 N_A_459_21#_c_162_n N_VGND_c_567_n 0.00431355f $X=4.38 $Y=1.16 $X2=0
+ $Y2=0
cc_221 N_A_459_21#_c_163_n N_VGND_c_567_n 0.0367019f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_222 N_A_459_21#_c_163_n N_VGND_c_569_n 0.0412732f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_223 N_A_459_21#_c_158_n N_VGND_c_572_n 0.00423334f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_224 N_A_459_21#_c_159_n N_VGND_c_572_n 0.00423261f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_225 N_A_459_21#_c_160_n N_VGND_c_574_n 0.00423334f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_226 N_A_459_21#_c_161_n N_VGND_c_574_n 0.00541359f $X=3.78 $Y=0.995 $X2=0
+ $Y2=0
cc_227 N_A_459_21#_c_163_n N_VGND_c_576_n 0.0231615f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_228 N_A_459_21#_M1012_s N_VGND_c_578_n 0.00225715f $X=4.445 $Y=0.235 $X2=0
+ $Y2=0
cc_229 N_A_459_21#_c_158_n N_VGND_c_578_n 0.00587047f $X=2.37 $Y=0.995 $X2=0
+ $Y2=0
cc_230 N_A_459_21#_c_159_n N_VGND_c_578_n 0.00609168f $X=2.84 $Y=0.995 $X2=0
+ $Y2=0
cc_231 N_A_459_21#_c_160_n N_VGND_c_578_n 0.00597024f $X=3.31 $Y=0.995 $X2=0
+ $Y2=0
cc_232 N_A_459_21#_c_161_n N_VGND_c_578_n 0.0110773f $X=3.78 $Y=0.995 $X2=0
+ $Y2=0
cc_233 N_A_459_21#_c_163_n N_VGND_c_578_n 0.0135821f $X=4.59 $Y=0.39 $X2=0 $Y2=0
cc_234 N_B_N_c_266_n N_VPWR_c_380_n 0.00913295f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_235 B_N N_VPWR_c_380_n 0.032799f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_236 N_B_N_c_265_n N_VPWR_c_380_n 0.0058213f $X=4.825 $Y=1.202 $X2=0 $Y2=0
cc_237 N_B_N_c_266_n N_VPWR_c_383_n 0.00673617f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B_N_c_266_n N_VPWR_c_376_n 0.0141776f $X=4.825 $Y=1.41 $X2=0 $Y2=0
cc_239 N_B_N_c_263_n N_VGND_c_567_n 0.00289784f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B_N_c_263_n N_VGND_c_569_n 0.00723785f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_241 B_N N_VGND_c_569_n 0.0239559f $X=5.2 $Y=1.105 $X2=0 $Y2=0
cc_242 N_B_N_c_265_n N_VGND_c_569_n 0.0063933f $X=4.825 $Y=1.202 $X2=0 $Y2=0
cc_243 N_B_N_c_263_n N_VGND_c_576_n 0.00541359f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_244 N_B_N_c_263_n N_VGND_c_578_n 0.0120732f $X=4.8 $Y=0.995 $X2=0 $Y2=0
cc_245 N_A_27_297#_c_290_n N_VPWR_M1002_d 0.00188315f $X=1.135 $Y=1.56 $X2=-0.19
+ $Y2=1.305
cc_246 N_A_27_297#_c_291_n N_VPWR_M1007_d 0.00184035f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_247 N_A_27_297#_c_289_n N_VPWR_c_377_n 0.0488071f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_248 N_A_27_297#_c_290_n N_VPWR_c_377_n 0.0212439f $X=1.135 $Y=1.56 $X2=0
+ $Y2=0
cc_249 N_A_27_297#_c_335_p N_VPWR_c_377_n 0.0385613f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_250 N_A_27_297#_c_335_p N_VPWR_c_378_n 0.0461742f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_251 N_A_27_297#_c_291_n N_VPWR_c_378_n 0.0194872f $X=1.945 $Y=1.56 $X2=0
+ $Y2=0
cc_252 N_A_27_297#_c_308_n N_VPWR_c_378_n 0.0496968f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_253 N_A_27_297#_c_289_n N_VPWR_c_381_n 0.0196165f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_254 N_A_27_297#_c_335_p N_VPWR_c_382_n 0.0118139f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_255 N_A_27_297#_c_308_n N_VPWR_c_383_n 0.0224921f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_256 N_A_27_297#_c_316_n N_VPWR_c_383_n 0.0317606f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_257 N_A_27_297#_c_318_n N_VPWR_c_383_n 0.0317606f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_258 N_A_27_297#_c_293_n N_VPWR_c_383_n 0.0260148f $X=4.025 $Y=2.295 $X2=0
+ $Y2=0
cc_259 N_A_27_297#_c_327_n N_VPWR_c_383_n 0.0220286f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_260 N_A_27_297#_M1002_s N_VPWR_c_376_n 0.00442207f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_261 N_A_27_297#_M1004_s N_VPWR_c_376_n 0.00647849f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_262 N_A_27_297#_M1013_s N_VPWR_c_376_n 0.00231261f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_263 N_A_27_297#_M1010_s N_VPWR_c_376_n 0.00231261f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_264 N_A_27_297#_M1017_s N_VPWR_c_376_n 0.00233913f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_265 N_A_27_297#_c_289_n N_VPWR_c_376_n 0.0107063f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_266 N_A_27_297#_c_335_p N_VPWR_c_376_n 0.00646998f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_267 N_A_27_297#_c_308_n N_VPWR_c_376_n 0.014078f $X=2.135 $Y=2.295 $X2=0
+ $Y2=0
cc_268 N_A_27_297#_c_316_n N_VPWR_c_376_n 0.0196262f $X=2.885 $Y=2.38 $X2=0
+ $Y2=0
cc_269 N_A_27_297#_c_318_n N_VPWR_c_376_n 0.0196262f $X=3.825 $Y=2.38 $X2=0
+ $Y2=0
cc_270 N_A_27_297#_c_293_n N_VPWR_c_376_n 0.0150121f $X=4.025 $Y=2.295 $X2=0
+ $Y2=0
cc_271 N_A_27_297#_c_327_n N_VPWR_c_376_n 0.0139179f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_272 N_A_27_297#_c_316_n N_Y_M1000_d 0.0034107f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_273 N_A_27_297#_c_318_n N_Y_M1015_d 0.0034107f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_274 N_A_27_297#_c_292_n N_Y_c_449_n 0.0132538f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_275 N_A_27_297#_c_308_n N_Y_c_511_n 0.0232292f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_276 N_A_27_297#_c_316_n N_Y_c_511_n 0.0128008f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_277 N_A_27_297#_c_327_n N_Y_c_511_n 0.0141845f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_278 N_A_27_297#_c_294_n N_Y_c_455_n 0.0142299f $X=4.04 $Y=1.66 $X2=0 $Y2=0
cc_279 N_A_27_297#_c_318_n N_Y_c_515_n 0.0128437f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_280 N_A_27_297#_c_294_n N_Y_c_515_n 0.0284474f $X=4.04 $Y=1.66 $X2=0 $Y2=0
cc_281 N_A_27_297#_c_327_n N_Y_c_515_n 0.0116296f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_282 N_A_27_297#_c_292_n N_Y_c_456_n 0.0150774f $X=2.135 $Y=1.665 $X2=0 $Y2=0
cc_283 N_A_27_297#_c_308_n N_Y_c_456_n 0.00543755f $X=2.135 $Y=2.295 $X2=0 $Y2=0
cc_284 N_A_27_297#_c_316_n N_Y_c_456_n 0.00296569f $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_285 N_A_27_297#_M1010_s N_Y_c_457_n 0.0020021f $X=2.955 $Y=1.485 $X2=0 $Y2=0
cc_286 N_A_27_297#_c_316_n N_Y_c_457_n 2.58037e-19 $X=2.885 $Y=2.38 $X2=0 $Y2=0
cc_287 N_A_27_297#_c_318_n N_Y_c_457_n 0.00438874f $X=3.825 $Y=2.38 $X2=0 $Y2=0
cc_288 N_A_27_297#_c_327_n N_Y_c_457_n 0.0197528f $X=3.1 $Y=2.02 $X2=0 $Y2=0
cc_289 N_A_27_297#_c_288_n N_VGND_c_562_n 0.0113923f $X=0.225 $Y=1.665 $X2=0
+ $Y2=0
cc_290 N_VPWR_c_376_n N_Y_M1000_d 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_291 N_VPWR_c_376_n N_Y_M1015_d 0.00232895f $X=5.29 $Y=2.72 $X2=0 $Y2=0
cc_292 N_Y_c_447_n N_VGND_M1008_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_293 N_Y_c_449_n N_VGND_M1016_d 0.00162089f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_294 N_Y_c_451_n N_VGND_M1005_d 0.00251047f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_295 N_Y_c_448_n N_VGND_c_562_n 0.00835667f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_296 N_Y_c_458_n N_VGND_c_563_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_297 N_Y_c_447_n N_VGND_c_563_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_298 N_Y_c_458_n N_VGND_c_564_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_299 N_Y_c_447_n N_VGND_c_564_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_300 N_Y_c_449_n N_VGND_c_565_n 0.0122559f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_301 N_Y_c_473_n N_VGND_c_566_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_302 N_Y_c_451_n N_VGND_c_566_n 0.0127273f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_303 N_Y_c_451_n N_VGND_c_567_n 0.0116109f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_304 N_Y_c_493_n N_VGND_c_567_n 0.0287371f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_305 N_Y_c_447_n N_VGND_c_570_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_306 N_Y_c_469_n N_VGND_c_570_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_307 N_Y_c_449_n N_VGND_c_570_n 0.00254521f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_308 N_Y_c_449_n N_VGND_c_572_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_309 N_Y_c_473_n N_VGND_c_572_n 0.0224037f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_310 N_Y_c_451_n N_VGND_c_572_n 0.00159127f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_311 N_Y_c_453_n N_VGND_c_572_n 0.00118043f $X=2.645 $Y=0.815 $X2=0 $Y2=0
cc_312 N_Y_c_451_n N_VGND_c_574_n 0.00198695f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_313 N_Y_c_493_n N_VGND_c_574_n 0.0223596f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_314 N_Y_M1003_s N_VGND_c_578_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_315 N_Y_M1009_s N_VGND_c_578_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_316 N_Y_M1001_s N_VGND_c_578_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_317 N_Y_M1006_s N_VGND_c_578_n 0.0025535f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_318 N_Y_c_458_n N_VGND_c_578_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_319 N_Y_c_447_n N_VGND_c_578_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_320 N_Y_c_469_n N_VGND_c_578_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_321 N_Y_c_449_n N_VGND_c_578_n 0.0094839f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_322 N_Y_c_473_n N_VGND_c_578_n 0.0141415f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_323 N_Y_c_451_n N_VGND_c_578_n 0.00800459f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_324 N_Y_c_493_n N_VGND_c_578_n 0.0141302f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_325 N_Y_c_453_n N_VGND_c_578_n 0.001841f $X=2.645 $Y=0.815 $X2=0 $Y2=0
