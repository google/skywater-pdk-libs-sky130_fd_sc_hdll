* File: sky130_fd_sc_hdll__xor2_4.pxi.spice
* Created: Thu Aug 27 19:29:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__XOR2_4%A N_A_c_158_n N_A_M1003_g N_A_c_169_n N_A_M1005_g
+ N_A_c_159_n N_A_M1014_g N_A_c_170_n N_A_M1012_g N_A_c_160_n N_A_M1030_g
+ N_A_c_171_n N_A_M1020_g N_A_c_172_n N_A_M1027_g N_A_c_161_n N_A_M1031_g
+ N_A_c_162_n N_A_M1004_g N_A_c_173_n N_A_M1001_g N_A_c_163_n N_A_M1008_g
+ N_A_c_174_n N_A_M1007_g N_A_c_164_n N_A_M1018_g N_A_c_175_n N_A_M1013_g
+ N_A_c_176_n N_A_M1015_g N_A_c_165_n N_A_M1032_g N_A_c_177_n N_A_c_178_n
+ N_A_c_184_p N_A_c_203_p N_A_c_179_n N_A_c_235_p N_A_c_166_n A N_A_c_167_n
+ N_A_c_168_n PM_SKY130_FD_SC_HDLL__XOR2_4%A
x_PM_SKY130_FD_SC_HDLL__XOR2_4%B N_B_c_386_n N_B_M1011_g N_B_c_398_n N_B_M1000_g
+ N_B_c_387_n N_B_M1025_g N_B_c_399_n N_B_M1006_g N_B_c_388_n N_B_M1026_g
+ N_B_c_400_n N_B_M1023_g N_B_c_389_n N_B_M1039_g N_B_c_401_n N_B_M1033_g
+ N_B_c_390_n N_B_c_391_n N_B_c_392_n N_B_M1002_g N_B_c_404_n N_B_M1009_g
+ N_B_c_393_n N_B_M1017_g N_B_c_405_n N_B_M1021_g N_B_c_394_n N_B_M1022_g
+ N_B_c_406_n N_B_M1028_g N_B_c_407_n N_B_M1035_g N_B_c_395_n N_B_M1037_g B
+ N_B_c_396_n N_B_c_397_n B PM_SKY130_FD_SC_HDLL__XOR2_4%B
x_PM_SKY130_FD_SC_HDLL__XOR2_4%A_112_47# N_A_112_47#_M1003_d N_A_112_47#_M1030_d
+ N_A_112_47#_M1011_s N_A_112_47#_M1026_s N_A_112_47#_M1000_s
+ N_A_112_47#_M1023_s N_A_112_47#_c_538_n N_A_112_47#_M1010_g
+ N_A_112_47#_c_555_n N_A_112_47#_M1016_g N_A_112_47#_c_539_n
+ N_A_112_47#_M1019_g N_A_112_47#_c_556_n N_A_112_47#_M1024_g
+ N_A_112_47#_c_540_n N_A_112_47#_M1036_g N_A_112_47#_c_557_n
+ N_A_112_47#_M1029_g N_A_112_47#_c_558_n N_A_112_47#_M1034_g
+ N_A_112_47#_c_541_n N_A_112_47#_M1038_g N_A_112_47#_c_542_n
+ N_A_112_47#_c_543_n N_A_112_47#_c_544_n N_A_112_47#_c_574_n
+ N_A_112_47#_c_545_n N_A_112_47#_c_581_n N_A_112_47#_c_546_n
+ N_A_112_47#_c_585_n N_A_112_47#_c_586_n N_A_112_47#_c_547_n
+ N_A_112_47#_c_640_n N_A_112_47#_c_548_n N_A_112_47#_c_549_n
+ N_A_112_47#_c_550_n N_A_112_47#_c_561_n N_A_112_47#_c_551_n
+ N_A_112_47#_c_552_n N_A_112_47#_c_553_n N_A_112_47#_c_562_n
+ N_A_112_47#_c_610_n N_A_112_47#_c_650_n N_A_112_47#_c_611_n
+ N_A_112_47#_c_563_n N_A_112_47#_c_564_n N_A_112_47#_c_565_n
+ N_A_112_47#_c_566_n N_A_112_47#_c_554_n PM_SKY130_FD_SC_HDLL__XOR2_4%A_112_47#
x_PM_SKY130_FD_SC_HDLL__XOR2_4%A_27_297# N_A_27_297#_M1005_s N_A_27_297#_M1012_s
+ N_A_27_297#_M1027_s N_A_27_297#_M1006_d N_A_27_297#_M1033_d
+ N_A_27_297#_c_822_n N_A_27_297#_c_824_n N_A_27_297#_c_839_n
+ N_A_27_297#_c_827_n N_A_27_297#_c_861_p N_A_27_297#_c_817_n
+ N_A_27_297#_c_826_n N_A_27_297#_c_818_n N_A_27_297#_c_850_n
+ N_A_27_297#_c_851_n PM_SKY130_FD_SC_HDLL__XOR2_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_4%VPWR N_VPWR_M1005_d N_VPWR_M1020_d N_VPWR_M1009_d
+ N_VPWR_M1028_d N_VPWR_M1001_d N_VPWR_M1013_d N_VPWR_c_882_n N_VPWR_c_883_n
+ N_VPWR_c_884_n N_VPWR_c_885_n N_VPWR_c_886_n N_VPWR_c_887_n N_VPWR_c_888_n
+ N_VPWR_c_889_n N_VPWR_c_890_n N_VPWR_c_891_n N_VPWR_c_892_n N_VPWR_c_893_n
+ N_VPWR_c_894_n N_VPWR_c_895_n N_VPWR_c_896_n VPWR N_VPWR_c_897_n
+ N_VPWR_c_881_n N_VPWR_c_899_n N_VPWR_c_900_n PM_SKY130_FD_SC_HDLL__XOR2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_297# N_A_886_297#_M1009_s
+ N_A_886_297#_M1021_s N_A_886_297#_M1035_s N_A_886_297#_M1007_s
+ N_A_886_297#_M1015_s N_A_886_297#_M1016_d N_A_886_297#_M1029_d
+ N_A_886_297#_c_1044_n N_A_886_297#_c_1045_n N_A_886_297#_c_1046_n
+ N_A_886_297#_c_1037_n N_A_886_297#_c_1056_n N_A_886_297#_c_1038_n
+ N_A_886_297#_c_1082_n N_A_886_297#_c_1039_n N_A_886_297#_c_1120_n
+ N_A_886_297#_c_1141_p N_A_886_297#_c_1084_n N_A_886_297#_c_1145_p
+ N_A_886_297#_c_1040_n N_A_886_297#_c_1061_n N_A_886_297#_c_1062_n
+ N_A_886_297#_c_1130_n N_A_886_297#_c_1132_n
+ PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_297#
x_PM_SKY130_FD_SC_HDLL__XOR2_4%X N_X_M1002_d N_X_M1022_d N_X_M1010_d N_X_M1036_d
+ N_X_M1016_s N_X_M1024_s N_X_M1034_s N_X_c_1157_n N_X_c_1158_n N_X_c_1159_n
+ N_X_c_1198_n N_X_c_1147_n N_X_c_1160_n N_X_c_1209_n N_X_c_1148_n N_X_c_1149_n
+ N_X_c_1150_n N_X_c_1151_n N_X_c_1162_n N_X_c_1152_n N_X_c_1163_n X
+ N_X_c_1176_n N_X_c_1153_n N_X_c_1154_n N_X_c_1155_n N_X_c_1156_n
+ PM_SKY130_FD_SC_HDLL__XOR2_4%X
x_PM_SKY130_FD_SC_HDLL__XOR2_4%VGND N_VGND_M1003_s N_VGND_M1014_s N_VGND_M1031_s
+ N_VGND_M1025_d N_VGND_M1039_d N_VGND_M1004_s N_VGND_M1018_s N_VGND_M1010_s
+ N_VGND_M1019_s N_VGND_M1038_s N_VGND_c_1306_n N_VGND_c_1307_n N_VGND_c_1308_n
+ N_VGND_c_1309_n N_VGND_c_1310_n N_VGND_c_1311_n N_VGND_c_1312_n
+ N_VGND_c_1313_n N_VGND_c_1314_n N_VGND_c_1315_n N_VGND_c_1316_n
+ N_VGND_c_1317_n N_VGND_c_1318_n N_VGND_c_1319_n N_VGND_c_1320_n
+ N_VGND_c_1321_n N_VGND_c_1322_n N_VGND_c_1323_n N_VGND_c_1324_n
+ N_VGND_c_1325_n N_VGND_c_1326_n N_VGND_c_1327_n N_VGND_c_1328_n
+ N_VGND_c_1329_n N_VGND_c_1330_n N_VGND_c_1331_n VGND N_VGND_c_1332_n
+ N_VGND_c_1333_n N_VGND_c_1334_n N_VGND_c_1335_n
+ PM_SKY130_FD_SC_HDLL__XOR2_4%VGND
x_PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_47# N_A_886_47#_M1002_s N_A_886_47#_M1017_s
+ N_A_886_47#_M1037_s N_A_886_47#_M1008_d N_A_886_47#_M1032_d
+ N_A_886_47#_c_1497_n N_A_886_47#_c_1503_n N_A_886_47#_c_1498_n
+ N_A_886_47#_c_1499_n N_A_886_47#_c_1513_n N_A_886_47#_c_1500_n
+ N_A_886_47#_c_1501_n N_A_886_47#_c_1502_n
+ PM_SKY130_FD_SC_HDLL__XOR2_4%A_886_47#
cc_1 VNB N_A_c_158_n 0.0197012f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_c_159_n 0.016761f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_A_c_160_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.425 $Y2=0.995
cc_4 VNB N_A_c_161_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=0.995
cc_5 VNB N_A_c_162_n 0.0162998f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=0.995
cc_6 VNB N_A_c_163_n 0.0165967f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=0.995
cc_7 VNB N_A_c_164_n 0.0170349f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.995
cc_8 VNB N_A_c_165_n 0.0220151f $X=-0.19 $Y=-0.24 $X2=8.105 $Y2=0.995
cc_9 VNB N_A_c_166_n 0.00467216f $X=-0.19 $Y=-0.24 $X2=2.88 $Y2=1.175
cc_10 VNB N_A_c_167_n 0.0767096f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.202
cc_11 VNB N_A_c_168_n 0.0803739f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.202
cc_12 VNB N_B_c_386_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_13 VNB N_B_c_387_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_14 VNB N_B_c_388_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.425 $Y2=0.995
cc_15 VNB N_B_c_389_n 0.0221076f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.41
cc_16 VNB N_B_c_390_n 0.0477207f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=0.995
cc_17 VNB N_B_c_391_n 0.0674992f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=0.56
cc_18 VNB N_B_c_392_n 0.0219752f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=0.56
cc_19 VNB N_B_c_393_n 0.0167438f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=0.56
cc_20 VNB N_B_c_394_n 0.0170767f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.56
cc_21 VNB N_B_c_395_n 0.0167925f $X=-0.19 $Y=-0.24 $X2=8.105 $Y2=0.56
cc_22 VNB N_B_c_396_n 0.00199342f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.202
cc_23 VNB N_B_c_397_n 0.0688016f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_24 VNB N_A_112_47#_c_538_n 0.0216918f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.41
cc_25 VNB N_A_112_47#_c_539_n 0.016763f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=0.995
cc_26 VNB N_A_112_47#_c_540_n 0.0171977f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=0.995
cc_27 VNB N_A_112_47#_c_541_n 0.0200668f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.41
cc_28 VNB N_A_112_47#_c_542_n 0.0190377f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.985
cc_29 VNB N_A_112_47#_c_543_n 0.00203902f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.985
cc_30 VNB N_A_112_47#_c_544_n 0.00773467f $X=-0.19 $Y=-0.24 $X2=8.105 $Y2=0.995
cc_31 VNB N_A_112_47#_c_545_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=6.595 $Y2=1.53
cc_32 VNB N_A_112_47#_c_546_n 0.00255474f $X=-0.19 $Y=-0.24 $X2=7.94 $Y2=1.16
cc_33 VNB N_A_112_47#_c_547_n 0.00525562f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_34 VNB N_A_112_47#_c_548_n 8.09078e-19 $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_35 VNB N_A_112_47#_c_549_n 0.00398328f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_36 VNB N_A_112_47#_c_550_n 0.0141968f $X=-0.19 $Y=-0.24 $X2=6.77 $Y2=1.202
cc_37 VNB N_A_112_47#_c_551_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.202
cc_38 VNB N_A_112_47#_c_552_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=7.94 $Y2=1.202
cc_39 VNB N_A_112_47#_c_553_n 0.0023781f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.202
cc_40 VNB N_A_112_47#_c_554_n 0.0827384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VPWR_c_881_n 0.459507f $X=-0.19 $Y=-0.24 $X2=6.77 $Y2=1.202
cc_42 VNB N_X_c_1147_n 0.00247032f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.985
cc_43 VNB N_X_c_1148_n 0.00963283f $X=-0.19 $Y=-0.24 $X2=8.105 $Y2=0.995
cc_44 VNB N_X_c_1149_n 0.0221179f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.275
cc_45 VNB N_X_c_1150_n 0.003375f $X=-0.19 $Y=-0.24 $X2=3.1 $Y2=1.53
cc_46 VNB N_X_c_1151_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=1.275
cc_47 VNB N_X_c_1152_n 0.00334519f $X=-0.19 $Y=-0.24 $X2=7.94 $Y2=1.175
cc_48 VNB N_X_c_1153_n 0.00228596f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_49 VNB N_X_c_1154_n 0.0126712f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_50 VNB N_X_c_1155_n 0.00621555f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_51 VNB N_X_c_1156_n 0.00311636f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.202
cc_52 VNB N_VGND_c_1306_n 0.0101714f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=0.995
cc_53 VNB N_VGND_c_1307_n 0.0182438f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=0.56
cc_54 VNB N_VGND_c_1308_n 0.019187f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.985
cc_55 VNB N_VGND_c_1309_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=0.56
cc_56 VNB N_VGND_c_1310_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.985
cc_57 VNB N_VGND_c_1311_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.985
cc_58 VNB N_VGND_c_1312_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.275
cc_59 VNB N_VGND_c_1313_n 0.0147986f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=1.275
cc_60 VNB N_VGND_c_1314_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=7.94 $Y2=1.16
cc_61 VNB N_VGND_c_1315_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=6.705 $Y2=1.175
cc_62 VNB N_VGND_c_1316_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_1317_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_64 VNB N_VGND_c_1318_n 0.0122507f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=1.202
cc_65 VNB N_VGND_c_1319_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=1.425 $Y2=1.202
cc_66 VNB N_VGND_c_1320_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_67 VNB N_VGND_c_1321_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.765 $Y2=1.16
cc_68 VNB N_VGND_c_1322_n 0.0200006f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=1.202
cc_69 VNB N_VGND_c_1323_n 0.00519339f $X=-0.19 $Y=-0.24 $X2=6.645 $Y2=1.202
cc_70 VNB N_VGND_c_1324_n 0.0604226f $X=-0.19 $Y=-0.24 $X2=6.77 $Y2=1.202
cc_71 VNB N_VGND_c_1325_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=7.115 $Y2=1.202
cc_72 VNB N_VGND_c_1326_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=7.585 $Y2=1.202
cc_73 VNB N_VGND_c_1327_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.202
cc_74 VNB N_VGND_c_1328_n 0.021605f $X=-0.19 $Y=-0.24 $X2=8.08 $Y2=1.202
cc_75 VNB N_VGND_c_1329_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=8.105 $Y2=1.202
cc_76 VNB N_VGND_c_1330_n 0.0191907f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1331_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.175
cc_78 VNB N_VGND_c_1332_n 0.019283f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1333_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1334_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1335_n 0.514676f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_A_886_47#_c_1497_n 0.00270572f $X=-0.19 $Y=-0.24 $X2=1.45 $Y2=1.41
cc_83 VNB N_A_886_47#_c_1498_n 0.00194195f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=0.56
cc_84 VNB N_A_886_47#_c_1499_n 0.00109126f $X=-0.19 $Y=-0.24 $X2=1.945 $Y2=0.56
cc_85 VNB N_A_886_47#_c_1500_n 0.00414013f $X=-0.19 $Y=-0.24 $X2=6.67 $Y2=1.985
cc_86 VNB N_A_886_47#_c_1501_n 0.00548011f $X=-0.19 $Y=-0.24 $X2=7.14 $Y2=1.41
cc_87 VNB N_A_886_47#_c_1502_n 0.00109312f $X=-0.19 $Y=-0.24 $X2=7.61 $Y2=1.41
cc_88 VPB N_A_c_169_n 0.0192002f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_89 VPB N_A_c_170_n 0.0158727f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_90 VPB N_A_c_171_n 0.0158196f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.41
cc_91 VPB N_A_c_172_n 0.0159269f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.41
cc_92 VPB N_A_c_173_n 0.0158458f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_93 VPB N_A_c_174_n 0.0160496f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.41
cc_94 VPB N_A_c_175_n 0.0159677f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.41
cc_95 VPB N_A_c_176_n 0.0191888f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.41
cc_96 VPB N_A_c_177_n 0.00115215f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.445
cc_97 VPB N_A_c_178_n 0.0277321f $X=-0.19 $Y=1.305 $X2=6.595 $Y2=1.53
cc_98 VPB N_A_c_179_n 0.00123098f $X=-0.19 $Y=1.305 $X2=6.705 $Y2=1.445
cc_99 VPB N_A_c_167_n 0.0455275f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.202
cc_100 VPB N_A_c_168_n 0.0487525f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.202
cc_101 VPB N_B_c_398_n 0.0157381f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_102 VPB N_B_c_399_n 0.0157419f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_103 VPB N_B_c_400_n 0.0158635f $X=-0.19 $Y=1.305 $X2=1.45 $Y2=1.41
cc_104 VPB N_B_c_401_n 0.0200905f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=0.995
cc_105 VPB N_B_c_390_n 0.0204896f $X=-0.19 $Y=1.305 $X2=6.645 $Y2=0.995
cc_106 VPB N_B_c_391_n 0.0481341f $X=-0.19 $Y=1.305 $X2=6.645 $Y2=0.56
cc_107 VPB N_B_c_404_n 0.0201091f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.985
cc_108 VPB N_B_c_405_n 0.0158911f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.985
cc_109 VPB N_B_c_406_n 0.0158911f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.985
cc_110 VPB N_B_c_407_n 0.0159807f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.985
cc_111 VPB N_B_c_397_n 0.0471806f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_112 VPB N_A_112_47#_c_555_n 0.0192809f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=0.995
cc_113 VPB N_A_112_47#_c_556_n 0.0158911f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_114 VPB N_A_112_47#_c_557_n 0.015872f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.41
cc_115 VPB N_A_112_47#_c_558_n 0.0191956f $X=-0.19 $Y=1.305 $X2=7.585 $Y2=0.995
cc_116 VPB N_A_112_47#_c_542_n 0.00689005f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.985
cc_117 VPB N_A_112_47#_c_548_n 0.00610017f $X=-0.19 $Y=1.305 $X2=1.765 $Y2=1.16
cc_118 VPB N_A_112_47#_c_561_n 0.00785262f $X=-0.19 $Y=1.305 $X2=7.585 $Y2=1.202
cc_119 VPB N_A_112_47#_c_562_n 0.0101831f $X=-0.19 $Y=1.305 $X2=8.105 $Y2=1.202
cc_120 VPB N_A_112_47#_c_563_n 0.00375306f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_112_47#_c_564_n 0.00168325f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_112_47#_c_565_n 0.00685629f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_112_47#_c_566_n 0.00173014f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_112_47#_c_554_n 0.046491f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_27_297#_c_817_n 0.00148837f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_126 VPB N_A_27_297#_c_818_n 0.0280239f $X=-0.19 $Y=1.305 $X2=7.14 $Y2=1.985
cc_127 VPB N_VPWR_c_882_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.945 $Y2=0.56
cc_128 VPB N_VPWR_c_883_n 0.0178757f $X=-0.19 $Y=1.305 $X2=6.645 $Y2=0.995
cc_129 VPB N_VPWR_c_884_n 0.00516582f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.985
cc_130 VPB N_VPWR_c_885_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.115 $Y2=0.56
cc_131 VPB N_VPWR_c_886_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.585 $Y2=0.995
cc_132 VPB N_VPWR_c_887_n 0.00516582f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.985
cc_133 VPB N_VPWR_c_888_n 0.00516582f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.985
cc_134 VPB N_VPWR_c_889_n 0.0736651f $X=-0.19 $Y=1.305 $X2=8.105 $Y2=0.56
cc_135 VPB N_VPWR_c_890_n 0.00478085f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.275
cc_136 VPB N_VPWR_c_891_n 0.0178757f $X=-0.19 $Y=1.305 $X2=6.595 $Y2=1.53
cc_137 VPB N_VPWR_c_892_n 0.00478085f $X=-0.19 $Y=1.305 $X2=3.1 $Y2=1.53
cc_138 VPB N_VPWR_c_893_n 0.0178757f $X=-0.19 $Y=1.305 $X2=6.705 $Y2=1.445
cc_139 VPB N_VPWR_c_894_n 0.00478085f $X=-0.19 $Y=1.305 $X2=6.815 $Y2=1.175
cc_140 VPB N_VPWR_c_895_n 0.0178757f $X=-0.19 $Y=1.305 $X2=7.94 $Y2=1.16
cc_141 VPB N_VPWR_c_896_n 0.00478085f $X=-0.19 $Y=1.305 $X2=7.94 $Y2=1.16
cc_142 VPB N_VPWR_c_897_n 0.0740728f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.202
cc_143 VPB N_VPWR_c_881_n 0.0589954f $X=-0.19 $Y=1.305 $X2=6.77 $Y2=1.202
cc_144 VPB N_VPWR_c_899_n 0.0228668f $X=-0.19 $Y=1.305 $X2=7.585 $Y2=1.202
cc_145 VPB N_VPWR_c_900_n 0.00478085f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.202
cc_146 VPB N_A_886_297#_c_1037_n 0.00214773f $X=-0.19 $Y=1.305 $X2=7.14
+ $Y2=1.985
cc_147 VPB N_A_886_297#_c_1038_n 0.00192772f $X=-0.19 $Y=1.305 $X2=7.61
+ $Y2=1.985
cc_148 VPB N_A_886_297#_c_1039_n 0.012098f $X=-0.19 $Y=1.305 $X2=8.08 $Y2=1.985
cc_149 VPB N_A_886_297#_c_1040_n 0.00199604f $X=-0.19 $Y=1.305 $X2=7.94 $Y2=1.16
cc_150 VPB N_X_c_1157_n 0.00429063f $X=-0.19 $Y=1.305 $X2=6.645 $Y2=0.56
cc_151 VPB N_X_c_1158_n 0.00510623f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.41
cc_152 VPB N_X_c_1159_n 0.00195599f $X=-0.19 $Y=1.305 $X2=6.67 $Y2=1.985
cc_153 VPB N_X_c_1160_n 0.00234077f $X=-0.19 $Y=1.305 $X2=7.61 $Y2=1.41
cc_154 VPB N_X_c_1149_n 0.00752017f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.275
cc_155 VPB N_X_c_1162_n 0.0014926f $X=-0.19 $Y=1.305 $X2=6.815 $Y2=1.175
cc_156 VPB N_X_c_1163_n 0.00873134f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB X 0.0352804f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=1.175
cc_158 N_A_c_161_n N_B_c_386_n 0.024433f $X=1.945 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_159 N_A_c_172_n N_B_c_398_n 0.0221449f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_160 N_A_c_184_p N_B_c_398_n 2.09341e-19 $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_161 N_A_c_177_n N_B_c_399_n 6.79361e-19 $X=2.99 $Y=1.445 $X2=0 $Y2=0
cc_162 N_A_c_184_p N_B_c_399_n 0.00510949f $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_163 N_A_c_177_n N_B_c_400_n 7.75865e-19 $X=2.99 $Y=1.445 $X2=0 $Y2=0
cc_164 N_A_c_178_n N_B_c_400_n 0.0122738f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_165 N_A_c_178_n N_B_c_401_n 0.0194073f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_c_178_n N_B_c_390_n 0.0192768f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_167 N_A_c_177_n N_B_c_391_n 0.0132286f $X=2.99 $Y=1.445 $X2=0 $Y2=0
cc_168 N_A_c_178_n N_B_c_391_n 0.0122503f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_169 N_A_c_166_n N_B_c_391_n 0.0374341f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_170 N_A_c_167_n N_B_c_391_n 0.024433f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_171 N_A_c_178_n N_B_c_404_n 0.0139099f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_172 N_A_c_178_n N_B_c_405_n 0.01191f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_173 N_A_c_178_n N_B_c_406_n 0.0118984f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_174 N_A_c_173_n N_B_c_407_n 0.0227665f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_178_n N_B_c_407_n 0.011855f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_176 N_A_c_179_n N_B_c_407_n 2.06453e-19 $X=6.705 $Y=1.445 $X2=0 $Y2=0
cc_177 N_A_c_162_n N_B_c_395_n 0.0174382f $X=6.645 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_178_n N_B_c_396_n 0.196476f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_179 N_A_c_203_p N_B_c_396_n 0.0110392f $X=6.705 $Y=1.275 $X2=0 $Y2=0
cc_180 N_A_c_166_n N_B_c_396_n 0.0167609f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_181 N_A_c_168_n N_B_c_396_n 0.00135129f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_182 N_A_c_178_n N_B_c_397_n 0.0231495f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_183 N_A_c_203_p N_B_c_397_n 4.0849e-19 $X=6.705 $Y=1.275 $X2=0 $Y2=0
cc_184 N_A_c_179_n N_B_c_397_n 8.78417e-19 $X=6.705 $Y=1.445 $X2=0 $Y2=0
cc_185 N_A_c_168_n N_B_c_397_n 0.0174382f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_186 N_A_c_178_n N_A_112_47#_M1023_s 0.00187091f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_187 N_A_c_158_n N_A_112_47#_c_542_n 0.0170306f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_188 N_A_c_169_n N_A_112_47#_c_542_n 0.00119489f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_166_n N_A_112_47#_c_542_n 0.015823f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_190 N_A_c_158_n N_A_112_47#_c_543_n 0.0101572f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_191 N_A_c_166_n N_A_112_47#_c_543_n 0.00717314f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_192 N_A_c_158_n N_A_112_47#_c_574_n 0.0107127f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_193 N_A_c_159_n N_A_112_47#_c_574_n 0.00686626f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_194 N_A_c_160_n N_A_112_47#_c_574_n 5.45498e-19 $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_195 N_A_c_159_n N_A_112_47#_c_545_n 0.00901745f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_196 N_A_c_160_n N_A_112_47#_c_545_n 0.00901745f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_197 N_A_c_166_n N_A_112_47#_c_545_n 0.0397461f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_198 N_A_c_167_n N_A_112_47#_c_545_n 0.00345541f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_199 N_A_c_159_n N_A_112_47#_c_581_n 5.24597e-19 $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_200 N_A_c_160_n N_A_112_47#_c_581_n 0.00651696f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_201 N_A_c_161_n N_A_112_47#_c_546_n 0.0106151f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A_c_166_n N_A_112_47#_c_546_n 0.0399644f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_203 N_A_c_161_n N_A_112_47#_c_585_n 5.32212e-19 $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A_c_178_n N_A_112_47#_c_586_n 0.0164917f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_205 N_A_c_184_p N_A_112_47#_c_586_n 0.011566f $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_206 N_A_c_166_n N_A_112_47#_c_586_n 0.00144764f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_207 N_A_c_178_n N_A_112_47#_c_547_n 0.00434751f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_208 N_A_c_166_n N_A_112_47#_c_547_n 0.0227112f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_209 N_A_c_176_n N_A_112_47#_c_548_n 0.00108129f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_168_n N_A_112_47#_c_548_n 0.00512058f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_211 N_A_c_235_p N_A_112_47#_c_549_n 0.0145272f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_c_168_n N_A_112_47#_c_549_n 0.00571708f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_213 N_A_c_158_n N_A_112_47#_c_551_n 0.00161382f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_159_n N_A_112_47#_c_551_n 0.00116636f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A_c_166_n N_A_112_47#_c_551_n 0.0306016f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_216 N_A_c_167_n N_A_112_47#_c_551_n 0.00358305f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_217 N_A_c_160_n N_A_112_47#_c_552_n 0.00119564f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_c_166_n N_A_112_47#_c_552_n 0.0307352f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_219 N_A_c_167_n N_A_112_47#_c_552_n 0.00486271f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_220 N_A_c_166_n N_A_112_47#_c_553_n 0.02961f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_221 N_A_c_169_n N_A_112_47#_c_562_n 0.0133681f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_170_n N_A_112_47#_c_562_n 0.01191f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_171_n N_A_112_47#_c_562_n 0.01191f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_172_n N_A_112_47#_c_562_n 0.011867f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_184_p N_A_112_47#_c_562_n 0.0098507f $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_226 N_A_c_166_n N_A_112_47#_c_562_n 0.157359f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_227 N_A_c_167_n N_A_112_47#_c_562_n 0.0231985f $X=1.92 $Y=1.202 $X2=0 $Y2=0
cc_228 N_A_c_166_n N_A_112_47#_c_610_n 8.215e-19 $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_229 N_A_c_178_n N_A_112_47#_c_611_n 0.012249f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_230 N_A_c_174_n N_A_112_47#_c_563_n 0.00496772f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_c_175_n N_A_112_47#_c_563_n 0.00496772f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_c_176_n N_A_112_47#_c_563_n 0.00125135f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_233 N_A_c_178_n N_A_112_47#_c_563_n 0.163768f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_234 N_A_c_184_p N_A_112_47#_c_563_n 0.0115163f $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_235 N_A_c_235_p N_A_112_47#_c_563_n 0.0142049f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_236 N_A_c_166_n N_A_112_47#_c_563_n 0.00737552f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_237 N_A_c_168_n N_A_112_47#_c_563_n 0.0110527f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_238 N_A_c_172_n N_A_112_47#_c_564_n 9.96005e-19 $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_177_n N_A_112_47#_c_564_n 8.95935e-19 $X=2.99 $Y=1.445 $X2=0 $Y2=0
cc_240 N_A_c_166_n N_A_112_47#_c_564_n 0.00776789f $X=2.88 $Y=1.175 $X2=0 $Y2=0
cc_241 N_A_c_176_n N_A_112_47#_c_565_n 0.00160344f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_c_175_n N_A_112_47#_c_566_n 7.23294e-19 $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_c_176_n N_A_112_47#_c_566_n 0.0124046f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_c_235_p N_A_112_47#_c_566_n 0.00660315f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_245 N_A_c_168_n N_A_112_47#_c_566_n 3.57927e-19 $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_246 N_A_c_178_n N_A_27_297#_M1006_d 8.73801e-19 $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_247 N_A_c_184_p N_A_27_297#_M1006_d 0.00102446f $X=3.1 $Y=1.53 $X2=0 $Y2=0
cc_248 N_A_c_178_n N_A_27_297#_M1033_d 0.00295094f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_249 N_A_c_169_n N_A_27_297#_c_822_n 0.0132707f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_250 N_A_c_170_n N_A_27_297#_c_822_n 0.0133261f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_c_171_n N_A_27_297#_c_824_n 0.0133261f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_c_172_n N_A_27_297#_c_824_n 0.0133261f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_178_n N_A_27_297#_c_826_n 0.0147221f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_254 N_A_c_178_n N_VPWR_M1009_d 0.00187547f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_255 N_A_c_178_n N_VPWR_M1028_d 0.00187547f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_256 N_A_c_169_n N_VPWR_c_882_n 0.00300743f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_c_170_n N_VPWR_c_882_n 0.00300743f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_c_170_n N_VPWR_c_883_n 0.00523784f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_259 N_A_c_171_n N_VPWR_c_883_n 0.00523784f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_260 N_A_c_171_n N_VPWR_c_884_n 0.00300743f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_c_172_n N_VPWR_c_884_n 0.00300743f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_c_173_n N_VPWR_c_887_n 0.00300743f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_c_174_n N_VPWR_c_887_n 0.00300743f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_c_175_n N_VPWR_c_888_n 0.00300743f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_265 N_A_c_176_n N_VPWR_c_888_n 0.00300743f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_266 N_A_c_172_n N_VPWR_c_889_n 0.00523784f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_c_173_n N_VPWR_c_893_n 0.00523784f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_268 N_A_c_174_n N_VPWR_c_895_n 0.00523784f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_c_175_n N_VPWR_c_895_n 0.00523784f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_270 N_A_c_176_n N_VPWR_c_897_n 0.00523784f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_c_169_n N_VPWR_c_881_n 0.00771171f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_c_170_n N_VPWR_c_881_n 0.00678659f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_c_171_n N_VPWR_c_881_n 0.00678659f $X=1.45 $Y=1.41 $X2=0 $Y2=0
cc_274 N_A_c_172_n N_VPWR_c_881_n 0.0068118f $X=1.92 $Y=1.41 $X2=0 $Y2=0
cc_275 N_A_c_173_n N_VPWR_c_881_n 0.0068118f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_276 N_A_c_174_n N_VPWR_c_881_n 0.00678659f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_277 N_A_c_175_n N_VPWR_c_881_n 0.00678659f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_278 N_A_c_176_n N_VPWR_c_881_n 0.00806894f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_279 N_A_c_169_n N_VPWR_c_899_n 0.00523784f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_280 N_A_c_178_n N_A_886_297#_M1009_s 0.00290685f $X=6.595 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_281 N_A_c_178_n N_A_886_297#_M1021_s 0.00187091f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_282 N_A_c_178_n N_A_886_297#_M1035_s 0.00187091f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_283 N_A_c_178_n N_A_886_297#_c_1044_n 0.0343218f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_284 N_A_c_178_n N_A_886_297#_c_1045_n 0.0343218f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_285 N_A_c_173_n N_A_886_297#_c_1046_n 0.0132167f $X=6.67 $Y=1.41 $X2=0 $Y2=0
cc_286 N_A_c_174_n N_A_886_297#_c_1046_n 0.014974f $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_287 N_A_c_178_n N_A_886_297#_c_1046_n 0.0123307f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_288 N_A_c_235_p N_A_886_297#_c_1046_n 0.00506447f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_c_168_n N_A_886_297#_c_1046_n 0.0042727f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_290 N_A_c_174_n N_A_886_297#_c_1037_n 6.72222e-19 $X=7.14 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A_c_175_n N_A_886_297#_c_1037_n 7.45525e-19 $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_c_178_n N_A_886_297#_c_1037_n 0.00248473f $X=6.595 $Y=1.53 $X2=0
+ $Y2=0
cc_293 N_A_c_235_p N_A_886_297#_c_1037_n 0.0169096f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_294 N_A_c_168_n N_A_886_297#_c_1037_n 0.00655264f $X=8.08 $Y=1.202 $X2=0
+ $Y2=0
cc_295 N_A_c_175_n N_A_886_297#_c_1056_n 0.014974f $X=7.61 $Y=1.41 $X2=0 $Y2=0
cc_296 N_A_c_176_n N_A_886_297#_c_1056_n 0.0134305f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_297 N_A_c_235_p N_A_886_297#_c_1056_n 0.00565689f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_298 N_A_c_168_n N_A_886_297#_c_1056_n 0.00489951f $X=8.08 $Y=1.202 $X2=0
+ $Y2=0
cc_299 N_A_c_178_n N_A_886_297#_c_1040_n 0.0155879f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_300 N_A_c_178_n N_A_886_297#_c_1061_n 0.0128801f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_301 N_A_c_178_n N_A_886_297#_c_1062_n 0.0128801f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_302 N_A_c_176_n N_X_c_1157_n 0.00213319f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_303 N_A_c_176_n N_X_c_1158_n 0.0028697f $X=8.08 $Y=1.41 $X2=0 $Y2=0
cc_304 N_A_c_165_n N_X_c_1150_n 2.57765e-19 $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_305 N_A_c_162_n N_X_c_1154_n 0.00167428f $X=6.645 $Y=0.995 $X2=0 $Y2=0
cc_306 N_A_c_163_n N_X_c_1154_n 0.00161901f $X=7.115 $Y=0.995 $X2=0 $Y2=0
cc_307 N_A_c_164_n N_X_c_1154_n 0.00163764f $X=7.585 $Y=0.995 $X2=0 $Y2=0
cc_308 N_A_c_165_n N_X_c_1154_n 0.00200111f $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_309 N_A_c_178_n N_X_c_1154_n 0.00261094f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_310 N_A_c_203_p N_X_c_1154_n 0.00232257f $X=6.705 $Y=1.275 $X2=0 $Y2=0
cc_311 N_A_c_235_p N_X_c_1154_n 0.0133778f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_312 N_A_c_168_n N_X_c_1154_n 0.00878068f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_313 N_A_c_158_n N_VGND_c_1307_n 0.00452312f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_314 N_A_c_158_n N_VGND_c_1308_n 0.00424416f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_315 N_A_c_159_n N_VGND_c_1308_n 0.00423334f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_316 N_A_c_159_n N_VGND_c_1309_n 0.00379224f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_317 N_A_c_160_n N_VGND_c_1309_n 0.00276126f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_318 N_A_c_160_n N_VGND_c_1310_n 0.00423334f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_319 N_A_c_161_n N_VGND_c_1310_n 0.00437852f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_320 N_A_c_161_n N_VGND_c_1311_n 0.00268723f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_321 N_A_c_162_n N_VGND_c_1314_n 0.00378935f $X=6.645 $Y=0.995 $X2=0 $Y2=0
cc_322 N_A_c_163_n N_VGND_c_1314_n 0.00276126f $X=7.115 $Y=0.995 $X2=0 $Y2=0
cc_323 N_A_c_164_n N_VGND_c_1315_n 0.00385467f $X=7.585 $Y=0.995 $X2=0 $Y2=0
cc_324 N_A_c_165_n N_VGND_c_1315_n 0.00365402f $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_325 N_A_c_165_n N_VGND_c_1316_n 0.00191367f $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_326 N_A_c_162_n N_VGND_c_1324_n 0.00421816f $X=6.645 $Y=0.995 $X2=0 $Y2=0
cc_327 N_A_c_163_n N_VGND_c_1326_n 0.00423334f $X=7.115 $Y=0.995 $X2=0 $Y2=0
cc_328 N_A_c_164_n N_VGND_c_1326_n 0.00423334f $X=7.585 $Y=0.995 $X2=0 $Y2=0
cc_329 N_A_c_165_n N_VGND_c_1328_n 0.00396605f $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_330 N_A_c_158_n N_VGND_c_1335_n 0.00683136f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_331 N_A_c_159_n N_VGND_c_1335_n 0.006093f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A_c_160_n N_VGND_c_1335_n 0.00608558f $X=1.425 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A_c_161_n N_VGND_c_1335_n 0.00615622f $X=1.945 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A_c_162_n N_VGND_c_1335_n 0.00569377f $X=6.645 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A_c_163_n N_VGND_c_1335_n 0.00566204f $X=7.115 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A_c_164_n N_VGND_c_1335_n 0.00590015f $X=7.585 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A_c_165_n N_VGND_c_1335_n 0.00692882f $X=8.105 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A_c_162_n N_A_886_47#_c_1503_n 0.00282739f $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_339 N_A_c_162_n N_A_886_47#_c_1498_n 0.00519746f $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_340 N_A_c_163_n N_A_886_47#_c_1498_n 4.74935e-19 $X=7.115 $Y=0.995 $X2=0
+ $Y2=0
cc_341 N_A_c_178_n N_A_886_47#_c_1498_n 0.00483984f $X=6.595 $Y=1.53 $X2=0 $Y2=0
cc_342 N_A_c_203_p N_A_886_47#_c_1498_n 3.31107e-19 $X=6.705 $Y=1.275 $X2=0
+ $Y2=0
cc_343 N_A_c_162_n N_A_886_47#_c_1499_n 0.00827789f $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_344 N_A_c_163_n N_A_886_47#_c_1499_n 0.00822505f $X=7.115 $Y=0.995 $X2=0
+ $Y2=0
cc_345 N_A_c_203_p N_A_886_47#_c_1499_n 0.0143048f $X=6.705 $Y=1.275 $X2=0 $Y2=0
cc_346 N_A_c_235_p N_A_886_47#_c_1499_n 0.021418f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_347 N_A_c_168_n N_A_886_47#_c_1499_n 0.00339144f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_348 N_A_c_162_n N_A_886_47#_c_1513_n 5.24597e-19 $X=6.645 $Y=0.995 $X2=0
+ $Y2=0
cc_349 N_A_c_163_n N_A_886_47#_c_1513_n 0.00651696f $X=7.115 $Y=0.995 $X2=0
+ $Y2=0
cc_350 N_A_c_164_n N_A_886_47#_c_1513_n 0.00693563f $X=7.585 $Y=0.995 $X2=0
+ $Y2=0
cc_351 N_A_c_165_n N_A_886_47#_c_1513_n 5.34196e-19 $X=8.105 $Y=0.995 $X2=0
+ $Y2=0
cc_352 N_A_c_164_n N_A_886_47#_c_1500_n 0.00855789f $X=7.585 $Y=0.995 $X2=0
+ $Y2=0
cc_353 N_A_c_165_n N_A_886_47#_c_1500_n 0.00901452f $X=8.105 $Y=0.995 $X2=0
+ $Y2=0
cc_354 N_A_c_235_p N_A_886_47#_c_1500_n 0.0360353f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_355 N_A_c_168_n N_A_886_47#_c_1500_n 0.00460274f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_356 N_A_c_164_n N_A_886_47#_c_1501_n 5.69266e-19 $X=7.585 $Y=0.995 $X2=0
+ $Y2=0
cc_357 N_A_c_165_n N_A_886_47#_c_1501_n 0.00857123f $X=8.105 $Y=0.995 $X2=0
+ $Y2=0
cc_358 N_A_c_163_n N_A_886_47#_c_1502_n 9.63332e-19 $X=7.115 $Y=0.995 $X2=0
+ $Y2=0
cc_359 N_A_c_164_n N_A_886_47#_c_1502_n 9.63332e-19 $X=7.585 $Y=0.995 $X2=0
+ $Y2=0
cc_360 N_A_c_235_p N_A_886_47#_c_1502_n 0.0245102f $X=7.94 $Y=1.16 $X2=0 $Y2=0
cc_361 N_A_c_168_n N_A_886_47#_c_1502_n 0.00344611f $X=8.08 $Y=1.202 $X2=0 $Y2=0
cc_362 N_B_c_386_n N_A_112_47#_c_546_n 0.00864834f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_363 N_B_c_386_n N_A_112_47#_c_585_n 0.00644736f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_364 N_B_c_387_n N_A_112_47#_c_585_n 0.00686626f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_365 N_B_c_388_n N_A_112_47#_c_585_n 5.45498e-19 $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_366 N_B_c_399_n N_A_112_47#_c_586_n 0.0117828f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_367 N_B_c_400_n N_A_112_47#_c_586_n 0.0107538f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_368 N_B_c_391_n N_A_112_47#_c_586_n 5.77563e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_369 N_B_c_387_n N_A_112_47#_c_547_n 0.00901006f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_370 N_B_c_388_n N_A_112_47#_c_547_n 0.0106213f $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_371 N_B_c_389_n N_A_112_47#_c_547_n 0.00324564f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_372 N_B_c_391_n N_A_112_47#_c_547_n 0.00721626f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_373 N_B_c_396_n N_A_112_47#_c_547_n 0.0349368f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_374 N_B_c_387_n N_A_112_47#_c_640_n 5.24597e-19 $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_375 N_B_c_388_n N_A_112_47#_c_640_n 0.00651696f $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_376 N_B_c_389_n N_A_112_47#_c_640_n 0.00599745f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_377 N_B_c_386_n N_A_112_47#_c_553_n 0.00110712f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_378 N_B_c_387_n N_A_112_47#_c_553_n 0.00116477f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_379 N_B_c_391_n N_A_112_47#_c_553_n 0.00358305f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_380 N_B_c_398_n N_A_112_47#_c_562_n 0.0137126f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_381 N_B_c_399_n N_A_112_47#_c_562_n 0.00114697f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_382 N_B_c_391_n N_A_112_47#_c_562_n 0.00521588f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_383 N_B_c_391_n N_A_112_47#_c_610_n 0.00158214f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_384 N_B_c_399_n N_A_112_47#_c_650_n 0.00376243f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_385 N_B_c_399_n N_A_112_47#_c_563_n 0.00297334f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_386 N_B_c_391_n N_A_112_47#_c_563_n 0.00285862f $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_387 N_B_c_396_n N_A_112_47#_c_563_n 0.0196467f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_388 N_B_c_398_n N_A_112_47#_c_564_n 0.00670553f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_389 N_B_c_391_n N_A_112_47#_c_564_n 3.26338e-19 $X=3.9 $Y=1.16 $X2=0 $Y2=0
cc_390 N_B_c_398_n N_A_27_297#_c_827_n 0.0143148f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_391 N_B_c_399_n N_A_27_297#_c_827_n 0.0100164f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_392 N_B_c_400_n N_A_27_297#_c_817_n 0.0100164f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_393 N_B_c_401_n N_A_27_297#_c_817_n 0.0143148f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_394 N_B_c_404_n N_VPWR_c_885_n 0.00300743f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_395 N_B_c_405_n N_VPWR_c_885_n 0.00300743f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_396 N_B_c_406_n N_VPWR_c_886_n 0.00300743f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_397 N_B_c_407_n N_VPWR_c_886_n 0.00300743f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_398 N_B_c_398_n N_VPWR_c_889_n 0.00429453f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_399 N_B_c_399_n N_VPWR_c_889_n 0.00429453f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_400 N_B_c_400_n N_VPWR_c_889_n 0.00429453f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_401 N_B_c_401_n N_VPWR_c_889_n 0.00429453f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_402 N_B_c_404_n N_VPWR_c_889_n 0.00523784f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_403 N_B_c_405_n N_VPWR_c_891_n 0.00523784f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_404 N_B_c_406_n N_VPWR_c_891_n 0.00523784f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_405 N_B_c_407_n N_VPWR_c_893_n 0.00523784f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_406 N_B_c_398_n N_VPWR_c_881_n 0.00609021f $X=2.39 $Y=1.41 $X2=0 $Y2=0
cc_407 N_B_c_399_n N_VPWR_c_881_n 0.00606499f $X=2.86 $Y=1.41 $X2=0 $Y2=0
cc_408 N_B_c_400_n N_VPWR_c_881_n 0.00606499f $X=3.33 $Y=1.41 $X2=0 $Y2=0
cc_409 N_B_c_401_n N_VPWR_c_881_n 0.00734734f $X=3.8 $Y=1.41 $X2=0 $Y2=0
cc_410 N_B_c_404_n N_VPWR_c_881_n 0.00806894f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_411 N_B_c_405_n N_VPWR_c_881_n 0.00678659f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_412 N_B_c_406_n N_VPWR_c_881_n 0.00678659f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_413 N_B_c_407_n N_VPWR_c_881_n 0.0068118f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_414 N_B_c_404_n N_A_886_297#_c_1044_n 0.0132364f $X=4.79 $Y=1.41 $X2=0 $Y2=0
cc_415 N_B_c_405_n N_A_886_297#_c_1044_n 0.0132364f $X=5.26 $Y=1.41 $X2=0 $Y2=0
cc_416 N_B_c_406_n N_A_886_297#_c_1045_n 0.0132364f $X=5.73 $Y=1.41 $X2=0 $Y2=0
cc_417 N_B_c_407_n N_A_886_297#_c_1045_n 0.0132364f $X=6.2 $Y=1.41 $X2=0 $Y2=0
cc_418 N_B_c_394_n N_X_c_1176_n 4.20042e-19 $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_419 N_B_c_396_n N_X_c_1176_n 0.00195803f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_420 N_B_c_395_n N_X_c_1154_n 0.00357687f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_421 N_B_c_396_n N_X_c_1154_n 0.00302344f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_422 N_B_c_390_n N_X_c_1155_n 8.71943e-19 $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_423 N_B_c_392_n N_X_c_1155_n 0.0123391f $X=4.765 $Y=0.995 $X2=0 $Y2=0
cc_424 N_B_c_393_n N_X_c_1155_n 0.0114353f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_425 N_B_c_394_n N_X_c_1155_n 0.00439082f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_426 N_B_c_396_n N_X_c_1155_n 0.0758521f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_427 N_B_c_397_n N_X_c_1155_n 0.00699375f $X=6.2 $Y=1.202 $X2=0 $Y2=0
cc_428 N_B_c_393_n N_X_c_1156_n 2.53296e-19 $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_429 N_B_c_394_n N_X_c_1156_n 0.00821074f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_430 N_B_c_395_n N_X_c_1156_n 0.0011756f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_431 N_B_c_396_n N_X_c_1156_n 0.0310846f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_432 N_B_c_397_n N_X_c_1156_n 0.00492344f $X=6.2 $Y=1.202 $X2=0 $Y2=0
cc_433 N_B_c_386_n N_VGND_c_1311_n 0.00268723f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_434 N_B_c_387_n N_VGND_c_1312_n 0.00379224f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_388_n N_VGND_c_1312_n 0.00276126f $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_436 N_B_c_389_n N_VGND_c_1313_n 0.00695442f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_390_n N_VGND_c_1313_n 0.00684795f $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_438 N_B_c_392_n N_VGND_c_1313_n 0.00685325f $X=4.765 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_396_n N_VGND_c_1313_n 0.0201588f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_440 N_B_c_386_n N_VGND_c_1320_n 0.00423334f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_387_n N_VGND_c_1320_n 0.00423334f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_388_n N_VGND_c_1322_n 0.00423334f $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_389_n N_VGND_c_1322_n 0.00541359f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_444 N_B_c_392_n N_VGND_c_1324_n 0.00357877f $X=4.765 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_393_n N_VGND_c_1324_n 0.00357877f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_446 N_B_c_394_n N_VGND_c_1324_n 0.00357877f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_c_395_n N_VGND_c_1324_n 0.00357877f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_448 N_B_c_386_n N_VGND_c_1335_n 0.00587047f $X=2.365 $Y=0.995 $X2=0 $Y2=0
cc_449 N_B_c_387_n N_VGND_c_1335_n 0.006093f $X=2.835 $Y=0.995 $X2=0 $Y2=0
cc_450 N_B_c_388_n N_VGND_c_1335_n 0.00597024f $X=3.305 $Y=0.995 $X2=0 $Y2=0
cc_451 N_B_c_389_n N_VGND_c_1335_n 0.0110773f $X=3.775 $Y=0.995 $X2=0 $Y2=0
cc_452 N_B_c_392_n N_VGND_c_1335_n 0.00668309f $X=4.765 $Y=0.995 $X2=0 $Y2=0
cc_453 N_B_c_393_n N_VGND_c_1335_n 0.00548399f $X=5.235 $Y=0.995 $X2=0 $Y2=0
cc_454 N_B_c_394_n N_VGND_c_1335_n 0.00547171f $X=5.705 $Y=0.995 $X2=0 $Y2=0
cc_455 N_B_c_395_n N_VGND_c_1335_n 0.00545144f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_456 N_B_c_390_n N_A_886_47#_c_1497_n 0.00316065f $X=4.69 $Y=1.16 $X2=0 $Y2=0
cc_457 N_B_c_392_n N_A_886_47#_c_1497_n 0.00931157f $X=4.765 $Y=0.995 $X2=0
+ $Y2=0
cc_458 N_B_c_393_n N_A_886_47#_c_1497_n 0.00931157f $X=5.235 $Y=0.995 $X2=0
+ $Y2=0
cc_459 N_B_c_394_n N_A_886_47#_c_1497_n 0.00958957f $X=5.705 $Y=0.995 $X2=0
+ $Y2=0
cc_460 N_B_c_395_n N_A_886_47#_c_1497_n 0.0114896f $X=6.225 $Y=0.995 $X2=0 $Y2=0
cc_461 N_B_c_396_n N_A_886_47#_c_1497_n 0.00645639f $X=5.285 $Y=1.16 $X2=0 $Y2=0
cc_462 N_B_c_395_n N_A_886_47#_c_1498_n 3.30353e-19 $X=6.225 $Y=0.995 $X2=0
+ $Y2=0
cc_463 N_A_112_47#_c_561_n N_A_27_297#_M1005_s 0.00208348f $X=0.255 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_464 N_A_112_47#_c_562_n N_A_27_297#_M1005_s 0.00113743f $X=2.5 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_465 N_A_112_47#_c_562_n N_A_27_297#_M1012_s 0.00187091f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_466 N_A_112_47#_c_562_n N_A_27_297#_M1027_s 0.00117265f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_467 N_A_112_47#_c_564_n N_A_27_297#_M1027_s 0.00256594f $X=2.415 $Y=1.53
+ $X2=0 $Y2=0
cc_468 N_A_112_47#_c_586_n N_A_27_297#_M1006_d 0.00332369f $X=3.44 $Y=1.87 $X2=0
+ $Y2=0
cc_469 N_A_112_47#_c_562_n N_A_27_297#_c_822_n 0.0378591f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_470 N_A_112_47#_c_562_n N_A_27_297#_c_824_n 0.0378591f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_471 N_A_112_47#_c_562_n N_A_27_297#_c_839_n 0.0137109f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_472 N_A_112_47#_c_564_n N_A_27_297#_c_839_n 0.0045571f $X=2.415 $Y=1.53 $X2=0
+ $Y2=0
cc_473 N_A_112_47#_M1000_s N_A_27_297#_c_827_n 0.00352392f $X=2.48 $Y=1.485
+ $X2=0 $Y2=0
cc_474 N_A_112_47#_c_586_n N_A_27_297#_c_827_n 0.00608347f $X=3.44 $Y=1.87 $X2=0
+ $Y2=0
cc_475 N_A_112_47#_c_610_n N_A_27_297#_c_827_n 0.0132435f $X=2.625 $Y=1.87 $X2=0
+ $Y2=0
cc_476 N_A_112_47#_M1023_s N_A_27_297#_c_817_n 0.00352392f $X=3.42 $Y=1.485
+ $X2=0 $Y2=0
cc_477 N_A_112_47#_c_586_n N_A_27_297#_c_817_n 0.00608347f $X=3.44 $Y=1.87 $X2=0
+ $Y2=0
cc_478 N_A_112_47#_c_611_n N_A_27_297#_c_817_n 0.0127274f $X=3.565 $Y=1.87 $X2=0
+ $Y2=0
cc_479 N_A_112_47#_c_563_n N_A_27_297#_c_826_n 0.00206914f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_480 N_A_112_47#_c_561_n N_A_27_297#_c_818_n 0.0154106f $X=0.255 $Y=1.53 $X2=0
+ $Y2=0
cc_481 N_A_112_47#_c_562_n N_A_27_297#_c_818_n 0.00875025f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_482 N_A_112_47#_c_562_n N_A_27_297#_c_850_n 0.0143191f $X=2.5 $Y=1.53 $X2=0
+ $Y2=0
cc_483 N_A_112_47#_c_586_n N_A_27_297#_c_851_n 0.0126843f $X=3.44 $Y=1.87 $X2=0
+ $Y2=0
cc_484 N_A_112_47#_c_562_n N_VPWR_M1005_d 0.00187547f $X=2.5 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_485 N_A_112_47#_c_562_n N_VPWR_M1020_d 0.00187547f $X=2.5 $Y=1.53 $X2=0 $Y2=0
cc_486 N_A_112_47#_c_563_n N_VPWR_M1001_d 0.00187762f $X=8.245 $Y=1.53 $X2=0
+ $Y2=0
cc_487 N_A_112_47#_c_563_n N_VPWR_M1013_d 0.00244296f $X=8.245 $Y=1.53 $X2=0
+ $Y2=0
cc_488 N_A_112_47#_c_555_n N_VPWR_c_897_n 0.00429453f $X=9.08 $Y=1.41 $X2=0
+ $Y2=0
cc_489 N_A_112_47#_c_556_n N_VPWR_c_897_n 0.00429453f $X=9.55 $Y=1.41 $X2=0
+ $Y2=0
cc_490 N_A_112_47#_c_557_n N_VPWR_c_897_n 0.00429453f $X=10.02 $Y=1.41 $X2=0
+ $Y2=0
cc_491 N_A_112_47#_c_558_n N_VPWR_c_897_n 0.00658436f $X=10.49 $Y=1.41 $X2=0
+ $Y2=0
cc_492 N_A_112_47#_M1000_s N_VPWR_c_881_n 0.00232092f $X=2.48 $Y=1.485 $X2=0
+ $Y2=0
cc_493 N_A_112_47#_M1023_s N_VPWR_c_881_n 0.00232092f $X=3.42 $Y=1.485 $X2=0
+ $Y2=0
cc_494 N_A_112_47#_c_555_n N_VPWR_c_881_n 0.00739666f $X=9.08 $Y=1.41 $X2=0
+ $Y2=0
cc_495 N_A_112_47#_c_556_n N_VPWR_c_881_n 0.00606499f $X=9.55 $Y=1.41 $X2=0
+ $Y2=0
cc_496 N_A_112_47#_c_557_n N_VPWR_c_881_n 0.00606499f $X=10.02 $Y=1.41 $X2=0
+ $Y2=0
cc_497 N_A_112_47#_c_558_n N_VPWR_c_881_n 0.0125304f $X=10.49 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_A_112_47#_c_586_n N_VPWR_c_881_n 0.00153883f $X=3.44 $Y=1.87 $X2=0
+ $Y2=0
cc_499 N_A_112_47#_c_563_n N_A_886_297#_M1007_s 2.88865e-19 $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_500 N_A_112_47#_c_548_n N_A_886_297#_M1015_s 9.93771e-19 $X=8.425 $Y=1.445
+ $X2=0 $Y2=0
cc_501 N_A_112_47#_c_565_n N_A_886_297#_M1015_s 0.00200743f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_502 N_A_112_47#_c_566_n N_A_886_297#_M1015_s 6.34336e-19 $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_503 N_A_112_47#_c_563_n N_A_886_297#_c_1044_n 0.00508579f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_504 N_A_112_47#_c_563_n N_A_886_297#_c_1045_n 0.00508579f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_505 N_A_112_47#_c_563_n N_A_886_297#_c_1046_n 0.0138242f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_506 N_A_112_47#_c_563_n N_A_886_297#_c_1037_n 0.0263618f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_507 N_A_112_47#_c_566_n N_A_886_297#_c_1037_n 0.00236413f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_508 N_A_112_47#_c_563_n N_A_886_297#_c_1056_n 0.0154279f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_509 N_A_112_47#_c_566_n N_A_886_297#_c_1056_n 0.00999959f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_510 N_A_112_47#_c_548_n N_A_886_297#_c_1038_n 0.00722003f $X=8.425 $Y=1.445
+ $X2=0 $Y2=0
cc_511 N_A_112_47#_c_563_n N_A_886_297#_c_1038_n 4.56591e-19 $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_512 N_A_112_47#_c_565_n N_A_886_297#_c_1038_n 0.00573091f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_513 N_A_112_47#_c_566_n N_A_886_297#_c_1038_n 0.00799355f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_514 N_A_112_47#_c_555_n N_A_886_297#_c_1082_n 0.00400988f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_515 N_A_112_47#_c_555_n N_A_886_297#_c_1039_n 0.0134508f $X=9.08 $Y=1.41
+ $X2=0 $Y2=0
cc_516 N_A_112_47#_c_556_n N_A_886_297#_c_1084_n 0.011451f $X=9.55 $Y=1.41 $X2=0
+ $Y2=0
cc_517 N_A_112_47#_c_557_n N_A_886_297#_c_1084_n 0.01161f $X=10.02 $Y=1.41 $X2=0
+ $Y2=0
cc_518 N_A_112_47#_c_563_n N_A_886_297#_c_1040_n 0.00209664f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_519 N_A_112_47#_c_563_n N_A_886_297#_c_1061_n 0.00209664f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_520 N_A_112_47#_c_563_n N_A_886_297#_c_1062_n 0.00209664f $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_521 N_A_112_47#_c_548_n N_X_c_1157_n 0.0126913f $X=8.425 $Y=1.445 $X2=0 $Y2=0
cc_522 N_A_112_47#_c_550_n N_X_c_1157_n 0.0238882f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_523 N_A_112_47#_c_565_n N_X_c_1157_n 0.00755503f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_524 N_A_112_47#_c_555_n N_X_c_1159_n 0.0146938f $X=9.08 $Y=1.41 $X2=0 $Y2=0
cc_525 N_A_112_47#_c_556_n N_X_c_1159_n 0.0143911f $X=9.55 $Y=1.41 $X2=0 $Y2=0
cc_526 N_A_112_47#_c_550_n N_X_c_1159_n 0.0494835f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_527 N_A_112_47#_c_554_n N_X_c_1159_n 0.00852346f $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_528 N_A_112_47#_c_538_n N_X_c_1198_n 0.00713548f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_529 N_A_112_47#_c_539_n N_X_c_1198_n 0.00686626f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_530 N_A_112_47#_c_540_n N_X_c_1198_n 5.45498e-19 $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_531 N_A_112_47#_c_539_n N_X_c_1147_n 0.00879805f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_532 N_A_112_47#_c_540_n N_X_c_1147_n 0.00879805f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_533 N_A_112_47#_c_550_n N_X_c_1147_n 0.0395697f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_534 N_A_112_47#_c_554_n N_X_c_1147_n 0.00345061f $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_535 N_A_112_47#_c_557_n N_X_c_1160_n 0.0133152f $X=10.02 $Y=1.41 $X2=0 $Y2=0
cc_536 N_A_112_47#_c_558_n N_X_c_1160_n 0.0150608f $X=10.49 $Y=1.41 $X2=0 $Y2=0
cc_537 N_A_112_47#_c_550_n N_X_c_1160_n 0.015279f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_538 N_A_112_47#_c_554_n N_X_c_1160_n 0.0091176f $X=10.49 $Y=1.202 $X2=0 $Y2=0
cc_539 N_A_112_47#_c_539_n N_X_c_1209_n 5.55006e-19 $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_540 N_A_112_47#_c_540_n N_X_c_1209_n 0.00670162f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_541 N_A_112_47#_c_541_n N_X_c_1148_n 0.0137257f $X=10.515 $Y=0.995 $X2=0
+ $Y2=0
cc_542 N_A_112_47#_c_558_n N_X_c_1149_n 0.00145198f $X=10.49 $Y=1.41 $X2=0 $Y2=0
cc_543 N_A_112_47#_c_541_n N_X_c_1149_n 0.0213159f $X=10.515 $Y=0.995 $X2=0
+ $Y2=0
cc_544 N_A_112_47#_c_550_n N_X_c_1149_n 0.00724749f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_545 N_A_112_47#_c_538_n N_X_c_1150_n 0.0101363f $X=9.055 $Y=0.995 $X2=0 $Y2=0
cc_546 N_A_112_47#_c_550_n N_X_c_1150_n 0.0300063f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_547 N_A_112_47#_c_538_n N_X_c_1151_n 0.00116636f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_548 N_A_112_47#_c_539_n N_X_c_1151_n 0.00132436f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_549 N_A_112_47#_c_550_n N_X_c_1151_n 0.0306016f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_550 N_A_112_47#_c_554_n N_X_c_1151_n 0.00358305f $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_551 N_A_112_47#_c_550_n N_X_c_1162_n 0.020385f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_552 N_A_112_47#_c_554_n N_X_c_1162_n 0.00663436f $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_553 N_A_112_47#_c_540_n N_X_c_1152_n 0.00116834f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_554 N_A_112_47#_c_550_n N_X_c_1152_n 0.00717779f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_555 N_A_112_47#_c_554_n N_X_c_1152_n 0.00600969f $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_556 N_A_112_47#_c_558_n N_X_c_1163_n 0.00207355f $X=10.49 $Y=1.41 $X2=0 $Y2=0
cc_557 N_A_112_47#_c_554_n N_X_c_1163_n 3.89106e-19 $X=10.49 $Y=1.202 $X2=0
+ $Y2=0
cc_558 N_A_112_47#_c_557_n X 5.75408e-19 $X=10.02 $Y=1.41 $X2=0 $Y2=0
cc_559 N_A_112_47#_c_558_n X 0.0111674f $X=10.49 $Y=1.41 $X2=0 $Y2=0
cc_560 N_A_112_47#_c_563_n N_X_c_1176_n 0.113372f $X=8.245 $Y=1.53 $X2=0 $Y2=0
cc_561 N_A_112_47#_c_538_n N_X_c_1153_n 0.00162656f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_562 N_A_112_47#_c_549_n N_X_c_1154_n 0.00268624f $X=8.51 $Y=1.175 $X2=0 $Y2=0
cc_563 N_A_112_47#_c_550_n N_X_c_1154_n 0.0157298f $X=9.945 $Y=1.16 $X2=0 $Y2=0
cc_564 N_A_112_47#_c_565_n N_X_c_1154_n 0.0145091f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_565 N_A_112_47#_c_566_n N_X_c_1154_n 0.00157657f $X=8.39 $Y=1.53 $X2=0 $Y2=0
cc_566 N_A_112_47#_c_543_n N_VGND_M1003_s 0.00100734f $X=0.53 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_567 N_A_112_47#_c_544_n N_VGND_M1003_s 0.002086f $X=0.255 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_568 N_A_112_47#_c_545_n N_VGND_M1014_s 0.00251047f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_569 N_A_112_47#_c_546_n N_VGND_M1031_s 0.00162089f $X=2.41 $Y=0.815 $X2=0
+ $Y2=0
cc_570 N_A_112_47#_c_547_n N_VGND_M1025_d 0.00251047f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_571 N_A_112_47#_c_543_n N_VGND_c_1307_n 0.00765622f $X=0.53 $Y=0.82 $X2=0
+ $Y2=0
cc_572 N_A_112_47#_c_544_n N_VGND_c_1307_n 0.0148186f $X=0.255 $Y=0.82 $X2=0
+ $Y2=0
cc_573 N_A_112_47#_c_543_n N_VGND_c_1308_n 0.00193763f $X=0.53 $Y=0.82 $X2=0
+ $Y2=0
cc_574 N_A_112_47#_c_574_n N_VGND_c_1308_n 0.0223596f $X=0.745 $Y=0.39 $X2=0
+ $Y2=0
cc_575 N_A_112_47#_c_545_n N_VGND_c_1308_n 0.00266636f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_576 N_A_112_47#_c_574_n N_VGND_c_1309_n 0.0183628f $X=0.745 $Y=0.39 $X2=0
+ $Y2=0
cc_577 N_A_112_47#_c_545_n N_VGND_c_1309_n 0.0127273f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_578 N_A_112_47#_c_545_n N_VGND_c_1310_n 0.00198695f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_579 N_A_112_47#_c_581_n N_VGND_c_1310_n 0.0231806f $X=1.685 $Y=0.39 $X2=0
+ $Y2=0
cc_580 N_A_112_47#_c_546_n N_VGND_c_1310_n 0.00254521f $X=2.41 $Y=0.815 $X2=0
+ $Y2=0
cc_581 N_A_112_47#_c_546_n N_VGND_c_1311_n 0.0122559f $X=2.41 $Y=0.815 $X2=0
+ $Y2=0
cc_582 N_A_112_47#_c_585_n N_VGND_c_1312_n 0.0183628f $X=2.625 $Y=0.39 $X2=0
+ $Y2=0
cc_583 N_A_112_47#_c_547_n N_VGND_c_1312_n 0.0127273f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_584 N_A_112_47#_c_547_n N_VGND_c_1313_n 0.0113219f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_585 N_A_112_47#_c_640_n N_VGND_c_1313_n 0.0297488f $X=3.565 $Y=0.39 $X2=0
+ $Y2=0
cc_586 N_A_112_47#_c_538_n N_VGND_c_1316_n 0.00438629f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_587 N_A_112_47#_c_539_n N_VGND_c_1317_n 0.00379224f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_588 N_A_112_47#_c_540_n N_VGND_c_1317_n 0.00276126f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_589 N_A_112_47#_c_541_n N_VGND_c_1319_n 0.00438629f $X=10.515 $Y=0.995 $X2=0
+ $Y2=0
cc_590 N_A_112_47#_c_546_n N_VGND_c_1320_n 0.00198695f $X=2.41 $Y=0.815 $X2=0
+ $Y2=0
cc_591 N_A_112_47#_c_585_n N_VGND_c_1320_n 0.0223596f $X=2.625 $Y=0.39 $X2=0
+ $Y2=0
cc_592 N_A_112_47#_c_547_n N_VGND_c_1320_n 0.00266636f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_593 N_A_112_47#_c_547_n N_VGND_c_1322_n 0.00198695f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_594 N_A_112_47#_c_640_n N_VGND_c_1322_n 0.0223596f $X=3.565 $Y=0.39 $X2=0
+ $Y2=0
cc_595 N_A_112_47#_c_538_n N_VGND_c_1330_n 0.00423334f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_596 N_A_112_47#_c_539_n N_VGND_c_1330_n 0.00424416f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_597 N_A_112_47#_c_540_n N_VGND_c_1332_n 0.00424416f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_598 N_A_112_47#_c_541_n N_VGND_c_1332_n 0.00439206f $X=10.515 $Y=0.995 $X2=0
+ $Y2=0
cc_599 N_A_112_47#_M1003_d N_VGND_c_1335_n 0.0025535f $X=0.56 $Y=0.235 $X2=0
+ $Y2=0
cc_600 N_A_112_47#_M1030_d N_VGND_c_1335_n 0.00304143f $X=1.5 $Y=0.235 $X2=0
+ $Y2=0
cc_601 N_A_112_47#_M1011_s N_VGND_c_1335_n 0.0025535f $X=2.44 $Y=0.235 $X2=0
+ $Y2=0
cc_602 N_A_112_47#_M1026_s N_VGND_c_1335_n 0.0025535f $X=3.38 $Y=0.235 $X2=0
+ $Y2=0
cc_603 N_A_112_47#_c_538_n N_VGND_c_1335_n 0.00712117f $X=9.055 $Y=0.995 $X2=0
+ $Y2=0
cc_604 N_A_112_47#_c_539_n N_VGND_c_1335_n 0.00611278f $X=9.525 $Y=0.995 $X2=0
+ $Y2=0
cc_605 N_A_112_47#_c_540_n N_VGND_c_1335_n 0.00610535f $X=9.995 $Y=0.995 $X2=0
+ $Y2=0
cc_606 N_A_112_47#_c_541_n N_VGND_c_1335_n 0.00715658f $X=10.515 $Y=0.995 $X2=0
+ $Y2=0
cc_607 N_A_112_47#_c_543_n N_VGND_c_1335_n 0.004202f $X=0.53 $Y=0.82 $X2=0 $Y2=0
cc_608 N_A_112_47#_c_544_n N_VGND_c_1335_n 7.18354e-19 $X=0.255 $Y=0.82 $X2=0
+ $Y2=0
cc_609 N_A_112_47#_c_574_n N_VGND_c_1335_n 0.0141302f $X=0.745 $Y=0.39 $X2=0
+ $Y2=0
cc_610 N_A_112_47#_c_545_n N_VGND_c_1335_n 0.00972452f $X=1.47 $Y=0.815 $X2=0
+ $Y2=0
cc_611 N_A_112_47#_c_581_n N_VGND_c_1335_n 0.0143352f $X=1.685 $Y=0.39 $X2=0
+ $Y2=0
cc_612 N_A_112_47#_c_546_n N_VGND_c_1335_n 0.0094839f $X=2.41 $Y=0.815 $X2=0
+ $Y2=0
cc_613 N_A_112_47#_c_585_n N_VGND_c_1335_n 0.0141302f $X=2.625 $Y=0.39 $X2=0
+ $Y2=0
cc_614 N_A_112_47#_c_547_n N_VGND_c_1335_n 0.00972452f $X=3.35 $Y=0.815 $X2=0
+ $Y2=0
cc_615 N_A_112_47#_c_640_n N_VGND_c_1335_n 0.0141302f $X=3.565 $Y=0.39 $X2=0
+ $Y2=0
cc_616 N_A_112_47#_c_563_n N_A_886_47#_c_1498_n 3.13965e-19 $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_617 N_A_112_47#_c_563_n N_A_886_47#_c_1499_n 2.18522e-19 $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_618 N_A_112_47#_c_538_n N_A_886_47#_c_1500_n 6.1243e-19 $X=9.055 $Y=0.995
+ $X2=0 $Y2=0
cc_619 N_A_112_47#_c_549_n N_A_886_47#_c_1500_n 0.0103246f $X=8.51 $Y=1.175
+ $X2=0 $Y2=0
cc_620 N_A_112_47#_c_563_n N_A_886_47#_c_1500_n 2.68676e-19 $X=8.245 $Y=1.53
+ $X2=0 $Y2=0
cc_621 N_A_112_47#_c_565_n N_A_886_47#_c_1500_n 5.83411e-19 $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_622 N_A_112_47#_c_566_n N_A_886_47#_c_1500_n 0.00414852f $X=8.39 $Y=1.53
+ $X2=0 $Y2=0
cc_623 N_A_112_47#_c_538_n N_A_886_47#_c_1501_n 0.0029957f $X=9.055 $Y=0.995
+ $X2=0 $Y2=0
cc_624 N_A_27_297#_c_822_n N_VPWR_M1005_d 0.00349582f $X=1.09 $Y=1.895 $X2=-0.19
+ $Y2=1.305
cc_625 N_A_27_297#_c_824_n N_VPWR_M1020_d 0.00349582f $X=2.03 $Y=1.895 $X2=0
+ $Y2=0
cc_626 N_A_27_297#_c_822_n N_VPWR_c_882_n 0.0139741f $X=1.09 $Y=1.895 $X2=0
+ $Y2=0
cc_627 N_A_27_297#_c_822_n N_VPWR_c_883_n 0.0028084f $X=1.09 $Y=1.895 $X2=0
+ $Y2=0
cc_628 N_A_27_297#_c_824_n N_VPWR_c_883_n 0.0028084f $X=2.03 $Y=1.895 $X2=0
+ $Y2=0
cc_629 N_A_27_297#_c_850_n N_VPWR_c_883_n 0.0149311f $X=1.215 $Y=1.96 $X2=0
+ $Y2=0
cc_630 N_A_27_297#_c_824_n N_VPWR_c_884_n 0.0139741f $X=2.03 $Y=1.895 $X2=0
+ $Y2=0
cc_631 N_A_27_297#_c_824_n N_VPWR_c_889_n 0.0028084f $X=2.03 $Y=1.895 $X2=0
+ $Y2=0
cc_632 N_A_27_297#_c_827_n N_VPWR_c_889_n 0.0386815f $X=2.97 $Y=2.38 $X2=0 $Y2=0
cc_633 N_A_27_297#_c_861_p N_VPWR_c_889_n 0.015002f $X=2.28 $Y=2.38 $X2=0 $Y2=0
cc_634 N_A_27_297#_c_817_n N_VPWR_c_889_n 0.0549564f $X=3.91 $Y=2.38 $X2=0 $Y2=0
cc_635 N_A_27_297#_c_851_n N_VPWR_c_889_n 0.014332f $X=3.095 $Y=2.3 $X2=0 $Y2=0
cc_636 N_A_27_297#_M1005_s N_VPWR_c_881_n 0.00238174f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_637 N_A_27_297#_M1012_s N_VPWR_c_881_n 0.0024798f $X=1.07 $Y=1.485 $X2=0
+ $Y2=0
cc_638 N_A_27_297#_M1027_s N_VPWR_c_881_n 0.00240425f $X=2.01 $Y=1.485 $X2=0
+ $Y2=0
cc_639 N_A_27_297#_M1006_d N_VPWR_c_881_n 0.00229658f $X=2.95 $Y=1.485 $X2=0
+ $Y2=0
cc_640 N_A_27_297#_M1033_d N_VPWR_c_881_n 0.00217519f $X=3.89 $Y=1.485 $X2=0
+ $Y2=0
cc_641 N_A_27_297#_c_822_n N_VPWR_c_881_n 0.0108264f $X=1.09 $Y=1.895 $X2=0
+ $Y2=0
cc_642 N_A_27_297#_c_824_n N_VPWR_c_881_n 0.0108264f $X=2.03 $Y=1.895 $X2=0
+ $Y2=0
cc_643 N_A_27_297#_c_827_n N_VPWR_c_881_n 0.0239144f $X=2.97 $Y=2.38 $X2=0 $Y2=0
cc_644 N_A_27_297#_c_861_p N_VPWR_c_881_n 0.00962794f $X=2.28 $Y=2.38 $X2=0
+ $Y2=0
cc_645 N_A_27_297#_c_817_n N_VPWR_c_881_n 0.0335426f $X=3.91 $Y=2.38 $X2=0 $Y2=0
cc_646 N_A_27_297#_c_818_n N_VPWR_c_881_n 0.0120542f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_647 N_A_27_297#_c_850_n N_VPWR_c_881_n 0.00955092f $X=1.215 $Y=1.96 $X2=0
+ $Y2=0
cc_648 N_A_27_297#_c_851_n N_VPWR_c_881_n 0.00938745f $X=3.095 $Y=2.3 $X2=0
+ $Y2=0
cc_649 N_A_27_297#_c_822_n N_VPWR_c_899_n 0.0028084f $X=1.09 $Y=1.895 $X2=0
+ $Y2=0
cc_650 N_A_27_297#_c_818_n N_VPWR_c_899_n 0.0208235f $X=0.275 $Y=1.96 $X2=0
+ $Y2=0
cc_651 N_A_27_297#_c_817_n N_A_886_297#_c_1040_n 0.0100846f $X=3.91 $Y=2.38
+ $X2=0 $Y2=0
cc_652 N_A_27_297#_c_826_n N_A_886_297#_c_1040_n 0.0282783f $X=4.035 $Y=1.96
+ $X2=0 $Y2=0
cc_653 N_VPWR_c_881_n N_A_886_297#_M1009_s 0.00225074f $X=10.81 $Y=2.72
+ $X2=-0.19 $Y2=-0.24
cc_654 N_VPWR_c_881_n N_A_886_297#_M1021_s 0.0024798f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_655 N_VPWR_c_881_n N_A_886_297#_M1035_s 0.0024798f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_656 N_VPWR_c_881_n N_A_886_297#_M1007_s 0.0024798f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_657 N_VPWR_c_881_n N_A_886_297#_M1015_s 0.0022668f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_658 N_VPWR_c_881_n N_A_886_297#_M1016_d 0.00231264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_659 N_VPWR_c_881_n N_A_886_297#_M1029_d 0.00297222f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_660 N_VPWR_M1009_d N_A_886_297#_c_1044_n 0.00334944f $X=4.88 $Y=1.485 $X2=0
+ $Y2=0
cc_661 N_VPWR_c_885_n N_A_886_297#_c_1044_n 0.0135607f $X=5.025 $Y=2.34 $X2=0
+ $Y2=0
cc_662 N_VPWR_c_889_n N_A_886_297#_c_1044_n 0.0028084f $X=4.9 $Y=2.72 $X2=0
+ $Y2=0
cc_663 N_VPWR_c_891_n N_A_886_297#_c_1044_n 0.0028084f $X=5.84 $Y=2.72 $X2=0
+ $Y2=0
cc_664 N_VPWR_c_881_n N_A_886_297#_c_1044_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_665 N_VPWR_M1028_d N_A_886_297#_c_1045_n 0.00334944f $X=5.82 $Y=1.485 $X2=0
+ $Y2=0
cc_666 N_VPWR_c_886_n N_A_886_297#_c_1045_n 0.0135607f $X=5.965 $Y=2.34 $X2=0
+ $Y2=0
cc_667 N_VPWR_c_891_n N_A_886_297#_c_1045_n 0.0028084f $X=5.84 $Y=2.72 $X2=0
+ $Y2=0
cc_668 N_VPWR_c_893_n N_A_886_297#_c_1045_n 0.0028084f $X=6.78 $Y=2.72 $X2=0
+ $Y2=0
cc_669 N_VPWR_c_881_n N_A_886_297#_c_1045_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_670 N_VPWR_M1001_d N_A_886_297#_c_1046_n 0.00412184f $X=6.76 $Y=1.485 $X2=0
+ $Y2=0
cc_671 N_VPWR_c_887_n N_A_886_297#_c_1046_n 0.0135607f $X=6.905 $Y=2.34 $X2=0
+ $Y2=0
cc_672 N_VPWR_c_893_n N_A_886_297#_c_1046_n 0.0028084f $X=6.78 $Y=2.72 $X2=0
+ $Y2=0
cc_673 N_VPWR_c_895_n N_A_886_297#_c_1046_n 0.0028084f $X=7.72 $Y=2.72 $X2=0
+ $Y2=0
cc_674 N_VPWR_c_881_n N_A_886_297#_c_1046_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_675 N_VPWR_M1013_d N_A_886_297#_c_1056_n 0.00412184f $X=7.7 $Y=1.485 $X2=0
+ $Y2=0
cc_676 N_VPWR_c_888_n N_A_886_297#_c_1056_n 0.0135607f $X=7.845 $Y=2.34 $X2=0
+ $Y2=0
cc_677 N_VPWR_c_895_n N_A_886_297#_c_1056_n 0.0028084f $X=7.72 $Y=2.72 $X2=0
+ $Y2=0
cc_678 N_VPWR_c_897_n N_A_886_297#_c_1056_n 0.0028084f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_679 N_VPWR_c_881_n N_A_886_297#_c_1056_n 0.0108264f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_680 N_VPWR_c_897_n N_A_886_297#_c_1039_n 0.0452646f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_681 N_VPWR_c_881_n N_A_886_297#_c_1039_n 0.0270376f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_682 N_VPWR_c_897_n N_A_886_297#_c_1120_n 0.0162911f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_683 N_VPWR_c_881_n N_A_886_297#_c_1120_n 0.00962794f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_684 N_VPWR_c_897_n N_A_886_297#_c_1084_n 0.0536701f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_685 N_VPWR_c_881_n N_A_886_297#_c_1084_n 0.0335386f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_686 N_VPWR_c_889_n N_A_886_297#_c_1040_n 0.0161853f $X=4.9 $Y=2.72 $X2=0
+ $Y2=0
cc_687 N_VPWR_c_881_n N_A_886_297#_c_1040_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_688 N_VPWR_c_891_n N_A_886_297#_c_1061_n 0.0149311f $X=5.84 $Y=2.72 $X2=0
+ $Y2=0
cc_689 N_VPWR_c_881_n N_A_886_297#_c_1061_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_690 N_VPWR_c_893_n N_A_886_297#_c_1062_n 0.0149311f $X=6.78 $Y=2.72 $X2=0
+ $Y2=0
cc_691 N_VPWR_c_881_n N_A_886_297#_c_1062_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_692 N_VPWR_c_895_n N_A_886_297#_c_1130_n 0.0149311f $X=7.72 $Y=2.72 $X2=0
+ $Y2=0
cc_693 N_VPWR_c_881_n N_A_886_297#_c_1130_n 0.00955092f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_694 N_VPWR_c_897_n N_A_886_297#_c_1132_n 0.014933f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_695 N_VPWR_c_881_n N_A_886_297#_c_1132_n 0.00960883f $X=10.81 $Y=2.72 $X2=0
+ $Y2=0
cc_696 N_VPWR_c_881_n N_X_M1016_s 0.00226545f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_697 N_VPWR_c_881_n N_X_M1024_s 0.00232895f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_698 N_VPWR_c_881_n N_X_M1034_s 0.00233913f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_699 N_VPWR_c_897_n X 0.0263741f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_700 N_VPWR_c_881_n X 0.0153152f $X=10.81 $Y=2.72 $X2=0 $Y2=0
cc_701 N_A_886_297#_c_1039_n N_X_M1016_s 0.00539485f $X=9.19 $Y=2.38 $X2=0 $Y2=0
cc_702 N_A_886_297#_c_1084_n N_X_M1024_s 0.00352392f $X=10.13 $Y=2.38 $X2=0
+ $Y2=0
cc_703 N_A_886_297#_c_1038_n N_X_c_1158_n 0.0147657f $X=8.315 $Y=2.005 $X2=0
+ $Y2=0
cc_704 N_A_886_297#_c_1082_n N_X_c_1158_n 0.00740215f $X=8.315 $Y=2.295 $X2=0
+ $Y2=0
cc_705 N_A_886_297#_c_1039_n N_X_c_1158_n 0.0192853f $X=9.19 $Y=2.38 $X2=0 $Y2=0
cc_706 N_A_886_297#_M1016_d N_X_c_1159_n 0.00188585f $X=9.17 $Y=1.485 $X2=0
+ $Y2=0
cc_707 N_A_886_297#_c_1039_n N_X_c_1159_n 0.00416884f $X=9.19 $Y=2.38 $X2=0
+ $Y2=0
cc_708 N_A_886_297#_c_1141_p N_X_c_1159_n 0.0144831f $X=9.315 $Y=2 $X2=0 $Y2=0
cc_709 N_A_886_297#_c_1084_n N_X_c_1159_n 0.00416884f $X=10.13 $Y=2.38 $X2=0
+ $Y2=0
cc_710 N_A_886_297#_M1029_d N_X_c_1160_n 0.00187422f $X=10.11 $Y=1.485 $X2=0
+ $Y2=0
cc_711 N_A_886_297#_c_1084_n N_X_c_1160_n 0.00387236f $X=10.13 $Y=2.38 $X2=0
+ $Y2=0
cc_712 N_A_886_297#_c_1145_p N_X_c_1160_n 0.0143571f $X=10.255 $Y=1.96 $X2=0
+ $Y2=0
cc_713 N_A_886_297#_c_1084_n N_X_c_1162_n 0.0134104f $X=10.13 $Y=2.38 $X2=0
+ $Y2=0
cc_714 N_X_c_1150_n N_VGND_M1010_s 0.00198367f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_715 N_X_c_1153_n N_VGND_M1010_s 0.00193855f $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_716 N_X_c_1147_n N_VGND_M1019_s 0.00255557f $X=10.04 $Y=0.82 $X2=0 $Y2=0
cc_717 N_X_c_1148_n N_VGND_M1038_s 0.00384351f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_718 N_X_c_1155_n N_VGND_c_1313_n 0.012822f $X=5.65 $Y=0.79 $X2=0 $Y2=0
cc_719 N_X_c_1154_n N_VGND_c_1314_n 7.99957e-19 $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_720 N_X_c_1154_n N_VGND_c_1315_n 7.99957e-19 $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_721 N_X_c_1150_n N_VGND_c_1316_n 0.0115042f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_722 N_X_c_1153_n N_VGND_c_1316_n 0.00198703f $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_723 N_X_c_1198_n N_VGND_c_1317_n 0.0183628f $X=9.315 $Y=0.39 $X2=0 $Y2=0
cc_724 N_X_c_1147_n N_VGND_c_1317_n 0.012101f $X=10.04 $Y=0.82 $X2=0 $Y2=0
cc_725 N_X_c_1148_n N_VGND_c_1318_n 0.00237165f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_726 N_X_c_1148_n N_VGND_c_1319_n 0.0133599f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_727 N_X_c_1150_n N_VGND_c_1328_n 0.00163475f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_728 N_X_c_1153_n N_VGND_c_1328_n 2.28408e-19 $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_729 N_X_c_1198_n N_VGND_c_1330_n 0.0223596f $X=9.315 $Y=0.39 $X2=0 $Y2=0
cc_730 N_X_c_1147_n N_VGND_c_1330_n 0.00260082f $X=10.04 $Y=0.82 $X2=0 $Y2=0
cc_731 N_X_c_1150_n N_VGND_c_1330_n 0.00216539f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_732 N_X_c_1153_n N_VGND_c_1330_n 2.58473e-19 $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_733 N_X_c_1147_n N_VGND_c_1332_n 0.00193763f $X=10.04 $Y=0.82 $X2=0 $Y2=0
cc_734 N_X_c_1209_n N_VGND_c_1332_n 0.0231806f $X=10.255 $Y=0.39 $X2=0 $Y2=0
cc_735 N_X_c_1148_n N_VGND_c_1332_n 0.00245178f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_736 N_X_M1002_d N_VGND_c_1335_n 0.00256987f $X=4.84 $Y=0.235 $X2=0 $Y2=0
cc_737 N_X_M1022_d N_VGND_c_1335_n 0.00237472f $X=5.78 $Y=0.235 $X2=0 $Y2=0
cc_738 N_X_M1010_d N_VGND_c_1335_n 0.0025535f $X=9.13 $Y=0.235 $X2=0 $Y2=0
cc_739 N_X_M1036_d N_VGND_c_1335_n 0.00304426f $X=10.07 $Y=0.235 $X2=0 $Y2=0
cc_740 N_X_c_1198_n N_VGND_c_1335_n 0.0141302f $X=9.315 $Y=0.39 $X2=0 $Y2=0
cc_741 N_X_c_1147_n N_VGND_c_1335_n 0.00962544f $X=10.04 $Y=0.82 $X2=0 $Y2=0
cc_742 N_X_c_1209_n N_VGND_c_1335_n 0.0143352f $X=10.255 $Y=0.39 $X2=0 $Y2=0
cc_743 N_X_c_1148_n N_VGND_c_1335_n 0.00976426f $X=10.635 $Y=0.82 $X2=0 $Y2=0
cc_744 N_X_c_1150_n N_VGND_c_1335_n 0.00369932f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_745 N_X_c_1176_n N_VGND_c_1335_n 0.0153719f $X=5.935 $Y=0.81 $X2=0 $Y2=0
cc_746 N_X_c_1153_n N_VGND_c_1335_n 0.0160771f $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_747 N_X_c_1154_n N_VGND_c_1335_n 0.126767f $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_748 N_X_c_1155_n N_A_886_47#_M1002_s 0.00441627f $X=5.65 $Y=0.79 $X2=-0.19
+ $Y2=-0.24
cc_749 N_X_c_1155_n N_A_886_47#_M1017_s 0.00214342f $X=5.65 $Y=0.79 $X2=0 $Y2=0
cc_750 N_X_c_1154_n N_A_886_47#_M1037_s 3.83238e-19 $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_751 N_X_M1002_d N_A_886_47#_c_1497_n 0.00400389f $X=4.84 $Y=0.235 $X2=0 $Y2=0
cc_752 N_X_M1022_d N_A_886_47#_c_1497_n 0.00491234f $X=5.78 $Y=0.235 $X2=0 $Y2=0
cc_753 N_X_c_1176_n N_A_886_47#_c_1497_n 0.001084f $X=5.935 $Y=0.81 $X2=0 $Y2=0
cc_754 N_X_c_1154_n N_A_886_47#_c_1497_n 0.00338403f $X=8.705 $Y=0.81 $X2=0
+ $Y2=0
cc_755 N_X_c_1155_n N_A_886_47#_c_1497_n 0.081737f $X=5.65 $Y=0.79 $X2=0 $Y2=0
cc_756 N_X_c_1176_n N_A_886_47#_c_1498_n 4.58815e-19 $X=5.935 $Y=0.81 $X2=0
+ $Y2=0
cc_757 N_X_c_1154_n N_A_886_47#_c_1498_n 0.014681f $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_758 N_X_c_1156_n N_A_886_47#_c_1498_n 0.00415537f $X=5.965 $Y=0.73 $X2=0
+ $Y2=0
cc_759 N_X_c_1154_n N_A_886_47#_c_1499_n 0.0181412f $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_760 N_X_c_1150_n N_A_886_47#_c_1500_n 0.01389f $X=9.1 $Y=0.815 $X2=0 $Y2=0
cc_761 N_X_c_1153_n N_A_886_47#_c_1500_n 3.95087e-19 $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_762 N_X_c_1154_n N_A_886_47#_c_1500_n 0.0379285f $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_763 N_X_c_1198_n N_A_886_47#_c_1501_n 0.00457692f $X=9.315 $Y=0.39 $X2=0
+ $Y2=0
cc_764 N_X_c_1153_n N_A_886_47#_c_1501_n 0.00100553f $X=8.85 $Y=0.81 $X2=0 $Y2=0
cc_765 N_X_c_1154_n N_A_886_47#_c_1502_n 0.0167328f $X=8.705 $Y=0.81 $X2=0 $Y2=0
cc_766 N_VGND_c_1335_n N_A_886_47#_M1002_s 0.00209344f $X=10.81 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_767 N_VGND_c_1335_n N_A_886_47#_M1017_s 0.00255381f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_768 N_VGND_c_1335_n N_A_886_47#_M1037_s 0.00177027f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_769 N_VGND_c_1335_n N_A_886_47#_M1008_d 0.00210051f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_770 N_VGND_c_1335_n N_A_886_47#_M1032_d 0.00172424f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_771 N_VGND_c_1313_n N_A_886_47#_c_1497_n 0.0190116f $X=4.035 $Y=0.39 $X2=0
+ $Y2=0
cc_772 N_VGND_c_1324_n N_A_886_47#_c_1497_n 0.112077f $X=6.82 $Y=0 $X2=0 $Y2=0
cc_773 N_VGND_c_1335_n N_A_886_47#_c_1497_n 0.0564526f $X=10.81 $Y=0 $X2=0 $Y2=0
cc_774 N_VGND_c_1314_n N_A_886_47#_c_1503_n 0.0141571f $X=6.905 $Y=0.39 $X2=0
+ $Y2=0
cc_775 N_VGND_c_1324_n N_A_886_47#_c_1503_n 0.0152108f $X=6.82 $Y=0 $X2=0 $Y2=0
cc_776 N_VGND_c_1335_n N_A_886_47#_c_1503_n 0.00447564f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_777 N_VGND_c_1314_n N_A_886_47#_c_1498_n 0.00471242f $X=6.905 $Y=0.39 $X2=0
+ $Y2=0
cc_778 N_VGND_M1004_s N_A_886_47#_c_1499_n 0.00251047f $X=6.72 $Y=0.235 $X2=0
+ $Y2=0
cc_779 N_VGND_c_1314_n N_A_886_47#_c_1499_n 0.0115286f $X=6.905 $Y=0.39 $X2=0
+ $Y2=0
cc_780 N_VGND_c_1324_n N_A_886_47#_c_1499_n 0.00266636f $X=6.82 $Y=0 $X2=0 $Y2=0
cc_781 N_VGND_c_1326_n N_A_886_47#_c_1499_n 0.00198695f $X=7.76 $Y=0 $X2=0 $Y2=0
cc_782 N_VGND_c_1335_n N_A_886_47#_c_1499_n 0.00428495f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_783 N_VGND_c_1315_n N_A_886_47#_c_1513_n 0.0183628f $X=7.845 $Y=0.39 $X2=0
+ $Y2=0
cc_784 N_VGND_c_1326_n N_A_886_47#_c_1513_n 0.0223596f $X=7.76 $Y=0 $X2=0 $Y2=0
cc_785 N_VGND_c_1335_n N_A_886_47#_c_1513_n 0.00672308f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_786 N_VGND_M1018_s N_A_886_47#_c_1500_n 0.00348805f $X=7.66 $Y=0.235 $X2=0
+ $Y2=0
cc_787 N_VGND_c_1315_n N_A_886_47#_c_1500_n 0.0119556f $X=7.845 $Y=0.39 $X2=0
+ $Y2=0
cc_788 N_VGND_c_1326_n N_A_886_47#_c_1500_n 0.00266636f $X=7.76 $Y=0 $X2=0 $Y2=0
cc_789 N_VGND_c_1328_n N_A_886_47#_c_1500_n 0.00199443f $X=8.76 $Y=0 $X2=0 $Y2=0
cc_790 N_VGND_c_1335_n N_A_886_47#_c_1500_n 0.00440626f $X=10.81 $Y=0 $X2=0
+ $Y2=0
cc_791 N_VGND_c_1315_n N_A_886_47#_c_1501_n 0.0223967f $X=7.845 $Y=0.39 $X2=0
+ $Y2=0
cc_792 N_VGND_c_1316_n N_A_886_47#_c_1501_n 0.0165694f $X=8.845 $Y=0.39 $X2=0
+ $Y2=0
cc_793 N_VGND_c_1328_n N_A_886_47#_c_1501_n 0.024373f $X=8.76 $Y=0 $X2=0 $Y2=0
cc_794 N_VGND_c_1335_n N_A_886_47#_c_1501_n 0.00671219f $X=10.81 $Y=0 $X2=0
+ $Y2=0
