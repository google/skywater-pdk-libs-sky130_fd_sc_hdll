* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb8to1_4 D[7] D[6] D[5] D[4] D[3] D[2] D[1] D[0] S[7]
+ S[6] S[5] S[4] S[3] S[2] S[1] S[0] VGND VNB VPB VPWR Z
X0 VGND D[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_1313_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND D[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_355_613# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_3797_297# a_4239_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X5 VPWR S[6] a_4239_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X6 a_1313_591# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VPWR D[2] a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 VPWR D[5] a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VPWR D[1] a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_4239_793# S[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_1755_793# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X12 a_2839_613# a_2626_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X13 VPWR D[7] a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 Z S[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X15 a_142_599# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X16 Z a_142_325# a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X17 a_1315_911# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND D[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Z a_2626_599# a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X20 a_2626_599# S[5] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 VPWR S[3] a_1755_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X22 a_3797_591# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X23 Z S[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X24 Z S[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X25 a_355_311# a_142_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X26 a_1313_297# a_1755_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X27 Z a_142_325# a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 Z a_4239_793# a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X29 a_1755_793# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X30 VGND S[2] a_1755_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X31 a_3799_911# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 a_142_325# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X33 a_405_66# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 a_3799_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X35 a_405_66# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 a_2839_311# a_2626_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X37 a_355_311# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 a_1315_911# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X39 a_355_311# a_142_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X40 a_3797_591# a_4239_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X41 a_3799_911# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X42 VPWR S[0] a_142_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 a_2839_613# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X44 VGND D[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X45 VPWR D[4] a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X46 a_1313_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X47 a_355_613# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 VPWR S[5] a_2626_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X49 a_3799_47# S[6] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X50 a_405_66# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X51 VPWR D[0] a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X52 VPWR D[6] a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X53 a_3799_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 VGND S[0] a_142_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X56 VPWR D[1] a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X57 VGND D[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X58 Z a_4239_265# a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X59 Z S[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 Z a_142_599# a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 a_3799_911# D[7] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X62 VGND D[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X63 VPWR D[7] a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X64 VPWR D[3] a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_3797_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 Z S[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X67 VPWR S[7] a_4239_793# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X68 a_355_613# a_142_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X69 a_1313_591# a_1755_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X70 Z a_142_599# a_355_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X71 Z a_2626_325# a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 VGND S[1] a_142_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X73 VGND S[5] a_2626_599# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X74 a_2839_613# a_2626_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X75 a_3799_911# S[7] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X76 a_2626_325# S[4] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X77 a_355_613# a_142_599# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X78 a_2839_311# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X79 a_1315_911# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X80 a_405_918# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X81 VGND S[3] a_1755_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X82 Z a_1755_265# a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X83 a_355_311# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X84 a_2626_325# S[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X85 a_405_918# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X86 a_2889_66# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X87 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X88 VGND D[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X89 a_142_599# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X90 a_1313_297# a_1755_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X91 VPWR D[0] a_355_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X92 Z a_4239_793# a_3797_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X93 VPWR D[6] a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X94 VPWR D[5] a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X95 VPWR D[2] a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X96 Z S[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X97 VPWR S[1] a_142_599# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X98 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X99 Z a_1755_265# a_1313_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X100 Z S[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X101 a_142_325# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X102 VGND D[0] a_405_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X103 a_4239_265# S[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X104 a_405_918# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X105 VGND D[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X106 VGND D[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X107 Z S[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X108 a_1755_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X109 a_2839_613# D[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X110 a_3797_297# a_4239_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X111 a_1315_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X112 VGND D[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X113 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X114 Z a_2626_599# a_2839_613# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X115 a_405_66# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X116 a_3797_591# D[7] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X117 a_1315_911# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X118 a_1313_591# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X119 a_405_918# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X120 VPWR S[2] a_1755_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X121 VGND S[7] a_4239_793# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X122 a_2889_918# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X123 Z a_1755_793# a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X124 a_2889_66# S[4] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X125 a_2889_918# S[5] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X126 VPWR D[3] a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X127 a_4239_265# S[6] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X128 a_2839_311# a_2626_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X129 a_2889_918# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X130 VGND D[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X131 VGND D[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X132 a_1755_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X133 a_1315_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X134 VGND D[2] a_1315_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X135 a_1313_591# a_1755_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X136 Z S[3] a_1315_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X137 a_2889_66# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X138 Z S[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X139 Z S[7] a_3799_911# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X140 Z S[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X141 VGND S[4] a_2626_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X142 VPWR D[4] a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X143 Z a_2626_325# a_2839_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X144 a_4239_793# S[7] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X145 VGND D[1] a_405_918# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X146 VPWR S[4] a_2626_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X147 Z a_1755_793# a_1313_591# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X148 Z S[4] a_2889_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X149 Z S[6] a_3799_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X150 a_3799_47# D[6] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X151 a_2839_311# D[4] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X152 a_2626_599# S[5] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X153 VGND S[6] a_4239_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X154 Z a_4239_265# a_3797_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X155 a_2889_918# D[5] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X156 a_3797_591# a_4239_793# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X157 Z S[5] a_2889_918# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X158 a_3797_297# D[6] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X159 a_2889_66# D[4] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
