* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
X0 VPWR B1 a_228_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VGND A2 a_230_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_27_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 a_230_47# B2 a_124_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_124_47# B1 a_230_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_27_297# C1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND a_27_297# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_297# A2 a_515_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_230_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_515_297# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 a_27_297# C1 a_124_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 a_228_297# B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
