* NGSPICE file created from sky130_fd_sc_hdll__o21ba_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
M1000 a_79_199# a_222_93# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=3e+11p pd=2.6e+06u as=9.257e+11p ps=7.95e+06u
M1001 a_222_93# B1_N VPWR VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1002 a_222_93# B1_N VGND VNB nshort w=420000u l=150000u
+  ad=1.302e+11p pd=1.46e+06u as=3.76e+11p ps=3.81e+06u
M1003 a_460_47# A1 VGND VNB nshort w=650000u l=150000u
+  ad=4.29e+11p pd=3.92e+06u as=0p ps=0u
M1004 VGND A2 a_460_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR a_79_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.7e+11p ps=2.54e+06u
M1006 VPWR A1 a_554_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1007 VGND a_79_199# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.69e+11p ps=1.82e+06u
M1008 a_554_297# A2 a_79_199# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_460_47# a_222_93# a_79_199# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.95e+11p ps=1.9e+06u
.ends

