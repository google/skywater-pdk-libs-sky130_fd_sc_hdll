* File: sky130_fd_sc_hdll__a211oi_2.spice
* Created: Thu Aug 27 18:51:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a211oi_2.pex.spice"
.subckt sky130_fd_sc_hdll__a211oi_2  VNB VPB C1 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1012 N_Y_M1012_d N_C1_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.20475 PD=0.98 PS=1.93 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1012_d N_C1_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.091 PD=0.98 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B1_M1001_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.091 PD=1.03 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1001_d N_B1_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.17225 PD=1.03 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_525_47#_M1002_d N_A1_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.17225 AS=0.1235 PD=1.83 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1007 N_A_525_47#_M1007_d N_A1_M1007_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.1235 PD=0.93 PS=1.03 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75000.7
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g N_A_525_47#_M1007_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.091 PD=1.03 PS=0.93 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1010 N_VGND_M1009_d N_A2_M1010_g N_A_525_47#_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.17225 PD=1.03 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_C1_M1004_g N_A_37_297#_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 N_Y_M1004_d N_C1_M1011_g N_A_37_297#_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1005 N_A_320_297#_M1005_d N_B1_M1005_g N_A_37_297#_M1011_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90001.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1013 N_A_320_297#_M1005_d N_B1_M1013_g N_A_37_297#_M1013_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1003 N_A_320_297#_M1003_d N_A1_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.275 PD=1.3 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1015 N_A_320_297#_M1003_d N_A1_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1015_s N_A2_M1000_g N_A_320_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A2_M1008_g N_A_320_297#_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX16_noxref VNB VPB NWDIODE A=8.7312 P=14.09
pX17_noxref noxref_13 B1 B1 PROBETYPE=1
pX18_noxref noxref_14 A1 A1 PROBETYPE=1
pX19_noxref noxref_15 A2 A2 PROBETYPE=1
c_38 VNB 0 1.83161e-19 $X=0.125 $Y=-0.085
*
.include "sky130_fd_sc_hdll__a211oi_2.pxi.spice"
*
.ends
*
*
