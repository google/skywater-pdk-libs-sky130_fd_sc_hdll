* NGSPICE file created from sky130_fd_sc_hdll__a32o_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
M1000 X a_21_199# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=1.01e+12p ps=8.02e+06u
M1001 VGND a_21_199# X VNB nshort w=650000u l=150000u
+  ad=8.5475e+11p pd=6.53e+06u as=2.08e+11p ps=1.94e+06u
M1002 VPWR A1 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.5e+11p ps=7.7e+06u
M1003 VPWR a_21_199# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_21_199# B1 a_382_47# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=2.3075e+11p ps=2.01e+06u
M1005 a_319_297# B1 a_21_199# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=2.9e+11p ps=2.58e+06u
M1006 VPWR A3 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_589_47# A1 a_21_199# VNB nshort w=650000u l=150000u
+  ad=3.445e+11p pd=2.36e+06u as=0p ps=0u
M1008 a_21_199# B2 a_319_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 X a_21_199# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1010 a_725_47# A2 a_589_47# VNB nshort w=650000u l=150000u
+  ad=1.755e+11p pd=1.84e+06u as=0p ps=0u
M1011 a_319_297# A2 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_382_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 VGND A3 a_725_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

