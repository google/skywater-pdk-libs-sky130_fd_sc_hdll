* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
X0 a_27_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X1 VGND a_184_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 VPWR a_27_47# a_184_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 VPWR a_184_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VGND a_184_21# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_184_21# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND A_N a_912_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 VPWR A_N a_912_21# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X8 VGND D a_606_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_836_47# a_912_21# a_184_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 X a_184_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 VPWR a_184_21# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_27_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 a_719_47# a_27_47# a_836_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 X a_184_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 X a_184_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 VPWR D a_184_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 X a_184_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 a_184_21# a_912_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_606_47# C a_719_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
