* File: sky130_fd_sc_hdll__or3_2.spice
* Created: Wed Sep  2 08:48:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or3_2.pex.spice"
.subckt sky130_fd_sc_hdll__or3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C_M1008_g N_A_30_53#_M1008_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.1302 PD=0.74 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.3 A=0.063 P=1.14 MULT=1
MM1004 N_A_30_53#_M1004_d N_B_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0672 AS=0.0672 PD=0.74 PS=0.74 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.7
+ SB=75001.9 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_30_53#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.128453 AS=0.0672 PD=0.926355 PS=0.74 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1000 N_VGND_M1002_d N_A_30_53#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.198797 AS=0.12025 PD=1.43364 PS=1.02 NRD=37.836 NRS=8.304 M=1 R=4.33333
+ SA=75001.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_30_53#_M1007_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.18525 AS=0.12025 PD=1.87 PS=1.02 NRD=3.684 NRS=8.304 M=1 R=4.33333
+ SA=75001.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 A_120_297# N_C_M1001_g N_A_30_53#_M1001_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0483 AS=0.1134 PD=0.65 PS=1.38 NRD=28.1316 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.4 A=0.0756 P=1.2 MULT=1
MM1009 A_202_297# N_B_M1009_g A_120_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0735
+ AS=0.0483 PD=0.77 PS=0.65 NRD=56.2829 NRS=28.1316 M=1 R=2.33333 SA=90000.6
+ SB=90002 A=0.0756 P=1.2 MULT=1
MM1006 N_VPWR_M1006_d N_A_M1006_g A_202_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.148094 AS=0.0735 PD=0.916901 PS=0.77 NRD=139.575 NRS=56.2829 M=1
+ R=2.33333 SA=90001.1 SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1003 N_VPWR_M1006_d N_A_30_53#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.352606 AS=0.145 PD=2.1831 PS=1.29 NRD=39.4 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_A_30_53#_M1005_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.325 AS=0.145 PD=2.65 PS=1.29 NRD=5.91 NRS=0.9653 M=1 R=5.55556 SA=90001.5
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
c_58 VPB 0 8.49032e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__or3_2.pxi.spice"
*
.ends
*
*
