* File: sky130_fd_sc_hdll__inv_4.pxi.spice
* Created: Wed Sep  2 08:33:11 2020
* 
x_PM_SKY130_FD_SC_HDLL__INV_4%A N_A_c_51_n N_A_M1000_g N_A_c_44_n N_A_M1002_g
+ N_A_c_52_n N_A_M1001_g N_A_c_45_n N_A_M1003_g N_A_c_53_n N_A_M1004_g
+ N_A_c_46_n N_A_M1005_g N_A_c_54_n N_A_M1007_g N_A_c_47_n N_A_M1006_g A A A A
+ N_A_c_48_n N_A_c_49_n N_A_c_50_n A A A PM_SKY130_FD_SC_HDLL__INV_4%A
x_PM_SKY130_FD_SC_HDLL__INV_4%VPWR N_VPWR_M1000_d N_VPWR_M1001_d N_VPWR_M1007_d
+ N_VPWR_c_123_n N_VPWR_c_124_n N_VPWR_c_125_n N_VPWR_c_126_n N_VPWR_c_127_n
+ N_VPWR_c_128_n N_VPWR_c_129_n N_VPWR_c_130_n VPWR N_VPWR_c_131_n
+ N_VPWR_c_122_n PM_SKY130_FD_SC_HDLL__INV_4%VPWR
x_PM_SKY130_FD_SC_HDLL__INV_4%Y N_Y_M1002_d N_Y_M1005_d N_Y_M1000_s N_Y_M1004_s
+ N_Y_c_172_n N_Y_c_173_n N_Y_c_177_n N_Y_c_164_n N_Y_c_165_n N_Y_c_187_n
+ N_Y_c_191_n N_Y_c_193_n N_Y_c_166_n N_Y_c_197_n N_Y_c_167_n N_Y_c_201_n Y Y Y
+ N_Y_c_169_n N_Y_c_171_n PM_SKY130_FD_SC_HDLL__INV_4%Y
x_PM_SKY130_FD_SC_HDLL__INV_4%VGND N_VGND_M1002_s N_VGND_M1003_s N_VGND_M1006_s
+ N_VGND_c_246_n N_VGND_c_247_n N_VGND_c_248_n N_VGND_c_249_n N_VGND_c_250_n
+ N_VGND_c_251_n N_VGND_c_252_n N_VGND_c_253_n VGND N_VGND_c_254_n
+ N_VGND_c_255_n PM_SKY130_FD_SC_HDLL__INV_4%VGND
cc_1 VNB N_A_c_44_n 0.0223575f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=0.995
cc_2 VNB N_A_c_45_n 0.0167673f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=0.995
cc_3 VNB N_A_c_46_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=0.995
cc_4 VNB N_A_c_47_n 0.01997f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=0.995
cc_5 VNB N_A_c_48_n 0.0338038f $X=-0.19 $Y=-0.24 $X2=0.445 $Y2=1.16
cc_6 VNB N_A_c_49_n 0.00932659f $X=-0.19 $Y=-0.24 $X2=1.72 $Y2=1.16
cc_7 VNB N_A_c_50_n 0.0746087f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.202
cc_8 VNB N_VPWR_c_122_n 0.117919f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=1.202
cc_9 VNB N_Y_c_164_n 0.00264748f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.985
cc_10 VNB N_Y_c_165_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=0.995
cc_11 VNB N_Y_c_166_n 0.00512972f $X=-0.19 $Y=-0.24 $X2=0.445 $Y2=1.16
cc_12 VNB N_Y_c_167_n 0.00232612f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.202
cc_13 VNB Y 0.0227262f $X=-0.19 $Y=-0.24 $X2=1.485 $Y2=1.202
cc_14 VNB N_Y_c_169_n 0.00970162f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_246_n 0.0114137f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=0.995
cc_16 VNB N_VGND_c_247_n 0.0175755f $X=-0.19 $Y=-0.24 $X2=1.04 $Y2=0.56
cc_17 VNB N_VGND_c_248_n 0.00468437f $X=-0.19 $Y=-0.24 $X2=1.51 $Y2=0.995
cc_18 VNB N_VGND_c_249_n 0.00518111f $X=-0.19 $Y=-0.24 $X2=1.955 $Y2=1.985
cc_19 VNB N_VGND_c_250_n 0.0199148f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=0.56
cc_20 VNB N_VGND_c_251_n 0.00323937f $X=-0.19 $Y=-0.24 $X2=1.98 $Y2=0.56
cc_21 VNB N_VGND_c_252_n 0.0192745f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.105
cc_22 VNB N_VGND_c_253_n 0.00478105f $X=-0.19 $Y=-0.24 $X2=1.055 $Y2=1.105
cc_23 VNB N_VGND_c_254_n 0.0138819f $X=-0.19 $Y=-0.24 $X2=0.545 $Y2=1.202
cc_24 VNB N_VGND_c_255_n 0.163897f $X=-0.19 $Y=-0.24 $X2=0.57 $Y2=1.202
cc_25 VPB N_A_c_51_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.545 $Y2=1.41
cc_26 VPB N_A_c_52_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.41
cc_27 VPB N_A_c_53_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.41
cc_28 VPB N_A_c_54_n 0.0194435f $X=-0.19 $Y=1.305 $X2=1.955 $Y2=1.41
cc_29 VPB N_A_c_48_n 0.0114928f $X=-0.19 $Y=1.305 $X2=0.445 $Y2=1.16
cc_30 VPB N_A_c_49_n 7.73822e-19 $X=-0.19 $Y=1.305 $X2=1.72 $Y2=1.16
cc_31 VPB N_A_c_50_n 0.0488711f $X=-0.19 $Y=1.305 $X2=1.955 $Y2=1.202
cc_32 VPB N_VPWR_c_123_n 0.0114158f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=0.995
cc_33 VPB N_VPWR_c_124_n 0.0433254f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=0.56
cc_34 VPB N_VPWR_c_125_n 0.00469739f $X=-0.19 $Y=1.305 $X2=1.51 $Y2=0.56
cc_35 VPB N_VPWR_c_126_n 0.00496839f $X=-0.19 $Y=1.305 $X2=1.98 $Y2=0.995
cc_36 VPB N_VPWR_c_127_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_37 VPB N_VPWR_c_128_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.105
cc_38 VPB N_VPWR_c_129_n 0.0206409f $X=-0.19 $Y=1.305 $X2=1.52 $Y2=1.105
cc_39 VPB N_VPWR_c_130_n 0.00401177f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_131_n 0.0163041f $X=-0.19 $Y=1.305 $X2=1.015 $Y2=1.202
cc_41 VPB N_VPWR_c_122_n 0.0490348f $X=-0.19 $Y=1.305 $X2=1.04 $Y2=1.202
cc_42 VPB Y 0.0107733f $X=-0.19 $Y=1.305 $X2=1.485 $Y2=1.202
cc_43 VPB N_Y_c_171_n 0.0127118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 N_A_c_51_n N_VPWR_c_124_n 0.00781009f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_45 N_A_c_48_n N_VPWR_c_124_n 0.00612676f $X=0.445 $Y=1.16 $X2=0 $Y2=0
cc_46 N_A_c_49_n N_VPWR_c_124_n 0.0214003f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A_c_52_n N_VPWR_c_125_n 0.0052072f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_48 N_A_c_53_n N_VPWR_c_125_n 0.004751f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_49 N_A_c_54_n N_VPWR_c_126_n 0.00583244f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A_c_51_n N_VPWR_c_127_n 0.00597712f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A_c_52_n N_VPWR_c_127_n 0.00673617f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_c_53_n N_VPWR_c_129_n 0.00597712f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A_c_54_n N_VPWR_c_129_n 0.00673617f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_54 N_A_c_51_n N_VPWR_c_122_n 0.0109493f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_55 N_A_c_52_n N_VPWR_c_122_n 0.0118438f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A_c_53_n N_VPWR_c_122_n 0.00999457f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A_c_54_n N_VPWR_c_122_n 0.0129427f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_58 N_A_c_44_n N_Y_c_172_n 0.0147385f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_59 N_A_c_51_n N_Y_c_173_n 0.00347232f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A_c_52_n N_Y_c_173_n 5.79575e-19 $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_61 N_A_c_49_n N_Y_c_173_n 0.0253353f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_62 N_A_c_50_n N_Y_c_173_n 0.00651614f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_63 N_A_c_51_n N_Y_c_177_n 0.0121679f $X=0.545 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A_c_52_n N_Y_c_177_n 0.0106248f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A_c_53_n N_Y_c_177_n 6.24653e-19 $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A_c_45_n N_Y_c_164_n 0.0131218f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A_c_46_n N_Y_c_164_n 0.00622594f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A_c_49_n N_Y_c_164_n 0.0404964f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_69 N_A_c_50_n N_Y_c_164_n 0.00345541f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_70 N_A_c_44_n N_Y_c_165_n 0.0128243f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A_c_49_n N_Y_c_165_n 0.030974f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A_c_50_n N_Y_c_165_n 0.00358305f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_73 N_A_c_52_n N_Y_c_187_n 0.0137916f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_74 N_A_c_53_n N_Y_c_187_n 0.0101048f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_c_49_n N_Y_c_187_n 0.0356113f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_76 N_A_c_50_n N_Y_c_187_n 0.00635951f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_77 N_A_c_45_n N_Y_c_191_n 6.12918e-19 $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_c_46_n N_Y_c_191_n 0.00982965f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_79 N_A_c_52_n N_Y_c_193_n 5.84907e-19 $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_80 N_A_c_53_n N_Y_c_193_n 0.0126343f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_c_54_n N_Y_c_193_n 0.0252512f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_c_47_n N_Y_c_166_n 0.0167901f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_c_54_n N_Y_c_197_n 0.018541f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_c_46_n N_Y_c_167_n 0.00489926f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_c_49_n N_Y_c_167_n 0.030974f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_c_50_n N_Y_c_167_n 0.00358305f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_87 N_A_c_53_n N_Y_c_201_n 0.00254223f $X=1.485 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_c_54_n N_Y_c_201_n 6.15357e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_c_49_n N_Y_c_201_n 0.0253353f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_90 N_A_c_50_n N_Y_c_201_n 0.00651614f $X=1.955 $Y=1.202 $X2=0 $Y2=0
cc_91 N_A_c_54_n Y 0.00255978f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A_c_47_n Y 0.0144736f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_c_49_n Y 0.00892144f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_c_44_n N_VGND_c_247_n 0.00530388f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_c_48_n N_VGND_c_247_n 0.00524994f $X=0.445 $Y=1.16 $X2=0 $Y2=0
cc_96 N_A_c_49_n N_VGND_c_247_n 0.00883493f $X=1.72 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A_c_45_n N_VGND_c_248_n 0.00276126f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_98 N_A_c_46_n N_VGND_c_248_n 0.0035663f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A_c_47_n N_VGND_c_249_n 0.0044954f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_c_44_n N_VGND_c_250_n 0.00465454f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_45_n N_VGND_c_250_n 0.00437852f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_c_46_n N_VGND_c_252_n 0.00396605f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_103 N_A_c_47_n N_VGND_c_252_n 0.00437852f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A_c_44_n N_VGND_c_255_n 0.00893928f $X=0.57 $Y=0.995 $X2=0 $Y2=0
cc_105 N_A_c_45_n N_VGND_c_255_n 0.00614065f $X=1.04 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_c_46_n N_VGND_c_255_n 0.00581484f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_c_47_n N_VGND_c_255_n 0.00716112f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_108 N_VPWR_c_122_n N_Y_M1000_s 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_109 N_VPWR_c_122_n N_Y_M1004_s 0.00231261f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_110 N_VPWR_c_124_n N_Y_c_173_n 0.0137878f $X=0.31 $Y=1.66 $X2=0 $Y2=0
cc_111 N_VPWR_c_124_n N_Y_c_177_n 0.0616825f $X=0.31 $Y=1.66 $X2=0 $Y2=0
cc_112 N_VPWR_c_125_n N_Y_c_177_n 0.0385613f $X=1.25 $Y=2 $X2=0 $Y2=0
cc_113 N_VPWR_c_127_n N_Y_c_177_n 0.0223557f $X=1.165 $Y=2.72 $X2=0 $Y2=0
cc_114 N_VPWR_c_122_n N_Y_c_177_n 0.0140101f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_M1001_d N_Y_c_187_n 0.00325884f $X=1.105 $Y=1.485 $X2=0 $Y2=0
cc_116 N_VPWR_c_125_n N_Y_c_187_n 0.0136682f $X=1.25 $Y=2 $X2=0 $Y2=0
cc_117 N_VPWR_c_125_n N_Y_c_193_n 0.0470327f $X=1.25 $Y=2 $X2=0 $Y2=0
cc_118 N_VPWR_c_126_n N_Y_c_193_n 0.0180305f $X=2.19 $Y=2.34 $X2=0 $Y2=0
cc_119 N_VPWR_c_129_n N_Y_c_193_n 0.0223557f $X=2.105 $Y=2.72 $X2=0 $Y2=0
cc_120 N_VPWR_c_122_n N_Y_c_193_n 0.0140101f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_121 N_VPWR_M1007_d N_Y_c_197_n 0.0139845f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_122 N_VPWR_c_126_n N_Y_c_197_n 0.00771958f $X=2.19 $Y=2.34 $X2=0 $Y2=0
cc_123 N_VPWR_M1007_d Y 2.09721e-19 $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_124 N_VPWR_M1007_d N_Y_c_171_n 0.00913336f $X=2.045 $Y=1.485 $X2=0 $Y2=0
cc_125 N_Y_c_164_n N_VGND_M1003_s 0.00255004f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_126 N_Y_c_166_n N_VGND_M1006_s 0.0046937f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_127 N_Y_c_169_n N_VGND_M1006_s 0.00478655f $X=2.53 $Y=0.905 $X2=0 $Y2=0
cc_128 N_Y_c_172_n N_VGND_c_247_n 0.0223739f $X=0.78 $Y=0.42 $X2=0 $Y2=0
cc_129 N_Y_c_164_n N_VGND_c_248_n 0.0121134f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_130 N_Y_c_191_n N_VGND_c_248_n 0.0216501f $X=1.72 $Y=0.42 $X2=0 $Y2=0
cc_131 N_Y_c_166_n N_VGND_c_249_n 0.0185426f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_132 N_Y_c_172_n N_VGND_c_250_n 0.023074f $X=0.78 $Y=0.42 $X2=0 $Y2=0
cc_133 N_Y_c_164_n N_VGND_c_250_n 0.00255089f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_134 N_Y_c_164_n N_VGND_c_252_n 0.00199443f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_135 N_Y_c_191_n N_VGND_c_252_n 0.023074f $X=1.72 $Y=0.42 $X2=0 $Y2=0
cc_136 N_Y_c_166_n N_VGND_c_252_n 0.00255089f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_137 N_Y_c_166_n N_VGND_c_254_n 5.66972e-19 $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_138 N_Y_c_169_n N_VGND_c_254_n 0.00443753f $X=2.53 $Y=0.905 $X2=0 $Y2=0
cc_139 N_Y_M1002_d N_VGND_c_255_n 0.00263993f $X=0.645 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_M1005_d N_VGND_c_255_n 0.00263993f $X=1.585 $Y=0.235 $X2=0 $Y2=0
cc_141 N_Y_c_172_n N_VGND_c_255_n 0.0141066f $X=0.78 $Y=0.42 $X2=0 $Y2=0
cc_142 N_Y_c_164_n N_VGND_c_255_n 0.0098008f $X=1.505 $Y=0.815 $X2=0 $Y2=0
cc_143 N_Y_c_191_n N_VGND_c_255_n 0.0141066f $X=1.72 $Y=0.42 $X2=0 $Y2=0
cc_144 N_Y_c_166_n N_VGND_c_255_n 0.00704533f $X=2.395 $Y=0.815 $X2=0 $Y2=0
cc_145 N_Y_c_169_n N_VGND_c_255_n 0.00760176f $X=2.53 $Y=0.905 $X2=0 $Y2=0
