* File: sky130_fd_sc_hdll__mux2_8.spice
* Created: Thu Aug 27 19:10:54 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2_8.pex.spice"
.subckt sky130_fd_sc_hdll__mux2_8  VNB VPB S A1 A0 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A0	A0
* A1	A1
* S	S
* VPB	VPB
* VNB	VNB
MM1006 N_X_M1006_d N_A_79_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75009.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1006_d N_A_79_21#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75009.2 A=0.0975 P=1.6 MULT=1
MM1010 N_X_M1010_d N_A_79_21#_M1010_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.1
+ SB=75008.8 A=0.0975 P=1.6 MULT=1
MM1020 N_X_M1010_d N_A_79_21#_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.6
+ SB=75008.3 A=0.0975 P=1.6 MULT=1
MM1026 N_X_M1026_d N_A_79_21#_M1026_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75007.8 A=0.0975 P=1.6 MULT=1
MM1027 N_X_M1026_d N_A_79_21#_M1027_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.5
+ SB=75007.4 A=0.0975 P=1.6 MULT=1
MM1029 N_X_M1029_d N_A_79_21#_M1029_g N_VGND_M1027_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003
+ SB=75006.9 A=0.0975 P=1.6 MULT=1
MM1030 N_X_M1029_d N_A_79_21#_M1030_g N_VGND_M1030_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.106066 PD=1.02 PS=0.982558 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75003.5 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1030_s N_S_M1007_g N_A_872_47#_M1007_s VNB NSHORT L=0.15 W=0.64
+ AD=0.104434 AS=0.0944 PD=0.967442 PS=0.935 NRD=9.372 NRS=3.744 M=1 R=4.26667
+ SA=75004 SB=75006 A=0.096 P=1.58 MULT=1
MM1003 N_A_79_21#_M1003_d N_A1_M1003_g N_A_872_47#_M1007_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.0944 PD=0.91 PS=0.935 NRD=0 NRS=0 M=1 R=4.26667
+ SA=75004.4 SB=75005.5 A=0.096 P=1.58 MULT=1
MM1005 N_A_79_21#_M1003_d N_A1_M1005_g N_A_872_47#_M1005_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0864 AS=0.384 PD=0.91 PS=1.84 NRD=0 NRS=0 M=1 R=4.26667 SA=75004.9
+ SB=75005.1 A=0.096 P=1.58 MULT=1
MM1023 N_VGND_M1023_d N_S_M1023_g N_A_872_47#_M1005_s VNB NSHORT L=0.15 W=0.64
+ AD=0.1232 AS=0.384 PD=1.025 PS=1.84 NRD=20.616 NRS=173.436 M=1 R=4.26667
+ SA=75006.2 SB=75003.8 A=0.096 P=1.58 MULT=1
MM1011 N_VGND_M1023_d N_A_1369_199#_M1011_g N_A_1422_47#_M1011_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.1232 AS=0.1552 PD=1.025 PS=1.125 NRD=0 NRS=16.872 M=1
+ R=4.26667 SA=75006.8 SB=75003.2 A=0.096 P=1.58 MULT=1
MM1017 N_A_79_21#_M1017_d N_A0_M1017_g N_A_1422_47#_M1011_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1184 AS=0.1552 PD=1.01 PS=1.125 NRD=8.436 NRS=21.552 M=1 R=4.26667
+ SA=75007.4 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1031 N_A_79_21#_M1017_d N_A0_M1031_g N_A_1422_47#_M1031_s VNB NSHORT L=0.15
+ W=0.64 AD=0.1184 AS=0.368 PD=1.01 PS=1.79 NRD=8.436 NRS=0 M=1 R=4.26667
+ SA=75007.9 SB=75002.1 A=0.096 P=1.58 MULT=1
MM1025 N_VGND_M1025_d N_A_1369_199#_M1025_g N_A_1422_47#_M1031_s VNB NSHORT
+ L=0.15 W=0.64 AD=0.128248 AS=0.368 PD=1.04186 PS=1.79 NRD=23.436 NRS=164.052
+ M=1 R=4.26667 SA=75009.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1032 N_A_1369_199#_M1032_d N_S_M1032_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.130252 PD=1.92 PS=1.05814 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75009.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90009.7 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_79_21#_M1001_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90009.3 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1001_d N_A_79_21#_M1004_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90008.8 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1008_d N_A_79_21#_M1008_g N_X_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90008.3 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1008_d N_A_79_21#_M1014_g N_X_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90007.9 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_79_21#_M1018_g N_X_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.5 SB=90007.4 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1018_d N_A_79_21#_M1021_g N_X_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90006.9 A=0.18 P=2.36 MULT=1
MM1028 N_VPWR_M1028_d N_A_79_21#_M1028_g N_X_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1475 AS=0.145 PD=1.295 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003.5 SB=90006.5 A=0.18 P=2.36 MULT=1
MM1022 N_A_870_297#_M1022_d N_S_M1022_g N_VPWR_M1028_d VPB PHIGHVT L=0.18 W=1
+ AD=0.5475 AS=0.1475 PD=2.095 PS=1.295 NRD=60.0653 NRS=1.9503 M=1 R=5.55556
+ SA=90003.9 SB=90006 A=0.18 P=2.36 MULT=1
MM1002 N_A_870_297#_M1022_d N_A0_M1002_g N_A_79_21#_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.5475 AS=0.145 PD=2.095 PS=1.29 NRD=100.45 NRS=0.9653 M=1 R=5.55556
+ SA=90005.2 SB=90004.7 A=0.18 P=2.36 MULT=1
MM1012 N_A_870_297#_M1012_d N_A0_M1012_g N_A_79_21#_M1002_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.7 SB=90004.2 A=0.18 P=2.36 MULT=1
MM1033 N_A_870_297#_M1012_d N_S_M1033_g N_VPWR_M1033_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1775 PD=1.29 PS=1.355 NRD=0.9653 NRS=10.8153 M=1 R=5.55556
+ SA=90006.2 SB=90003.8 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1033_s N_A_1369_199#_M1013_g N_A_1420_297#_M1013_s VPB PHIGHVT
+ L=0.18 W=1 AD=0.1775 AS=0.6925 PD=1.355 PS=2.385 NRD=3.9203 NRS=0.9653 M=1
+ R=5.55556 SA=90006.7 SB=90003.2 A=0.18 P=2.36 MULT=1
MM1016 N_A_1420_297#_M1013_s N_A1_M1016_g N_A_79_21#_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.6925 AS=0.145 PD=2.385 PS=1.29 NRD=216.68 NRS=0.9653 M=1 R=5.55556
+ SA=90008.3 SB=90001.7 A=0.18 P=2.36 MULT=1
MM1024 N_A_1420_297#_M1024_d N_A1_M1024_g N_A_79_21#_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90008.7 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_1369_199#_M1015_g N_A_1420_297#_M1024_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.185 AS=0.145 PD=1.37 PS=1.29 NRD=16.7253 NRS=0.9653 M=1
+ R=5.55556 SA=90009.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_A_1369_199#_M1019_d N_S_M1019_g N_VPWR_M1015_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.185 PD=2.54 PS=1.37 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90009.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX34_noxref VNB VPB NWDIODE A=17.5908 P=25.13
*
.include "sky130_fd_sc_hdll__mux2_8.pxi.spice"
*
.ends
*
*
