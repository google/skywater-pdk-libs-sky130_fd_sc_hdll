* File: sky130_fd_sc_hdll__o22ai_1.spice
* Created: Wed Sep  2 08:45:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o22ai_1  VNB VPB B1 B2 A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1005 N_Y_M1005_d N_B1_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128375 AS=0.2015 PD=1.045 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1003 N_A_27_47#_M1003_d N_B2_M1003_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.128375 PD=1.19 PS=1.045 NRD=32.304 NRS=22.152 M=1 R=4.33333
+ SA=75000.8 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1000_d N_A2_M1000_g N_A_27_47#_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.1755 PD=0.96 PS=1.19 NRD=0.912 NRS=15.684 M=1 R=4.33333
+ SA=75001.5 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_27_47#_M1006_d N_A1_M1006_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.208 AS=0.10075 PD=1.94 PS=0.96 NRD=10.152 NRS=4.608 M=1 R=4.33333
+ SA=75001.9 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1004 A_117_297# N_B1_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1 AD=0.2075
+ AS=0.27 PD=1.415 PS=2.54 NRD=30.0228 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.9 A=0.18 P=2.36 MULT=1
MM1007 N_Y_M1007_d N_B2_M1007_g A_117_297# VPB PHIGHVT L=0.18 W=1 AD=0.28
+ AS=0.2075 PD=1.56 PS=1.415 NRD=15.7403 NRS=30.0228 M=1 R=5.55556 SA=90000.8
+ SB=90001.3 A=0.18 P=2.36 MULT=1
MM1002 A_384_297# N_A2_M1002_g N_Y_M1007_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.28 PD=1.23 PS=1.56 NRD=11.8003 NRS=39.4 M=1 R=5.55556 SA=90001.5
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g A_384_297# VPB PHIGHVT L=0.18 W=1 AD=0.28
+ AS=0.115 PD=2.56 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90001.9
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.0397 P=9.49
pX9_noxref noxref_13 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o22ai_1.pxi.spice"
*
.ends
*
*
