* File: sky130_fd_sc_hdll__ebufn_1.spice
* Created: Wed Sep  2 08:30:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__ebufn_1.pex.spice"
.subckt sky130_fd_sc_hdll__ebufn_1  VNB VPB A TE_B VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* TE_B	TE_B
* A	A
* VPB	VPB
* VNB	VNB
MM1005 N_VGND_M1005_d N_A_M1005_g N_A_27_47#_M1005_s VNB NSHORT L=0.15 W=0.42
+ AD=0.098125 AS=0.1302 PD=1.005 PS=1.46 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1006 N_A_211_369#_M1006_d N_TE_B_M1006_g N_VGND_M1005_d VNB NSHORT L=0.15
+ W=0.42 AD=0.2814 AS=0.098125 PD=2.18 PS=1.005 NRD=109.992 NRS=51.036 M=1 R=2.8
+ SA=75000.4 SB=75000.6 A=0.063 P=1.14 MULT=1
MM1002 A_543_47# N_A_211_369#_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.06825 AS=0.169 PD=0.86 PS=1.82 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1000 N_Z_M1000_d N_A_27_47#_M1000_g A_543_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.3055 AS=0.06825 PD=2.24 PS=0.86 NRD=37.836 NRS=9.228 M=1 R=4.33333
+ SA=75000.5 SB=75000.4 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_A_27_47#_M1001_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0928 AS=0.1728 PD=0.93 PS=1.82 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90000.6 A=0.1152 P=1.64 MULT=1
MM1007 N_A_211_369#_M1007_d N_TE_B_M1007_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.1728 AS=0.0928 PD=1.82 PS=0.93 NRD=1.5366 NRS=1.5366 M=1 R=3.55556
+ SA=90000.6 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1003 A_411_297# N_TE_B_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.44
+ AS=0.28 PD=1.88 PS=2.56 NRD=75.8253 NRS=2.9353 M=1 R=5.55556 SA=90000.2
+ SB=90001.4 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_27_47#_M1004_g A_411_297# VPB PHIGHVT L=0.18 W=1 AD=0.395
+ AS=0.44 PD=2.79 PS=1.88 NRD=25.5903 NRS=75.8253 M=1 R=5.55556 SA=90001.2
+ SB=90000.3 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__ebufn_1.pxi.spice"
*
.ends
*
*
