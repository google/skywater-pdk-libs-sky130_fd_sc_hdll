* File: sky130_fd_sc_hdll__o21bai_1.pex.spice
* Created: Wed Sep  2 08:44:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%B1_N 2 5 6 7 11 17 18 20 23
c41 11 0 3.08172e-19 $X=0.935 $Y=1.97
r42 18 24 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.475 $Y2=1.325
r43 18 23 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.475 $Y=1.16
+ $X2=0.475 $Y2=0.995
r44 17 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.45
+ $Y=1.16 $X2=0.45 $Y2=1.16
r45 14 20 8.35926 $w=2.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.22 $Y=1.345
+ $X2=0.22 $Y2=1.53
r46 13 17 7.5732 $w=3.48e-07 $l=2.3e-07 $layer=LI1_cond $X=0.22 $Y=1.17 $X2=0.45
+ $Y2=1.17
r47 13 14 2.25943 $w=2.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.22 $Y=1.17
+ $X2=0.22 $Y2=1.345
r48 8 11 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.935 $Y=1.685
+ $X2=0.935 $Y2=1.97
r49 6 8 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=0.845 $Y=1.61
+ $X2=0.935 $Y2=1.685
r50 6 7 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=0.845 $Y=1.61
+ $X2=0.635 $Y2=1.61
r51 5 23 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.56 $Y=0.675
+ $X2=0.56 $Y2=0.995
r52 2 7 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=0.535 $Y=1.535
+ $X2=0.635 $Y2=1.61
r53 2 24 69.6312 $w=2e-07 $l=2.1e-07 $layer=POLY_cond $X=0.535 $Y=1.535
+ $X2=0.535 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%A_105_352# 1 2 7 9 10 12 13 14 17 21 22
+ 24 31 34
c59 22 0 1.47323e-19 $X=0.917 $Y=1.535
c60 17 0 1.60849e-19 $X=0.7 $Y=1.96
r61 33 34 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=0.855 $Y=0.825
+ $X2=0.855 $Y2=0.995
r62 31 33 8.65224 $w=2.63e-07 $l=1.65e-07 $layer=LI1_cond $X=0.807 $Y=0.66
+ $X2=0.807 $Y2=0.825
r63 24 25 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.98
+ $Y=1.16 $X2=0.98 $Y2=1.16
r64 22 24 14.6497 $w=2.93e-07 $l=3.75e-07 $layer=LI1_cond $X=0.917 $Y=1.535
+ $X2=0.917 $Y2=1.16
r65 21 34 7.79447 $w=2.93e-07 $l=1.47e-07 $layer=LI1_cond $X=0.917 $Y=1.142
+ $X2=0.917 $Y2=0.995
r66 21 24 0.703186 $w=2.93e-07 $l=1.8e-08 $layer=LI1_cond $X=0.917 $Y=1.142
+ $X2=0.917 $Y2=1.16
r67 15 22 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=0.687 $Y=1.62
+ $X2=0.917 $Y2=1.62
r68 15 17 9.04224 $w=3.23e-07 $l=2.55e-07 $layer=LI1_cond $X=0.687 $Y=1.705
+ $X2=0.687 $Y2=1.96
r69 13 25 79.5619 $w=3.3e-07 $l=4.55e-07 $layer=POLY_cond $X=1.435 $Y=1.16
+ $X2=0.98 $Y2=1.16
r70 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.435 $Y=1.16
+ $X2=1.535 $Y2=1.202
r71 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.56 $Y=0.995
+ $X2=1.535 $Y2=1.202
r72 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.56 $Y=0.995
+ $X2=1.56 $Y2=0.56
r73 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.202
r74 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.985
r75 2 17 600 $w=1.7e-07 $l=2.73861e-07 $layer=licon1_PDIFF $count=1 $X=0.525
+ $Y=1.76 $X2=0.7 $Y2=1.96
r76 1 31 182 $w=1.7e-07 $l=2.55588e-07 $layer=licon1_NDIFF $count=1 $X=0.635
+ $Y=0.465 $X2=0.775 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%A2 1 3 4 6 7 15
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2 $Y=1.16
+ $X2=2 $Y2=1.16
r31 7 15 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=1.76 $Y=1.175 $X2=2
+ $Y2=1.175
r32 4 10 39.1718 $w=2.59e-07 $l=1.93959e-07 $layer=POLY_cond $X=2.06 $Y=0.995
+ $X2=1.997 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.06 $Y=0.995 $X2=2.06
+ $Y2=0.56
r34 1 10 51.0578 $w=2.59e-07 $l=2.68328e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=1.997 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.035 $Y=1.41
+ $X2=2.035 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%A1 1 3 4 6 7 14
r21 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.53
+ $Y=1.16 $X2=2.53 $Y2=1.16
r22 7 14 13.2035 $w=2.08e-07 $l=2.5e-07 $layer=LI1_cond $X=2.78 $Y=1.18 $X2=2.53
+ $Y2=1.18
r23 4 10 39.2931 $w=2.55e-07 $l=1.69926e-07 $layer=POLY_cond $X=2.54 $Y=0.995
+ $X2=2.53 $Y2=1.16
r24 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.54 $Y=0.995 $X2=2.54
+ $Y2=0.56
r25 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.53 $Y2=1.16
r26 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.495 $Y=1.41
+ $X2=2.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%VPWR 1 2 9 13 15 19 21 26 32 36
r33 36 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 35 38 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r35 35 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r36 32 33 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 30 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 30 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r39 29 30 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r40 27 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=2.72
+ $X2=1.235 $Y2=2.72
r41 27 29 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.4 $Y=2.72 $X2=1.61
+ $Y2=2.72
r42 26 35 6.92095 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=2.47 $Y=2.72
+ $X2=2.845 $Y2=2.72
r43 26 29 56.107 $w=1.68e-07 $l=8.6e-07 $layer=LI1_cond $X=2.47 $Y=2.72 $X2=1.61
+ $Y2=2.72
r44 21 32 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=1.235 $Y2=2.72
r45 21 23 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=1.07 $Y=2.72
+ $X2=0.23 $Y2=2.72
r46 19 33 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r47 19 23 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r48 15 18 13.7853 $w=5.88e-07 $l=6.8e-07 $layer=LI1_cond $X=2.765 $Y=1.62
+ $X2=2.765 $Y2=2.3
r49 13 35 3.04522 $w=5.9e-07 $l=1.18427e-07 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.845 $Y2=2.72
r50 13 18 6.79129 $w=5.88e-07 $l=3.35e-07 $layer=LI1_cond $X=2.765 $Y=2.635
+ $X2=2.765 $Y2=2.3
r51 9 12 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.235 $Y=1.96
+ $X2=1.235 $Y2=2.3
r52 7 32 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=2.635
+ $X2=1.235 $Y2=2.72
r53 7 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.235 $Y=2.635
+ $X2=1.235 $Y2=2.3
r54 2 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.485 $X2=2.73 $Y2=2.3
r55 2 15 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.585
+ $Y=1.485 $X2=2.73 $Y2=1.62
r56 1 12 600 $w=1.7e-07 $l=6.36396e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.76 $X2=1.235 $Y2=2.3
r57 1 9 600 $w=1.7e-07 $l=2.93428e-07 $layer=licon1_PDIFF $count=1 $X=1.025
+ $Y=1.76 $X2=1.235 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%Y 1 2 9 16 18
r32 18 24 2.07014 $w=5.18e-07 $l=9e-08 $layer=LI1_cond $X=1.895 $Y=2.21
+ $X2=1.895 $Y2=2.3
r33 16 18 13.4559 $w=5.18e-07 $l=5.85e-07 $layer=LI1_cond $X=1.895 $Y=1.625
+ $X2=1.895 $Y2=2.21
r34 14 16 5.85354 $w=1.78e-07 $l=9.5e-08 $layer=LI1_cond $X=1.8 $Y=1.535
+ $X2=1.895 $Y2=1.535
r35 7 14 28.0354 $w=1.78e-07 $l=4.55e-07 $layer=LI1_cond $X=1.345 $Y=1.535
+ $X2=1.8 $Y2=1.535
r36 7 9 47.1454 $w=2.18e-07 $l=9e-07 $layer=LI1_cond $X=1.345 $Y=1.445 $X2=1.345
+ $Y2=0.545
r37 2 24 400 $w=1.7e-07 $l=8.98248e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.485 $X2=1.8 $Y2=2.3
r38 2 14 400 $w=1.7e-07 $l=2.32916e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.485 $X2=1.8 $Y2=1.62
r39 1 9 182 $w=1.7e-07 $l=3.8775e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.35 $Y2=0.545
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%VGND 1 2 7 9 13 16 17 18 28 29
r37 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r38 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r39 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r40 23 26 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r41 22 25 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r42 22 23 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r43 20 32 4.29305 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.18
+ $Y2=0
r44 20 22 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=0.36 $Y=0 $X2=0.69
+ $Y2=0
r45 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r46 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r47 16 25 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.07
+ $Y2=0
r48 16 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=0 $X2=2.28
+ $Y2=0
r49 15 28 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.99
+ $Y2=0
r50 15 17 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.365 $Y=0 $X2=2.28
+ $Y2=0
r51 11 17 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0
r52 11 13 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.28 $Y=0.085
+ $X2=2.28 $Y2=0.39
r53 7 32 3.02899 $w=2.75e-07 $l=1.03899e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.18 $Y2=0
r54 7 9 24.0965 $w=2.73e-07 $l=5.75e-07 $layer=LI1_cond $X=0.222 $Y=0.085
+ $X2=0.222 $Y2=0.66
r55 2 13 182 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=1 $X=2.135
+ $Y=0.235 $X2=2.28 $Y2=0.39
r56 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21BAI_1%A_327_47# 1 2 9 11 12 15
r28 13 15 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.725 $Y=0.735
+ $X2=2.725 $Y2=0.39
r29 11 13 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=2.535 $Y=0.82
+ $X2=2.725 $Y2=0.735
r30 11 12 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=2.535 $Y=0.82
+ $X2=1.97 $Y2=0.82
r31 7 12 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=1.805 $Y=0.735
+ $X2=1.97 $Y2=0.82
r32 7 9 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=1.805 $Y=0.735
+ $X2=1.805 $Y2=0.4
r33 2 15 91 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=2 $X=2.615
+ $Y=0.235 $X2=2.75 $Y2=0.39
r34 1 9 91 $w=1.7e-07 $l=2.38642e-07 $layer=licon1_NDIFF $count=2 $X=1.635
+ $Y=0.235 $X2=1.805 $Y2=0.4
.ends

