* File: sky130_fd_sc_hdll__xnor3_2.spice
* Created: Wed Sep  2 08:54:07 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__xnor3_2.pex.spice"
.subckt sky130_fd_sc_hdll__xnor3_2  VNB VPB C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_79_21#_M1002_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75000.2
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1023 N_VGND_M1023_d N_A_79_21#_M1023_g N_X_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.157336 AS=0.12025 PD=1.30607 PS=1.02 NRD=6.456 NRS=4.608 M=1 R=4.33333
+ SA=75000.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_A_328_93#_M1009_d N_C_M1009_g N_VGND_M1023_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1995 AS=0.101664 PD=1.79 PS=0.843925 NRD=54.276 NRS=53.436 M=1 R=2.8
+ SA=75001.3 SB=75000.4 A=0.063 P=1.14 MULT=1
MM1007 N_A_79_21#_M1007_d N_C_M1007_g N_A_477_49#_M1007_s VNB NSHORT L=0.15
+ W=0.64 AD=0.0928 AS=0.2048 PD=0.93 PS=1.92 NRD=0.936 NRS=8.436 M=1 R=4.26667
+ SA=75000.2 SB=75000.8 A=0.096 P=1.58 MULT=1
MM1008 N_A_453_325#_M1008_d N_A_328_93#_M1008_g N_A_79_21#_M1007_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.256 AS=0.0928 PD=2.08 PS=0.93 NRD=21.552 NRS=0.936 M=1
+ R=4.26667 SA=75000.7 SB=75000.3 A=0.096 P=1.58 MULT=1
MM1022 N_A_885_297#_M1022_d N_B_M1022_g N_VGND_M1022_s VNB NSHORT L=0.15 W=0.65
+ AD=0.16515 AS=0.2535 PD=1.82 PS=2.08 NRD=0 NRS=17.532 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_A_453_325#_M1015_d N_B_M1015_g N_A_1003_297#_M1015_s VNB NSHORT L=0.15
+ W=0.64 AD=0.232513 AS=0.19475 PD=1.56377 PS=1.9 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75000.2 SB=75002.6 A=0.096 P=1.58 MULT=1
MM1001 N_A_1286_297#_M1001_d N_A_885_297#_M1001_g N_A_453_325#_M1015_d VNB
+ NSHORT L=0.15 W=0.42 AD=0.152666 AS=0.152587 PD=1.0183 PS=1.02623 NRD=88.14
+ NRS=108.564 M=1 R=2.8 SA=75001 SB=75002.9 A=0.063 P=1.14 MULT=1
MM1004 N_A_477_49#_M1004_d N_B_M1004_g N_A_1286_297#_M1001_d VNB NSHORT L=0.15
+ W=0.64 AD=0.175819 AS=0.232634 PD=1.23355 PS=1.5517 NRD=10.308 NRS=12.18 M=1
+ R=4.26667 SA=75001.4 SB=75002 A=0.096 P=1.58 MULT=1
MM1012 N_A_1003_297#_M1012_d N_A_885_297#_M1012_g N_A_477_49#_M1004_d VNB NSHORT
+ L=0.15 W=0.6 AD=0.123387 AS=0.164831 PD=1.01129 PS=1.15645 NRD=15.996
+ NRS=41.988 M=1 R=4 SA=75002.1 SB=75001.4 A=0.09 P=1.5 MULT=1
MM1021 N_VGND_M1021_d N_A_M1021_g N_A_1003_297#_M1012_d VNB NSHORT L=0.15 W=0.64
+ AD=0.0864 AS=0.131613 PD=0.91 PS=1.07871 NRD=0 NRS=8.436 M=1 R=4.26667
+ SA=75002.5 SB=75000.9 A=0.096 P=1.58 MULT=1
MM1020 N_A_1286_297#_M1020_d N_A_1003_297#_M1020_g N_VGND_M1021_d VNB NSHORT
+ L=0.15 W=0.64 AD=0.3296 AS=0.0864 PD=2.31 PS=0.91 NRD=42.18 NRS=0 M=1
+ R=4.26667 SA=75002.9 SB=75000.4 A=0.096 P=1.58 MULT=1
MM1013 N_X_M1013_d N_A_79_21#_M1013_g N_VPWR_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.27 PD=1.31 PS=2.54 NRD=4.9053 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1019 N_X_M1013_d N_A_79_21#_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.240488 PD=1.31 PS=1.7378 NRD=0.9653 NRS=9.8303 M=1 R=5.55556
+ SA=90000.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_A_328_93#_M1003_d N_C_M1003_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1856 AS=0.153912 PD=1.86 PS=1.1122 NRD=1.5366 NRS=57.0906 M=1 R=3.55556
+ SA=90001.3 SB=90000.2 A=0.1152 P=1.64 MULT=1
MM1016 N_A_79_21#_M1016_d N_C_M1016_g N_A_453_325#_M1016_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.16135 AS=0.2814 PD=1.335 PS=2.35 NRD=1.1623 NRS=1.1623 M=1
+ R=4.66667 SA=90000.2 SB=90000.7 A=0.1512 P=2.04 MULT=1
MM1000 N_A_477_49#_M1000_d N_A_328_93#_M1000_g N_A_79_21#_M1016_d VPB PHIGHVT
+ L=0.18 W=0.84 AD=0.33075 AS=0.16135 PD=2.47 PS=1.335 NRD=25.7873 NRS=17.5724
+ M=1 R=4.66667 SA=90000.7 SB=90000.3 A=0.1512 P=2.04 MULT=1
MM1005 N_A_885_297#_M1005_d N_B_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.32 AS=0.26655 PD=2.64 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1010 N_A_477_49#_M1010_d N_B_M1010_g N_A_1003_297#_M1010_s VPB PHIGHVT L=0.18
+ W=0.84 AD=0.284351 AS=0.3612 PD=1.66297 PS=2.54 NRD=48.068 NRS=38.6908 M=1
+ R=4.66667 SA=90000.3 SB=90002.4 A=0.1512 P=2.04 MULT=1
MM1017 N_A_1286_297#_M1017_d N_A_885_297#_M1017_g N_A_477_49#_M1010_d VPB
+ PHIGHVT L=0.18 W=0.64 AD=0.2268 AS=0.216649 PD=1.465 PS=1.26703 NRD=95.4071
+ NRS=43.0839 M=1 R=3.55556 SA=90001.1 SB=90002.3 A=0.1152 P=1.64 MULT=1
MM1006 N_A_453_325#_M1006_d N_B_M1006_g N_A_1286_297#_M1017_d VPB PHIGHVT L=0.18
+ W=0.64 AD=0.154638 AS=0.2268 PD=1.12865 PS=1.465 NRD=57.4255 NRS=3.0732 M=1
+ R=3.55556 SA=90001.6 SB=90002.1 A=0.1152 P=1.64 MULT=1
MM1014 N_A_1003_297#_M1014_d N_A_885_297#_M1014_g N_A_453_325#_M1006_d VPB
+ PHIGHVT L=0.18 W=0.84 AD=0.164987 AS=0.202962 PD=1.25543 PS=1.48135
+ NRD=33.1551 NRS=0 M=1 R=4.66667 SA=90001.7 SB=90001.4 A=0.1512 P=2.04 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_A_1003_297#_M1014_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.196413 PD=1.29 PS=1.49457 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1011 N_A_1286_297#_M1011_d N_A_1003_297#_M1011_g N_VPWR_M1018_d VPB PHIGHVT
+ L=0.18 W=1 AD=0.475 AS=0.145 PD=2.95 PS=1.29 NRD=37.9225 NRS=0.9653 M=1
+ R=5.55556 SA=90002.4 SB=90000.4 A=0.18 P=2.36 MULT=1
DX24_noxref VNB VPB NWDIODE A=16.1142 P=23.29
*
.include "sky130_fd_sc_hdll__xnor3_2.pxi.spice"
*
.ends
*
*
