* File: sky130_fd_sc_hdll__nor3_2.pex.spice
* Created: Thu Aug 27 19:16:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%A 1 3 4 6 7 9 10 12 13 14 22 27
c37 14 0 1.93357e-19 $X=0.66 $Y=1.105
r38 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.01 $Y2=1.202
r39 20 22 43.1263 $w=3.8e-07 $l=3.4e-07 $layer=POLY_cond $X=0.645 $Y=1.202
+ $X2=0.985 $Y2=1.202
r40 20 27 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.645
+ $Y=1.16 $X2=0.645 $Y2=1.16
r41 18 20 16.4895 $w=3.8e-07 $l=1.3e-07 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.645 $Y2=1.202
r42 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.49 $Y=1.202
+ $X2=0.515 $Y2=1.202
r43 14 27 5.28139 $w=2.08e-07 $l=1e-07 $layer=LI1_cond $X=0.745 $Y=1.18
+ $X2=0.645 $Y2=1.18
r44 13 27 21.6537 $w=2.08e-07 $l=4.1e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.645 $Y2=1.18
r45 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=1.202
r46 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.01 $Y=0.995
+ $X2=1.01 $Y2=0.56
r47 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r48 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r49 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r50 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
r51 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.49 $Y=0.995
+ $X2=0.49 $Y2=1.202
r52 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.49 $Y=0.995 $X2=0.49
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%B 1 3 4 6 7 9 10 12 13 14 22 25
c42 22 0 1.93357e-19 $X=1.925 $Y=1.202
r43 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.925 $Y=1.202
+ $X2=1.95 $Y2=1.202
r44 20 22 31.7105 $w=3.8e-07 $l=2.5e-07 $layer=POLY_cond $X=1.675 $Y=1.202
+ $X2=1.925 $Y2=1.202
r45 18 20 27.9053 $w=3.8e-07 $l=2.2e-07 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.675 $Y2=1.202
r46 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.43 $Y=1.202
+ $X2=1.455 $Y2=1.202
r47 13 14 23.7662 $w=2.08e-07 $l=4.5e-07 $layer=LI1_cond $X=1.62 $Y=1.18
+ $X2=2.07 $Y2=1.18
r48 13 25 0.264069 $w=2.08e-07 $l=5e-09 $layer=LI1_cond $X=1.62 $Y=1.18
+ $X2=1.615 $Y2=1.18
r49 13 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.675
+ $Y=1.16 $X2=1.675 $Y2=1.16
r50 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.202
r51 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=0.56
r52 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.202
r53 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.925 $Y=1.41
+ $X2=1.925 $Y2=1.985
r54 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r55 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r56 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.43 $Y=0.995
+ $X2=1.43 $Y2=1.202
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.43 $Y=0.995 $X2=1.43
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%C 1 3 4 6 7 9 10 12 15 18 19 25 27
c43 4 0 1.50204e-19 $X=3.03 $Y=1.41
r44 25 26 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.5 $Y=1.202
+ $X2=3.525 $Y2=1.202
r45 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.005 $Y=1.202
+ $X2=3.03 $Y2=1.202
r46 18 19 8.29932 $w=4.88e-07 $l=3.4e-07 $layer=LI1_cond $X=2.69 $Y=1.19
+ $X2=2.69 $Y2=1.53
r47 18 27 0.244098 $w=4.88e-07 $l=1e-08 $layer=LI1_cond $X=2.69 $Y=1.19 $X2=2.69
+ $Y2=1.18
r48 16 25 51.3711 $w=3.8e-07 $l=4.05e-07 $layer=POLY_cond $X=3.095 $Y=1.202
+ $X2=3.5 $Y2=1.202
r49 16 23 8.24474 $w=3.8e-07 $l=6.5e-08 $layer=POLY_cond $X=3.095 $Y=1.202
+ $X2=3.03 $Y2=1.202
r50 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.095
+ $Y=1.16 $X2=3.095 $Y2=1.16
r51 13 27 5.72758 $w=2.1e-07 $l=2.45e-07 $layer=LI1_cond $X=2.935 $Y=1.18
+ $X2=2.69 $Y2=1.18
r52 13 15 8.45022 $w=2.08e-07 $l=1.6e-07 $layer=LI1_cond $X=2.935 $Y=1.18
+ $X2=3.095 $Y2=1.18
r53 10 26 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.525 $Y=0.995
+ $X2=3.525 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.525 $Y=0.995
+ $X2=3.525 $Y2=0.56
r55 7 25 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.5 $Y=1.41 $X2=3.5
+ $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.5 $Y=1.41 $X2=3.5
+ $Y2=1.985
r57 4 23 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.03 $Y=1.41
+ $X2=3.03 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.03 $Y=1.41 $X2=3.03
+ $Y2=1.985
r59 1 22 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.005 $Y=0.995
+ $X2=3.005 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%A_27_297# 1 2 3 10 12 14 18 20 27 29
r35 21 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=1.54
+ $X2=1.22 $Y2=1.54
r36 20 29 4.1433 $w=1.7e-07 $l=1.2e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=2.155 $Y2=1.54
r37 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.035 $Y=1.54
+ $X2=1.345 $Y2=1.54
r38 16 27 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=1.54
r39 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=1.22 $Y=1.625
+ $X2=1.22 $Y2=2.3
r40 15 25 4.31308 $w=1.7e-07 $l=1.28e-07 $layer=LI1_cond $X=0.405 $Y=1.54
+ $X2=0.277 $Y2=1.54
r41 14 27 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=1.22 $Y2=1.54
r42 14 15 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.095 $Y=1.54
+ $X2=0.405 $Y2=1.54
r43 10 25 2.86415 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=1.54
r44 10 12 30.5058 $w=2.53e-07 $l=6.75e-07 $layer=LI1_cond $X=0.277 $Y=1.625
+ $X2=0.277 $Y2=2.3
r45 3 29 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=2.015
+ $Y=1.485 $X2=2.16 $Y2=1.62
r46 2 27 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=1.62
r47 2 18 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r48 1 25 400 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.62
r49 1 12 400 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%VPWR 1 8 10 17 18 21
r40 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 17 18 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r42 15 18 0.785335 $w=4.8e-07 $l=2.76e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r43 15 22 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 14 17 180.064 $w=1.68e-07 $l=2.76e-06 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=3.91 $Y2=2.72
r45 14 15 2.65714 $w=1.7e-07 $l=5.95e-07 $layer=mcon $count=3 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r46 12 21 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=0.75 $Y2=2.72
r47 12 14 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=0.875 $Y=2.72
+ $X2=1.15 $Y2=2.72
r48 10 22 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 6 21 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=2.635
+ $X2=0.75 $Y2=2.72
r50 6 8 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.75 $Y=2.635 $X2=0.75
+ $Y2=1.96
r51 1 8 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%A_309_297# 1 2 3 12 14 15 18 20 24 26
r31 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=3.735 $Y=2.295
+ $X2=3.735 $Y2=1.96
r32 21 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.92 $Y=2.38
+ $X2=2.815 $Y2=2.38
r33 20 22 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=3.61 $Y=2.38
+ $X2=3.735 $Y2=2.295
r34 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=3.61 $Y=2.38 $X2=2.92
+ $Y2=2.38
r35 16 26 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=2.815 $Y=2.295
+ $X2=2.815 $Y2=2.38
r36 16 18 17.6926 $w=2.08e-07 $l=3.35e-07 $layer=LI1_cond $X=2.815 $Y=2.295
+ $X2=2.815 $Y2=1.96
r37 14 26 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=2.71 $Y=2.38
+ $X2=2.815 $Y2=2.38
r38 14 15 58.3904 $w=1.68e-07 $l=8.95e-07 $layer=LI1_cond $X=2.71 $Y=2.38
+ $X2=1.815 $Y2=2.38
r39 10 15 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=1.69 $Y=2.295
+ $X2=1.815 $Y2=2.38
r40 10 12 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.69 $Y=2.295
+ $X2=1.69 $Y2=1.96
r41 3 24 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.59
+ $Y=1.485 $X2=3.735 $Y2=1.96
r42 2 18 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=2.67
+ $Y=1.485 $X2=2.795 $Y2=1.96
r43 1 12 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%Y 1 2 3 4 15 17 18 21 23 27 31 34 36 42 45
c69 36 0 1.50204e-19 $X=3.785 $Y=1.445
r70 42 45 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=3.265 $Y=1.54
+ $X2=3.57 $Y2=1.54
r71 39 45 10.8952 $w=1.68e-07 $l=1.67e-07 $layer=LI1_cond $X=3.737 $Y=1.54
+ $X2=3.57 $Y2=1.54
r72 36 39 8.677 $w=1.68e-07 $l=1.33e-07 $layer=LI1_cond $X=3.87 $Y=1.54
+ $X2=3.737 $Y2=1.54
r73 36 39 0.116124 $w=5.13e-07 $l=5e-09 $layer=LI1_cond $X=3.737 $Y=1.45
+ $X2=3.737 $Y2=1.455
r74 34 36 12.6575 $w=5.13e-07 $l=5.45e-07 $layer=LI1_cond $X=3.737 $Y=0.905
+ $X2=3.737 $Y2=1.45
r75 25 34 30.6232 $w=1.78e-07 $l=4.97e-07 $layer=LI1_cond $X=3.24 $Y=0.815
+ $X2=3.737 $Y2=0.815
r76 25 27 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.24 $Y=0.725
+ $X2=3.24 $Y2=0.39
r77 24 31 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.855 $Y=0.815
+ $X2=1.665 $Y2=0.815
r78 23 25 11.7071 $w=1.78e-07 $l=1.9e-07 $layer=LI1_cond $X=3.05 $Y=0.815
+ $X2=3.24 $Y2=0.815
r79 23 24 73.6313 $w=1.78e-07 $l=1.195e-06 $layer=LI1_cond $X=3.05 $Y=0.815
+ $X2=1.855 $Y2=0.815
r80 19 31 1.15089 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.815
r81 19 21 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.665 $Y=0.725
+ $X2=1.665 $Y2=0.39
r82 17 31 9.12476 $w=1.8e-07 $l=1.9e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=1.665 $Y2=0.815
r83 17 18 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=1.475 $Y=0.815
+ $X2=0.915 $Y2=0.815
r84 13 18 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.915 $Y2=0.815
r85 13 15 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.725 $Y=0.725
+ $X2=0.725 $Y2=0.39
r86 4 42 300 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=2 $X=3.12
+ $Y=1.485 $X2=3.265 $Y2=1.62
r87 3 27 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=3.08
+ $Y=0.235 $X2=3.265 $Y2=0.39
r88 2 21 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.505
+ $Y=0.235 $X2=1.69 $Y2=0.39
r89 1 15 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=0.565
+ $Y=0.235 $X2=0.75 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR3_2%VGND 1 2 3 4 5 16 18 20 24 26 28 30 37 46
+ 50 56 59
r55 58 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r56 55 56 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.795 $Y=0.235
+ $X2=2.88 $Y2=0.235
r57 52 55 4.95251 $w=6.38e-07 $l=2.65e-07 $layer=LI1_cond $X=2.53 $Y=0.235
+ $X2=2.795 $Y2=0.235
r58 52 53 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r59 49 52 6.91483 $w=6.38e-07 $l=3.7e-07 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.53 $Y2=0.235
r60 49 50 8.92176 $w=6.38e-07 $l=8.5e-08 $layer=LI1_cond $X=2.16 $Y=0.235
+ $X2=2.075 $Y2=0.235
r61 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 41 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r63 41 53 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r64 40 56 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.45 $Y=0 $X2=2.88
+ $Y2=0
r65 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r66 37 58 4.23784 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.895
+ $Y2=0
r67 37 40 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=3.65 $Y=0 $X2=3.45
+ $Y2=0
r68 36 53 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r69 36 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r70 35 50 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.07 $Y=0 $X2=2.075
+ $Y2=0
r71 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r72 33 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=0 $X2=1.22
+ $Y2=0
r73 33 35 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=1.305 $Y=0 $X2=2.07
+ $Y2=0
r74 30 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r75 30 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 26 58 3.2 $w=2.9e-07 $l=1.36015e-07 $layer=LI1_cond $X=3.795 $Y=0.085
+ $X2=3.895 $Y2=0
r77 26 28 12.1205 $w=2.88e-07 $l=3.05e-07 $layer=LI1_cond $X=3.795 $Y=0.085
+ $X2=3.795 $Y2=0.39
r78 22 46 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r79 22 24 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.39
r80 21 43 4.28094 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r81 20 46 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.135 $Y=0 $X2=1.22
+ $Y2=0
r82 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.135 $Y=0 $X2=0.365
+ $Y2=0
r83 16 43 3.0411 $w=2.75e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.182 $Y2=0
r84 16 18 12.7816 $w=2.73e-07 $l=3.05e-07 $layer=LI1_cond $X=0.227 $Y=0.085
+ $X2=0.227 $Y2=0.39
r85 5 28 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.6
+ $Y=0.235 $X2=3.735 $Y2=0.39
r86 4 55 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.67
+ $Y=0.235 $X2=2.795 $Y2=0.39
r87 3 49 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.16 $Y2=0.39
r88 2 24 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.085
+ $Y=0.235 $X2=1.22 $Y2=0.39
r89 1 18 91 $w=1.7e-07 $l=2.13834e-07 $layer=licon1_NDIFF $count=2 $X=0.14
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

