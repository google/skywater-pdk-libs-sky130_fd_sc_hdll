* File: sky130_fd_sc_hdll__einvn_4.pex.spice
* Created: Thu Aug 27 19:07:35 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%TE_B 1 3 4 6 7 8 9 11 12 14 16 17 19 21 22
+ 24 26 27 30 31 32
c80 31 0 7.37964e-20 $X=1.96 $Y=1.395
c81 30 0 7.37964e-20 $X=1.49 $Y=1.395
c82 22 0 2.39076e-19 $X=2.34 $Y=1.395
c83 17 0 1.65302e-19 $X=1.87 $Y=1.395
c84 4 0 1.15275e-19 $X=0.495 $Y=1.41
r85 37 38 3.48266 $w=3.46e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.202
+ $X2=0.495 $Y2=1.202
r86 35 37 31.3439 $w=3.46e-07 $l=2.25e-07 $layer=POLY_cond $X=0.245 $Y=1.202
+ $X2=0.47 $Y2=1.202
r87 32 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.245
+ $Y=1.16 $X2=0.245 $Y2=1.16
r88 27 29 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=1.02 $Y=1.25 $X2=1.02
+ $Y2=1.395
r89 24 26 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=2.43 $Y=1.47
+ $X2=2.43 $Y2=2.015
r90 23 31 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=2.05 $Y=1.395 $X2=1.96
+ $Y2=1.395
r91 22 24 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=2.34 $Y=1.395
+ $X2=2.43 $Y2=1.47
r92 22 23 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=2.34 $Y=1.395
+ $X2=2.05 $Y2=1.395
r93 19 31 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.96 $Y=1.47 $X2=1.96
+ $Y2=1.395
r94 19 21 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.96 $Y=1.47
+ $X2=1.96 $Y2=2.015
r95 18 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.58 $Y=1.395 $X2=1.49
+ $Y2=1.395
r96 17 31 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.87 $Y=1.395 $X2=1.96
+ $Y2=1.395
r97 17 18 148.702 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=1.87 $Y=1.395
+ $X2=1.58 $Y2=1.395
r98 14 30 2.7459 $w=1.8e-07 $l=7.5e-08 $layer=POLY_cond $X=1.49 $Y=1.47 $X2=1.49
+ $Y2=1.395
r99 14 16 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.49 $Y=1.47
+ $X2=1.49 $Y2=2.015
r100 13 29 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=1.12 $Y=1.395
+ $X2=1.02 $Y2=1.395
r101 12 30 23.6879 $w=1.5e-07 $l=9e-08 $layer=POLY_cond $X=1.4 $Y=1.395 $X2=1.49
+ $Y2=1.395
r102 12 13 143.574 $w=1.5e-07 $l=2.8e-07 $layer=POLY_cond $X=1.4 $Y=1.395
+ $X2=1.12 $Y2=1.395
r103 9 29 25.676 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=1.02 $Y=1.47 $X2=1.02
+ $Y2=1.395
r104 9 11 145.939 $w=1.8e-07 $l=5.45e-07 $layer=POLY_cond $X=1.02 $Y=1.47
+ $X2=1.02 $Y2=2.015
r105 8 38 29.6845 $w=3.46e-07 $l=1.21655e-07 $layer=POLY_cond $X=0.595 $Y=1.25
+ $X2=0.495 $Y2=1.202
r106 7 27 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=0.92 $Y=1.25 $X2=1.02
+ $Y2=1.25
r107 7 8 166.649 $w=1.5e-07 $l=3.25e-07 $layer=POLY_cond $X=0.92 $Y=1.25
+ $X2=0.595 $Y2=1.25
r108 4 38 18.0377 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r109 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r110 1 37 22.3532 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=1.202
r111 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.47 $Y=0.995
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%A_27_47# 1 2 7 9 10 11 12 14 15 17 19 20
+ 22 24 25 26 27 30 32 36 40
c97 25 0 1.07001e-19 $X=1.98 $Y=1.035
c98 15 0 3.80504e-19 $X=2.375 $Y=1.035
c99 10 0 1.17964e-19 $X=1.905 $Y=1.035
r100 37 40 19.2492 $w=3.13e-07 $l=1.25e-07 $layer=POLY_cond $X=2.9 $Y=1.16
+ $X2=2.9 $Y2=1.035
r101 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.875
+ $Y=1.16 $X2=2.875 $Y2=1.16
r102 34 39 3.44264 $w=3.3e-07 $l=3.8e-07 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=0.515 $Y2=1.16
r103 34 36 69.1466 $w=3.28e-07 $l=1.98e-06 $layer=LI1_cond $X=0.895 $Y=1.16
+ $X2=2.875 $Y2=1.16
r104 30 39 14.8547 $w=5.24e-07 $l=6.37593e-07 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.515 $Y2=1.16
r105 30 32 6.64871 $w=2.58e-07 $l=1.5e-07 $layer=LI1_cond $X=0.215 $Y=1.665
+ $X2=0.215 $Y2=1.815
r106 27 39 14.8547 $w=5.24e-07 $l=6.37593e-07 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.515 $Y2=1.16
r107 27 29 4.45769 $w=2.6e-07 $l=9.5e-08 $layer=LI1_cond $X=0.215 $Y=0.655
+ $X2=0.215 $Y2=0.56
r108 22 40 24.674 $w=3.13e-07 $l=8.44097e-08 $layer=POLY_cond $X=2.92 $Y=0.96
+ $X2=2.9 $Y2=1.035
r109 22 24 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.92 $Y=0.96 $X2=2.92
+ $Y2=0.56
r110 21 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.525 $Y=1.035
+ $X2=2.45 $Y2=1.035
r111 20 40 19.9686 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=2.74 $Y=1.035
+ $X2=2.9 $Y2=1.035
r112 20 21 110.245 $w=1.5e-07 $l=2.15e-07 $layer=POLY_cond $X=2.74 $Y=1.035
+ $X2=2.525 $Y2=1.035
r113 17 26 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.45 $Y=0.96
+ $X2=2.45 $Y2=1.035
r114 17 19 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.45 $Y=0.96 $X2=2.45
+ $Y2=0.56
r115 16 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.055 $Y=1.035
+ $X2=1.98 $Y2=1.035
r116 15 26 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=2.375 $Y=1.035
+ $X2=2.45 $Y2=1.035
r117 15 16 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.375 $Y=1.035
+ $X2=2.055 $Y2=1.035
r118 12 25 5.30422 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.98 $Y=0.96
+ $X2=1.98 $Y2=1.035
r119 12 14 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.98 $Y=0.96 $X2=1.98
+ $Y2=0.56
r120 10 25 20.4101 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=1.905 $Y=1.035
+ $X2=1.98 $Y2=1.035
r121 10 11 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.905 $Y=1.035
+ $X2=1.585 $Y2=1.035
r122 7 11 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=1.51 $Y=0.96
+ $X2=1.585 $Y2=1.035
r123 7 9 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=1.51 $Y=0.96 $X2=1.51
+ $Y2=0.56
r124 2 32 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.815
r125 1 29 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%A 1 3 4 6 7 9 10 12 13 15 16 18 19 21 22
+ 24 25 26 36
r67 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.145
+ $Y=1.16 $X2=5.145 $Y2=1.16
r68 36 38 34.9945 $w=3.65e-07 $l=2.65e-07 $layer=POLY_cond $X=4.88 $Y=1.202
+ $X2=5.145 $Y2=1.202
r69 35 36 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.855 $Y=1.202
+ $X2=4.88 $Y2=1.202
r70 34 35 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=4.41 $Y=1.202
+ $X2=4.855 $Y2=1.202
r71 33 34 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=4.385 $Y=1.202
+ $X2=4.41 $Y2=1.202
r72 32 33 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=3.94 $Y=1.202
+ $X2=4.385 $Y2=1.202
r73 31 32 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.915 $Y=1.202
+ $X2=3.94 $Y2=1.202
r74 30 31 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=3.47 $Y=1.202
+ $X2=3.915 $Y2=1.202
r75 29 30 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.445 $Y=1.202
+ $X2=3.47 $Y2=1.202
r76 26 39 0.794788 $w=4.33e-07 $l=3e-08 $layer=LI1_cond $X=5.197 $Y=1.19
+ $X2=5.197 $Y2=1.16
r77 25 39 8.21281 $w=4.33e-07 $l=3.1e-07 $layer=LI1_cond $X=5.197 $Y=0.85
+ $X2=5.197 $Y2=1.16
r78 22 36 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.88 $Y=1.41
+ $X2=4.88 $Y2=1.202
r79 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.88 $Y=1.41
+ $X2=4.88 $Y2=1.985
r80 19 35 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=1.202
r81 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.855 $Y=0.995
+ $X2=4.855 $Y2=0.56
r82 16 34 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.41 $Y=1.41
+ $X2=4.41 $Y2=1.202
r83 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.41 $Y=1.41
+ $X2=4.41 $Y2=1.985
r84 13 33 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=1.202
r85 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.385 $Y=0.995
+ $X2=4.385 $Y2=0.56
r86 10 32 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.94 $Y=1.41
+ $X2=3.94 $Y2=1.202
r87 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.94 $Y=1.41
+ $X2=3.94 $Y2=1.985
r88 7 31 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.915 $Y=0.995
+ $X2=3.915 $Y2=1.202
r89 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.915 $Y=0.995
+ $X2=3.915 $Y2=0.56
r90 4 30 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.202
r91 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.47 $Y=1.41 $X2=3.47
+ $Y2=1.985
r92 1 29 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=1.202
r93 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.445 $Y=0.995
+ $X2=3.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%VPWR 1 2 3 12 16 18 22 24 26 31 41 42 45
+ 48 51
r74 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r75 49 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r76 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r77 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r78 41 42 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 39 42 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r80 39 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 38 41 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r82 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r83 36 51 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.89 $Y=2.72 $X2=2.67
+ $Y2=2.72
r84 36 38 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=2.89 $Y=2.72 $X2=2.99
+ $Y2=2.72
r85 35 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r86 35 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r87 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r88 32 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r89 32 34 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r90 31 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.51 $Y=2.72 $X2=1.7
+ $Y2=2.72
r91 31 34 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=1.51 $Y=2.72
+ $X2=1.15 $Y2=2.72
r92 26 45 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r93 26 28 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r94 24 46 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r95 24 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r96 20 51 1.73497 $w=4.4e-07 $l=8.5e-08 $layer=LI1_cond $X=2.67 $Y=2.635
+ $X2=2.67 $Y2=2.72
r97 20 22 16.6318 $w=4.38e-07 $l=6.35e-07 $layer=LI1_cond $X=2.67 $Y=2.635
+ $X2=2.67 $Y2=2
r98 19 48 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.89 $Y=2.72 $X2=1.7
+ $Y2=2.72
r99 18 51 10.4332 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=2.45 $Y=2.72 $X2=2.67
+ $Y2=2.72
r100 18 19 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.45 $Y=2.72
+ $X2=1.89 $Y2=2.72
r101 14 48 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.7 $Y=2.635 $X2=1.7
+ $Y2=2.72
r102 14 16 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=1.7 $Y=2.635
+ $X2=1.7 $Y2=2.02
r103 10 45 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r104 10 12 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.02
r105 3 22 300 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=2 $X=2.52
+ $Y=1.545 $X2=2.665 $Y2=2
r106 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.58
+ $Y=1.545 $X2=1.725 $Y2=2.02
r107 1 12 300 $w=1.7e-07 $l=6.03158e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.02
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%A_222_309# 1 2 3 4 5 18 20 21 24 26 31 32
+ 33 36 38 42 44 45
c72 44 0 1.83817e-19 $X=2.195 $Y=1.58
c73 21 0 1.15275e-19 $X=1.34 $Y=1.58
c74 20 0 2.24965e-19 $X=2.11 $Y=1.58
r75 40 42 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=5.115 $Y=2.295
+ $X2=5.115 $Y2=1.815
r76 39 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.26 $Y=2.38
+ $X2=4.175 $Y2=2.38
r77 38 40 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.03 $Y=2.38
+ $X2=5.115 $Y2=2.295
r78 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.03 $Y=2.38
+ $X2=4.26 $Y2=2.38
r79 34 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.175 $Y=2.295
+ $X2=4.175 $Y2=2.38
r80 34 36 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=4.175 $Y=2.295
+ $X2=4.175 $Y2=1.815
r81 32 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=2.38
+ $X2=4.175 $Y2=2.38
r82 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=4.09 $Y=2.38
+ $X2=3.32 $Y2=2.38
r83 29 33 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.215 $Y=2.295
+ $X2=3.32 $Y2=2.38
r84 29 31 25.3506 $w=2.08e-07 $l=4.8e-07 $layer=LI1_cond $X=3.215 $Y=2.295
+ $X2=3.215 $Y2=1.815
r85 28 31 7.92208 $w=2.08e-07 $l=1.5e-07 $layer=LI1_cond $X=3.215 $Y=1.665
+ $X2=3.215 $Y2=1.815
r86 27 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.28 $Y=1.58
+ $X2=2.195 $Y2=1.58
r87 26 28 6.91519 $w=1.7e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.11 $Y=1.58
+ $X2=3.215 $Y2=1.665
r88 26 27 54.1497 $w=1.68e-07 $l=8.3e-07 $layer=LI1_cond $X=3.11 $Y=1.58
+ $X2=2.28 $Y2=1.58
r89 22 44 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.58
r90 22 24 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.195 $Y=1.665
+ $X2=2.195 $Y2=1.815
r91 20 44 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.11 $Y=1.58
+ $X2=2.195 $Y2=1.58
r92 20 21 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.11 $Y=1.58
+ $X2=1.34 $Y2=1.58
r93 16 21 7.32204 $w=1.7e-07 $l=1.75425e-07 $layer=LI1_cond $X=1.202 $Y=1.665
+ $X2=1.34 $Y2=1.58
r94 16 18 6.28605 $w=2.73e-07 $l=1.5e-07 $layer=LI1_cond $X=1.202 $Y=1.665
+ $X2=1.202 $Y2=1.815
r95 5 42 300 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=2 $X=4.97
+ $Y=1.485 $X2=5.115 $Y2=1.815
r96 4 36 300 $w=1.7e-07 $l=3.95917e-07 $layer=licon1_PDIFF $count=2 $X=4.03
+ $Y=1.485 $X2=4.175 $Y2=1.815
r97 3 31 300 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=2 $X=3.11
+ $Y=1.485 $X2=3.235 $Y2=1.815
r98 2 24 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=2.05
+ $Y=1.545 $X2=2.195 $Y2=1.815
r99 1 18 300 $w=1.7e-07 $l=3.34739e-07 $layer=licon1_PDIFF $count=2 $X=1.11
+ $Y=1.545 $X2=1.255 $Y2=1.815
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%Z 1 2 3 4 15 19 21 23 34 38 43
r44 41 43 0.354651 $w=8.58e-07 $l=2.5e-08 $layer=LI1_cond $X=4.62 $Y=1.05
+ $X2=4.645 $Y2=1.05
r45 32 34 2.83721 $w=8.58e-07 $l=2e-07 $layer=LI1_cond $X=3.705 $Y=1.05
+ $X2=3.905 $Y2=1.05
r46 29 32 0.354651 $w=8.58e-07 $l=2.5e-08 $layer=LI1_cond $X=3.68 $Y=1.05
+ $X2=3.705 $Y2=1.05
r47 23 41 3.47558 $w=8.58e-07 $l=2.45e-07 $layer=LI1_cond $X=4.375 $Y=1.05
+ $X2=4.62 $Y2=1.05
r48 23 38 0.14186 $w=8.58e-07 $l=1e-08 $layer=LI1_cond $X=4.375 $Y=1.05
+ $X2=4.365 $Y2=1.05
r49 21 38 6.38372 $w=8.58e-07 $l=4.5e-07 $layer=LI1_cond $X=3.915 $Y=1.05
+ $X2=4.365 $Y2=1.05
r50 21 34 0.14186 $w=8.58e-07 $l=1e-08 $layer=LI1_cond $X=3.915 $Y=1.05
+ $X2=3.905 $Y2=1.05
r51 17 41 5.54258 $w=3.8e-07 $l=4.3e-07 $layer=LI1_cond $X=4.62 $Y=1.48 $X2=4.62
+ $Y2=1.05
r52 17 19 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=4.62 $Y=1.48
+ $X2=4.62 $Y2=1.61
r53 13 29 5.54258 $w=3.8e-07 $l=4.3e-07 $layer=LI1_cond $X=3.68 $Y=1.48 $X2=3.68
+ $Y2=1.05
r54 13 15 3.94257 $w=3.78e-07 $l=1.3e-07 $layer=LI1_cond $X=3.68 $Y=1.48
+ $X2=3.68 $Y2=1.61
r55 4 19 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=4.5
+ $Y=1.485 $X2=4.645 $Y2=1.61
r56 3 15 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.485 $X2=3.705 $Y2=1.61
r57 2 43 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=4.46
+ $Y=0.235 $X2=4.645 $Y2=0.74
r58 1 32 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.52
+ $Y=0.235 $X2=3.705 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%VGND 1 2 3 12 14 18 22 25 26 27 29 42 43
+ 46 49
r74 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r75 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r76 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r77 42 43 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r78 40 43 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r79 39 42 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r80 39 40 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r81 37 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r82 37 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=1.61
+ $Y2=0
r83 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r84 34 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=1.77
+ $Y2=0
r85 34 36 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=1.935 $Y=0 $X2=2.53
+ $Y2=0
r86 29 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r87 29 31 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r88 27 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r89 27 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r90 25 36 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.53
+ $Y2=0
r91 25 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.545 $Y=0 $X2=2.71
+ $Y2=0
r92 24 39 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.99
+ $Y2=0
r93 24 26 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.875 $Y=0 $X2=2.71
+ $Y2=0
r94 20 26 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0
r95 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.71 $Y=0.085
+ $X2=2.71 $Y2=0.36
r96 16 49 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0
r97 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.77 $Y=0.085
+ $X2=1.77 $Y2=0.36
r98 15 46 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r99 14 49 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.605 $Y=0 $X2=1.77
+ $Y2=0
r100 14 15 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=1.605 $Y=0
+ $X2=0.895 $Y2=0
r101 10 46 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0
r102 10 12 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=0.705 $Y=0.085
+ $X2=0.705 $Y2=0.38
r103 3 22 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.71 $Y2=0.36
r104 2 18 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.77 $Y2=0.36
r105 1 12 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__EINVN_4%A_235_47# 1 2 3 4 5 16 19 20 21 24 29 30
+ 34 36
c65 36 0 9.85391e-20 $X=2.24 $Y=0.74
c66 24 0 7.41152e-20 $X=3.125 $Y=0.74
c67 19 0 5.76004e-19 $X=2.155 $Y=0.74
r68 32 34 53.4639 $w=1.93e-07 $l=9.4e-07 $layer=LI1_cond $X=4.175 $Y=0.352
+ $X2=5.115 $Y2=0.352
r69 30 32 50.0513 $w=1.93e-07 $l=8.8e-07 $layer=LI1_cond $X=3.295 $Y=0.352
+ $X2=4.175 $Y2=0.352
r70 27 29 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=3.21 $Y=0.655
+ $X2=3.21 $Y2=0.56
r71 26 30 6.85817 $w=1.95e-07 $l=1.33918e-07 $layer=LI1_cond $X=3.21 $Y=0.45
+ $X2=3.295 $Y2=0.352
r72 26 29 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=3.21 $Y=0.45
+ $X2=3.21 $Y2=0.56
r73 25 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.325 $Y=0.74
+ $X2=2.24 $Y2=0.74
r74 24 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.125 $Y=0.74
+ $X2=3.21 $Y2=0.655
r75 24 25 52.1925 $w=1.68e-07 $l=8e-07 $layer=LI1_cond $X=3.125 $Y=0.74
+ $X2=2.325 $Y2=0.74
r76 21 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.24 $Y=0.655
+ $X2=2.24 $Y2=0.74
r77 21 23 6.81765 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=2.24 $Y=0.655
+ $X2=2.24 $Y2=0.56
r78 19 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=0.74
+ $X2=2.24 $Y2=0.74
r79 19 20 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.155 $Y=0.74
+ $X2=1.385 $Y2=0.74
r80 16 20 7.68211 $w=1.7e-07 $l=1.9799e-07 $layer=LI1_cond $X=1.225 $Y=0.655
+ $X2=1.385 $Y2=0.74
r81 16 18 3.62188 $w=3.2e-07 $l=9.5e-08 $layer=LI1_cond $X=1.225 $Y=0.655
+ $X2=1.225 $Y2=0.56
r82 5 34 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=4.93
+ $Y=0.235 $X2=5.115 $Y2=0.365
r83 4 32 182 $w=1.7e-07 $l=2.41402e-07 $layer=licon1_NDIFF $count=1 $X=3.99
+ $Y=0.235 $X2=4.175 $Y2=0.365
r84 3 29 182 $w=1.7e-07 $l=4.18927e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.21 $Y2=0.56
r85 2 23 182 $w=1.7e-07 $l=4.07124e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.24 $Y2=0.56
r86 1 18 182 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.56
.ends

