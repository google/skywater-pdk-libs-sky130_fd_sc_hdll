* File: sky130_fd_sc_hdll__or3b_1.pex.spice
* Created: Wed Sep  2 08:48:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%C_N 1 3 4 6 7 12 15
c23 7 0 1.51781e-19 $X=0.15 $Y=1.105
r24 12 13 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r25 10 12 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=0.26 $Y=1.202
+ $X2=0.495 $Y2=1.202
r26 7 15 0.230489 $w=2.48e-07 $l=5e-09 $layer=LI1_cond $X=0.235 $Y=1.2 $X2=0.23
+ $Y2=1.2
r27 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.26
+ $Y=1.16 $X2=0.26 $Y2=1.16
r28 4 13 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r29 4 6 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.675
r30 1 12 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r31 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%A_117_297# 1 2 7 9 12 14 15 16 18
c42 16 0 1.80681e-19 $X=0.73 $Y=1.325
c43 14 0 1.51781e-19 $X=1.385 $Y=1.16
r44 23 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.185
+ $Y=1.16 $X2=1.185 $Y2=1.16
r45 21 23 11.0909 $w=4.62e-07 $l=4.2e-07 $layer=LI1_cond $X=0.892 $Y=0.74
+ $X2=0.892 $Y2=1.16
r46 16 23 9.47731 $w=4.62e-07 $l=2.32282e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.892 $Y2=1.16
r47 16 18 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.73 $Y=1.325
+ $X2=0.73 $Y2=1.63
r48 14 24 34.9723 $w=3.3e-07 $l=2e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.185 $Y2=1.16
r49 14 15 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.485 $Y2=1.202
r50 10 15 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.485 $Y2=1.202
r51 10 12 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.51 $Y2=0.475
r52 7 15 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.202
r53 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.695
r54 2 18 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r55 1 21 182 $w=1.7e-07 $l=3.35783e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.465 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%B 1 2 3 4 6 9 10 11 12 13 19 21 25 28
c40 2 0 2.65584e-19 $X=1.905 $Y=1.31
r41 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.94
+ $Y=2.31 $X2=1.94 $Y2=2.31
r42 13 19 8.03218 $w=3.28e-07 $l=2.3e-07 $layer=LI1_cond $X=1.71 $Y=2.29
+ $X2=1.94 $Y2=2.29
r43 13 28 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=2.29 $X2=1.61
+ $Y2=2.29
r44 12 28 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=1.2 $Y=2.29 $X2=1.61
+ $Y2=2.29
r45 12 25 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=2.29 $X2=1.15
+ $Y2=2.29
r46 11 25 14.3182 $w=3.28e-07 $l=4.1e-07 $layer=LI1_cond $X=0.74 $Y=2.29
+ $X2=1.15 $Y2=2.29
r47 11 21 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=0.74 $Y=2.29 $X2=0.69
+ $Y2=2.29
r48 9 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=1.93 $Y=0.475 $X2=1.93
+ $Y2=0.76
r49 4 18 56.6054 $w=2.52e-07 $l=2.91976e-07 $layer=POLY_cond $X=1.905 $Y=2.035
+ $X2=1.94 $Y2=2.31
r50 4 6 132.161 $w=1.8e-07 $l=3.4e-07 $layer=POLY_cond $X=1.905 $Y=2.035
+ $X2=1.905 $Y2=1.695
r51 3 6 110.782 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.695
r52 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.905 $Y=1.31 $X2=1.905
+ $Y2=1.41
r53 1 10 37.4512 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.905 $Y=0.86 $X2=1.905
+ $Y2=0.76
r54 1 2 149.21 $w=2e-07 $l=4.5e-07 $layer=POLY_cond $X=1.905 $Y=0.86 $X2=1.905
+ $Y2=1.31
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%A 1 3 6 8 9 10 16 17 23
r49 21 23 10.4768 $w=3.28e-07 $l=3e-07 $layer=LI1_cond $X=1.77 $Y=1.16 $X2=2.07
+ $Y2=1.16
r50 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.38
+ $Y=1.16 $X2=2.38 $Y2=1.16
r51 10 16 5.5876 $w=3.28e-07 $l=1.6e-07 $layer=LI1_cond $X=2.22 $Y=1.16 $X2=2.38
+ $Y2=1.16
r52 10 23 5.23838 $w=3.28e-07 $l=1.5e-07 $layer=LI1_cond $X=2.22 $Y=1.16
+ $X2=2.07 $Y2=1.16
r53 9 17 9.64289 $w=2.43e-07 $l=2.05e-07 $layer=LI1_cond $X=1.647 $Y=1.53
+ $X2=1.647 $Y2=1.325
r54 8 17 4.01731 $w=2.45e-07 $l=1.65e-07 $layer=LI1_cond $X=1.647 $Y=1.16
+ $X2=1.647 $Y2=1.325
r55 8 21 2.99472 $w=3.3e-07 $l=1.23e-07 $layer=LI1_cond $X=1.647 $Y=1.16
+ $X2=1.77 $Y2=1.16
r56 4 15 39.1718 $w=2.59e-07 $l=1.93959e-07 $layer=POLY_cond $X=2.445 $Y=0.995
+ $X2=2.382 $Y2=1.16
r57 4 6 266.638 $w=1.5e-07 $l=5.2e-07 $layer=POLY_cond $X=2.445 $Y=0.995
+ $X2=2.445 $Y2=0.475
r58 1 15 51.0578 $w=2.59e-07 $l=2.68328e-07 $layer=POLY_cond $X=2.42 $Y=1.41
+ $X2=2.382 $Y2=1.16
r59 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.42 $Y=1.41 $X2=2.42
+ $Y2=1.695
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%A_225_53# 1 2 3 10 12 13 15 18 22 24 25 26
+ 27 30 32 34 39 40 41 46 48
c93 46 0 1.33059e-19 $X=2.91 $Y=1.16
c94 39 0 1.07404e-19 $X=2.805 $Y=1.495
r95 46 49 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.857 $Y=1.16
+ $X2=2.857 $Y2=1.325
r96 46 48 8.58424 $w=2.73e-07 $l=1.65e-07 $layer=LI1_cond $X=2.857 $Y=1.16
+ $X2=2.857 $Y2=0.995
r97 46 47 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.16 $X2=2.91 $Y2=1.16
r98 41 43 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=2.265 $Y=1.58
+ $X2=2.265 $Y2=1.87
r99 39 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.805 $Y=1.495
+ $X2=2.805 $Y2=1.325
r100 36 48 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.805 $Y=0.825
+ $X2=2.805 $Y2=0.995
r101 35 41 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.35 $Y=1.58
+ $X2=2.265 $Y2=1.58
r102 34 39 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=1.58
+ $X2=2.805 $Y2=1.495
r103 34 35 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=2.72 $Y=1.58
+ $X2=2.35 $Y2=1.58
r104 33 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=0.74
+ $X2=2.19 $Y2=0.74
r105 32 36 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.72 $Y=0.74
+ $X2=2.805 $Y2=0.825
r106 32 33 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=2.72 $Y=0.74
+ $X2=2.275 $Y2=0.74
r107 28 40 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.655
+ $X2=2.19 $Y2=0.74
r108 28 30 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.19 $Y=0.655
+ $X2=2.19 $Y2=0.47
r109 26 43 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=1.87
+ $X2=2.265 $Y2=1.87
r110 26 27 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=2.18 $Y=1.87
+ $X2=1.335 $Y2=1.87
r111 24 40 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=2.19 $Y2=0.74
r112 24 25 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.105 $Y=0.74
+ $X2=1.335 $Y2=0.74
r113 20 27 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.205 $Y=1.785
+ $X2=1.335 $Y2=1.87
r114 20 22 4.43247 $w=2.58e-07 $l=1e-07 $layer=LI1_cond $X=1.205 $Y=1.785
+ $X2=1.205 $Y2=1.685
r115 16 25 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=1.205 $Y=0.655
+ $X2=1.335 $Y2=0.74
r116 16 18 10.4163 $w=2.58e-07 $l=2.35e-07 $layer=LI1_cond $X=1.205 $Y=0.655
+ $X2=1.205 $Y2=0.42
r117 13 47 38.9672 $w=2.67e-07 $l=1.96074e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.917 $Y2=1.16
r118 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.985 $Y=0.995
+ $X2=2.985 $Y2=0.56
r119 10 47 50.2707 $w=2.67e-07 $l=2.70647e-07 $layer=POLY_cond $X=2.96 $Y=1.41
+ $X2=2.917 $Y2=1.16
r120 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.96 $Y=1.41
+ $X2=2.96 $Y2=1.985
r121 3 22 600 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.685
r122 2 30 182 $w=1.7e-07 $l=2.82754e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.265 $X2=2.19 $Y2=0.47
r123 1 18 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.265 $X2=1.25 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%VPWR 1 2 7 9 13 16 17 18 28 29
c33 9 0 1.56946e-19 $X=0.26 $Y=1.66
c34 2 0 1.07404e-19 $X=2.51 $Y=1.485
r35 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r36 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r37 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 23 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r39 22 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=2.72
+ $X2=2.53 $Y2=2.72
r40 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r41 20 32 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r42 20 22 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.69 $Y2=2.72
r43 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r45 16 25 2.60963 $w=1.68e-07 $l=4e-08 $layer=LI1_cond $X=2.57 $Y=2.72 $X2=2.53
+ $Y2=2.72
r46 16 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.57 $Y=2.72 $X2=2.71
+ $Y2=2.72
r47 15 28 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=2.85 $Y=2.72 $X2=3.45
+ $Y2=2.72
r48 15 17 7.6511 $w=1.7e-07 $l=1.4e-07 $layer=LI1_cond $X=2.85 $Y=2.72 $X2=2.71
+ $Y2=2.72
r49 11 17 0.375625 $w=2.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2.72
r50 11 13 26.1358 $w=2.78e-07 $l=6.35e-07 $layer=LI1_cond $X=2.71 $Y=2.635
+ $X2=2.71 $Y2=2
r51 7 32 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.172 $Y2=2.72
r52 7 9 43.2166 $w=2.58e-07 $l=9.75e-07 $layer=LI1_cond $X=0.215 $Y=2.635
+ $X2=0.215 $Y2=1.66
r53 2 13 300 $w=1.7e-07 $l=6.11044e-07 $layer=licon1_PDIFF $count=2 $X=2.51
+ $Y=1.485 $X2=2.72 $Y2=2
r54 1 9 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%X 1 2 10 13 14 15
r18 13 15 3.74205 $w=4.23e-07 $l=1.38e-07 $layer=LI1_cond $X=3.322 $Y=1.707
+ $X2=3.322 $Y2=1.845
r19 13 14 6.47855 $w=4.23e-07 $l=2.12e-07 $layer=LI1_cond $X=3.322 $Y=1.707
+ $X2=3.322 $Y2=1.495
r20 12 14 26.4702 $w=3.18e-07 $l=7.35e-07 $layer=LI1_cond $X=3.375 $Y=0.76
+ $X2=3.375 $Y2=1.495
r21 10 12 5.33966 $w=4.23e-07 $l=1.7e-07 $layer=LI1_cond $X=3.322 $Y=0.59
+ $X2=3.322 $Y2=0.76
r22 2 15 300 $w=1.7e-07 $l=4.2638e-07 $layer=licon1_PDIFF $count=2 $X=3.05
+ $Y=1.485 $X2=3.195 $Y2=1.845
r23 1 10 182 $w=1.7e-07 $l=4.17073e-07 $layer=licon1_NDIFF $count=1 $X=3.06
+ $Y=0.235 $X2=3.195 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR3B_1%VGND 1 2 3 10 12 16 18 20 25 32 33 39
c47 12 0 1.56946e-19 $X=0.26 $Y=0.73
r48 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r49 33 44 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r50 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r51 30 32 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.87 $Y=0 $X2=3.45
+ $Y2=0
r52 29 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r53 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r54 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r55 26 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=1.695
+ $Y2=0
r56 26 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=1.885 $Y=0 $X2=2.07
+ $Y2=0
r57 25 46 10.8465 $w=4.23e-07 $l=4e-07 $layer=LI1_cond $X=2.657 $Y=0 $X2=2.657
+ $Y2=0.4
r58 25 30 6.14847 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=2.657 $Y=0 $X2=2.87
+ $Y2=0
r59 25 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r60 25 28 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.445 $Y=0 $X2=2.07
+ $Y2=0
r61 24 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=1.61
+ $Y2=0
r62 23 24 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r63 21 36 4.14523 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r64 21 23 52.5187 $w=1.68e-07 $l=8.05e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=1.15
+ $Y2=0
r65 20 39 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.695
+ $Y2=0
r66 20 23 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.505 $Y=0 $X2=1.15
+ $Y2=0
r67 18 24 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r68 18 36 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r69 14 39 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0
r70 14 16 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=1.695 $Y=0.085
+ $X2=1.695 $Y2=0.4
r71 10 36 3.06699 $w=2.6e-07 $l=1.04307e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.172 $Y2=0
r72 10 12 28.5895 $w=2.58e-07 $l=6.45e-07 $layer=LI1_cond $X=0.215 $Y=0.085
+ $X2=0.215 $Y2=0.73
r73 3 46 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=2.52
+ $Y=0.265 $X2=2.705 $Y2=0.4
r74 2 16 182 $w=1.7e-07 $l=1.90919e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.265 $X2=1.72 $Y2=0.4
r75 1 12 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.465 $X2=0.26 $Y2=0.73
.ends

