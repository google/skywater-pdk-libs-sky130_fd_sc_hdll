* File: sky130_fd_sc_hdll__mux2_4.pxi.spice
* Created: Thu Aug 27 19:10:48 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2_4%S N_S_c_80_n N_S_M1004_g N_S_c_81_n N_S_M1010_g
+ N_S_c_88_n N_S_M1012_g N_S_c_82_n N_S_M1008_g N_S_c_83_n N_S_c_93_p
+ N_S_c_157_p N_S_c_84_n N_S_c_85_n S N_S_c_86_n N_S_c_125_p
+ PM_SKY130_FD_SC_HDLL__MUX2_4%S
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A_27_47# N_A_27_47#_M1010_s N_A_27_47#_M1004_s
+ N_A_27_47#_c_174_n N_A_27_47#_M1016_g N_A_27_47#_c_175_n N_A_27_47#_M1015_g
+ N_A_27_47#_c_176_n N_A_27_47#_c_181_n N_A_27_47#_c_195_n N_A_27_47#_c_177_n
+ N_A_27_47#_c_178_n N_A_27_47#_c_183_n PM_SKY130_FD_SC_HDLL__MUX2_4%A_27_47#
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A0 N_A0_c_228_n N_A0_M1001_g N_A0_c_224_n
+ N_A0_M1011_g N_A0_c_225_n N_A0_c_226_n A0 A0 N_A0_c_227_n
+ PM_SKY130_FD_SC_HDLL__MUX2_4%A0
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A1 N_A1_c_257_n N_A1_M1014_g N_A1_c_258_n
+ N_A1_M1006_g A1 N_A1_c_259_n A1 PM_SKY130_FD_SC_HDLL__MUX2_4%A1
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A_424_297# N_A_424_297#_M1011_d
+ N_A_424_297#_M1001_d N_A_424_297#_c_296_n N_A_424_297#_M1000_g
+ N_A_424_297#_c_288_n N_A_424_297#_M1003_g N_A_424_297#_c_297_n
+ N_A_424_297#_M1002_g N_A_424_297#_c_289_n N_A_424_297#_M1005_g
+ N_A_424_297#_c_298_n N_A_424_297#_M1007_g N_A_424_297#_c_290_n
+ N_A_424_297#_M1009_g N_A_424_297#_c_299_n N_A_424_297#_M1013_g
+ N_A_424_297#_c_291_n N_A_424_297#_M1017_g N_A_424_297#_c_306_n
+ N_A_424_297#_c_300_n N_A_424_297#_c_314_n N_A_424_297#_c_316_n
+ N_A_424_297#_c_319_n N_A_424_297#_c_292_n N_A_424_297#_c_293_n
+ N_A_424_297#_c_369_p N_A_424_297#_c_294_n N_A_424_297#_c_295_n
+ PM_SKY130_FD_SC_HDLL__MUX2_4%A_424_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_4%VPWR N_VPWR_M1004_d N_VPWR_M1012_d N_VPWR_M1002_d
+ N_VPWR_M1013_d N_VPWR_c_425_n N_VPWR_c_426_n N_VPWR_c_427_n N_VPWR_c_428_n
+ VPWR N_VPWR_c_429_n N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n N_VPWR_c_424_n
+ PM_SKY130_FD_SC_HDLL__MUX2_4%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A_222_297# N_A_222_297#_M1016_d
+ N_A_222_297#_M1014_d N_A_222_297#_c_507_n N_A_222_297#_c_508_n
+ PM_SKY130_FD_SC_HDLL__MUX2_4%A_222_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_4%A_334_297# N_A_334_297#_M1001_s
+ N_A_334_297#_M1012_s N_A_334_297#_c_530_n N_A_334_297#_c_538_n
+ PM_SKY130_FD_SC_HDLL__MUX2_4%A_334_297#
x_PM_SKY130_FD_SC_HDLL__MUX2_4%X N_X_M1003_d N_X_M1009_d N_X_M1000_s N_X_M1007_s
+ N_X_c_558_n N_X_c_559_n N_X_c_562_n N_X_c_566_n N_X_c_568_n N_X_c_572_n
+ N_X_c_577_n N_X_c_578_n N_X_c_580_n N_X_c_583_n N_X_c_585_n N_X_c_587_n X X X
+ N_X_c_554_n N_X_c_556_n X X PM_SKY130_FD_SC_HDLL__MUX2_4%X
x_PM_SKY130_FD_SC_HDLL__MUX2_4%VGND N_VGND_M1010_d N_VGND_M1008_d N_VGND_M1005_s
+ N_VGND_M1017_s VGND N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n
+ N_VGND_c_633_n N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n N_VGND_c_637_n
+ N_VGND_c_638_n PM_SKY130_FD_SC_HDLL__MUX2_4%VGND
cc_1 VNB N_S_c_80_n 0.0275228f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_S_c_81_n 0.0199123f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_S_c_82_n 0.0200245f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.995
cc_4 VNB N_S_c_83_n 0.00213724f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.995
cc_5 VNB N_S_c_84_n 0.00479919f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=0.995
cc_6 VNB N_S_c_85_n 0.00209372f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=1.16
cc_7 VNB N_S_c_86_n 0.0461754f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.16
cc_8 VNB N_A_27_47#_c_174_n 0.0268667f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_27_47#_c_175_n 0.0231693f $X=-0.19 $Y=-0.24 $X2=3.595 $Y2=1.985
cc_10 VNB N_A_27_47#_c_176_n 0.0288959f $X=-0.19 $Y=-0.24 $X2=3.62 $Y2=0.56
cc_11 VNB N_A_27_47#_c_177_n 6.63473e-19 $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_12 VNB N_A_27_47#_c_178_n 0.0127969f $X=-0.19 $Y=-0.24 $X2=2.905 $Y2=1.105
cc_13 VNB N_A0_c_224_n 0.0231022f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_14 VNB N_A0_c_225_n 0.0260952f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A0_c_226_n 0.0113974f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A0_c_227_n 0.00558613f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.805
cc_17 VNB N_A1_c_257_n 0.0250499f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_18 VNB N_A1_c_258_n 0.0204934f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_19 VNB N_A1_c_259_n 0.00226885f $X=-0.19 $Y=-0.24 $X2=3.595 $Y2=1.985
cc_20 VNB N_A_424_297#_c_288_n 0.0171395f $X=-0.19 $Y=-0.24 $X2=3.595 $Y2=1.985
cc_21 VNB N_A_424_297#_c_289_n 0.0164573f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.995
cc_22 VNB N_A_424_297#_c_290_n 0.0169682f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.16
cc_23 VNB N_A_424_297#_c_291_n 0.0185183f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_424_297#_c_292_n 0.00278721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_424_297#_c_293_n 3.7607e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_424_297#_c_294_n 0.00110875f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_424_297#_c_295_n 0.0796931f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VPWR_c_424_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_554_n 0.00760977f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.0245332f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_630_n 0.0153048f $X=-0.19 $Y=-0.24 $X2=0.705 $Y2=0.805
cc_32 VNB N_VGND_c_631_n 0.067702f $X=-0.19 $Y=-0.24 $X2=2.965 $Y2=0.995
cc_33 VNB N_VGND_c_632_n 0.0144191f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_633_n 0.0134014f $X=-0.19 $Y=-0.24 $X2=3.51 $Y2=1.16
cc_35 VNB N_VGND_c_634_n 0.00860652f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_635_n 0.00792095f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_636_n 0.00781721f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_637_n 0.0233724f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_638_n 0.296928f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VPB N_S_c_80_n 0.0295121f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB N_S_c_88_n 0.0207519f $X=-0.19 $Y=1.305 $X2=3.595 $Y2=1.41
cc_42 VPB N_S_c_84_n 0.00204496f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=0.995
cc_43 VPB N_S_c_85_n 9.49428e-19 $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_44 VPB N_S_c_86_n 0.022001f $X=-0.19 $Y=1.305 $X2=3.51 $Y2=1.16
cc_45 VPB N_A_27_47#_c_174_n 0.0317842f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_A_27_47#_c_176_n 0.00902809f $X=-0.19 $Y=1.305 $X2=3.62 $Y2=0.56
cc_47 VPB N_A_27_47#_c_181_n 0.0304719f $X=-0.19 $Y=1.305 $X2=2.88 $Y2=0.72
cc_48 VPB N_A_27_47#_c_177_n 0.00175591f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_49 VPB N_A_27_47#_c_183_n 0.00720662f $X=-0.19 $Y=1.305 $X2=0.54 $Y2=1.16
cc_50 VPB N_A0_c_228_n 0.0197564f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_A0_c_225_n 0.0117723f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A0_c_226_n 0.00678725f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A0_c_227_n 0.008477f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=0.805
cc_54 VPB N_A1_c_257_n 0.0342837f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB N_A1_c_259_n 0.00259849f $X=-0.19 $Y=1.305 $X2=3.595 $Y2=1.985
cc_56 VPB N_A_424_297#_c_296_n 0.0157797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A_424_297#_c_297_n 0.0158087f $X=-0.19 $Y=1.305 $X2=3.62 $Y2=0.56
cc_58 VPB N_A_424_297#_c_298_n 0.01609f $X=-0.19 $Y=1.305 $X2=2.965 $Y2=0.805
cc_59 VPB N_A_424_297#_c_299_n 0.0180323f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=1.16
cc_60 VPB N_A_424_297#_c_300_n 0.00678936f $X=-0.19 $Y=1.305 $X2=3.062 $Y2=1.16
cc_61 VPB N_A_424_297#_c_293_n 0.00162451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_424_297#_c_295_n 0.04826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_VPWR_c_425_n 0.00269553f $X=-0.19 $Y=1.305 $X2=0.705 $Y2=0.805
cc_64 VPB N_VPWR_c_426_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=2.965 $Y2=0.805
cc_65 VPB N_VPWR_c_427_n 0.0112517f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_66 VPB N_VPWR_c_428_n 0.0254666f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.16
cc_67 VPB N_VPWR_c_429_n 0.0151047f $X=-0.19 $Y=1.305 $X2=2.905 $Y2=1.105
cc_68 VPB N_VPWR_c_430_n 0.0658349f $X=-0.19 $Y=1.305 $X2=3.51 $Y2=1.16
cc_69 VPB N_VPWR_c_431_n 0.0141085f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_432_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_433_n 0.00532298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_434_n 0.0054644f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_435_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_VPWR_c_424_n 0.0502731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_A_222_297#_c_507_n 0.00919862f $X=-0.19 $Y=1.305 $X2=3.595 $Y2=1.41
cc_76 VPB N_A_222_297#_c_508_n 0.00666098f $X=-0.19 $Y=1.305 $X2=3.62 $Y2=0.995
cc_77 VPB N_A_334_297#_c_530_n 0.00979017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_X_c_556_n 0.00777576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB X 0.0126538f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 N_S_c_80_n N_A_27_47#_c_174_n 0.051602f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_81 N_S_c_93_p N_A_27_47#_c_174_n 0.00309954f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_82 N_S_c_85_n N_A_27_47#_c_174_n 0.00205493f $X=0.705 $Y=1.16 $X2=0 $Y2=0
cc_83 N_S_c_81_n N_A_27_47#_c_175_n 0.0189841f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_84 N_S_c_83_n N_A_27_47#_c_175_n 0.0040103f $X=0.705 $Y=0.995 $X2=0 $Y2=0
cc_85 N_S_c_93_p N_A_27_47#_c_175_n 0.0142909f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_86 N_S_c_80_n N_A_27_47#_c_176_n 0.0139665f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_87 N_S_c_81_n N_A_27_47#_c_176_n 0.00729071f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_88 N_S_c_83_n N_A_27_47#_c_176_n 0.0065627f $X=0.705 $Y=0.995 $X2=0 $Y2=0
cc_89 N_S_c_85_n N_A_27_47#_c_176_n 0.0249363f $X=0.705 $Y=1.16 $X2=0 $Y2=0
cc_90 N_S_c_80_n N_A_27_47#_c_181_n 0.00751475f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_91 N_S_c_80_n N_A_27_47#_c_195_n 0.0198562f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_S_c_85_n N_A_27_47#_c_195_n 0.0245059f $X=0.705 $Y=1.16 $X2=0 $Y2=0
cc_93 N_S_c_80_n N_A_27_47#_c_177_n 0.00129325f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_S_c_93_p N_A_27_47#_c_177_n 0.0130468f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_95 N_S_c_85_n N_A_27_47#_c_177_n 0.0255193f $X=0.705 $Y=1.16 $X2=0 $Y2=0
cc_96 N_S_c_93_p N_A0_c_224_n 0.0139486f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_97 N_S_c_93_p N_A0_c_225_n 0.00752321f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_98 N_S_c_93_p N_A0_c_227_n 0.0251041f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_99 N_S_c_93_p N_A1_c_257_n 0.00301939f $X=2.88 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_100 N_S_c_84_n N_A1_c_257_n 0.00313448f $X=2.965 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_101 N_S_c_86_n N_A1_c_257_n 0.0105163f $X=3.51 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_102 N_S_c_93_p N_A1_c_258_n 0.0145387f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_103 N_S_c_84_n N_A1_c_258_n 0.00605028f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_104 N_S_c_93_p N_A1_c_259_n 0.0381081f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_105 N_S_c_84_n N_A1_c_259_n 0.0192835f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_106 N_S_c_86_n N_A1_c_259_n 2.90987e-19 $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_107 N_S_c_93_p N_A_424_297#_M1011_d 0.0053912f $X=2.88 $Y=0.72 $X2=-0.19
+ $Y2=-0.24
cc_108 N_S_c_88_n N_A_424_297#_c_296_n 0.0368018f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_109 N_S_c_82_n N_A_424_297#_c_288_n 0.00992053f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_110 N_S_c_82_n N_A_424_297#_c_306_n 0.00367848f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_111 N_S_c_93_p N_A_424_297#_c_306_n 0.0557657f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_112 N_S_c_86_n N_A_424_297#_c_306_n 0.00362358f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_113 N_S_c_125_p N_A_424_297#_c_306_n 0.00635313f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_114 N_S_c_88_n N_A_424_297#_c_300_n 0.0210969f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_115 N_S_c_84_n N_A_424_297#_c_300_n 0.0102322f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_116 N_S_c_86_n N_A_424_297#_c_300_n 0.00926207f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_117 N_S_c_125_p N_A_424_297#_c_300_n 0.0267348f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_118 N_S_c_82_n N_A_424_297#_c_314_n 0.00686832f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_119 N_S_c_93_p N_A_424_297#_c_314_n 0.00135923f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_120 N_S_c_82_n N_A_424_297#_c_316_n 0.015448f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_121 N_S_c_86_n N_A_424_297#_c_316_n 0.00259935f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_122 N_S_c_125_p N_A_424_297#_c_316_n 0.00991814f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_123 N_S_c_93_p N_A_424_297#_c_319_n 0.011546f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_124 N_S_c_84_n N_A_424_297#_c_319_n 0.00135923f $X=2.965 $Y=0.995 $X2=0 $Y2=0
cc_125 N_S_c_86_n N_A_424_297#_c_319_n 0.00392529f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_126 N_S_c_125_p N_A_424_297#_c_319_n 0.0137618f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_127 N_S_c_82_n N_A_424_297#_c_292_n 0.00444676f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_128 N_S_c_125_p N_A_424_297#_c_292_n 0.00518297f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_129 N_S_c_88_n N_A_424_297#_c_293_n 0.00404704f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_130 N_S_c_86_n N_A_424_297#_c_293_n 0.0025078f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_131 N_S_c_125_p N_A_424_297#_c_293_n 0.00518297f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_132 N_S_c_86_n N_A_424_297#_c_294_n 0.00147534f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_133 N_S_c_125_p N_A_424_297#_c_294_n 0.0125165f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_134 N_S_c_86_n N_A_424_297#_c_295_n 0.0303434f $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_135 N_S_c_125_p N_A_424_297#_c_295_n 2.67853e-19 $X=3.51 $Y=1.16 $X2=0 $Y2=0
cc_136 N_S_c_80_n N_VPWR_c_425_n 0.0170292f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_137 N_S_c_80_n N_VPWR_c_429_n 0.00427505f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_S_c_88_n N_VPWR_c_430_n 0.00429282f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_139 N_S_c_88_n N_VPWR_c_434_n 0.0117752f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_140 N_S_c_80_n N_VPWR_c_424_n 0.0082412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_141 N_S_c_88_n N_VPWR_c_424_n 0.00861216f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_142 N_S_c_88_n N_A_334_297#_c_530_n 0.00801661f $X=3.595 $Y=1.41 $X2=0 $Y2=0
cc_143 N_S_c_83_n N_VGND_M1010_d 0.00100437f $X=0.705 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_144 N_S_c_93_p N_VGND_M1010_d 0.00631878f $X=2.88 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_145 N_S_c_157_p N_VGND_M1010_d 0.0026614f $X=0.79 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_146 N_S_c_81_n N_VGND_c_630_n 0.00273179f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_147 N_S_c_82_n N_VGND_c_631_n 0.00199743f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_148 N_S_c_93_p N_VGND_c_631_n 0.0190549f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_149 N_S_c_80_n N_VGND_c_634_n 2.41877e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_150 N_S_c_81_n N_VGND_c_634_n 0.0137315f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_151 N_S_c_93_p N_VGND_c_634_n 0.00790208f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_152 N_S_c_157_p N_VGND_c_634_n 0.0111292f $X=0.79 $Y=0.72 $X2=0 $Y2=0
cc_153 N_S_c_85_n N_VGND_c_634_n 0.00282478f $X=0.705 $Y=1.16 $X2=0 $Y2=0
cc_154 N_S_c_82_n N_VGND_c_635_n 0.0127089f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_155 N_S_c_81_n N_VGND_c_638_n 0.00600638f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_156 N_S_c_82_n N_VGND_c_638_n 0.00403341f $X=3.62 $Y=0.995 $X2=0 $Y2=0
cc_157 N_S_c_93_p N_VGND_c_638_n 0.0341968f $X=2.88 $Y=0.72 $X2=0 $Y2=0
cc_158 N_S_c_157_p N_VGND_c_638_n 8.07506e-19 $X=0.79 $Y=0.72 $X2=0 $Y2=0
cc_159 N_S_c_93_p A_226_47# 0.0311516f $X=2.88 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_160 N_S_c_93_p A_530_47# 0.0140052f $X=2.88 $Y=0.72 $X2=-0.19 $Y2=-0.24
cc_161 N_S_c_84_n A_530_47# 0.00214639f $X=2.965 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_162 N_A_27_47#_c_174_n N_A0_c_225_n 0.0107922f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_177_n N_A0_c_225_n 3.2841e-19 $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_164 N_A_27_47#_c_174_n N_A0_c_227_n 0.00436693f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_195_n N_A0_c_227_n 0.00747957f $X=0.96 $Y=1.58 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_177_n N_A0_c_227_n 0.0280061f $X=1.045 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_195_n N_VPWR_M1004_d 0.00701377f $X=0.96 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_168 N_A_27_47#_c_174_n N_VPWR_c_425_n 0.0111859f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_181_n N_VPWR_c_425_n 0.0482148f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_195_n N_VPWR_c_425_n 0.0236824f $X=0.96 $Y=1.58 $X2=0 $Y2=0
cc_171 N_A_27_47#_c_181_n N_VPWR_c_429_n 0.0178516f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_172 N_A_27_47#_c_174_n N_VPWR_c_430_n 0.00599625f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_27_47#_M1004_s N_VPWR_c_424_n 0.00425811f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_174 N_A_27_47#_c_174_n N_VPWR_c_424_n 0.0115131f $X=1.02 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_27_47#_c_181_n N_VPWR_c_424_n 0.00974347f $X=0.26 $Y=1.96 $X2=0 $Y2=0
cc_176 N_A_27_47#_c_195_n N_A_222_297#_M1016_d 0.00406385f $X=0.96 $Y=1.58
+ $X2=-0.19 $Y2=-0.24
cc_177 N_A_27_47#_c_174_n N_A_222_297#_c_508_n 0.0105606f $X=1.02 $Y=1.41 $X2=0
+ $Y2=0
cc_178 N_A_27_47#_c_195_n N_A_222_297#_c_508_n 0.00468399f $X=0.96 $Y=1.58 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_178_n N_VGND_c_630_n 0.013968f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_180 N_A_27_47#_c_175_n N_VGND_c_631_n 0.00425094f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_175_n N_VGND_c_634_n 0.00927917f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_178_n N_VGND_c_634_n 0.0130779f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_183 N_A_27_47#_M1010_s N_VGND_c_638_n 0.0060609f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_175_n N_VGND_c_638_n 0.00751371f $X=1.055 $Y=0.995 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_178_n N_VGND_c_638_n 0.00948668f $X=0.26 $Y=0.46 $X2=0 $Y2=0
cc_186 N_A0_c_228_n N_A1_c_257_n 0.0319991f $X=2.03 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_187 N_A0_c_226_n N_A1_c_257_n 0.0223839f $X=2.03 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_188 N_A0_c_224_n N_A1_c_258_n 0.0258905f $X=2.055 $Y=0.995 $X2=0 $Y2=0
cc_189 N_A0_c_226_n N_A1_c_259_n 0.0200725f $X=2.03 $Y=1.202 $X2=0 $Y2=0
cc_190 N_A0_c_227_n N_A1_c_259_n 0.0260741f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_191 N_A0_c_224_n N_A_424_297#_c_306_n 0.00961348f $X=2.055 $Y=0.995 $X2=0
+ $Y2=0
cc_192 N_A0_c_228_n N_VPWR_c_430_n 0.00434439f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A0_c_228_n N_VPWR_c_424_n 0.00758895f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A0_c_228_n N_A_222_297#_c_507_n 0.0131041f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A0_c_227_n N_A_222_297#_c_507_n 0.00580313f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_196 N_A0_c_228_n N_A_222_297#_c_508_n 0.00371926f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A0_c_227_n N_A_334_297#_M1001_s 0.00419359f $X=1.71 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_198 N_A0_c_228_n N_A_334_297#_c_530_n 0.0128741f $X=2.03 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A0_c_225_n N_A_334_297#_c_530_n 0.00331088f $X=1.93 $Y=1.16 $X2=0 $Y2=0
cc_200 N_A0_c_227_n N_A_334_297#_c_530_n 0.00843607f $X=1.71 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A0_c_224_n N_VGND_c_631_n 0.00403467f $X=2.055 $Y=0.995 $X2=0 $Y2=0
cc_202 N_A0_c_224_n N_VGND_c_638_n 0.00724919f $X=2.055 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_258_n N_A_424_297#_c_306_n 0.0124698f $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_204 N_A1_c_257_n N_A_424_297#_c_300_n 0.0156075f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A1_c_259_n N_A_424_297#_c_300_n 0.0215402f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_206 N_A1_c_258_n N_A_424_297#_c_314_n 0.00374734f $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_207 N_A1_c_258_n N_A_424_297#_c_319_n 5.84083e-19 $X=2.575 $Y=0.995 $X2=0
+ $Y2=0
cc_208 N_A1_c_257_n N_VPWR_c_430_n 0.00434439f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A1_c_257_n N_VPWR_c_424_n 0.00749869f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A1_c_257_n N_A_222_297#_c_507_n 0.00928151f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_211 N_A1_c_257_n N_A_334_297#_c_530_n 0.0141061f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_212 N_A1_c_259_n N_A_334_297#_c_530_n 0.00397174f $X=2.5 $Y=1.16 $X2=0 $Y2=0
cc_213 N_A1_c_257_n N_A_334_297#_c_538_n 0.00247568f $X=2.55 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A1_c_258_n N_VGND_c_631_n 0.00366111f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A1_c_258_n N_VGND_c_638_n 0.00691926f $X=2.575 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_424_297#_c_300_n N_VPWR_M1012_d 0.00593905f $X=3.815 $Y=1.68 $X2=0
+ $Y2=0
cc_217 N_A_424_297#_c_293_n N_VPWR_M1012_d 0.00123403f $X=3.9 $Y=1.595 $X2=0
+ $Y2=0
cc_218 N_A_424_297#_c_296_n N_VPWR_c_426_n 6.33692e-19 $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_424_297#_c_297_n N_VPWR_c_426_n 0.0141913f $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_424_297#_c_298_n N_VPWR_c_426_n 0.0107665f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_424_297#_c_299_n N_VPWR_c_426_n 5.96427e-19 $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_424_297#_c_298_n N_VPWR_c_428_n 6.33692e-19 $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_424_297#_c_299_n N_VPWR_c_428_n 0.0152179f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_424_297#_c_296_n N_VPWR_c_431_n 0.0062441f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_424_297#_c_297_n N_VPWR_c_431_n 0.00427505f $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_424_297#_c_298_n N_VPWR_c_432_n 0.00622633f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_424_297#_c_299_n N_VPWR_c_432_n 0.00427505f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_424_297#_c_296_n N_VPWR_c_434_n 0.00716348f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_229 N_A_424_297#_c_297_n N_VPWR_c_434_n 4.88209e-19 $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_424_297#_c_300_n N_VPWR_c_434_n 0.00924749f $X=3.815 $Y=1.68 $X2=0
+ $Y2=0
cc_231 N_A_424_297#_M1001_d N_VPWR_c_424_n 0.00274149f $X=2.12 $Y=1.485 $X2=0
+ $Y2=0
cc_232 N_A_424_297#_c_296_n N_VPWR_c_424_n 0.0104012f $X=4.065 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A_424_297#_c_297_n N_VPWR_c_424_n 0.00732977f $X=4.535 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_424_297#_c_298_n N_VPWR_c_424_n 0.0104011f $X=5.005 $Y=1.41 $X2=0
+ $Y2=0
cc_235 N_A_424_297#_c_299_n N_VPWR_c_424_n 0.00732977f $X=5.475 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_424_297#_c_300_n N_A_222_297#_M1014_d 0.0118051f $X=3.815 $Y=1.68
+ $X2=0 $Y2=0
cc_237 N_A_424_297#_M1001_d N_A_222_297#_c_507_n 0.00462568f $X=2.12 $Y=1.485
+ $X2=0 $Y2=0
cc_238 N_A_424_297#_c_300_n N_A_334_297#_M1012_s 0.00530375f $X=3.815 $Y=1.68
+ $X2=0 $Y2=0
cc_239 N_A_424_297#_M1001_d N_A_334_297#_c_530_n 0.00468216f $X=2.12 $Y=1.485
+ $X2=0 $Y2=0
cc_240 N_A_424_297#_c_300_n N_A_334_297#_c_530_n 0.084845f $X=3.815 $Y=1.68
+ $X2=0 $Y2=0
cc_241 N_A_424_297#_c_289_n N_X_c_558_n 0.00377939f $X=4.56 $Y=0.995 $X2=0 $Y2=0
cc_242 N_A_424_297#_c_296_n N_X_c_559_n 0.0104664f $X=4.065 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_424_297#_c_297_n N_X_c_559_n 0.00490547f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_244 N_A_424_297#_c_300_n N_X_c_559_n 0.00121446f $X=3.815 $Y=1.68 $X2=0 $Y2=0
cc_245 N_A_424_297#_c_289_n N_X_c_562_n 0.0117298f $X=4.56 $Y=0.995 $X2=0 $Y2=0
cc_246 N_A_424_297#_c_290_n N_X_c_562_n 0.0129187f $X=5.03 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_424_297#_c_369_p N_X_c_562_n 0.0314633f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_424_297#_c_295_n N_X_c_562_n 0.00344781f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_249 N_A_424_297#_c_369_p N_X_c_566_n 0.00902757f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_424_297#_c_295_n N_X_c_566_n 0.00312289f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_251 N_A_424_297#_c_297_n N_X_c_568_n 0.0158817f $X=4.535 $Y=1.41 $X2=0 $Y2=0
cc_252 N_A_424_297#_c_298_n N_X_c_568_n 0.0178551f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_424_297#_c_369_p N_X_c_568_n 0.0264366f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_424_297#_c_295_n N_X_c_568_n 0.00608435f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_255 N_A_424_297#_c_296_n N_X_c_572_n 0.0016148f $X=4.065 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_424_297#_c_300_n N_X_c_572_n 0.0103688f $X=3.815 $Y=1.68 $X2=0 $Y2=0
cc_257 N_A_424_297#_c_293_n N_X_c_572_n 0.00122453f $X=3.9 $Y=1.595 $X2=0 $Y2=0
cc_258 N_A_424_297#_c_369_p N_X_c_572_n 0.00806945f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_424_297#_c_295_n N_X_c_572_n 0.00411408f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_260 N_A_424_297#_c_291_n N_X_c_577_n 0.00377652f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_424_297#_c_298_n N_X_c_578_n 0.00530373f $X=5.005 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_424_297#_c_299_n N_X_c_578_n 0.00490547f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_424_297#_c_291_n N_X_c_580_n 0.0171722f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_424_297#_c_369_p N_X_c_580_n 0.00366099f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_265 N_A_424_297#_c_295_n N_X_c_580_n 2.26856e-19 $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_266 N_A_424_297#_c_299_n N_X_c_583_n 0.0210405f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_424_297#_c_369_p N_X_c_583_n 0.00298838f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_424_297#_c_369_p N_X_c_585_n 0.00902757f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_269 N_A_424_297#_c_295_n N_X_c_585_n 0.00312289f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_270 N_A_424_297#_c_369_p N_X_c_587_n 0.00806945f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_271 N_A_424_297#_c_295_n N_X_c_587_n 0.00411408f $X=5.475 $Y=1.202 $X2=0
+ $Y2=0
cc_272 N_A_424_297#_c_299_n X 0.006513f $X=5.475 $Y=1.41 $X2=0 $Y2=0
cc_273 N_A_424_297#_c_291_n X 0.0236794f $X=5.5 $Y=0.995 $X2=0 $Y2=0
cc_274 N_A_424_297#_c_369_p X 0.0112927f $X=5.265 $Y=1.16 $X2=0 $Y2=0
cc_275 N_A_424_297#_c_316_n N_VGND_M1008_d 0.00541165f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_276 N_A_424_297#_c_292_n N_VGND_M1008_d 7.5176e-19 $X=3.9 $Y=1.075 $X2=0
+ $Y2=0
cc_277 N_A_424_297#_c_306_n N_VGND_c_631_n 0.065108f $X=3.26 $Y=0.38 $X2=0 $Y2=0
cc_278 N_A_424_297#_c_316_n N_VGND_c_631_n 0.00258755f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_279 N_A_424_297#_c_288_n N_VGND_c_632_n 0.00585385f $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_424_297#_c_289_n N_VGND_c_632_n 0.00198377f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_424_297#_c_290_n N_VGND_c_633_n 0.00425094f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_282 N_A_424_297#_c_291_n N_VGND_c_633_n 0.00197669f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_424_297#_c_288_n N_VGND_c_635_n 0.00162962f $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_424_297#_c_306_n N_VGND_c_635_n 0.0132795f $X=3.26 $Y=0.38 $X2=0
+ $Y2=0
cc_285 N_A_424_297#_c_316_n N_VGND_c_635_n 0.0203912f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_286 N_A_424_297#_c_288_n N_VGND_c_636_n 5.64511e-19 $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_287 N_A_424_297#_c_289_n N_VGND_c_636_n 0.00960147f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_288 N_A_424_297#_c_290_n N_VGND_c_636_n 0.0016282f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_289 N_A_424_297#_c_290_n N_VGND_c_637_n 5.65297e-19 $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_290 N_A_424_297#_c_291_n N_VGND_c_637_n 0.0107903f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_291 N_A_424_297#_M1011_d N_VGND_c_638_n 0.00299627f $X=2.13 $Y=0.235 $X2=0
+ $Y2=0
cc_292 N_A_424_297#_c_288_n N_VGND_c_638_n 0.0107343f $X=4.09 $Y=0.995 $X2=0
+ $Y2=0
cc_293 N_A_424_297#_c_289_n N_VGND_c_638_n 0.00271758f $X=4.56 $Y=0.995 $X2=0
+ $Y2=0
cc_294 N_A_424_297#_c_290_n N_VGND_c_638_n 0.00584696f $X=5.03 $Y=0.995 $X2=0
+ $Y2=0
cc_295 N_A_424_297#_c_291_n N_VGND_c_638_n 0.00270442f $X=5.5 $Y=0.995 $X2=0
+ $Y2=0
cc_296 N_A_424_297#_c_306_n N_VGND_c_638_n 0.0484074f $X=3.26 $Y=0.38 $X2=0
+ $Y2=0
cc_297 N_A_424_297#_c_316_n N_VGND_c_638_n 0.00657122f $X=3.815 $Y=0.74 $X2=0
+ $Y2=0
cc_298 N_A_424_297#_c_306_n A_530_47# 0.021461f $X=3.26 $Y=0.38 $X2=-0.19
+ $Y2=-0.24
cc_299 N_A_424_297#_c_314_n A_530_47# 0.00627734f $X=3.345 $Y=0.655 $X2=-0.19
+ $Y2=-0.24
cc_300 N_A_424_297#_c_316_n A_530_47# 0.00149403f $X=3.815 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_301 N_A_424_297#_c_319_n A_530_47# 0.00427672f $X=3.43 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_302 N_VPWR_c_424_n N_A_222_297#_M1016_d 0.00234812f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_303 N_VPWR_c_424_n N_A_222_297#_M1014_d 0.00251338f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_304 N_VPWR_c_430_n N_A_222_297#_c_507_n 0.0800446f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_305 N_VPWR_c_424_n N_A_222_297#_c_507_n 0.0545762f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_306 N_VPWR_c_425_n N_A_222_297#_c_508_n 0.0403842f $X=0.73 $Y=2 $X2=0 $Y2=0
cc_307 N_VPWR_c_430_n N_A_222_297#_c_508_n 0.0225051f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_308 N_VPWR_c_424_n N_A_222_297#_c_508_n 0.0146699f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_309 N_VPWR_c_424_n N_A_334_297#_M1001_s 0.00219219f $X=5.75 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_310 N_VPWR_c_424_n N_A_334_297#_M1012_s 0.00438456f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_311 N_VPWR_c_430_n N_A_334_297#_c_530_n 0.00578029f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_312 N_VPWR_c_424_n N_A_334_297#_c_530_n 0.01133f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_313 N_VPWR_c_430_n N_A_334_297#_c_538_n 0.0116015f $X=3.615 $Y=2.72 $X2=0
+ $Y2=0
cc_314 N_VPWR_c_434_n N_A_334_297#_c_538_n 0.0156776f $X=3.83 $Y=2.34 $X2=0
+ $Y2=0
cc_315 N_VPWR_c_424_n N_A_334_297#_c_538_n 0.00642843f $X=5.75 $Y=2.72 $X2=0
+ $Y2=0
cc_316 N_VPWR_c_424_n N_X_M1000_s 0.00647849f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_317 N_VPWR_c_424_n N_X_M1007_s 0.00647849f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_426_n N_X_c_559_n 0.0410603f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_319 N_VPWR_c_431_n N_X_c_559_n 0.0118139f $X=4.555 $Y=2.72 $X2=0 $Y2=0
cc_320 N_VPWR_c_434_n N_X_c_559_n 0.0128538f $X=3.83 $Y=2.34 $X2=0 $Y2=0
cc_321 N_VPWR_c_424_n N_X_c_559_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_M1002_d N_X_c_568_n 0.00386757f $X=4.625 $Y=1.485 $X2=0 $Y2=0
cc_323 N_VPWR_c_426_n N_X_c_568_n 0.0209383f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_324 N_VPWR_c_426_n N_X_c_578_n 0.0336646f $X=4.77 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_c_428_n N_X_c_578_n 0.0410603f $X=5.71 $Y=2 $X2=0 $Y2=0
cc_326 N_VPWR_c_432_n N_X_c_578_n 0.0118139f $X=5.495 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_424_n N_X_c_578_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_M1013_d N_X_c_583_n 0.00131722f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_329 N_VPWR_c_428_n N_X_c_583_n 0.00745553f $X=5.71 $Y=2 $X2=0 $Y2=0
cc_330 N_VPWR_M1013_d N_X_c_556_n 0.00288305f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_331 N_VPWR_c_428_n N_X_c_556_n 0.0202891f $X=5.71 $Y=2 $X2=0 $Y2=0
cc_332 N_VPWR_M1013_d X 0.00146706f $X=5.565 $Y=1.485 $X2=0 $Y2=0
cc_333 N_A_222_297#_c_507_n N_A_334_297#_M1001_s 0.00519649f $X=2.805 $Y=2.36
+ $X2=-0.19 $Y2=1.305
cc_334 N_A_222_297#_M1014_d N_A_334_297#_c_530_n 0.00648816f $X=2.64 $Y=1.485
+ $X2=0 $Y2=0
cc_335 N_A_222_297#_c_507_n N_A_334_297#_c_530_n 0.074805f $X=2.805 $Y=2.36
+ $X2=0 $Y2=0
cc_336 N_A_222_297#_c_508_n N_A_334_297#_c_530_n 0.0139281f $X=1.275 $Y=2.02
+ $X2=0 $Y2=0
cc_337 N_A_222_297#_c_507_n N_A_334_297#_c_538_n 0.00919609f $X=2.805 $Y=2.36
+ $X2=0 $Y2=0
cc_338 N_X_c_562_n N_VGND_M1005_s 0.00439476f $X=5.155 $Y=0.72 $X2=0 $Y2=0
cc_339 N_X_c_580_n N_VGND_M1017_s 8.22501e-19 $X=5.65 $Y=0.72 $X2=0 $Y2=0
cc_340 N_X_c_554_n N_VGND_M1017_s 0.00272217f $X=5.765 $Y=0.805 $X2=0 $Y2=0
cc_341 X N_VGND_M1017_s 0.00125528f $X=5.755 $Y=0.85 $X2=0 $Y2=0
cc_342 N_X_c_558_n N_VGND_c_632_n 0.01143f $X=4.3 $Y=0.42 $X2=0 $Y2=0
cc_343 N_X_c_562_n N_VGND_c_632_n 0.00244812f $X=5.155 $Y=0.72 $X2=0 $Y2=0
cc_344 N_X_c_562_n N_VGND_c_633_n 0.00313948f $X=5.155 $Y=0.72 $X2=0 $Y2=0
cc_345 N_X_c_577_n N_VGND_c_633_n 0.01143f $X=5.24 $Y=0.42 $X2=0 $Y2=0
cc_346 N_X_c_580_n N_VGND_c_633_n 0.00243833f $X=5.65 $Y=0.72 $X2=0 $Y2=0
cc_347 N_X_c_558_n N_VGND_c_636_n 0.0156777f $X=4.3 $Y=0.42 $X2=0 $Y2=0
cc_348 N_X_c_562_n N_VGND_c_636_n 0.0213178f $X=5.155 $Y=0.72 $X2=0 $Y2=0
cc_349 N_X_c_577_n N_VGND_c_637_n 0.015756f $X=5.24 $Y=0.42 $X2=0 $Y2=0
cc_350 N_X_c_580_n N_VGND_c_637_n 0.00701254f $X=5.65 $Y=0.72 $X2=0 $Y2=0
cc_351 N_X_c_554_n N_VGND_c_637_n 0.0191948f $X=5.765 $Y=0.805 $X2=0 $Y2=0
cc_352 N_X_M1003_d N_VGND_c_638_n 0.00466109f $X=4.165 $Y=0.235 $X2=0 $Y2=0
cc_353 N_X_M1009_d N_VGND_c_638_n 0.00309587f $X=5.105 $Y=0.235 $X2=0 $Y2=0
cc_354 N_X_c_558_n N_VGND_c_638_n 0.00643448f $X=4.3 $Y=0.42 $X2=0 $Y2=0
cc_355 N_X_c_562_n N_VGND_c_638_n 0.0114934f $X=5.155 $Y=0.72 $X2=0 $Y2=0
cc_356 N_X_c_577_n N_VGND_c_638_n 0.00643448f $X=5.24 $Y=0.42 $X2=0 $Y2=0
cc_357 N_X_c_580_n N_VGND_c_638_n 0.00507606f $X=5.65 $Y=0.72 $X2=0 $Y2=0
cc_358 N_X_c_554_n N_VGND_c_638_n 0.00128469f $X=5.765 $Y=0.805 $X2=0 $Y2=0
cc_359 N_VGND_c_638_n A_226_47# 0.0100088f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
cc_360 N_VGND_c_638_n A_530_47# 0.00782464f $X=5.75 $Y=0 $X2=-0.19 $Y2=-0.24
