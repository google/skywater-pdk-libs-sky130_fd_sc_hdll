* File: sky130_fd_sc_hdll__a21o_2.spice
* Created: Thu Aug 27 18:52:50 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21o_2.pex.spice"
.subckt sky130_fd_sc_hdll__a21o_2  VNB VPB B1 A1 A2 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1003 N_X_M1003_d N_A_80_21#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13975 AS=0.17225 PD=1.08 PS=1.83 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1007 N_X_M1003_d N_A_80_21#_M1007_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13975 AS=0.2405 PD=1.08 PS=1.39 NRD=18.456 NRS=40.608 M=1 R=4.33333
+ SA=75000.8 SB=75002.3 A=0.0975 P=1.6 MULT=1
MM1006 N_A_80_21#_M1006_d N_B1_M1006_g N_VGND_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.15925 AS=0.2405 PD=1.14 PS=1.39 NRD=0 NRS=44.304 M=1 R=4.33333 SA=75001.7
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1008 A_532_47# N_A1_M1008_g N_A_80_21#_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.118625 AS=0.15925 PD=1.015 PS=1.14 NRD=23.532 NRS=39.684 M=1 R=4.33333
+ SA=75002.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_VGND_M1009_d N_A2_M1009_g A_532_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.118625 PD=1.92 PS=1.015 NRD=8.304 NRS=23.532 M=1 R=4.33333 SA=75002.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_X_M1002_d N_A_80_21#_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.275 PD=1.35 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90000.8 A=0.18 P=2.36 MULT=1
MM1005 N_X_M1002_d N_A_80_21#_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.325 PD=1.35 PS=2.65 NRD=11.8003 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_A_444_297#_M1004_d N_B1_M1004_g N_A_80_21#_M1004_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.325 PD=1.3 PS=2.65 NRD=1.9503 NRS=11.8003 M=1 R=5.55556
+ SA=90000.2 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_444_297#_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1675 AS=0.15 PD=1.335 PS=1.3 NRD=5.8903 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1000 N_A_444_297#_M1000_d N_A2_M1000_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.1675 PD=2.54 PS=1.335 NRD=0.9653 NRS=4.9053 M=1 R=5.55556
+ SA=90001.2 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_48 VPB 0 8.49032e-20 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__a21o_2.pxi.spice"
*
.ends
*
*
