* File: sky130_fd_sc_hdll__and4b_2.pxi.spice
* Created: Thu Aug 27 18:59:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__AND4B_2%A_N N_A_N_c_86_n N_A_N_c_87_n N_A_N_M1001_g
+ N_A_N_M1008_g A_N A_N A_N N_A_N_c_85_n PM_SKY130_FD_SC_HDLL__AND4B_2%A_N
x_PM_SKY130_FD_SC_HDLL__AND4B_2%A_27_413# N_A_27_413#_M1008_d
+ N_A_27_413#_M1001_s N_A_27_413#_c_116_n N_A_27_413#_c_122_n
+ N_A_27_413#_c_123_n N_A_27_413#_M1011_g N_A_27_413#_c_117_n
+ N_A_27_413#_c_118_n N_A_27_413#_M1010_g N_A_27_413#_c_124_n
+ N_A_27_413#_c_125_n N_A_27_413#_c_126_n N_A_27_413#_c_119_n
+ N_A_27_413#_c_127_n N_A_27_413#_c_162_p N_A_27_413#_c_120_n
+ PM_SKY130_FD_SC_HDLL__AND4B_2%A_27_413#
x_PM_SKY130_FD_SC_HDLL__AND4B_2%B N_B_M1005_g N_B_c_186_n N_B_c_187_n
+ N_B_M1006_g N_B_c_183_n N_B_c_188_n B B B B N_B_c_185_n
+ PM_SKY130_FD_SC_HDLL__AND4B_2%B
x_PM_SKY130_FD_SC_HDLL__AND4B_2%C N_C_c_224_n N_C_c_225_n N_C_M1009_g
+ N_C_M1013_g C C C C N_C_c_223_n PM_SKY130_FD_SC_HDLL__AND4B_2%C
x_PM_SKY130_FD_SC_HDLL__AND4B_2%D N_D_c_267_n N_D_c_268_n N_D_M1000_g
+ N_D_M1002_g D D D N_D_c_266_n PM_SKY130_FD_SC_HDLL__AND4B_2%D
x_PM_SKY130_FD_SC_HDLL__AND4B_2%A_211_413# N_A_211_413#_M1010_s
+ N_A_211_413#_M1011_d N_A_211_413#_M1009_d N_A_211_413#_c_316_n
+ N_A_211_413#_M1004_g N_A_211_413#_c_311_n N_A_211_413#_M1003_g
+ N_A_211_413#_c_317_n N_A_211_413#_M1007_g N_A_211_413#_c_312_n
+ N_A_211_413#_M1012_g N_A_211_413#_c_340_n N_A_211_413#_c_318_n
+ N_A_211_413#_c_319_n N_A_211_413#_c_352_n N_A_211_413#_c_320_n
+ N_A_211_413#_c_321_n N_A_211_413#_c_322_n N_A_211_413#_c_313_n
+ N_A_211_413#_c_338_n N_A_211_413#_c_314_n N_A_211_413#_c_315_n
+ PM_SKY130_FD_SC_HDLL__AND4B_2%A_211_413#
x_PM_SKY130_FD_SC_HDLL__AND4B_2%VPWR N_VPWR_M1001_d N_VPWR_M1006_d
+ N_VPWR_M1000_d N_VPWR_M1007_s N_VPWR_c_430_n N_VPWR_c_431_n N_VPWR_c_432_n
+ N_VPWR_c_433_n N_VPWR_c_434_n N_VPWR_c_435_n VPWR N_VPWR_c_436_n
+ N_VPWR_c_437_n N_VPWR_c_438_n N_VPWR_c_439_n N_VPWR_c_440_n N_VPWR_c_429_n
+ PM_SKY130_FD_SC_HDLL__AND4B_2%VPWR
x_PM_SKY130_FD_SC_HDLL__AND4B_2%X N_X_M1003_s N_X_M1004_d X X X X X X
+ N_X_c_506_n X X PM_SKY130_FD_SC_HDLL__AND4B_2%X
x_PM_SKY130_FD_SC_HDLL__AND4B_2%VGND N_VGND_M1008_s N_VGND_M1002_d
+ N_VGND_M1012_d N_VGND_c_544_n N_VGND_c_545_n N_VGND_c_546_n N_VGND_c_547_n
+ VGND N_VGND_c_548_n N_VGND_c_549_n N_VGND_c_550_n
+ PM_SKY130_FD_SC_HDLL__AND4B_2%VGND
cc_1 VNB N_A_N_M1008_g 0.0378956f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB A_N 0.0134551f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_3 VNB N_A_N_c_85_n 0.0480964f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.16
cc_4 VNB N_A_27_413#_c_116_n 0.0503595f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_5 VNB N_A_27_413#_c_117_n 0.0385264f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_6 VNB N_A_27_413#_c_118_n 0.0173533f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_27_413#_c_119_n 0.00683076f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_27_413#_c_120_n 0.00268127f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_B_M1005_g 0.0358917f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.99
cc_10 VNB N_B_c_183_n 0.0129562f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_11 VNB B 0.00441215f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B_c_185_n 0.00663656f $X=-0.19 $Y=-0.24 $X2=0.235 $Y2=0.85
cc_13 VNB N_C_M1013_g 0.0289822f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_14 VNB C 0.0066282f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_C_c_223_n 0.0222981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_D_M1002_g 0.0277529f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_17 VNB D 0.00949239f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_18 VNB N_D_c_266_n 0.0193485f $X=-0.19 $Y=-0.24 $X2=0.245 $Y2=1.16
cc_19 VNB N_A_211_413#_c_311_n 0.018087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_211_413#_c_312_n 0.0190959f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_211_413#_c_313_n 0.00985932f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_211_413#_c_314_n 0.00253552f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_211_413#_c_315_n 0.0509391f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VPWR_c_429_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB X 0.00825301f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_26 VNB X 0.0227136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_544_n 0.0115458f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_28 VNB N_VGND_c_545_n 0.0153468f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_29 VNB N_VGND_c_546_n 0.00801182f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_547_n 0.0728129f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_548_n 0.0163621f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_549_n 0.0250796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_550_n 0.247547f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VPB N_A_N_c_86_n 0.0401646f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_35 VPB N_A_N_c_87_n 0.0256644f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_36 VPB A_N 0.0170388f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_37 VPB N_A_N_c_85_n 0.0112694f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_38 VPB N_A_27_413#_c_116_n 0.00646937f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_39 VPB N_A_27_413#_c_122_n 0.0351488f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_40 VPB N_A_27_413#_c_123_n 0.0259078f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_A_27_413#_c_124_n 0.00287295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_A_27_413#_c_125_n 0.0085818f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_43 VPB N_A_27_413#_c_126_n 0.00854499f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB N_A_27_413#_c_127_n 0.00956739f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_45 VPB N_A_27_413#_c_120_n 4.83739e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_B_c_186_n 0.0101188f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_47 VPB N_B_c_187_n 0.0254007f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.445
cc_48 VPB N_B_c_188_n 0.0115151f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB B 0.00451303f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_B_c_185_n 0.021433f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=0.85
cc_51 VPB N_C_c_224_n 0.0309012f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_52 VPB N_C_c_225_n 0.0222667f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_53 VPB C 0.00440836f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_C_c_223_n 0.00331124f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_D_c_267_n 0.0310219f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.89
cc_56 VPB N_D_c_268_n 0.0235304f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.99
cc_57 VPB D 0.00520047f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_58 VPB N_D_c_266_n 0.00301727f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_59 VPB N_A_211_413#_c_316_n 0.0165946f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_60 VPB N_A_211_413#_c_317_n 0.0195644f $X=-0.19 $Y=1.305 $X2=0.245 $Y2=1.16
cc_61 VPB N_A_211_413#_c_318_n 0.0261056f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.53
cc_62 VPB N_A_211_413#_c_319_n 0.00763843f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_211_413#_c_320_n 0.00445452f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_211_413#_c_321_n 0.00110566f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_211_413#_c_322_n 0.0157754f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_211_413#_c_313_n 0.00852237f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_211_413#_c_314_n 2.30056e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_211_413#_c_315_n 0.0268914f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_430_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_431_n 0.00287347f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_432_n 0.0117623f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=1.16
cc_72 VPB N_VPWR_c_433_n 0.0300471f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=0.85
cc_73 VPB N_VPWR_c_434_n 0.0177825f $X=-0.19 $Y=1.305 $X2=0.235 $Y2=1.16
cc_74 VPB N_VPWR_c_435_n 0.00513434f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_VPWR_c_436_n 0.0152577f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_VPWR_c_437_n 0.0189775f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_438_n 0.00503031f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_78 VPB N_VPWR_c_439_n 0.0210304f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_440_n 0.0118622f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_429_n 0.0478595f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB X 0.00614618f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_82 VPB X 0.011463f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 N_A_N_M1008_g N_A_27_413#_c_116_n 0.00790114f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_84 A_N N_A_27_413#_c_116_n 2.48101e-19 $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_85 N_A_N_c_85_n N_A_27_413#_c_116_n 0.0210246f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_N_c_86_n N_A_27_413#_c_122_n 0.0131033f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_87 N_A_N_c_87_n N_A_27_413#_c_123_n 0.0251464f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_88 N_A_N_c_87_n N_A_27_413#_c_124_n 0.00662f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_89 N_A_N_c_86_n N_A_27_413#_c_125_n 0.0115768f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_90 N_A_N_c_87_n N_A_27_413#_c_125_n 0.00913427f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_91 N_A_N_c_85_n N_A_27_413#_c_125_n 0.00130998f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_92 A_N N_A_27_413#_c_126_n 0.0132061f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_93 N_A_N_c_85_n N_A_27_413#_c_126_n 9.93381e-19 $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_94 N_A_N_M1008_g N_A_27_413#_c_119_n 0.00747831f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_95 A_N N_A_27_413#_c_119_n 0.0117563f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_96 N_A_N_c_86_n N_A_27_413#_c_127_n 0.00730207f $X=0.495 $Y=1.89 $X2=0 $Y2=0
cc_97 A_N N_A_27_413#_c_127_n 0.014058f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_98 A_N N_A_27_413#_c_120_n 0.0148927f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_99 N_A_N_c_85_n N_A_27_413#_c_120_n 0.00324847f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_100 N_A_N_c_87_n N_VPWR_c_430_n 0.011944f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_101 N_A_N_c_87_n N_VPWR_c_436_n 0.00323276f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_102 N_A_N_c_87_n N_VPWR_c_429_n 0.00477569f $X=0.495 $Y=1.99 $X2=0 $Y2=0
cc_103 N_A_N_M1008_g N_VGND_c_545_n 0.00482545f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_104 A_N N_VGND_c_545_n 0.0114029f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_105 N_A_N_c_85_n N_VGND_c_545_n 0.00382627f $X=0.52 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_N_M1008_g N_VGND_c_547_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_107 N_A_N_M1008_g N_VGND_c_550_n 0.0127868f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_108 A_N N_VGND_c_550_n 0.00107484f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_109 N_A_27_413#_c_116_n N_B_M1005_g 0.00424142f $X=0.965 $Y=1.325 $X2=0 $Y2=0
cc_110 N_A_27_413#_c_118_n N_B_M1005_g 0.0373108f $X=1.51 $Y=0.73 $X2=0 $Y2=0
cc_111 N_A_27_413#_c_118_n B 0.00167921f $X=1.51 $Y=0.73 $X2=0 $Y2=0
cc_112 N_A_27_413#_c_116_n N_A_211_413#_c_322_n 3.57503e-19 $X=0.965 $Y=1.325
+ $X2=0 $Y2=0
cc_113 N_A_27_413#_c_122_n N_A_211_413#_c_322_n 0.00831163f $X=0.965 $Y=1.89
+ $X2=0 $Y2=0
cc_114 N_A_27_413#_c_123_n N_A_211_413#_c_322_n 0.00727211f $X=0.965 $Y=1.99
+ $X2=0 $Y2=0
cc_115 N_A_27_413#_c_125_n N_A_211_413#_c_322_n 0.0110751f $X=0.685 $Y=1.915
+ $X2=0 $Y2=0
cc_116 N_A_27_413#_c_127_n N_A_211_413#_c_322_n 0.00990573f $X=0.77 $Y=1.83
+ $X2=0 $Y2=0
cc_117 N_A_27_413#_c_116_n N_A_211_413#_c_313_n 0.00553331f $X=0.965 $Y=1.325
+ $X2=0 $Y2=0
cc_118 N_A_27_413#_c_122_n N_A_211_413#_c_313_n 0.00746912f $X=0.965 $Y=1.89
+ $X2=0 $Y2=0
cc_119 N_A_27_413#_c_117_n N_A_211_413#_c_313_n 0.0150624f $X=1.435 $Y=0.805
+ $X2=0 $Y2=0
cc_120 N_A_27_413#_c_118_n N_A_211_413#_c_313_n 0.00281191f $X=1.51 $Y=0.73
+ $X2=0 $Y2=0
cc_121 N_A_27_413#_c_119_n N_A_211_413#_c_313_n 0.0165286f $X=0.77 $Y=0.995
+ $X2=0 $Y2=0
cc_122 N_A_27_413#_c_127_n N_A_211_413#_c_313_n 0.0141267f $X=0.77 $Y=1.83 $X2=0
+ $Y2=0
cc_123 N_A_27_413#_c_120_n N_A_211_413#_c_313_n 0.02509f $X=0.94 $Y=1.16 $X2=0
+ $Y2=0
cc_124 N_A_27_413#_c_117_n N_A_211_413#_c_338_n 0.00187101f $X=1.435 $Y=0.805
+ $X2=0 $Y2=0
cc_125 N_A_27_413#_c_162_p N_A_211_413#_c_338_n 0.0149168f $X=0.73 $Y=0.42 $X2=0
+ $Y2=0
cc_126 N_A_27_413#_c_123_n N_VPWR_c_430_n 0.00973767f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_127 N_A_27_413#_c_124_n N_VPWR_c_430_n 0.0201569f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_128 N_A_27_413#_c_125_n N_VPWR_c_430_n 0.0209571f $X=0.685 $Y=1.915 $X2=0
+ $Y2=0
cc_129 N_A_27_413#_c_124_n N_VPWR_c_436_n 0.0117547f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_130 N_A_27_413#_c_125_n N_VPWR_c_436_n 0.00239659f $X=0.685 $Y=1.915 $X2=0
+ $Y2=0
cc_131 N_A_27_413#_c_123_n N_VPWR_c_439_n 0.00643335f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_132 N_A_27_413#_c_123_n N_VPWR_c_440_n 0.00255931f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_133 N_A_27_413#_M1001_s N_VPWR_c_429_n 0.0038794f $X=0.135 $Y=2.065 $X2=0
+ $Y2=0
cc_134 N_A_27_413#_c_123_n N_VPWR_c_429_n 0.0119419f $X=0.965 $Y=1.99 $X2=0
+ $Y2=0
cc_135 N_A_27_413#_c_124_n N_VPWR_c_429_n 0.00645836f $X=0.26 $Y=2.3 $X2=0 $Y2=0
cc_136 N_A_27_413#_c_125_n N_VPWR_c_429_n 0.0053989f $X=0.685 $Y=1.915 $X2=0
+ $Y2=0
cc_137 N_A_27_413#_c_116_n N_VGND_c_547_n 0.00528256f $X=0.965 $Y=1.325 $X2=0
+ $Y2=0
cc_138 N_A_27_413#_c_117_n N_VGND_c_547_n 7.2576e-19 $X=1.435 $Y=0.805 $X2=0
+ $Y2=0
cc_139 N_A_27_413#_c_118_n N_VGND_c_547_n 0.00585385f $X=1.51 $Y=0.73 $X2=0
+ $Y2=0
cc_140 N_A_27_413#_c_162_p N_VGND_c_547_n 0.0143008f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_141 N_A_27_413#_M1008_d N_VGND_c_550_n 0.00382094f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_142 N_A_27_413#_c_116_n N_VGND_c_550_n 0.00733702f $X=0.965 $Y=1.325 $X2=0
+ $Y2=0
cc_143 N_A_27_413#_c_118_n N_VGND_c_550_n 0.0120642f $X=1.51 $Y=0.73 $X2=0 $Y2=0
cc_144 N_A_27_413#_c_162_p N_VGND_c_550_n 0.00798371f $X=0.73 $Y=0.42 $X2=0
+ $Y2=0
cc_145 N_B_c_186_n N_C_c_224_n 0.00467623f $X=1.945 $Y=1.89 $X2=0 $Y2=0
cc_146 B N_C_c_224_n 0.00370141f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_147 N_B_c_185_n N_C_c_224_n 0.0185442f $X=1.98 $Y=1.24 $X2=0 $Y2=0
cc_148 N_B_c_187_n N_C_c_225_n 0.0191617f $X=1.945 $Y=1.99 $X2=0 $Y2=0
cc_149 N_B_M1005_g N_C_M1013_g 0.0230566f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_150 B N_C_M1013_g 0.0019513f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_151 N_B_M1005_g C 0.00166657f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_152 N_B_c_183_n C 2.71585e-19 $X=1.98 $Y=1.21 $X2=0 $Y2=0
cc_153 B C 0.0775767f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_154 N_B_c_185_n C 9.32012e-19 $X=1.98 $Y=1.24 $X2=0 $Y2=0
cc_155 N_B_M1005_g N_C_c_223_n 0.0026834f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_156 N_B_c_183_n N_C_c_223_n 0.0153546f $X=1.98 $Y=1.21 $X2=0 $Y2=0
cc_157 B N_C_c_223_n 0.00209969f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_158 N_B_c_187_n N_A_211_413#_c_340_n 0.00486536f $X=1.945 $Y=1.99 $X2=0 $Y2=0
cc_159 N_B_c_187_n N_A_211_413#_c_318_n 0.01606f $X=1.945 $Y=1.99 $X2=0 $Y2=0
cc_160 N_B_c_188_n N_A_211_413#_c_318_n 4.87475e-19 $X=1.98 $Y=1.745 $X2=0 $Y2=0
cc_161 B N_A_211_413#_c_318_n 0.0202382f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_162 N_B_c_187_n N_A_211_413#_c_322_n 4.35297e-19 $X=1.945 $Y=1.99 $X2=0 $Y2=0
cc_163 N_B_c_188_n N_A_211_413#_c_322_n 0.00814131f $X=1.98 $Y=1.745 $X2=0 $Y2=0
cc_164 N_B_M1005_g N_A_211_413#_c_313_n 0.00853411f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_165 B N_A_211_413#_c_313_n 0.0400781f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_166 N_B_c_187_n N_VPWR_c_440_n 0.0234005f $X=1.945 $Y=1.99 $X2=0 $Y2=0
cc_167 N_B_M1005_g N_VGND_c_547_n 0.00456292f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_168 B N_VGND_c_547_n 0.00765038f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_169 N_B_M1005_g N_VGND_c_550_n 0.00767831f $X=1.92 $Y=0.445 $X2=0 $Y2=0
cc_170 B N_VGND_c_550_n 0.00854438f $X=1.94 $Y=0.425 $X2=0 $Y2=0
cc_171 B A_399_47# 0.00368299f $X=1.94 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_172 N_C_c_224_n N_D_c_267_n 0.0144696f $X=2.495 $Y=1.89 $X2=0 $Y2=0
cc_173 C N_D_c_267_n 7.61769e-19 $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_174 N_C_c_225_n N_D_c_268_n 0.0240947f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_175 N_C_M1013_g N_D_M1002_g 0.030986f $X=2.52 $Y=0.445 $X2=0 $Y2=0
cc_176 C N_D_M1002_g 8.37536e-19 $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_177 N_C_M1013_g D 0.0032739f $X=2.52 $Y=0.445 $X2=0 $Y2=0
cc_178 C D 0.0783954f $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_179 C N_D_c_266_n 9.58467e-19 $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_180 N_C_c_223_n N_D_c_266_n 0.0196168f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_181 N_C_c_225_n N_A_211_413#_c_318_n 0.0151847f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_182 C N_A_211_413#_c_318_n 0.0118144f $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_183 N_C_c_223_n N_A_211_413#_c_318_n 0.00130845f $X=2.46 $Y=1.16 $X2=0 $Y2=0
cc_184 N_C_c_224_n N_A_211_413#_c_319_n 0.0036668f $X=2.495 $Y=1.89 $X2=0 $Y2=0
cc_185 N_C_c_225_n N_A_211_413#_c_352_n 0.00418471f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_186 N_C_c_225_n N_VPWR_c_434_n 0.00456002f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_187 N_C_c_225_n N_VPWR_c_440_n 0.00834198f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_188 N_C_c_225_n N_VPWR_c_429_n 0.00520553f $X=2.495 $Y=1.99 $X2=0 $Y2=0
cc_189 N_C_M1013_g N_VGND_c_546_n 0.00206181f $X=2.52 $Y=0.445 $X2=0 $Y2=0
cc_190 N_C_M1013_g N_VGND_c_547_n 0.0038979f $X=2.52 $Y=0.445 $X2=0 $Y2=0
cc_191 C N_VGND_c_547_n 0.00659474f $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_192 N_C_M1013_g N_VGND_c_550_n 0.0060513f $X=2.52 $Y=0.445 $X2=0 $Y2=0
cc_193 C N_VGND_c_550_n 0.00759195f $X=2.425 $Y=0.425 $X2=0 $Y2=0
cc_194 C A_399_47# 0.00255245f $X=2.425 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_195 N_D_c_267_n N_A_211_413#_c_316_n 0.0182228f $X=2.99 $Y=1.89 $X2=0 $Y2=0
cc_196 N_D_c_268_n N_A_211_413#_c_316_n 0.0135715f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_197 D N_A_211_413#_c_316_n 5.43348e-19 $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_198 N_D_M1002_g N_A_211_413#_c_311_n 0.0196542f $X=3.015 $Y=0.445 $X2=0 $Y2=0
cc_199 D N_A_211_413#_c_311_n 0.00276322f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_200 N_D_c_268_n N_A_211_413#_c_319_n 0.00336482f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_201 D N_A_211_413#_c_319_n 0.00664914f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_202 N_D_c_267_n N_A_211_413#_c_320_n 0.00671928f $X=2.99 $Y=1.89 $X2=0 $Y2=0
cc_203 N_D_c_268_n N_A_211_413#_c_320_n 0.00830855f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_204 D N_A_211_413#_c_320_n 0.0188919f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_205 N_D_c_267_n N_A_211_413#_c_321_n 0.00466672f $X=2.99 $Y=1.89 $X2=0 $Y2=0
cc_206 D N_A_211_413#_c_321_n 0.0219044f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_207 D N_A_211_413#_c_314_n 0.0258756f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_208 N_D_c_266_n N_A_211_413#_c_314_n 0.0010244f $X=2.955 $Y=1.16 $X2=0 $Y2=0
cc_209 N_D_c_267_n N_A_211_413#_c_315_n 0.00284235f $X=2.99 $Y=1.89 $X2=0 $Y2=0
cc_210 D N_A_211_413#_c_315_n 0.00125042f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_211 N_D_c_266_n N_A_211_413#_c_315_n 0.0177661f $X=2.955 $Y=1.16 $X2=0 $Y2=0
cc_212 N_D_c_268_n N_VPWR_c_431_n 0.00632419f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_213 N_D_c_268_n N_VPWR_c_434_n 0.00563419f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_214 N_D_c_268_n N_VPWR_c_440_n 0.00108755f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_215 N_D_c_268_n N_VPWR_c_429_n 0.00787625f $X=2.99 $Y=1.99 $X2=0 $Y2=0
cc_216 D X 0.00707525f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_217 N_D_M1002_g N_X_c_506_n 6.16236e-19 $X=3.015 $Y=0.445 $X2=0 $Y2=0
cc_218 D X 0.00567546f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_219 N_D_M1002_g N_VGND_c_546_n 0.0128076f $X=3.015 $Y=0.445 $X2=0 $Y2=0
cc_220 D N_VGND_c_546_n 0.00589357f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_221 N_D_M1002_g N_VGND_c_547_n 0.00198995f $X=3.015 $Y=0.445 $X2=0 $Y2=0
cc_222 D N_VGND_c_547_n 0.00360847f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_223 N_D_M1002_g N_VGND_c_550_n 0.00285201f $X=3.015 $Y=0.445 $X2=0 $Y2=0
cc_224 D N_VGND_c_550_n 0.00685945f $X=2.79 $Y=0.765 $X2=0 $Y2=0
cc_225 D A_519_47# 0.00188003f $X=2.79 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_226 N_A_211_413#_c_318_n N_VPWR_M1006_d 0.00262418f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_227 N_A_211_413#_c_320_n N_VPWR_M1000_d 0.00664488f $X=3.295 $Y=1.88 $X2=0
+ $Y2=0
cc_228 N_A_211_413#_c_321_n N_VPWR_M1000_d 0.00325377f $X=3.38 $Y=1.795 $X2=0
+ $Y2=0
cc_229 N_A_211_413#_c_340_n N_VPWR_c_430_n 0.0165263f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_230 N_A_211_413#_c_316_n N_VPWR_c_431_n 0.00855809f $X=3.54 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_211_413#_c_317_n N_VPWR_c_431_n 9.49425e-19 $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_232 N_A_211_413#_c_320_n N_VPWR_c_431_n 0.0166758f $X=3.295 $Y=1.88 $X2=0
+ $Y2=0
cc_233 N_A_211_413#_c_317_n N_VPWR_c_433_n 0.00704965f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_211_413#_c_318_n N_VPWR_c_434_n 0.0036485f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_235 N_A_211_413#_c_352_n N_VPWR_c_434_n 0.0126306f $X=2.755 $Y=2.3 $X2=0
+ $Y2=0
cc_236 N_A_211_413#_c_320_n N_VPWR_c_434_n 0.00365041f $X=3.295 $Y=1.88 $X2=0
+ $Y2=0
cc_237 N_A_211_413#_c_316_n N_VPWR_c_437_n 0.00622633f $X=3.54 $Y=1.41 $X2=0
+ $Y2=0
cc_238 N_A_211_413#_c_317_n N_VPWR_c_437_n 0.00643255f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_239 N_A_211_413#_c_340_n N_VPWR_c_439_n 0.0118139f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_240 N_A_211_413#_c_318_n N_VPWR_c_439_n 0.00506621f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_241 N_A_211_413#_c_322_n N_VPWR_c_439_n 0.00249276f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_242 N_A_211_413#_M1011_d N_VPWR_c_440_n 0.00466001f $X=1.055 $Y=2.065 $X2=0
+ $Y2=0
cc_243 N_A_211_413#_c_340_n N_VPWR_c_440_n 0.00875114f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_244 N_A_211_413#_c_318_n N_VPWR_c_440_n 0.0406458f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_245 N_A_211_413#_c_352_n N_VPWR_c_440_n 0.0125331f $X=2.755 $Y=2.3 $X2=0
+ $Y2=0
cc_246 N_A_211_413#_M1011_d N_VPWR_c_429_n 0.00865828f $X=1.055 $Y=2.065 $X2=0
+ $Y2=0
cc_247 N_A_211_413#_M1009_d N_VPWR_c_429_n 0.0030151f $X=2.585 $Y=2.065 $X2=0
+ $Y2=0
cc_248 N_A_211_413#_c_316_n N_VPWR_c_429_n 0.0104879f $X=3.54 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_211_413#_c_317_n N_VPWR_c_429_n 0.0121535f $X=4.045 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_211_413#_c_340_n N_VPWR_c_429_n 0.00646998f $X=1.2 $Y=2.3 $X2=0 $Y2=0
cc_251 N_A_211_413#_c_318_n N_VPWR_c_429_n 0.0174406f $X=2.67 $Y=2 $X2=0 $Y2=0
cc_252 N_A_211_413#_c_352_n N_VPWR_c_429_n 0.00723365f $X=2.755 $Y=2.3 $X2=0
+ $Y2=0
cc_253 N_A_211_413#_c_320_n N_VPWR_c_429_n 0.00774161f $X=3.295 $Y=1.88 $X2=0
+ $Y2=0
cc_254 N_A_211_413#_c_322_n N_VPWR_c_429_n 0.00388138f $X=1.265 $Y=2 $X2=0 $Y2=0
cc_255 N_A_211_413#_c_317_n X 0.0172663f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_211_413#_c_320_n X 0.0112115f $X=3.295 $Y=1.88 $X2=0 $Y2=0
cc_257 N_A_211_413#_c_311_n X 0.0104255f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A_211_413#_c_312_n X 0.0118029f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_211_413#_c_315_n X 0.00194336f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_260 N_A_211_413#_c_316_n X 0.00920579f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_211_413#_c_317_n X 0.0135312f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_211_413#_c_321_n X 0.015893f $X=3.38 $Y=1.795 $X2=0 $Y2=0
cc_263 N_A_211_413#_c_315_n X 0.00372299f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_264 N_A_211_413#_c_311_n N_X_c_506_n 0.00807166f $X=3.565 $Y=0.995 $X2=0
+ $Y2=0
cc_265 N_A_211_413#_c_312_n N_X_c_506_n 0.0045409f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_211_413#_c_316_n X 0.00119264f $X=3.54 $Y=1.41 $X2=0 $Y2=0
cc_267 N_A_211_413#_c_311_n X 0.00248829f $X=3.565 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_211_413#_c_317_n X 0.0057162f $X=4.045 $Y=1.41 $X2=0 $Y2=0
cc_269 N_A_211_413#_c_312_n X 0.00755537f $X=4.07 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_211_413#_c_321_n X 0.0106754f $X=3.38 $Y=1.795 $X2=0 $Y2=0
cc_271 N_A_211_413#_c_314_n X 0.0209276f $X=3.47 $Y=1.16 $X2=0 $Y2=0
cc_272 N_A_211_413#_c_315_n X 0.0360858f $X=4.045 $Y=1.202 $X2=0 $Y2=0
cc_273 N_A_211_413#_c_311_n N_VGND_c_546_n 0.00355157f $X=3.565 $Y=0.995 $X2=0
+ $Y2=0
cc_274 N_A_211_413#_c_314_n N_VGND_c_546_n 0.0033107f $X=3.47 $Y=1.16 $X2=0
+ $Y2=0
cc_275 N_A_211_413#_c_315_n N_VGND_c_546_n 9.74653e-19 $X=4.045 $Y=1.202 $X2=0
+ $Y2=0
cc_276 N_A_211_413#_c_338_n N_VGND_c_547_n 0.0139021f $X=1.3 $Y=0.42 $X2=0 $Y2=0
cc_277 N_A_211_413#_c_311_n N_VGND_c_548_n 0.00465454f $X=3.565 $Y=0.995 $X2=0
+ $Y2=0
cc_278 N_A_211_413#_c_312_n N_VGND_c_548_n 0.0019794f $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_279 N_A_211_413#_c_311_n N_VGND_c_549_n 5.24816e-19 $X=3.565 $Y=0.995 $X2=0
+ $Y2=0
cc_280 N_A_211_413#_c_312_n N_VGND_c_549_n 0.0110987f $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_281 N_A_211_413#_M1010_s N_VGND_c_550_n 0.00256467f $X=1.175 $Y=0.235 $X2=0
+ $Y2=0
cc_282 N_A_211_413#_c_311_n N_VGND_c_550_n 0.00838544f $X=3.565 $Y=0.995 $X2=0
+ $Y2=0
cc_283 N_A_211_413#_c_312_n N_VGND_c_550_n 0.00279076f $X=4.07 $Y=0.995 $X2=0
+ $Y2=0
cc_284 N_A_211_413#_c_338_n N_VGND_c_550_n 0.00836197f $X=1.3 $Y=0.42 $X2=0
+ $Y2=0
cc_285 N_VPWR_c_429_n N_X_M1004_d 0.0046766f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_c_431_n X 0.017087f $X=3.305 $Y=2.34 $X2=0 $Y2=0
cc_287 N_VPWR_c_433_n X 0.042057f $X=4.28 $Y=2 $X2=0 $Y2=0
cc_288 N_VPWR_c_437_n X 0.0192051f $X=4.195 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_429_n X 0.0114183f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_M1007_s X 0.00293f $X=4.135 $Y=1.485 $X2=0 $Y2=0
cc_291 N_VPWR_c_433_n X 0.0229665f $X=4.28 $Y=2 $X2=0 $Y2=0
cc_292 N_VPWR_M1007_s X 2.16973e-19 $X=4.135 $Y=1.485 $X2=0 $Y2=0
cc_293 X N_VGND_M1012_d 0.00300766f $X=4.22 $Y=0.765 $X2=0 $Y2=0
cc_294 X N_VGND_M1012_d 2.61253e-19 $X=3.905 $Y=0.85 $X2=0 $Y2=0
cc_295 N_X_c_506_n N_VGND_c_546_n 0.0164985f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_296 X N_VGND_c_548_n 0.00260748f $X=4.22 $Y=0.765 $X2=0 $Y2=0
cc_297 N_X_c_506_n N_VGND_c_548_n 0.0210913f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_298 X N_VGND_c_549_n 0.0266648f $X=4.22 $Y=0.765 $X2=0 $Y2=0
cc_299 N_X_c_506_n N_VGND_c_549_n 0.0165902f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_300 N_X_M1003_s N_VGND_c_550_n 0.00321778f $X=3.64 $Y=0.235 $X2=0 $Y2=0
cc_301 X N_VGND_c_550_n 0.0066116f $X=4.22 $Y=0.765 $X2=0 $Y2=0
cc_302 N_X_c_506_n N_VGND_c_550_n 0.0123534f $X=3.81 $Y=0.42 $X2=0 $Y2=0
cc_303 N_VGND_c_550_n A_317_47# 0.0111139f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_304 N_VGND_c_550_n A_399_47# 0.0115473f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_305 N_VGND_c_550_n A_519_47# 0.00936378f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
