* File: sky130_fd_sc_hdll__o32ai_4.pex.spice
* Created: Wed Sep  2 08:47:20 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%B2 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 46 47 55
r73 47 48 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.212
+ $X2=1.93 $Y2=1.212
r74 45 47 33.9132 $w=3.34e-07 $l=2.35e-07 $layer=POLY_cond $X=1.67 $Y=1.212
+ $X2=1.905 $Y2=1.212
r75 45 46 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=1.67
+ $Y=1.16 $X2=1.67 $Y2=1.16
r76 43 45 30.3054 $w=3.34e-07 $l=2.1e-07 $layer=POLY_cond $X=1.46 $Y=1.212
+ $X2=1.67 $Y2=1.212
r77 42 43 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.212
+ $X2=1.46 $Y2=1.212
r78 41 42 64.2186 $w=3.34e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.212
+ $X2=1.435 $Y2=1.212
r79 40 41 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.212
+ $X2=0.99 $Y2=1.212
r80 39 40 64.2186 $w=3.34e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.212
+ $X2=0.965 $Y2=1.212
r81 38 39 3.60778 $w=3.34e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.212
+ $X2=0.52 $Y2=1.212
r82 36 38 31.7485 $w=3.34e-07 $l=2.2e-07 $layer=POLY_cond $X=0.275 $Y=1.212
+ $X2=0.495 $Y2=1.212
r83 31 46 28.0045 $w=1.98e-07 $l=5.05e-07 $layer=LI1_cond $X=1.165 $Y=1.175
+ $X2=1.67 $Y2=1.175
r84 31 55 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=1.165 $Y=1.175
+ $X2=1.155 $Y2=1.175
r85 30 55 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.695 $Y=1.175
+ $X2=1.155 $Y2=1.175
r86 29 30 25.5091 $w=1.98e-07 $l=4.6e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.695 $Y2=1.175
r87 29 36 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.275
+ $Y=1.16 $X2=0.275 $Y2=1.16
r88 25 48 21.5099 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.93 $Y=1.015
+ $X2=1.93 $Y2=1.212
r89 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.93 $Y=1.015
+ $X2=1.93 $Y2=0.56
r90 22 47 17.2128 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.212
r91 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r92 18 43 21.5099 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=1.46 $Y=1.015
+ $X2=1.46 $Y2=1.212
r93 18 20 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=1.46 $Y=1.015
+ $X2=1.46 $Y2=0.56
r94 15 42 17.2128 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.212
r95 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r96 11 41 21.5099 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.99 $Y=1.015
+ $X2=0.99 $Y2=1.212
r97 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.99 $Y=1.015
+ $X2=0.99 $Y2=0.56
r98 8 40 17.2128 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.212
r99 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r100 4 39 21.5099 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=1.212
r101 4 6 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.52 $Y=1.015
+ $X2=0.52 $Y2=0.56
r102 1 38 17.2128 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.212
r103 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%B1 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 46 47 52 55 58
c68 27 0 1.98558e-19 $X=3.825 $Y=0.56
r69 47 48 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=3.8 $Y=1.212
+ $X2=3.825 $Y2=1.212
r70 46 58 6.1 $w=1.98e-07 $l=1.1e-07 $layer=LI1_cond $X=3.565 $Y=1.175 $X2=3.455
+ $Y2=1.175
r71 45 47 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=3.565 $Y=1.212
+ $X2=3.8 $Y2=1.212
r72 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.565
+ $Y=1.16 $X2=3.565 $Y2=1.16
r73 43 45 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=3.33 $Y=1.212
+ $X2=3.565 $Y2=1.212
r74 42 43 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=3.305 $Y=1.212
+ $X2=3.33 $Y2=1.212
r75 41 42 62.7164 $w=3.42e-07 $l=4.45e-07 $layer=POLY_cond $X=2.86 $Y=1.212
+ $X2=3.305 $Y2=1.212
r76 40 41 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=2.835 $Y=1.212
+ $X2=2.86 $Y2=1.212
r77 38 40 30.3012 $w=3.42e-07 $l=2.15e-07 $layer=POLY_cond $X=2.62 $Y=1.212
+ $X2=2.835 $Y2=1.212
r78 38 52 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.62
+ $Y=1.16 $X2=2.62 $Y2=1.16
r79 36 38 32.4152 $w=3.42e-07 $l=2.3e-07 $layer=POLY_cond $X=2.39 $Y=1.212
+ $X2=2.62 $Y2=1.212
r80 35 36 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=2.365 $Y=1.212
+ $X2=2.39 $Y2=1.212
r81 31 58 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.175
+ $X2=3.455 $Y2=1.175
r82 31 55 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=3.45 $Y=1.175
+ $X2=2.995 $Y2=1.175
r83 30 55 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.99 $Y=1.175
+ $X2=2.995 $Y2=1.175
r84 30 52 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=2.99 $Y=1.175
+ $X2=2.535 $Y2=1.175
r85 29 52 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.175
+ $X2=2.535 $Y2=1.175
r86 25 48 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=3.825 $Y=1.015
+ $X2=3.825 $Y2=1.212
r87 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.825 $Y=1.015
+ $X2=3.825 $Y2=0.56
r88 22 47 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=3.8 $Y=1.41 $X2=3.8
+ $Y2=1.212
r89 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.8 $Y=1.41 $X2=3.8
+ $Y2=1.985
r90 19 43 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=3.33 $Y=1.41
+ $X2=3.33 $Y2=1.212
r91 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.33 $Y=1.41
+ $X2=3.33 $Y2=1.985
r92 15 42 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=3.305 $Y=1.015
+ $X2=3.305 $Y2=1.212
r93 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=3.305 $Y=1.015
+ $X2=3.305 $Y2=0.56
r94 12 41 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=2.86 $Y=1.41
+ $X2=2.86 $Y2=1.212
r95 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.86 $Y=1.41
+ $X2=2.86 $Y2=1.985
r96 8 40 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=2.835 $Y=1.015
+ $X2=2.835 $Y2=1.212
r97 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.835 $Y=1.015
+ $X2=2.835 $Y2=0.56
r98 5 36 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=2.39 $Y=1.41
+ $X2=2.39 $Y2=1.212
r99 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.39 $Y=1.41 $X2=2.39
+ $Y2=1.985
r100 1 35 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=2.365 $Y=1.015
+ $X2=2.365 $Y2=1.212
r101 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=2.365 $Y=1.015
+ $X2=2.365 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A3 3 7 9 11 14 16 18 19 21 24 26 28 29 30
+ 31 32 33 38 50 55 58 61 63
c87 33 0 1.52421e-19 $X=5.675 $Y=1.105
r88 61 63 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=5.295 $Y=1.175
+ $X2=5.745 $Y2=1.175
r89 50 51 54.5794 $w=3.4e-07 $l=3.85e-07 $layer=POLY_cond $X=5.815 $Y=1.212
+ $X2=6.2 $Y2=1.212
r90 48 50 9.92353 $w=3.4e-07 $l=7e-08 $layer=POLY_cond $X=5.745 $Y=1.212
+ $X2=5.815 $Y2=1.212
r91 48 63 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.745
+ $Y=1.16 $X2=5.745 $Y2=1.16
r92 46 48 2.12647 $w=3.4e-07 $l=1.5e-08 $layer=POLY_cond $X=5.73 $Y=1.212
+ $X2=5.745 $Y2=1.212
r93 45 46 66.6294 $w=3.4e-07 $l=4.7e-07 $layer=POLY_cond $X=5.26 $Y=1.212
+ $X2=5.73 $Y2=1.212
r94 44 45 10.6324 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=5.185 $Y=1.212
+ $X2=5.26 $Y2=1.212
r95 43 44 55.9971 $w=3.4e-07 $l=3.95e-07 $layer=POLY_cond $X=4.79 $Y=1.212
+ $X2=5.185 $Y2=1.212
r96 42 43 10.6324 $w=3.4e-07 $l=7.5e-08 $layer=POLY_cond $X=4.715 $Y=1.212
+ $X2=4.79 $Y2=1.212
r97 38 42 11.8119 $w=3.4e-07 $l=9.75961e-08 $layer=POLY_cond $X=4.64 $Y=1.16
+ $X2=4.715 $Y2=1.212
r98 38 40 63.0897 $w=2.9e-07 $l=3.05e-07 $layer=POLY_cond $X=4.64 $Y=1.16
+ $X2=4.335 $Y2=1.16
r99 33 63 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=5.76 $Y=1.175
+ $X2=5.745 $Y2=1.175
r100 32 61 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=5.27 $Y=1.175
+ $X2=5.295 $Y2=1.175
r101 32 58 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=5.27 $Y=1.175
+ $X2=4.835 $Y2=1.175
r102 31 58 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=4.825 $Y=1.175
+ $X2=4.835 $Y2=1.175
r103 31 55 24.9545 $w=1.98e-07 $l=4.5e-07 $layer=LI1_cond $X=4.825 $Y=1.175
+ $X2=4.375 $Y2=1.175
r104 30 55 2.21818 $w=1.98e-07 $l=4e-08 $layer=LI1_cond $X=4.335 $Y=1.175
+ $X2=4.375 $Y2=1.175
r105 30 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.335
+ $Y=1.16 $X2=4.335 $Y2=1.16
r106 29 40 3.10277 $w=2.9e-07 $l=1.5e-08 $layer=POLY_cond $X=4.32 $Y=1.16
+ $X2=4.335 $Y2=1.16
r107 26 51 17.6285 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.212
r108 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.2 $Y=1.41
+ $X2=6.2 $Y2=1.985
r109 22 50 21.9347 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.815 $Y=1.015
+ $X2=5.815 $Y2=1.212
r110 22 24 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.815 $Y=1.015
+ $X2=5.815 $Y2=0.56
r111 19 46 17.6285 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.212
r112 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.73 $Y=1.41
+ $X2=5.73 $Y2=1.985
r113 16 45 17.6285 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.212
r114 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.985
r115 12 44 21.9347 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.185 $Y=1.015
+ $X2=5.185 $Y2=1.212
r116 12 14 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.185 $Y=1.015
+ $X2=5.185 $Y2=0.56
r117 9 43 17.6285 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.212
r118 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.985
r119 5 42 21.9347 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=4.715 $Y=1.015
+ $X2=4.715 $Y2=1.212
r120 5 7 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.715 $Y=1.015
+ $X2=4.715 $Y2=0.56
r121 1 29 30.6382 $w=2.9e-07 $l=1.78606e-07 $layer=POLY_cond $X=4.245 $Y=1.015
+ $X2=4.32 $Y2=1.16
r122 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=4.245 $Y=1.015
+ $X2=4.245 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A2 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 46 47 52 56 58
c77 47 0 1.52421e-19 $X=8.08 $Y=1.212
r78 56 58 23.8455 $w=1.98e-07 $l=4.3e-07 $layer=LI1_cond $X=7.135 $Y=1.175
+ $X2=7.565 $Y2=1.175
r79 47 48 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=8.08 $Y=1.212
+ $X2=8.105 $Y2=1.212
r80 45 47 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=7.845 $Y=1.212
+ $X2=8.08 $Y2=1.212
r81 45 46 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=7.845
+ $Y=1.16 $X2=7.845 $Y2=1.16
r82 43 45 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=7.61 $Y=1.212
+ $X2=7.845 $Y2=1.212
r83 42 43 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=7.585 $Y=1.212
+ $X2=7.61 $Y2=1.212
r84 41 42 62.7164 $w=3.42e-07 $l=4.45e-07 $layer=POLY_cond $X=7.14 $Y=1.212
+ $X2=7.585 $Y2=1.212
r85 40 41 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=7.115 $Y=1.212
+ $X2=7.14 $Y2=1.212
r86 39 52 12.7545 $w=1.98e-07 $l=2.3e-07 $layer=LI1_cond $X=6.905 $Y=1.175
+ $X2=6.675 $Y2=1.175
r87 38 40 29.5965 $w=3.42e-07 $l=2.1e-07 $layer=POLY_cond $X=6.905 $Y=1.212
+ $X2=7.115 $Y2=1.212
r88 38 39 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=6.905
+ $Y=1.16 $X2=6.905 $Y2=1.16
r89 36 38 33.1199 $w=3.42e-07 $l=2.35e-07 $layer=POLY_cond $X=6.67 $Y=1.212
+ $X2=6.905 $Y2=1.212
r90 35 36 3.52339 $w=3.42e-07 $l=2.5e-08 $layer=POLY_cond $X=6.645 $Y=1.212
+ $X2=6.67 $Y2=1.212
r91 31 46 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=7.58 $Y=1.175
+ $X2=7.845 $Y2=1.175
r92 31 58 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=7.58 $Y=1.175
+ $X2=7.565 $Y2=1.175
r93 30 56 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=7.125 $Y=1.175
+ $X2=7.135 $Y2=1.175
r94 30 39 12.2 $w=1.98e-07 $l=2.2e-07 $layer=LI1_cond $X=7.125 $Y=1.175
+ $X2=6.905 $Y2=1.175
r95 29 52 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=6.665 $Y=1.175
+ $X2=6.675 $Y2=1.175
r96 25 48 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=8.105 $Y=1.015
+ $X2=8.105 $Y2=1.212
r97 25 27 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=8.105 $Y=1.015
+ $X2=8.105 $Y2=0.56
r98 22 47 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=8.08 $Y=1.41
+ $X2=8.08 $Y2=1.212
r99 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.08 $Y=1.41
+ $X2=8.08 $Y2=1.985
r100 19 43 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.212
r101 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.61 $Y=1.41
+ $X2=7.61 $Y2=1.985
r102 15 42 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=7.585 $Y=1.015
+ $X2=7.585 $Y2=1.212
r103 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.585 $Y=1.015
+ $X2=7.585 $Y2=0.56
r104 12 41 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.212
r105 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.14 $Y=1.41
+ $X2=7.14 $Y2=1.985
r106 8 40 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=7.115 $Y=1.015
+ $X2=7.115 $Y2=1.212
r107 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=7.115 $Y=1.015
+ $X2=7.115 $Y2=0.56
r108 5 36 17.7656 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.212
r109 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.67 $Y=1.41
+ $X2=6.67 $Y2=1.985
r110 1 35 22.0749 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=6.645 $Y=1.015
+ $X2=6.645 $Y2=1.212
r111 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=6.645 $Y=1.015
+ $X2=6.645 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A1 3 5 7 10 12 14 17 19 21 22 23 26 28 30
+ 31 32 33 34 49 57 60 63
r78 52 63 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=10.615 $Y=1.175
+ $X2=10.35 $Y2=1.175
r79 51 52 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=10.615
+ $Y=1.16 $X2=10.615 $Y2=1.16
r80 49 51 12.7214 $w=3.41e-07 $l=9e-08 $layer=POLY_cond $X=10.525 $Y=1.212
+ $X2=10.615 $Y2=1.212
r81 48 49 3.53372 $w=3.41e-07 $l=2.5e-08 $layer=POLY_cond $X=10.5 $Y=1.212
+ $X2=10.525 $Y2=1.212
r82 46 47 3.49275 $w=3.45e-07 $l=2.5e-08 $layer=POLY_cond $X=9.985 $Y=1.212
+ $X2=10.01 $Y2=1.212
r83 45 46 62.171 $w=3.45e-07 $l=4.45e-07 $layer=POLY_cond $X=9.54 $Y=1.212
+ $X2=9.985 $Y2=1.212
r84 44 45 3.49275 $w=3.45e-07 $l=2.5e-08 $layer=POLY_cond $X=9.515 $Y=1.212
+ $X2=9.54 $Y2=1.212
r85 42 44 29.3391 $w=3.45e-07 $l=2.1e-07 $layer=POLY_cond $X=9.305 $Y=1.212
+ $X2=9.515 $Y2=1.212
r86 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=9.305
+ $Y=1.16 $X2=9.305 $Y2=1.16
r87 40 42 32.8319 $w=3.45e-07 $l=2.35e-07 $layer=POLY_cond $X=9.07 $Y=1.212
+ $X2=9.305 $Y2=1.212
r88 39 40 3.49275 $w=3.45e-07 $l=2.5e-08 $layer=POLY_cond $X=9.045 $Y=1.212
+ $X2=9.07 $Y2=1.212
r89 34 52 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=10.805 $Y=1.175
+ $X2=10.615 $Y2=1.175
r90 33 63 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=10.345 $Y=1.175
+ $X2=10.35 $Y2=1.175
r91 33 60 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=10.345 $Y=1.175
+ $X2=9.91 $Y2=1.175
r92 32 60 0.831818 $w=1.98e-07 $l=1.5e-08 $layer=LI1_cond $X=9.895 $Y=1.175
+ $X2=9.91 $Y2=1.175
r93 32 57 24.4 $w=1.98e-07 $l=4.4e-07 $layer=LI1_cond $X=9.895 $Y=1.175
+ $X2=9.455 $Y2=1.175
r94 31 57 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=9.43 $Y=1.175
+ $X2=9.455 $Y2=1.175
r95 31 43 6.93182 $w=1.98e-07 $l=1.25e-07 $layer=LI1_cond $X=9.43 $Y=1.175
+ $X2=9.305 $Y2=1.175
r96 28 49 17.6972 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=10.525 $Y=1.41
+ $X2=10.525 $Y2=1.212
r97 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.525 $Y=1.41
+ $X2=10.525 $Y2=1.985
r98 24 48 22.0049 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=10.5 $Y=1.015
+ $X2=10.5 $Y2=1.212
r99 24 26 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=10.5 $Y=1.015
+ $X2=10.5 $Y2=0.56
r100 23 47 15.3369 $w=3.45e-07 $l=1.23288e-07 $layer=POLY_cond $X=10.11 $Y=1.16
+ $X2=10.01 $Y2=1.212
r101 22 48 11.8174 $w=3.41e-07 $l=9.75961e-08 $layer=POLY_cond $X=10.425 $Y=1.16
+ $X2=10.5 $Y2=1.212
r102 22 23 65.1582 $w=2.9e-07 $l=3.15e-07 $layer=POLY_cond $X=10.425 $Y=1.16
+ $X2=10.11 $Y2=1.16
r103 19 47 17.97 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.212
r104 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.985
r105 15 46 22.2839 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=9.985 $Y=1.015
+ $X2=9.985 $Y2=1.212
r106 15 17 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.985 $Y=1.015
+ $X2=9.985 $Y2=0.56
r107 12 45 17.97 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.212
r108 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.985
r109 8 44 22.2839 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=9.515 $Y=1.015
+ $X2=9.515 $Y2=1.212
r110 8 10 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.515 $Y=1.015
+ $X2=9.515 $Y2=0.56
r111 5 40 17.97 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=9.07 $Y=1.41 $X2=9.07
+ $Y2=1.212
r112 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.07 $Y=1.41
+ $X2=9.07 $Y2=1.985
r113 1 39 22.2839 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=1.212
r114 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=9.045 $Y=1.015
+ $X2=9.045 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_297# 1 2 3 4 5 16 18 20 24 26 31 32
+ 33 36 38 40 42 47 49
c77 3 0 3.29093e-19 $X=1.995 $Y=1.485
r78 40 51 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=2.005
+ $X2=4.075 $Y2=1.92
r79 40 42 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.075 $Y=2.005
+ $X2=4.075 $Y2=2.26
r80 39 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=1.92
+ $X2=3.095 $Y2=1.92
r81 38 51 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=3.95 $Y=1.92
+ $X2=4.075 $Y2=1.92
r82 38 39 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.95 $Y=1.92
+ $X2=3.18 $Y2=1.92
r83 34 49 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.095 $Y=2.005
+ $X2=3.095 $Y2=1.92
r84 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=3.095 $Y=2.005
+ $X2=3.095 $Y2=2.26
r85 32 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.01 $Y=1.92
+ $X2=3.095 $Y2=1.92
r86 32 33 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=3.01 $Y=1.92
+ $X2=2.24 $Y2=1.92
r87 29 31 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.155 $Y=2.255
+ $X2=2.155 $Y2=2.17
r88 28 33 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.155 $Y=2.005
+ $X2=2.24 $Y2=1.92
r89 28 31 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=2.155 $Y=2.005
+ $X2=2.155 $Y2=2.17
r90 27 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.36 $X2=1.2
+ $Y2=2.36
r91 26 29 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.07 $Y=2.36
+ $X2=2.155 $Y2=2.255
r92 26 27 41.4589 $w=2.08e-07 $l=7.85e-07 $layer=LI1_cond $X=2.07 $Y=2.36
+ $X2=1.285 $Y2=2.36
r93 22 47 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=1.2 $Y=2.255 $X2=1.2
+ $Y2=2.36
r94 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=1.2 $Y=2.255
+ $X2=1.2 $Y2=2
r95 21 45 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=2.36
+ $X2=0.217 $Y2=2.36
r96 20 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.36 $X2=1.2
+ $Y2=2.36
r97 20 21 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.36
+ $X2=0.345 $Y2=2.36
r98 16 45 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.217 $Y=2.255
+ $X2=0.217 $Y2=2.36
r99 16 18 26.8903 $w=2.53e-07 $l=5.95e-07 $layer=LI1_cond $X=0.217 $Y=2.255
+ $X2=0.217 $Y2=1.66
r100 5 51 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.485 $X2=4.035 $Y2=1.92
r101 5 42 600 $w=1.7e-07 $l=8.44393e-07 $layer=licon1_PDIFF $count=1 $X=3.89
+ $Y=1.485 $X2=4.035 $Y2=2.26
r102 4 49 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.485 $X2=3.095 $Y2=1.92
r103 4 36 600 $w=1.7e-07 $l=8.44393e-07 $layer=licon1_PDIFF $count=1 $X=2.95
+ $Y=1.485 $X2=3.095 $Y2=2.26
r104 3 31 600 $w=1.7e-07 $l=7.60805e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.155 $Y2=2.17
r105 2 47 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2.34
r106 2 24 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r107 1 45 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r108 1 18 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%Y 1 2 3 4 5 6 7 8 25 33 35 38 43 45 49 54
+ 57 58 59 61 63 64
c129 45 0 1.29579e-19 $X=4.86 $Y=1.58
c130 38 0 1.99513e-19 $X=2.145 $Y=1.495
r131 55 64 5.98103 $w=3.93e-07 $l=2.05e-07 $layer=LI1_cond $X=1.652 $Y=1.665
+ $X2=1.652 $Y2=1.87
r132 55 57 1.43204 $w=3.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.652 $Y=1.665
+ $X2=1.652 $Y2=1.58
r133 50 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.19 $Y=1.58
+ $X2=5.025 $Y2=1.58
r134 49 63 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.75 $Y=1.58
+ $X2=5.94 $Y2=1.58
r135 49 50 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.75 $Y=1.58
+ $X2=5.19 $Y2=1.58
r136 46 59 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.235 $Y=1.58
+ $X2=2.145 $Y2=1.58
r137 45 61 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.86 $Y=1.58
+ $X2=5.025 $Y2=1.58
r138 45 46 171.257 $w=1.68e-07 $l=2.625e-06 $layer=LI1_cond $X=4.86 $Y=1.58
+ $X2=2.235 $Y2=1.58
r139 41 43 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=2.625 $Y=0.78
+ $X2=3.565 $Y2=0.78
r140 39 58 3.89906 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.235 $Y=0.78
+ $X2=2.145 $Y2=0.78
r141 39 41 17.9781 $w=2.48e-07 $l=3.9e-07 $layer=LI1_cond $X=2.235 $Y=0.78
+ $X2=2.625 $Y2=0.78
r142 38 59 1.13756 $w=1.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.145 $Y=1.495
+ $X2=2.145 $Y2=1.58
r143 37 58 2.54814 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=2.145 $Y=0.905
+ $X2=2.145 $Y2=0.78
r144 37 38 36.3535 $w=1.78e-07 $l=5.9e-07 $layer=LI1_cond $X=2.145 $Y=0.905
+ $X2=2.145 $Y2=1.495
r145 36 57 9.73034 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=1.85 $Y=1.58
+ $X2=1.652 $Y2=1.58
r146 35 59 5.41628 $w=1.7e-07 $l=9e-08 $layer=LI1_cond $X=2.055 $Y=1.58
+ $X2=2.145 $Y2=1.58
r147 35 36 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.055 $Y=1.58
+ $X2=1.85 $Y2=1.58
r148 34 54 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=1.58
+ $X2=0.705 $Y2=1.58
r149 33 57 9.73034 $w=1.7e-07 $l=1.97e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=1.652 $Y2=1.58
r150 33 34 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.58
+ $X2=0.895 $Y2=1.58
r151 27 30 43.3319 $w=2.48e-07 $l=9.4e-07 $layer=LI1_cond $X=0.73 $Y=0.78
+ $X2=1.67 $Y2=0.78
r152 25 58 3.89906 $w=2.5e-07 $l=9e-08 $layer=LI1_cond $X=2.055 $Y=0.78
+ $X2=2.145 $Y2=0.78
r153 25 30 17.7476 $w=2.48e-07 $l=3.85e-07 $layer=LI1_cond $X=2.055 $Y=0.78
+ $X2=1.67 $Y2=0.78
r154 8 63 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=5.82
+ $Y=1.485 $X2=5.965 $Y2=1.66
r155 7 61 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.485 $X2=5.025 $Y2=1.66
r156 6 57 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.66
r157 5 54 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
r158 4 43 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.38
+ $Y=0.235 $X2=3.565 $Y2=0.74
r159 3 41 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=2.44
+ $Y=0.235 $X2=2.625 $Y2=0.74
r160 2 30 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.74
r161 1 27 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%VPWR 1 2 3 4 5 18 22 26 30 32 34 39 40 42
+ 43 44 46 54 69 74 77 81
r149 80 81 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r150 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r151 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r152 72 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r153 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r154 69 80 4.01252 $w=1.7e-07 $l=1.82e-07 $layer=LI1_cond $X=10.675 $Y=2.72
+ $X2=10.857 $Y2=2.72
r155 69 71 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=10.675 $Y=2.72
+ $X2=10.35 $Y2=2.72
r156 68 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r157 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r158 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r159 64 65 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r160 62 65 1.30889 $w=4.8e-07 $l=4.6e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=8.51 $Y2=2.72
r161 62 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=3.45 $Y2=2.72
r162 61 64 300.107 $w=1.68e-07 $l=4.6e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=8.51 $Y2=2.72
r163 61 62 1.69091 $w=1.7e-07 $l=9.35e-07 $layer=mcon $count=5 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r164 59 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.54 $Y2=2.72
r165 59 61 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=3.73 $Y=2.72
+ $X2=3.91 $Y2=2.72
r166 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r167 58 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r168 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r169 55 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.79 $Y=2.72 $X2=2.6
+ $Y2=2.72
r170 55 57 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=2.79 $Y=2.72 $X2=2.99
+ $Y2=2.72
r171 54 77 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.35 $Y=2.72
+ $X2=3.54 $Y2=2.72
r172 54 57 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=3.35 $Y=2.72
+ $X2=2.99 $Y2=2.72
r173 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r174 52 53 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r175 48 52 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r176 46 74 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.41 $Y=2.72 $X2=2.6
+ $Y2=2.72
r177 46 52 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=2.41 $Y=2.72
+ $X2=2.07 $Y2=2.72
r178 44 53 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r179 44 48 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r180 42 67 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.43 $Y2=2.72
r181 42 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.775 $Y2=2.72
r182 41 71 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=10.35 $Y2=2.72
r183 41 43 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=9.775 $Y2=2.72
r184 39 64 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=8.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r185 39 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.67 $Y=2.72
+ $X2=8.795 $Y2=2.72
r186 38 67 33.2727 $w=1.68e-07 $l=5.1e-07 $layer=LI1_cond $X=8.92 $Y=2.72
+ $X2=9.43 $Y2=2.72
r187 38 40 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=8.92 $Y=2.72
+ $X2=8.795 $Y2=2.72
r188 34 37 31.3464 $w=2.48e-07 $l=6.8e-07 $layer=LI1_cond $X=10.8 $Y=1.66
+ $X2=10.8 $Y2=2.34
r189 32 80 3.13065 $w=2.5e-07 $l=1.09864e-07 $layer=LI1_cond $X=10.8 $Y=2.635
+ $X2=10.857 $Y2=2.72
r190 32 37 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=10.8 $Y=2.635
+ $X2=10.8 $Y2=2.34
r191 28 43 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=2.72
r192 28 30 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=2
r193 24 40 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.795 $Y=2.635
+ $X2=8.795 $Y2=2.72
r194 24 26 29.2721 $w=2.48e-07 $l=6.35e-07 $layer=LI1_cond $X=8.795 $Y=2.635
+ $X2=8.795 $Y2=2
r195 20 77 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=3.54 $Y=2.635
+ $X2=3.54 $Y2=2.72
r196 20 22 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=3.54 $Y=2.635
+ $X2=3.54 $Y2=2.34
r197 16 74 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.6 $Y=2.635 $X2=2.6
+ $Y2=2.72
r198 16 18 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.6 $Y=2.635
+ $X2=2.6 $Y2=2.34
r199 5 37 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.485 $X2=10.76 $Y2=2.34
r200 5 34 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.615
+ $Y=1.485 $X2=10.76 $Y2=1.66
r201 4 30 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.63
+ $Y=1.485 $X2=9.775 $Y2=2
r202 3 26 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=8.71
+ $Y=1.485 $X2=8.835 $Y2=2
r203 2 22 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.42
+ $Y=1.485 $X2=3.565 $Y2=2.34
r204 1 18 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.48
+ $Y=1.485 $X2=2.625 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A_886_297# 1 2 3 4 5 16 18 20 24 26 30 32
+ 36 38 40 42 47 49 51
r70 40 53 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=8.355 $Y=2.255
+ $X2=8.355 $Y2=2.36
r71 40 42 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=8.355 $Y=2.255
+ $X2=8.355 $Y2=2
r72 39 51 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.46 $Y=2.36 $X2=7.375
+ $Y2=2.36
r73 38 53 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=8.23 $Y=2.36
+ $X2=8.355 $Y2=2.36
r74 38 39 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=8.23 $Y=2.36
+ $X2=7.46 $Y2=2.36
r75 34 51 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=7.375 $Y=2.255
+ $X2=7.375 $Y2=2.36
r76 34 36 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.375 $Y=2.255
+ $X2=7.375 $Y2=2
r77 33 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.36 $X2=6.435
+ $Y2=2.36
r78 32 51 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=7.29 $Y=2.36 $X2=7.375
+ $Y2=2.36
r79 32 33 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=7.29 $Y=2.36
+ $X2=6.52 $Y2=2.36
r80 28 49 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.435 $Y=2.255
+ $X2=6.435 $Y2=2.36
r81 28 30 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=6.435 $Y=2.255
+ $X2=6.435 $Y2=2
r82 27 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.58 $Y=2.36 $X2=5.495
+ $Y2=2.36
r83 26 49 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.35 $Y=2.36 $X2=6.435
+ $Y2=2.36
r84 26 27 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=6.35 $Y=2.36
+ $X2=5.58 $Y2=2.36
r85 22 47 2.11342 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.495 $Y=2.255
+ $X2=5.495 $Y2=2.36
r86 22 24 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=5.495 $Y=2.255
+ $X2=5.495 $Y2=2
r87 21 45 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=4.64 $Y=2.36
+ $X2=4.515 $Y2=2.36
r88 20 47 4.3182 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=5.41 $Y=2.36 $X2=5.495
+ $Y2=2.36
r89 20 21 40.6667 $w=2.08e-07 $l=7.7e-07 $layer=LI1_cond $X=5.41 $Y=2.36
+ $X2=4.64 $Y2=2.36
r90 16 45 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.515 $Y=2.255
+ $X2=4.515 $Y2=2.36
r91 16 18 11.7549 $w=2.48e-07 $l=2.55e-07 $layer=LI1_cond $X=4.515 $Y=2.255
+ $X2=4.515 $Y2=2
r92 5 53 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=8.17
+ $Y=1.485 $X2=8.315 $Y2=2.34
r93 5 42 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=8.17
+ $Y=1.485 $X2=8.315 $Y2=2
r94 4 51 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=2.34
r95 4 36 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=7.23
+ $Y=1.485 $X2=7.375 $Y2=2
r96 3 49 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.485 $X2=6.435 $Y2=2.34
r97 3 30 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=6.29
+ $Y=1.485 $X2=6.435 $Y2=2
r98 2 47 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.485 $X2=5.495 $Y2=2.34
r99 2 24 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=5.35
+ $Y=1.485 $X2=5.495 $Y2=2
r100 1 45 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.485 $X2=4.555 $Y2=2.34
r101 1 18 600 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=1 $X=4.43
+ $Y=1.485 $X2=4.555 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A_1352_297# 1 2 3 4 15 19 23 25 27 29 32
+ 34 36
r66 27 38 2.53352 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.22 $Y=1.665
+ $X2=10.22 $Y2=1.58
r67 27 29 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=10.22 $Y=1.665
+ $X2=10.22 $Y2=2.34
r68 26 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.47 $Y=1.58 $X2=9.28
+ $Y2=1.58
r69 25 38 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.03 $Y=1.58
+ $X2=10.22 $Y2=1.58
r70 25 26 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=10.03 $Y=1.58
+ $X2=9.47 $Y2=1.58
r71 21 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.28 $Y=1.665
+ $X2=9.28 $Y2=1.58
r72 21 23 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=9.28 $Y=1.665
+ $X2=9.28 $Y2=2.34
r73 20 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.01 $Y=1.58 $X2=7.82
+ $Y2=1.58
r74 19 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.09 $Y=1.58 $X2=9.28
+ $Y2=1.58
r75 19 20 70.4599 $w=1.68e-07 $l=1.08e-06 $layer=LI1_cond $X=9.09 $Y=1.58
+ $X2=8.01 $Y2=1.58
r76 16 32 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.07 $Y=1.58 $X2=6.88
+ $Y2=1.58
r77 15 34 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.63 $Y=1.58 $X2=7.82
+ $Y2=1.58
r78 15 16 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.63 $Y=1.58
+ $X2=7.07 $Y2=1.58
r79 4 38 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=1.66
r80 4 29 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=2.34
r81 3 36 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.485 $X2=9.305 $Y2=1.66
r82 3 23 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=9.16
+ $Y=1.485 $X2=9.305 $Y2=2.34
r83 2 34 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=7.7
+ $Y=1.485 $X2=7.845 $Y2=1.66
r84 1 32 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=6.76
+ $Y=1.485 $X2=6.905 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%A_27_47# 1 2 3 4 5 6 7 8 9 10 11 34 36 38
+ 46 47 48 52 56 60 64 68 70 74 82 85 86 87 90 91 92
c172 47 0 1.98558e-19 $X=4.075 $Y=0.735
r173 89 91 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.675 $Y=0.58
+ $X2=8.84 $Y2=0.58
r174 89 90 18.0264 $w=6.48e-07 $l=5.75e-07 $layer=LI1_cond $X=8.675 $Y=0.58
+ $X2=8.1 $Y2=0.58
r175 84 86 10.4819 $w=6.48e-07 $l=1.65e-07 $layer=LI1_cond $X=6.415 $Y=0.58
+ $X2=6.58 $Y2=0.58
r176 84 85 16.7383 $w=6.48e-07 $l=5.05e-07 $layer=LI1_cond $X=6.415 $Y=0.58
+ $X2=5.91 $Y2=0.58
r177 72 74 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=10.735 $Y=0.735
+ $X2=10.735 $Y2=0.38
r178 71 92 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.94 $Y=0.82
+ $X2=9.75 $Y2=0.82
r179 70 72 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=10.545 $Y=0.82
+ $X2=10.735 $Y2=0.735
r180 70 71 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=10.545 $Y=0.82
+ $X2=9.94 $Y2=0.82
r181 66 92 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.75 $Y=0.735
+ $X2=9.75 $Y2=0.82
r182 66 68 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=9.75 $Y=0.735
+ $X2=9.75 $Y2=0.38
r183 64 92 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.56 $Y=0.82
+ $X2=9.75 $Y2=0.82
r184 64 91 46.9733 $w=1.68e-07 $l=7.2e-07 $layer=LI1_cond $X=9.56 $Y=0.82
+ $X2=8.84 $Y2=0.82
r185 63 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.54 $Y=0.82
+ $X2=7.35 $Y2=0.82
r186 63 90 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.54 $Y=0.82
+ $X2=8.1 $Y2=0.82
r187 58 87 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.35 $Y=0.735
+ $X2=7.35 $Y2=0.82
r188 58 60 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=7.35 $Y=0.735
+ $X2=7.35 $Y2=0.38
r189 56 87 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.16 $Y=0.82
+ $X2=7.35 $Y2=0.82
r190 56 86 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=7.16 $Y=0.82
+ $X2=6.58 $Y2=0.82
r191 55 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.14 $Y=0.82
+ $X2=4.95 $Y2=0.82
r192 55 85 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=5.14 $Y=0.82
+ $X2=5.91 $Y2=0.82
r193 50 82 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.95 $Y=0.735
+ $X2=4.95 $Y2=0.82
r194 50 52 10.7662 $w=3.78e-07 $l=3.55e-07 $layer=LI1_cond $X=4.95 $Y=0.735
+ $X2=4.95 $Y2=0.38
r195 49 81 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.2 $Y=0.82
+ $X2=4.075 $Y2=0.82
r196 48 82 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.76 $Y=0.82
+ $X2=4.95 $Y2=0.82
r197 48 49 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.76 $Y=0.82
+ $X2=4.2 $Y2=0.82
r198 47 81 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.075 $Y=0.735
+ $X2=4.075 $Y2=0.82
r199 46 79 3.14258 $w=2.5e-07 $l=1.05e-07 $layer=LI1_cond $X=4.075 $Y=0.465
+ $X2=4.075 $Y2=0.36
r200 46 47 12.4464 $w=2.48e-07 $l=2.7e-07 $layer=LI1_cond $X=4.075 $Y=0.465
+ $X2=4.075 $Y2=0.735
r201 43 45 50.4372 $w=2.08e-07 $l=9.55e-07 $layer=LI1_cond $X=2.14 $Y=0.36
+ $X2=3.095 $Y2=0.36
r202 41 43 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=1.2 $Y=0.36 $X2=2.14
+ $Y2=0.36
r203 39 77 3.79048 $w=2.1e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=0.217 $Y2=0.36
r204 39 41 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=0.36
+ $X2=1.2 $Y2=0.36
r205 38 79 3.74117 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=3.95 $Y=0.36
+ $X2=4.075 $Y2=0.36
r206 38 45 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=3.95 $Y=0.36
+ $X2=3.095 $Y2=0.36
r207 34 77 3.10938 $w=2.55e-07 $l=1.05e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.36
r208 34 36 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.217 $Y=0.465
+ $X2=0.217 $Y2=0.72
r209 11 74 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=10.575
+ $Y=0.235 $X2=10.76 $Y2=0.38
r210 10 68 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=9.59
+ $Y=0.235 $X2=9.775 $Y2=0.38
r211 9 89 45.5 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_NDIFF $count=4 $X=8.18
+ $Y=0.235 $X2=8.675 $Y2=0.38
r212 8 60 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=7.19
+ $Y=0.235 $X2=7.375 $Y2=0.38
r213 7 84 45.5 $w=1.7e-07 $l=5.93085e-07 $layer=licon1_NDIFF $count=4 $X=5.89
+ $Y=0.235 $X2=6.415 $Y2=0.38
r214 6 52 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=4.79
+ $Y=0.235 $X2=4.975 $Y2=0.38
r215 5 81 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.035 $Y2=0.74
r216 5 79 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.035 $Y2=0.38
r217 4 45 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=2.91
+ $Y=0.235 $X2=3.095 $Y2=0.38
r218 3 43 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r219 2 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r220 1 77 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
r221 1 36 182 $w=1.7e-07 $l=5.43921e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__O32AI_4%VGND 1 2 3 4 5 6 21 25 29 33 37 41 44 45
+ 47 48 50 51 53 54 56 57 59 60 61 92 93
r143 92 93 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r144 90 93 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.89 $Y=0
+ $X2=10.81 $Y2=0
r145 89 90 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.89 $Y=0 $X2=9.89
+ $Y2=0
r146 87 90 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=0 $X2=9.89
+ $Y2=0
r147 86 87 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=0 $X2=8.97
+ $Y2=0
r148 84 87 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r149 83 86 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.05 $Y=0 $X2=8.97
+ $Y2=0
r150 83 84 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.05 $Y=0 $X2=8.05
+ $Y2=0
r151 81 84 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.59 $Y=0 $X2=8.05
+ $Y2=0
r152 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r153 78 81 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0 $X2=7.59
+ $Y2=0
r154 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r155 75 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r156 74 77 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=5.75 $Y=0 $X2=6.67
+ $Y2=0
r157 74 75 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r158 72 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=5.75
+ $Y2=0
r159 71 72 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r160 69 72 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r161 68 69 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r162 64 68 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=0.23 $Y=0 $X2=4.37
+ $Y2=0
r163 61 69 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=0.23 $Y=0 $X2=4.37
+ $Y2=0
r164 61 64 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r165 59 89 17.615 $w=1.68e-07 $l=2.7e-07 $layer=LI1_cond $X=10.16 $Y=0 $X2=9.89
+ $Y2=0
r166 59 60 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=10.16 $Y=0
+ $X2=10.267 $Y2=0
r167 58 92 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=10.375 $Y=0
+ $X2=10.81 $Y2=0
r168 58 60 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=10.375 $Y=0
+ $X2=10.267 $Y2=0
r169 56 86 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=9.22 $Y=0 $X2=8.97
+ $Y2=0
r170 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.22 $Y=0 $X2=9.305
+ $Y2=0
r171 55 89 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=9.39 $Y=0 $X2=9.89
+ $Y2=0
r172 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.39 $Y=0 $X2=9.305
+ $Y2=0
r173 53 80 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.59
+ $Y2=0
r174 53 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.76 $Y=0 $X2=7.845
+ $Y2=0
r175 52 83 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.93 $Y=0 $X2=8.05
+ $Y2=0
r176 52 54 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.93 $Y=0 $X2=7.845
+ $Y2=0
r177 50 77 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.67
+ $Y2=0
r178 50 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.82 $Y=0 $X2=6.905
+ $Y2=0
r179 49 80 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.99 $Y=0 $X2=7.59
+ $Y2=0
r180 49 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.99 $Y=0 $X2=6.905
+ $Y2=0
r181 47 71 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.29
+ $Y2=0
r182 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.36 $Y=0 $X2=5.525
+ $Y2=0
r183 46 74 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.75
+ $Y2=0
r184 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.69 $Y=0 $X2=5.525
+ $Y2=0
r185 44 68 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.37
+ $Y2=0
r186 44 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.42 $Y=0 $X2=4.505
+ $Y2=0
r187 43 71 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=4.59 $Y=0 $X2=5.29
+ $Y2=0
r188 43 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.59 $Y=0 $X2=4.505
+ $Y2=0
r189 39 60 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=10.267 $Y=0.085
+ $X2=10.267 $Y2=0
r190 39 41 15.8126 $w=2.13e-07 $l=2.95e-07 $layer=LI1_cond $X=10.267 $Y=0.085
+ $X2=10.267 $Y2=0.38
r191 35 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.305 $Y=0.085
+ $X2=9.305 $Y2=0
r192 35 37 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=9.305 $Y=0.085
+ $X2=9.305 $Y2=0.38
r193 31 54 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.845 $Y=0.085
+ $X2=7.845 $Y2=0
r194 31 33 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=7.845 $Y=0.085
+ $X2=7.845 $Y2=0.38
r195 27 51 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0
r196 27 29 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.905 $Y=0.085
+ $X2=6.905 $Y2=0.38
r197 23 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.525 $Y=0.085
+ $X2=5.525 $Y2=0
r198 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.525 $Y=0.085
+ $X2=5.525 $Y2=0.38
r199 19 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.505 $Y=0.085
+ $X2=4.505 $Y2=0
r200 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.505 $Y=0.085
+ $X2=4.505 $Y2=0.38
r201 6 41 182 $w=1.7e-07 $l=2.93684e-07 $layer=licon1_NDIFF $count=1 $X=10.06
+ $Y=0.235 $X2=10.29 $Y2=0.38
r202 5 37 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=9.12
+ $Y=0.235 $X2=9.305 $Y2=0.38
r203 4 33 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=7.66
+ $Y=0.235 $X2=7.845 $Y2=0.38
r204 3 29 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=6.72
+ $Y=0.235 $X2=6.905 $Y2=0.38
r205 2 25 182 $w=1.7e-07 $l=3.29621e-07 $layer=licon1_NDIFF $count=1 $X=5.26
+ $Y=0.235 $X2=5.525 $Y2=0.38
r206 1 21 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=4.32
+ $Y=0.235 $X2=4.505 $Y2=0.38
.ends

