* File: sky130_fd_sc_hdll__nor4_4.pxi.spice
* Created: Thu Aug 27 19:17:07 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4_4%A N_A_c_121_n N_A_M1003_g N_A_c_127_n N_A_M1002_g
+ N_A_c_122_n N_A_M1015_g N_A_c_128_n N_A_M1008_g N_A_c_123_n N_A_M1016_g
+ N_A_c_129_n N_A_M1013_g N_A_c_130_n N_A_M1020_g N_A_c_124_n N_A_M1025_g A
+ N_A_c_125_n N_A_c_126_n A PM_SKY130_FD_SC_HDLL__NOR4_4%A
x_PM_SKY130_FD_SC_HDLL__NOR4_4%B N_B_c_193_n N_B_M1011_g N_B_c_199_n N_B_M1000_g
+ N_B_c_194_n N_B_M1012_g N_B_c_200_n N_B_M1017_g N_B_c_195_n N_B_M1022_g
+ N_B_c_201_n N_B_M1024_g N_B_c_202_n N_B_M1030_g N_B_c_196_n N_B_M1028_g B B B
+ N_B_c_198_n B B PM_SKY130_FD_SC_HDLL__NOR4_4%B
x_PM_SKY130_FD_SC_HDLL__NOR4_4%C N_C_c_269_n N_C_M1005_g N_C_c_275_n N_C_M1004_g
+ N_C_c_270_n N_C_M1006_g N_C_c_276_n N_C_M1014_g N_C_c_271_n N_C_M1019_g
+ N_C_c_277_n N_C_M1021_g N_C_c_278_n N_C_M1027_g N_C_c_272_n N_C_M1023_g C
+ N_C_c_273_n N_C_c_274_n C PM_SKY130_FD_SC_HDLL__NOR4_4%C
x_PM_SKY130_FD_SC_HDLL__NOR4_4%D N_D_c_345_n N_D_M1007_g N_D_c_351_n N_D_M1001_g
+ N_D_c_346_n N_D_M1018_g N_D_c_352_n N_D_M1009_g N_D_c_347_n N_D_M1026_g
+ N_D_c_353_n N_D_M1010_g N_D_c_354_n N_D_M1031_g N_D_c_348_n N_D_M1029_g D
+ N_D_c_349_n N_D_c_350_n D PM_SKY130_FD_SC_HDLL__NOR4_4%D
x_PM_SKY130_FD_SC_HDLL__NOR4_4%A_27_297# N_A_27_297#_M1002_s N_A_27_297#_M1008_s
+ N_A_27_297#_M1020_s N_A_27_297#_M1017_s N_A_27_297#_M1030_s
+ N_A_27_297#_c_422_n N_A_27_297#_c_423_n N_A_27_297#_c_424_n
+ N_A_27_297#_c_449_p N_A_27_297#_c_425_n N_A_27_297#_c_426_n
+ N_A_27_297#_c_451_p N_A_27_297#_c_442_n N_A_27_297#_c_471_p
+ N_A_27_297#_c_427_n N_A_27_297#_c_428_n N_A_27_297#_c_429_n
+ N_A_27_297#_c_454_p PM_SKY130_FD_SC_HDLL__NOR4_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_4%VPWR N_VPWR_M1002_d N_VPWR_M1013_d N_VPWR_c_485_n
+ N_VPWR_c_486_n N_VPWR_c_487_n VPWR N_VPWR_c_488_n N_VPWR_c_484_n
+ N_VPWR_c_490_n N_VPWR_c_491_n PM_SKY130_FD_SC_HDLL__NOR4_4%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4_4%A_497_297# N_A_497_297#_M1000_d
+ N_A_497_297#_M1024_d N_A_497_297#_M1004_d N_A_497_297#_M1021_d
+ N_A_497_297#_c_576_n N_A_497_297#_c_577_n N_A_497_297#_c_578_n
+ N_A_497_297#_c_579_n N_A_497_297#_c_580_n N_A_497_297#_c_581_n
+ N_A_497_297#_c_582_n PM_SKY130_FD_SC_HDLL__NOR4_4%A_497_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_4%A_887_297# N_A_887_297#_M1004_s
+ N_A_887_297#_M1014_s N_A_887_297#_M1027_s N_A_887_297#_M1009_d
+ N_A_887_297#_M1031_d N_A_887_297#_c_635_n N_A_887_297#_c_638_n
+ N_A_887_297#_c_636_n N_A_887_297#_c_677_n N_A_887_297#_c_640_n
+ N_A_887_297#_c_642_n N_A_887_297#_c_643_n N_A_887_297#_c_685_p
+ N_A_887_297#_c_637_n N_A_887_297#_c_689_p N_A_887_297#_c_664_n
+ N_A_887_297#_c_666_n N_A_887_297#_c_668_n
+ PM_SKY130_FD_SC_HDLL__NOR4_4%A_887_297#
x_PM_SKY130_FD_SC_HDLL__NOR4_4%Y N_Y_M1003_s N_Y_M1016_s N_Y_M1011_d N_Y_M1022_d
+ N_Y_M1005_d N_Y_M1019_d N_Y_M1007_s N_Y_M1026_s N_Y_M1001_s N_Y_M1010_s
+ N_Y_c_715_n N_Y_c_692_n N_Y_c_693_n N_Y_c_726_n N_Y_c_694_n N_Y_c_730_n
+ N_Y_c_695_n N_Y_c_743_n N_Y_c_696_n N_Y_c_756_n N_Y_c_697_n N_Y_c_763_n
+ N_Y_c_698_n N_Y_c_767_n N_Y_c_710_n N_Y_c_699_n N_Y_c_788_n N_Y_c_711_n
+ N_Y_c_700_n N_Y_c_701_n N_Y_c_702_n N_Y_c_703_n N_Y_c_704_n N_Y_c_705_n
+ N_Y_c_706_n N_Y_c_712_n N_Y_c_707_n N_Y_c_713_n Y N_Y_c_709_n
+ PM_SKY130_FD_SC_HDLL__NOR4_4%Y
x_PM_SKY130_FD_SC_HDLL__NOR4_4%VGND N_VGND_M1003_d N_VGND_M1015_d N_VGND_M1025_d
+ N_VGND_M1012_s N_VGND_M1028_s N_VGND_M1006_s N_VGND_M1023_s N_VGND_M1018_d
+ N_VGND_M1029_d N_VGND_c_898_n N_VGND_c_899_n N_VGND_c_900_n N_VGND_c_901_n
+ N_VGND_c_902_n N_VGND_c_903_n N_VGND_c_904_n N_VGND_c_905_n N_VGND_c_906_n
+ N_VGND_c_907_n N_VGND_c_908_n N_VGND_c_909_n N_VGND_c_910_n N_VGND_c_911_n
+ N_VGND_c_912_n N_VGND_c_913_n N_VGND_c_914_n N_VGND_c_915_n N_VGND_c_916_n
+ N_VGND_c_917_n N_VGND_c_918_n N_VGND_c_919_n VGND N_VGND_c_920_n
+ N_VGND_c_921_n N_VGND_c_922_n N_VGND_c_923_n N_VGND_c_924_n
+ PM_SKY130_FD_SC_HDLL__NOR4_4%VGND
cc_1 VNB N_A_c_121_n 0.0218461f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_2 VNB N_A_c_122_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_3 VNB N_A_c_123_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_4 VNB N_A_c_124_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_5 VNB N_A_c_125_n 0.0161158f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_6 VNB N_A_c_126_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_7 VNB N_B_c_193_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_8 VNB N_B_c_194_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_9 VNB N_B_c_195_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_10 VNB N_B_c_196_n 0.0224149f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_11 VNB B 0.0163812f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_12 VNB N_B_c_198_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.18
cc_13 VNB N_C_c_269_n 0.021971f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_14 VNB N_C_c_270_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_15 VNB N_C_c_271_n 0.0172026f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_16 VNB N_C_c_272_n 0.0169382f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_17 VNB N_C_c_273_n 0.00349977f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_18 VNB N_C_c_274_n 0.0801694f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_19 VNB N_D_c_345_n 0.0164943f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=0.995
cc_20 VNB N_D_c_346_n 0.0167631f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=0.995
cc_21 VNB N_D_c_347_n 0.0172006f $X=-0.19 $Y=-0.24 $X2=1.43 $Y2=0.995
cc_22 VNB N_D_c_348_n 0.0201672f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=0.995
cc_23 VNB N_D_c_349_n 0.00389209f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.16
cc_24 VNB N_D_c_350_n 0.0767323f $X=-0.19 $Y=-0.24 $X2=1.925 $Y2=1.202
cc_25 VNB N_VPWR_c_484_n 0.364621f $X=-0.19 $Y=-0.24 $X2=0.49 $Y2=1.202
cc_26 VNB N_Y_c_692_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.455 $Y2=1.202
cc_27 VNB N_Y_c_693_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.202
cc_28 VNB N_Y_c_694_n 0.00447396f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.18
cc_29 VNB N_Y_c_695_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.18
cc_30 VNB N_Y_c_696_n 0.00909655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_Y_c_697_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_Y_c_698_n 0.00697564f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_Y_c_699_n 0.00247276f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_Y_c_700_n 0.00250594f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_Y_c_701_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_Y_c_702_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_703_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_704_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_Y_c_705_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_Y_c_706_n 0.00252317f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_Y_c_707_n 0.00262404f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB Y 0.0219386f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_Y_c_709_n 0.011352f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_898_n 0.0103581f $X=-0.19 $Y=-0.24 $X2=0.515 $Y2=1.202
cc_45 VNB N_VGND_c_899_n 0.0340224f $X=-0.19 $Y=-0.24 $X2=0.58 $Y2=1.16
cc_46 VNB N_VGND_c_900_n 0.0198149f $X=-0.19 $Y=-0.24 $X2=0.96 $Y2=1.202
cc_47 VNB N_VGND_c_901_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.75 $Y2=1.202
cc_48 VNB N_VGND_c_902_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=1.95 $Y2=1.202
cc_49 VNB N_VGND_c_903_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.19
cc_50 VNB N_VGND_c_904_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_905_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_906_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_907_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_908_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_909_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_910_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_911_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_912_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_913_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_914_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_915_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_916_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_917_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_918_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_919_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_920_n 0.0119703f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_921_n 0.41131f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_922_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_923_n 0.0192911f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_VGND_c_924_n 0.0208752f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VPB N_A_c_127_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_72 VPB N_A_c_128_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_73 VPB N_A_c_129_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_74 VPB N_A_c_130_n 0.0161064f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_75 VPB N_A_c_126_n 0.048391f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_76 VPB N_B_c_199_n 0.0164231f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_77 VPB N_B_c_200_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_78 VPB N_B_c_201_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_79 VPB N_B_c_202_n 0.0203443f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_80 VPB N_B_c_198_n 0.0492916f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.18
cc_81 VPB N_C_c_275_n 0.0203443f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_82 VPB N_C_c_276_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_83 VPB N_C_c_277_n 0.0159747f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_84 VPB N_C_c_278_n 0.0164331f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_85 VPB N_C_c_274_n 0.0492916f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_86 VPB N_D_c_351_n 0.0164331f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.41
cc_87 VPB N_D_c_352_n 0.0159747f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.41
cc_88 VPB N_D_c_353_n 0.0159562f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_89 VPB N_D_c_354_n 0.0191939f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_90 VPB N_D_c_350_n 0.0465457f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.202
cc_91 VPB N_A_27_297#_c_422_n 0.0108308f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.41
cc_92 VPB N_A_27_297#_c_423_n 0.0327764f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_93 VPB N_A_27_297#_c_424_n 0.00196267f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.985
cc_94 VPB N_A_27_297#_c_425_n 0.00201678f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_A_27_297#_c_426_n 0.00416269f $X=-0.19 $Y=1.305 $X2=0.515 $Y2=1.202
cc_96 VPB N_A_27_297#_c_427_n 0.0019907f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.202
cc_97 VPB N_A_27_297#_c_428_n 0.00518462f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=1.202
cc_98 VPB N_A_27_297#_c_429_n 0.00151002f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_485_n 0.00516582f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.985
cc_100 VPB N_VPWR_c_486_n 0.0195604f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.995
cc_101 VPB N_VPWR_c_487_n 0.00516582f $X=-0.19 $Y=1.305 $X2=1.455 $Y2=1.985
cc_102 VPB N_VPWR_c_488_n 0.162315f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_484_n 0.061448f $X=-0.19 $Y=1.305 $X2=0.49 $Y2=1.202
cc_104 VPB N_VPWR_c_490_n 0.0238702f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_105 VPB N_VPWR_c_491_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0.985 $Y2=1.202
cc_106 VPB N_A_497_297#_c_576_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=0.56
cc_107 VPB N_A_497_297#_c_577_n 0.0179977f $X=-0.19 $Y=1.305 $X2=1.925 $Y2=1.41
cc_108 VPB N_A_497_297#_c_578_n 0.00193318f $X=-0.19 $Y=1.305 $X2=1.95 $Y2=0.56
cc_109 VPB N_A_497_297#_c_579_n 0.00174485f $X=-0.19 $Y=1.305 $X2=0.515
+ $Y2=1.202
cc_110 VPB N_A_497_297#_c_580_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0.58 $Y2=1.16
cc_111 VPB N_A_497_297#_c_581_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0.96 $Y2=1.202
cc_112 VPB N_A_497_297#_c_582_n 0.00187638f $X=-0.19 $Y=1.305 $X2=1.43 $Y2=1.202
cc_113 VPB N_A_887_297#_c_635_n 0.00452881f $X=-0.19 $Y=1.305 $X2=1.455
+ $Y2=1.985
cc_114 VPB N_A_887_297#_c_636_n 0.00166712f $X=-0.19 $Y=1.305 $X2=1.925
+ $Y2=1.985
cc_115 VPB N_A_887_297#_c_637_n 0.00692367f $X=-0.19 $Y=1.305 $X2=1.75 $Y2=1.16
cc_116 VPB N_Y_c_710_n 0.00193318f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_Y_c_711_n 0.0181949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_Y_c_712_n 0.00187638f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_Y_c_713_n 0.00149756f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB Y 0.00841712f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 N_A_c_124_n N_B_c_193_n 0.0243397f $X=1.95 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_122 N_A_c_130_n N_B_c_199_n 0.00971598f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_c_125_n B 0.0121231f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_124 N_A_c_126_n B 2.62535e-19 $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_125 N_A_c_125_n N_B_c_198_n 2.62535e-19 $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A_c_126_n N_B_c_198_n 0.0243397f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_127 N_A_c_125_n N_A_27_297#_c_422_n 0.0192812f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_128 N_A_c_127_n N_A_27_297#_c_424_n 0.0158609f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_c_128_n N_A_27_297#_c_424_n 0.0156273f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_125_n N_A_27_297#_c_424_n 0.0487385f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_c_126_n N_A_27_297#_c_424_n 0.00837544f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_132 N_A_c_129_n N_A_27_297#_c_425_n 0.0156273f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_133 N_A_c_130_n N_A_27_297#_c_425_n 0.0155666f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_125_n N_A_27_297#_c_425_n 0.0480109f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_c_126_n N_A_27_297#_c_425_n 0.00816971f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_136 N_A_c_125_n N_A_27_297#_c_429_n 0.0204509f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_137 N_A_c_126_n N_A_27_297#_c_429_n 0.00656533f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_138 N_A_c_127_n N_VPWR_c_485_n 0.00300743f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_128_n N_VPWR_c_485_n 0.00300743f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_128_n N_VPWR_c_486_n 0.00702461f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_129_n N_VPWR_c_486_n 0.00702461f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_129_n N_VPWR_c_487_n 0.00300743f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_130_n N_VPWR_c_487_n 0.00300743f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_130_n N_VPWR_c_488_n 0.00702461f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_127_n N_VPWR_c_484_n 0.0133387f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_128_n N_VPWR_c_484_n 0.0124092f $X=0.985 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_c_129_n N_VPWR_c_484_n 0.0124092f $X=1.455 $Y=1.41 $X2=0 $Y2=0
cc_148 N_A_c_130_n N_VPWR_c_484_n 0.0124344f $X=1.925 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A_c_127_n N_VPWR_c_490_n 0.00702461f $X=0.515 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A_c_121_n N_Y_c_715_n 0.00539651f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_c_122_n N_Y_c_715_n 0.00686626f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A_c_123_n N_Y_c_715_n 5.45498e-19 $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A_c_122_n N_Y_c_692_n 0.00901745f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A_c_123_n N_Y_c_692_n 0.00901745f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_155 N_A_c_125_n N_Y_c_692_n 0.0398926f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_156 N_A_c_126_n N_Y_c_692_n 0.00345541f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_157 N_A_c_121_n N_Y_c_693_n 0.00266157f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_158 N_A_c_122_n N_Y_c_693_n 0.00116636f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_159 N_A_c_125_n N_Y_c_693_n 0.0307014f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_160 N_A_c_126_n N_Y_c_693_n 0.00358305f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_161 N_A_c_122_n N_Y_c_726_n 5.24597e-19 $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_162 N_A_c_123_n N_Y_c_726_n 0.00651696f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_c_124_n N_Y_c_694_n 0.0106151f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_164 N_A_c_125_n N_Y_c_694_n 0.0118017f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_c_124_n N_Y_c_730_n 5.32212e-19 $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_166 N_A_c_123_n N_Y_c_701_n 0.00119564f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_167 N_A_c_125_n N_Y_c_701_n 0.030835f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_168 N_A_c_126_n N_Y_c_701_n 0.00486271f $X=1.925 $Y=1.202 $X2=0 $Y2=0
cc_169 N_A_c_121_n N_VGND_c_899_n 0.00496762f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_170 N_A_c_125_n N_VGND_c_899_n 0.0157677f $X=1.75 $Y=1.16 $X2=0 $Y2=0
cc_171 N_A_c_121_n N_VGND_c_900_n 0.00541359f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_172 N_A_c_122_n N_VGND_c_900_n 0.00423334f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_173 N_A_c_122_n N_VGND_c_901_n 0.00379224f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_c_123_n N_VGND_c_901_n 0.00276126f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_175 N_A_c_124_n N_VGND_c_902_n 0.00268723f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_176 N_A_c_123_n N_VGND_c_908_n 0.00423334f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_177 N_A_c_124_n N_VGND_c_908_n 0.00437852f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_178 N_A_c_121_n N_VGND_c_921_n 0.0106014f $X=0.49 $Y=0.995 $X2=0 $Y2=0
cc_179 N_A_c_122_n N_VGND_c_921_n 0.006093f $X=0.96 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A_c_123_n N_VGND_c_921_n 0.00608558f $X=1.43 $Y=0.995 $X2=0 $Y2=0
cc_181 N_A_c_124_n N_VGND_c_921_n 0.00615622f $X=1.95 $Y=0.995 $X2=0 $Y2=0
cc_182 B N_C_c_273_n 0.0150083f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_183 B N_C_c_274_n 0.00157386f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_184 N_B_c_199_n N_A_27_297#_c_426_n 2.98195e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B_c_199_n N_A_27_297#_c_442_n 0.0143578f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_200_n N_A_27_297#_c_442_n 0.01161f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_201_n N_A_27_297#_c_427_n 0.01161f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_202_n N_A_27_297#_c_427_n 0.01161f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B_c_199_n N_VPWR_c_488_n 0.00429453f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_200_n N_VPWR_c_488_n 0.00429453f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_201_n N_VPWR_c_488_n 0.00429453f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B_c_202_n N_VPWR_c_488_n 0.00429453f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_c_199_n N_VPWR_c_484_n 0.00609021f $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B_c_200_n N_VPWR_c_484_n 0.00606499f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B_c_201_n N_VPWR_c_484_n 0.00606499f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_202_n N_VPWR_c_484_n 0.00734734f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_200_n N_A_497_297#_c_576_n 0.0128188f $X=2.865 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B_c_201_n N_A_497_297#_c_576_n 0.0128795f $X=3.335 $Y=1.41 $X2=0 $Y2=0
cc_199 B N_A_497_297#_c_576_n 0.0486996f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_200 N_B_c_198_n N_A_497_297#_c_576_n 0.00864922f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_201 N_B_c_202_n N_A_497_297#_c_577_n 0.0148794f $X=3.805 $Y=1.41 $X2=0 $Y2=0
cc_202 B N_A_497_297#_c_577_n 0.0577826f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_203 N_B_c_198_n N_A_497_297#_c_577_n 8.84531e-19 $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_204 N_B_c_199_n N_A_497_297#_c_579_n 2.98195e-19 $X=2.395 $Y=1.41 $X2=0 $Y2=0
cc_205 B N_A_497_297#_c_579_n 0.0204252f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_206 N_B_c_198_n N_A_497_297#_c_579_n 0.00655199f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_207 B N_A_497_297#_c_580_n 0.0204252f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_208 N_B_c_198_n N_A_497_297#_c_580_n 0.00634604f $X=3.805 $Y=1.202 $X2=0
+ $Y2=0
cc_209 N_B_c_193_n N_Y_c_694_n 0.00865686f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_210 B N_Y_c_694_n 0.00826974f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_211 N_B_c_193_n N_Y_c_730_n 0.00644736f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_212 N_B_c_194_n N_Y_c_730_n 0.00686626f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_213 N_B_c_195_n N_Y_c_730_n 5.45498e-19 $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_214 N_B_c_194_n N_Y_c_695_n 0.00901745f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_215 N_B_c_195_n N_Y_c_695_n 0.00901745f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_216 B N_Y_c_695_n 0.0398926f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_217 N_B_c_198_n N_Y_c_695_n 0.00345541f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_218 N_B_c_194_n N_Y_c_743_n 5.24597e-19 $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_219 N_B_c_195_n N_Y_c_743_n 0.00651696f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_220 N_B_c_196_n N_Y_c_696_n 0.01289f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_221 B N_Y_c_696_n 0.0552267f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_222 N_B_c_193_n N_Y_c_702_n 0.00116636f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_223 N_B_c_194_n N_Y_c_702_n 0.00116636f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_224 B N_Y_c_702_n 0.0307014f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_225 N_B_c_198_n N_Y_c_702_n 0.00358305f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_226 N_B_c_195_n N_Y_c_703_n 0.00119564f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_227 B N_Y_c_703_n 0.030835f $X=4.23 $Y=1.105 $X2=0 $Y2=0
cc_228 N_B_c_198_n N_Y_c_703_n 0.00486271f $X=3.805 $Y=1.202 $X2=0 $Y2=0
cc_229 N_B_c_193_n N_VGND_c_902_n 0.00268723f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_230 N_B_c_194_n N_VGND_c_903_n 0.00379224f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_231 N_B_c_195_n N_VGND_c_903_n 0.00276126f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_232 N_B_c_193_n N_VGND_c_910_n 0.00423334f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_233 N_B_c_194_n N_VGND_c_910_n 0.00423334f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_234 N_B_c_193_n N_VGND_c_921_n 0.00587047f $X=2.37 $Y=0.995 $X2=0 $Y2=0
cc_235 N_B_c_194_n N_VGND_c_921_n 0.006093f $X=2.84 $Y=0.995 $X2=0 $Y2=0
cc_236 N_B_c_195_n N_VGND_c_921_n 0.00608558f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_237 N_B_c_196_n N_VGND_c_921_n 0.00745263f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_238 N_B_c_195_n N_VGND_c_923_n 0.00423334f $X=3.31 $Y=0.995 $X2=0 $Y2=0
cc_239 N_B_c_196_n N_VGND_c_923_n 0.00437852f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_240 N_B_c_196_n N_VGND_c_924_n 0.00481673f $X=3.83 $Y=0.995 $X2=0 $Y2=0
cc_241 N_C_c_272_n N_D_c_345_n 0.0243397f $X=6.23 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_242 N_C_c_278_n N_D_c_351_n 0.0213499f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_243 N_C_c_273_n N_D_c_349_n 0.0185441f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_244 N_C_c_274_n N_D_c_349_n 8.21108e-19 $X=6.205 $Y=1.202 $X2=0 $Y2=0
cc_245 N_C_c_273_n N_D_c_350_n 2.16854e-19 $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_246 N_C_c_274_n N_D_c_350_n 0.0243397f $X=6.205 $Y=1.202 $X2=0 $Y2=0
cc_247 N_C_c_275_n N_VPWR_c_488_n 0.00429453f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_248 N_C_c_276_n N_VPWR_c_488_n 0.00429453f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_249 N_C_c_277_n N_VPWR_c_488_n 0.00429453f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_250 N_C_c_278_n N_VPWR_c_488_n 0.00429453f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_251 N_C_c_275_n N_VPWR_c_484_n 0.00734734f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_252 N_C_c_276_n N_VPWR_c_484_n 0.00606499f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_253 N_C_c_277_n N_VPWR_c_484_n 0.00606499f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_254 N_C_c_278_n N_VPWR_c_484_n 0.00609021f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_255 N_C_c_275_n N_A_497_297#_c_577_n 0.0148794f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_256 N_C_c_273_n N_A_497_297#_c_577_n 0.0145434f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_257 N_C_c_274_n N_A_497_297#_c_577_n 8.84531e-19 $X=6.205 $Y=1.202 $X2=0
+ $Y2=0
cc_258 N_C_c_276_n N_A_497_297#_c_578_n 0.0128795f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_259 N_C_c_277_n N_A_497_297#_c_578_n 0.0128188f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_260 N_C_c_273_n N_A_497_297#_c_578_n 0.0486996f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_261 N_C_c_274_n N_A_497_297#_c_578_n 0.00864922f $X=6.205 $Y=1.202 $X2=0
+ $Y2=0
cc_262 N_C_c_273_n N_A_497_297#_c_581_n 0.0204252f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_263 N_C_c_274_n N_A_497_297#_c_581_n 0.00655199f $X=6.205 $Y=1.202 $X2=0
+ $Y2=0
cc_264 N_C_c_278_n N_A_497_297#_c_582_n 9.73013e-19 $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_265 N_C_c_273_n N_A_497_297#_c_582_n 0.0204252f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_266 N_C_c_274_n N_A_497_297#_c_582_n 0.00634604f $X=6.205 $Y=1.202 $X2=0
+ $Y2=0
cc_267 N_C_c_275_n N_A_887_297#_c_638_n 0.01161f $X=4.795 $Y=1.41 $X2=0 $Y2=0
cc_268 N_C_c_276_n N_A_887_297#_c_638_n 0.01161f $X=5.265 $Y=1.41 $X2=0 $Y2=0
cc_269 N_C_c_277_n N_A_887_297#_c_640_n 0.01161f $X=5.735 $Y=1.41 $X2=0 $Y2=0
cc_270 N_C_c_278_n N_A_887_297#_c_640_n 0.0143578f $X=6.205 $Y=1.41 $X2=0 $Y2=0
cc_271 N_C_c_269_n N_Y_c_696_n 0.0109318f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_272 N_C_c_273_n N_Y_c_696_n 0.00826974f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_273 N_C_c_269_n N_Y_c_756_n 0.0110728f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_274 N_C_c_270_n N_Y_c_756_n 0.00686626f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_275 N_C_c_271_n N_Y_c_756_n 5.45498e-19 $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_276 N_C_c_270_n N_Y_c_697_n 0.00901745f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_277 N_C_c_271_n N_Y_c_697_n 0.00901745f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_278 N_C_c_273_n N_Y_c_697_n 0.0398926f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_279 N_C_c_274_n N_Y_c_697_n 0.00345541f $X=6.205 $Y=1.202 $X2=0 $Y2=0
cc_280 N_C_c_270_n N_Y_c_763_n 5.24597e-19 $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_281 N_C_c_271_n N_Y_c_763_n 0.00651696f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_282 N_C_c_272_n N_Y_c_698_n 0.0106151f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_283 N_C_c_273_n N_Y_c_698_n 0.0118017f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_284 N_C_c_272_n N_Y_c_767_n 5.32212e-19 $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_285 N_C_c_269_n N_Y_c_704_n 0.00116636f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_286 N_C_c_270_n N_Y_c_704_n 0.00116636f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_287 N_C_c_273_n N_Y_c_704_n 0.0307014f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_288 N_C_c_274_n N_Y_c_704_n 0.00358305f $X=6.205 $Y=1.202 $X2=0 $Y2=0
cc_289 N_C_c_271_n N_Y_c_705_n 0.00119564f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_290 N_C_c_273_n N_Y_c_705_n 0.030835f $X=6.03 $Y=1.16 $X2=0 $Y2=0
cc_291 N_C_c_274_n N_Y_c_705_n 0.00486271f $X=6.205 $Y=1.202 $X2=0 $Y2=0
cc_292 N_C_c_270_n N_VGND_c_904_n 0.00379224f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_293 N_C_c_271_n N_VGND_c_904_n 0.00276126f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_294 N_C_c_272_n N_VGND_c_905_n 0.00268723f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_295 N_C_c_269_n N_VGND_c_912_n 0.00423334f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_296 N_C_c_270_n N_VGND_c_912_n 0.00423334f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_297 N_C_c_271_n N_VGND_c_914_n 0.00423334f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_298 N_C_c_272_n N_VGND_c_914_n 0.00437852f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_299 N_C_c_269_n N_VGND_c_921_n 0.00716687f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_300 N_C_c_270_n N_VGND_c_921_n 0.006093f $X=5.24 $Y=0.995 $X2=0 $Y2=0
cc_301 N_C_c_271_n N_VGND_c_921_n 0.00608558f $X=5.71 $Y=0.995 $X2=0 $Y2=0
cc_302 N_C_c_272_n N_VGND_c_921_n 0.00615622f $X=6.23 $Y=0.995 $X2=0 $Y2=0
cc_303 N_C_c_269_n N_VGND_c_924_n 0.00481673f $X=4.77 $Y=0.995 $X2=0 $Y2=0
cc_304 N_D_c_351_n N_VPWR_c_488_n 0.00429453f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_305 N_D_c_352_n N_VPWR_c_488_n 0.00429453f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_306 N_D_c_353_n N_VPWR_c_488_n 0.00429453f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_307 N_D_c_354_n N_VPWR_c_488_n 0.00429453f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_308 N_D_c_351_n N_VPWR_c_484_n 0.00609021f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_309 N_D_c_352_n N_VPWR_c_484_n 0.00606499f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_310 N_D_c_353_n N_VPWR_c_484_n 0.00606499f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_311 N_D_c_354_n N_VPWR_c_484_n 0.0070948f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_312 N_D_c_349_n N_A_887_297#_c_642_n 0.00266826f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_313 N_D_c_351_n N_A_887_297#_c_643_n 0.0143578f $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_314 N_D_c_352_n N_A_887_297#_c_643_n 0.01161f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_315 N_D_c_353_n N_A_887_297#_c_637_n 0.01161f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_316 N_D_c_354_n N_A_887_297#_c_637_n 0.01161f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_317 N_D_c_345_n N_Y_c_698_n 0.00865686f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_318 N_D_c_349_n N_Y_c_698_n 0.0159556f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_319 N_D_c_345_n N_Y_c_767_n 0.00644736f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_320 N_D_c_346_n N_Y_c_767_n 0.00686626f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_321 N_D_c_347_n N_Y_c_767_n 5.45498e-19 $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_322 N_D_c_352_n N_Y_c_710_n 0.0128188f $X=7.145 $Y=1.41 $X2=0 $Y2=0
cc_323 N_D_c_353_n N_Y_c_710_n 0.0128795f $X=7.615 $Y=1.41 $X2=0 $Y2=0
cc_324 N_D_c_349_n N_Y_c_710_n 0.0486996f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_325 N_D_c_350_n N_Y_c_710_n 0.00864922f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_326 N_D_c_346_n N_Y_c_699_n 0.00901745f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_327 N_D_c_347_n N_Y_c_699_n 0.00901745f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_328 N_D_c_349_n N_Y_c_699_n 0.0398926f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_329 N_D_c_350_n N_Y_c_699_n 0.00345541f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_330 N_D_c_346_n N_Y_c_788_n 5.24597e-19 $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_331 N_D_c_347_n N_Y_c_788_n 0.00651696f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_332 N_D_c_354_n N_Y_c_711_n 0.0160435f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_333 N_D_c_349_n N_Y_c_711_n 0.0048601f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_334 N_D_c_350_n N_Y_c_711_n 9.33689e-19 $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_335 N_D_c_348_n N_Y_c_700_n 0.0141313f $X=8.11 $Y=0.995 $X2=0 $Y2=0
cc_336 N_D_c_349_n N_Y_c_700_n 0.00211379f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_337 N_D_c_345_n N_Y_c_706_n 0.00116636f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_338 N_D_c_346_n N_Y_c_706_n 0.00116636f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_339 N_D_c_349_n N_Y_c_706_n 0.0307014f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_340 N_D_c_350_n N_Y_c_706_n 0.00358305f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_341 N_D_c_351_n N_Y_c_712_n 9.73013e-19 $X=6.675 $Y=1.41 $X2=0 $Y2=0
cc_342 N_D_c_349_n N_Y_c_712_n 0.0204252f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_343 N_D_c_350_n N_Y_c_712_n 0.00655199f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_344 N_D_c_347_n N_Y_c_707_n 0.00119564f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_345 N_D_c_349_n N_Y_c_707_n 0.030835f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_346 N_D_c_350_n N_Y_c_707_n 0.00486271f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_347 N_D_c_349_n N_Y_c_713_n 0.0204252f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_348 N_D_c_350_n N_Y_c_713_n 0.00634604f $X=8.085 $Y=1.202 $X2=0 $Y2=0
cc_349 N_D_c_354_n Y 0.00159768f $X=8.085 $Y=1.41 $X2=0 $Y2=0
cc_350 N_D_c_348_n Y 0.0175063f $X=8.11 $Y=0.995 $X2=0 $Y2=0
cc_351 N_D_c_349_n Y 0.0108179f $X=7.88 $Y=1.16 $X2=0 $Y2=0
cc_352 N_D_c_345_n N_VGND_c_905_n 0.00268723f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_353 N_D_c_346_n N_VGND_c_906_n 0.00379224f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_354 N_D_c_347_n N_VGND_c_906_n 0.00276126f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_355 N_D_c_348_n N_VGND_c_907_n 0.00438629f $X=8.11 $Y=0.995 $X2=0 $Y2=0
cc_356 N_D_c_345_n N_VGND_c_916_n 0.00423334f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_357 N_D_c_346_n N_VGND_c_916_n 0.00423334f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_358 N_D_c_347_n N_VGND_c_918_n 0.00423334f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_359 N_D_c_348_n N_VGND_c_918_n 0.00437852f $X=8.11 $Y=0.995 $X2=0 $Y2=0
cc_360 N_D_c_345_n N_VGND_c_921_n 0.00587047f $X=6.65 $Y=0.995 $X2=0 $Y2=0
cc_361 N_D_c_346_n N_VGND_c_921_n 0.006093f $X=7.12 $Y=0.995 $X2=0 $Y2=0
cc_362 N_D_c_347_n N_VGND_c_921_n 0.00608558f $X=7.59 $Y=0.995 $X2=0 $Y2=0
cc_363 N_D_c_348_n N_VGND_c_921_n 0.00720525f $X=8.11 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A_27_297#_c_424_n N_VPWR_M1002_d 0.00187091f $X=1.095 $Y=1.54 $X2=-0.19
+ $Y2=1.305
cc_365 N_A_27_297#_c_425_n N_VPWR_M1013_d 0.00187091f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_366 N_A_27_297#_c_424_n N_VPWR_c_485_n 0.0143191f $X=1.095 $Y=1.54 $X2=0
+ $Y2=0
cc_367 N_A_27_297#_c_449_p N_VPWR_c_486_n 0.0149311f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_368 N_A_27_297#_c_425_n N_VPWR_c_487_n 0.0143191f $X=2.035 $Y=1.54 $X2=0
+ $Y2=0
cc_369 N_A_27_297#_c_451_p N_VPWR_c_488_n 0.015002f $X=2.16 $Y=2.295 $X2=0 $Y2=0
cc_370 N_A_27_297#_c_442_n N_VPWR_c_488_n 0.0386815f $X=2.975 $Y=2.38 $X2=0
+ $Y2=0
cc_371 N_A_27_297#_c_427_n N_VPWR_c_488_n 0.0588952f $X=3.915 $Y=2.38 $X2=0
+ $Y2=0
cc_372 N_A_27_297#_c_454_p N_VPWR_c_488_n 0.0149886f $X=3.1 $Y=2.38 $X2=0 $Y2=0
cc_373 N_A_27_297#_M1002_s N_VPWR_c_484_n 0.00303344f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_374 N_A_27_297#_M1008_s N_VPWR_c_484_n 0.00370124f $X=1.075 $Y=1.485 $X2=0
+ $Y2=0
cc_375 N_A_27_297#_M1020_s N_VPWR_c_484_n 0.00297222f $X=2.015 $Y=1.485 $X2=0
+ $Y2=0
cc_376 N_A_27_297#_M1017_s N_VPWR_c_484_n 0.00231264f $X=2.955 $Y=1.485 $X2=0
+ $Y2=0
cc_377 N_A_27_297#_M1030_s N_VPWR_c_484_n 0.00217519f $X=3.895 $Y=1.485 $X2=0
+ $Y2=0
cc_378 N_A_27_297#_c_423_n N_VPWR_c_484_n 0.0120542f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_379 N_A_27_297#_c_449_p N_VPWR_c_484_n 0.00955092f $X=1.22 $Y=2.3 $X2=0 $Y2=0
cc_380 N_A_27_297#_c_451_p N_VPWR_c_484_n 0.00962794f $X=2.16 $Y=2.295 $X2=0
+ $Y2=0
cc_381 N_A_27_297#_c_442_n N_VPWR_c_484_n 0.0239144f $X=2.975 $Y=2.38 $X2=0
+ $Y2=0
cc_382 N_A_27_297#_c_427_n N_VPWR_c_484_n 0.035656f $X=3.915 $Y=2.38 $X2=0 $Y2=0
cc_383 N_A_27_297#_c_454_p N_VPWR_c_484_n 0.00962421f $X=3.1 $Y=2.38 $X2=0 $Y2=0
cc_384 N_A_27_297#_c_423_n N_VPWR_c_490_n 0.0208166f $X=0.28 $Y=2.3 $X2=0 $Y2=0
cc_385 N_A_27_297#_c_442_n N_A_497_297#_M1000_d 0.00352392f $X=2.975 $Y=2.38
+ $X2=-0.19 $Y2=1.305
cc_386 N_A_27_297#_c_427_n N_A_497_297#_M1024_d 0.00352392f $X=3.915 $Y=2.38
+ $X2=0 $Y2=0
cc_387 N_A_27_297#_M1017_s N_A_497_297#_c_576_n 0.00187091f $X=2.955 $Y=1.485
+ $X2=0 $Y2=0
cc_388 N_A_27_297#_c_442_n N_A_497_297#_c_576_n 0.00385532f $X=2.975 $Y=2.38
+ $X2=0 $Y2=0
cc_389 N_A_27_297#_c_471_p N_A_497_297#_c_576_n 0.0143018f $X=3.1 $Y=1.96 $X2=0
+ $Y2=0
cc_390 N_A_27_297#_c_427_n N_A_497_297#_c_576_n 0.00385532f $X=3.915 $Y=2.38
+ $X2=0 $Y2=0
cc_391 N_A_27_297#_M1030_s N_A_497_297#_c_577_n 0.00295666f $X=3.895 $Y=1.485
+ $X2=0 $Y2=0
cc_392 N_A_27_297#_c_427_n N_A_497_297#_c_577_n 0.00385532f $X=3.915 $Y=2.38
+ $X2=0 $Y2=0
cc_393 N_A_27_297#_c_428_n N_A_497_297#_c_577_n 0.0218636f $X=4.04 $Y=1.96 $X2=0
+ $Y2=0
cc_394 N_A_27_297#_c_426_n N_A_497_297#_c_579_n 0.00226124f $X=2.16 $Y=1.625
+ $X2=0 $Y2=0
cc_395 N_A_27_297#_c_442_n N_A_497_297#_c_579_n 0.013395f $X=2.975 $Y=2.38 $X2=0
+ $Y2=0
cc_396 N_A_27_297#_c_427_n N_A_497_297#_c_580_n 0.013395f $X=3.915 $Y=2.38 $X2=0
+ $Y2=0
cc_397 N_A_27_297#_c_428_n N_A_887_297#_c_635_n 0.0384367f $X=4.04 $Y=1.96 $X2=0
+ $Y2=0
cc_398 N_A_27_297#_c_427_n N_A_887_297#_c_636_n 0.0149967f $X=3.915 $Y=2.38
+ $X2=0 $Y2=0
cc_399 N_A_27_297#_c_425_n N_Y_c_694_n 3.18413e-19 $X=2.035 $Y=1.54 $X2=0 $Y2=0
cc_400 N_A_27_297#_c_426_n N_Y_c_694_n 0.00936521f $X=2.16 $Y=1.625 $X2=0 $Y2=0
cc_401 N_A_27_297#_c_422_n N_VGND_c_899_n 0.00367361f $X=0.247 $Y=1.625 $X2=0
+ $Y2=0
cc_402 N_VPWR_c_484_n N_A_497_297#_M1000_d 0.00232895f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_403 N_VPWR_c_484_n N_A_497_297#_M1024_d 0.00232895f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_404 N_VPWR_c_484_n N_A_497_297#_M1004_d 0.00232895f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_405 N_VPWR_c_484_n N_A_497_297#_M1021_d 0.00232895f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_406 N_VPWR_c_484_n N_A_887_297#_M1004_s 0.00217519f $X=8.51 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_407 N_VPWR_c_484_n N_A_887_297#_M1014_s 0.00231264f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_408 N_VPWR_c_484_n N_A_887_297#_M1027_s 0.00231264f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_409 N_VPWR_c_484_n N_A_887_297#_M1009_d 0.00231264f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_410 N_VPWR_c_484_n N_A_887_297#_M1031_d 0.00217519f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_411 N_VPWR_c_488_n N_A_887_297#_c_638_n 0.0386815f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_412 N_VPWR_c_484_n N_A_887_297#_c_638_n 0.0239144f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_413 N_VPWR_c_488_n N_A_887_297#_c_636_n 0.0184233f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_414 N_VPWR_c_484_n N_A_887_297#_c_636_n 0.0107791f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_415 N_VPWR_c_488_n N_A_887_297#_c_640_n 0.0386815f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_416 N_VPWR_c_484_n N_A_887_297#_c_640_n 0.0239144f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_417 N_VPWR_c_488_n N_A_887_297#_c_643_n 0.0386815f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_418 N_VPWR_c_484_n N_A_887_297#_c_643_n 0.0239144f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_419 N_VPWR_c_488_n N_A_887_297#_c_637_n 0.0549564f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_420 N_VPWR_c_484_n N_A_887_297#_c_637_n 0.0335386f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_421 N_VPWR_c_488_n N_A_887_297#_c_664_n 0.0149886f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_422 N_VPWR_c_484_n N_A_887_297#_c_664_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_423 N_VPWR_c_488_n N_A_887_297#_c_666_n 0.0149886f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_424 N_VPWR_c_484_n N_A_887_297#_c_666_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_425 N_VPWR_c_488_n N_A_887_297#_c_668_n 0.0149886f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_426 N_VPWR_c_484_n N_A_887_297#_c_668_n 0.00962421f $X=8.51 $Y=2.72 $X2=0
+ $Y2=0
cc_427 N_VPWR_c_484_n N_Y_M1001_s 0.00232895f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_428 N_VPWR_c_484_n N_Y_M1010_s 0.00232895f $X=8.51 $Y=2.72 $X2=0 $Y2=0
cc_429 N_A_497_297#_c_577_n N_A_887_297#_M1004_s 0.00295666f $X=4.905 $Y=1.54
+ $X2=-0.19 $Y2=1.305
cc_430 N_A_497_297#_c_578_n N_A_887_297#_M1014_s 0.00187091f $X=5.845 $Y=1.54
+ $X2=0 $Y2=0
cc_431 N_A_497_297#_c_577_n N_A_887_297#_c_635_n 0.0197547f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_432 N_A_497_297#_M1004_d N_A_887_297#_c_638_n 0.00352392f $X=4.885 $Y=1.485
+ $X2=0 $Y2=0
cc_433 N_A_497_297#_c_577_n N_A_887_297#_c_638_n 0.00385532f $X=4.905 $Y=1.54
+ $X2=0 $Y2=0
cc_434 N_A_497_297#_c_578_n N_A_887_297#_c_638_n 0.00385532f $X=5.845 $Y=1.54
+ $X2=0 $Y2=0
cc_435 N_A_497_297#_c_581_n N_A_887_297#_c_638_n 0.013395f $X=5.03 $Y=1.62 $X2=0
+ $Y2=0
cc_436 N_A_497_297#_c_578_n N_A_887_297#_c_677_n 0.0143018f $X=5.845 $Y=1.54
+ $X2=0 $Y2=0
cc_437 N_A_497_297#_M1021_d N_A_887_297#_c_640_n 0.00352392f $X=5.825 $Y=1.485
+ $X2=0 $Y2=0
cc_438 N_A_497_297#_c_578_n N_A_887_297#_c_640_n 0.00385532f $X=5.845 $Y=1.54
+ $X2=0 $Y2=0
cc_439 N_A_497_297#_c_582_n N_A_887_297#_c_640_n 0.013395f $X=5.97 $Y=1.62 $X2=0
+ $Y2=0
cc_440 N_A_497_297#_c_577_n N_Y_c_696_n 0.00753964f $X=4.905 $Y=1.54 $X2=0 $Y2=0
cc_441 N_A_887_297#_c_643_n N_Y_M1001_s 0.00352392f $X=7.255 $Y=2.38 $X2=0 $Y2=0
cc_442 N_A_887_297#_c_637_n N_Y_M1010_s 0.00352392f $X=8.195 $Y=2.38 $X2=0 $Y2=0
cc_443 N_A_887_297#_M1009_d N_Y_c_710_n 0.00187091f $X=7.235 $Y=1.485 $X2=0
+ $Y2=0
cc_444 N_A_887_297#_c_643_n N_Y_c_710_n 0.00385532f $X=7.255 $Y=2.38 $X2=0 $Y2=0
cc_445 N_A_887_297#_c_685_p N_Y_c_710_n 0.0143018f $X=7.38 $Y=1.96 $X2=0 $Y2=0
cc_446 N_A_887_297#_c_637_n N_Y_c_710_n 0.00385532f $X=8.195 $Y=2.38 $X2=0 $Y2=0
cc_447 N_A_887_297#_M1031_d N_Y_c_711_n 0.00296904f $X=8.175 $Y=1.485 $X2=0
+ $Y2=0
cc_448 N_A_887_297#_c_637_n N_Y_c_711_n 0.00385532f $X=8.195 $Y=2.38 $X2=0 $Y2=0
cc_449 N_A_887_297#_c_689_p N_Y_c_711_n 0.0179301f $X=8.32 $Y=1.96 $X2=0 $Y2=0
cc_450 N_A_887_297#_c_643_n N_Y_c_712_n 0.013395f $X=7.255 $Y=2.38 $X2=0 $Y2=0
cc_451 N_A_887_297#_c_637_n N_Y_c_713_n 0.013395f $X=8.195 $Y=2.38 $X2=0 $Y2=0
cc_452 N_Y_c_692_n N_VGND_M1015_d 0.00251047f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_453 N_Y_c_694_n N_VGND_M1025_d 0.00162089f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_454 N_Y_c_695_n N_VGND_M1012_s 0.00251047f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_455 N_Y_c_696_n N_VGND_M1028_s 0.0108248f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_456 N_Y_c_697_n N_VGND_M1006_s 0.00251047f $X=5.755 $Y=0.815 $X2=0 $Y2=0
cc_457 N_Y_c_698_n N_VGND_M1023_s 0.00162089f $X=6.695 $Y=0.815 $X2=0 $Y2=0
cc_458 N_Y_c_699_n N_VGND_M1018_d 0.00251047f $X=7.635 $Y=0.815 $X2=0 $Y2=0
cc_459 N_Y_c_700_n N_VGND_M1029_d 0.00121567f $X=8.36 $Y=0.815 $X2=0 $Y2=0
cc_460 N_Y_c_709_n N_VGND_M1029_d 0.00198968f $X=8.495 $Y=0.905 $X2=0 $Y2=0
cc_461 N_Y_c_693_n N_VGND_c_899_n 0.00835456f $X=0.915 $Y=0.815 $X2=0 $Y2=0
cc_462 N_Y_c_715_n N_VGND_c_900_n 0.0223596f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_463 N_Y_c_692_n N_VGND_c_900_n 0.00266636f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_464 N_Y_c_715_n N_VGND_c_901_n 0.0183628f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_465 N_Y_c_692_n N_VGND_c_901_n 0.0127273f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_466 N_Y_c_694_n N_VGND_c_902_n 0.0122559f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_467 N_Y_c_730_n N_VGND_c_903_n 0.0183628f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_468 N_Y_c_695_n N_VGND_c_903_n 0.0127273f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_469 N_Y_c_756_n N_VGND_c_904_n 0.0183628f $X=5.03 $Y=0.39 $X2=0 $Y2=0
cc_470 N_Y_c_697_n N_VGND_c_904_n 0.0127273f $X=5.755 $Y=0.815 $X2=0 $Y2=0
cc_471 N_Y_c_698_n N_VGND_c_905_n 0.0122559f $X=6.695 $Y=0.815 $X2=0 $Y2=0
cc_472 N_Y_c_767_n N_VGND_c_906_n 0.0183628f $X=6.91 $Y=0.39 $X2=0 $Y2=0
cc_473 N_Y_c_699_n N_VGND_c_906_n 0.0127273f $X=7.635 $Y=0.815 $X2=0 $Y2=0
cc_474 N_Y_c_700_n N_VGND_c_907_n 0.00923644f $X=8.36 $Y=0.815 $X2=0 $Y2=0
cc_475 N_Y_c_709_n N_VGND_c_907_n 0.00380511f $X=8.495 $Y=0.905 $X2=0 $Y2=0
cc_476 N_Y_c_692_n N_VGND_c_908_n 0.00198695f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_477 N_Y_c_726_n N_VGND_c_908_n 0.0231806f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_478 N_Y_c_694_n N_VGND_c_908_n 0.00254521f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_479 N_Y_c_694_n N_VGND_c_910_n 0.00198695f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_480 N_Y_c_730_n N_VGND_c_910_n 0.0223596f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_481 N_Y_c_695_n N_VGND_c_910_n 0.00266636f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_482 N_Y_c_696_n N_VGND_c_912_n 0.00198695f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_483 N_Y_c_756_n N_VGND_c_912_n 0.0223596f $X=5.03 $Y=0.39 $X2=0 $Y2=0
cc_484 N_Y_c_697_n N_VGND_c_912_n 0.00266636f $X=5.755 $Y=0.815 $X2=0 $Y2=0
cc_485 N_Y_c_697_n N_VGND_c_914_n 0.00198695f $X=5.755 $Y=0.815 $X2=0 $Y2=0
cc_486 N_Y_c_763_n N_VGND_c_914_n 0.0231806f $X=5.97 $Y=0.39 $X2=0 $Y2=0
cc_487 N_Y_c_698_n N_VGND_c_914_n 0.00254521f $X=6.695 $Y=0.815 $X2=0 $Y2=0
cc_488 N_Y_c_698_n N_VGND_c_916_n 0.00198695f $X=6.695 $Y=0.815 $X2=0 $Y2=0
cc_489 N_Y_c_767_n N_VGND_c_916_n 0.0223596f $X=6.91 $Y=0.39 $X2=0 $Y2=0
cc_490 N_Y_c_699_n N_VGND_c_916_n 0.00266636f $X=7.635 $Y=0.815 $X2=0 $Y2=0
cc_491 N_Y_c_699_n N_VGND_c_918_n 0.00198695f $X=7.635 $Y=0.815 $X2=0 $Y2=0
cc_492 N_Y_c_788_n N_VGND_c_918_n 0.0231806f $X=7.85 $Y=0.39 $X2=0 $Y2=0
cc_493 N_Y_c_700_n N_VGND_c_918_n 0.00254521f $X=8.36 $Y=0.815 $X2=0 $Y2=0
cc_494 N_Y_c_709_n N_VGND_c_920_n 0.00378405f $X=8.495 $Y=0.905 $X2=0 $Y2=0
cc_495 N_Y_M1003_s N_VGND_c_921_n 0.0025535f $X=0.565 $Y=0.235 $X2=0 $Y2=0
cc_496 N_Y_M1016_s N_VGND_c_921_n 0.00304143f $X=1.505 $Y=0.235 $X2=0 $Y2=0
cc_497 N_Y_M1011_d N_VGND_c_921_n 0.0025535f $X=2.445 $Y=0.235 $X2=0 $Y2=0
cc_498 N_Y_M1022_d N_VGND_c_921_n 0.00304143f $X=3.385 $Y=0.235 $X2=0 $Y2=0
cc_499 N_Y_M1005_d N_VGND_c_921_n 0.0025535f $X=4.845 $Y=0.235 $X2=0 $Y2=0
cc_500 N_Y_M1019_d N_VGND_c_921_n 0.00304143f $X=5.785 $Y=0.235 $X2=0 $Y2=0
cc_501 N_Y_M1007_s N_VGND_c_921_n 0.0025535f $X=6.725 $Y=0.235 $X2=0 $Y2=0
cc_502 N_Y_M1026_s N_VGND_c_921_n 0.00304143f $X=7.665 $Y=0.235 $X2=0 $Y2=0
cc_503 N_Y_c_715_n N_VGND_c_921_n 0.0141302f $X=0.75 $Y=0.39 $X2=0 $Y2=0
cc_504 N_Y_c_692_n N_VGND_c_921_n 0.00972452f $X=1.475 $Y=0.815 $X2=0 $Y2=0
cc_505 N_Y_c_726_n N_VGND_c_921_n 0.0143352f $X=1.69 $Y=0.39 $X2=0 $Y2=0
cc_506 N_Y_c_694_n N_VGND_c_921_n 0.0094839f $X=2.415 $Y=0.815 $X2=0 $Y2=0
cc_507 N_Y_c_730_n N_VGND_c_921_n 0.0141302f $X=2.63 $Y=0.39 $X2=0 $Y2=0
cc_508 N_Y_c_695_n N_VGND_c_921_n 0.00972452f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_509 N_Y_c_743_n N_VGND_c_921_n 0.0143352f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_510 N_Y_c_696_n N_VGND_c_921_n 0.0114512f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_511 N_Y_c_756_n N_VGND_c_921_n 0.0141302f $X=5.03 $Y=0.39 $X2=0 $Y2=0
cc_512 N_Y_c_697_n N_VGND_c_921_n 0.00972452f $X=5.755 $Y=0.815 $X2=0 $Y2=0
cc_513 N_Y_c_763_n N_VGND_c_921_n 0.0143352f $X=5.97 $Y=0.39 $X2=0 $Y2=0
cc_514 N_Y_c_698_n N_VGND_c_921_n 0.0094839f $X=6.695 $Y=0.815 $X2=0 $Y2=0
cc_515 N_Y_c_767_n N_VGND_c_921_n 0.0141302f $X=6.91 $Y=0.39 $X2=0 $Y2=0
cc_516 N_Y_c_699_n N_VGND_c_921_n 0.00972452f $X=7.635 $Y=0.815 $X2=0 $Y2=0
cc_517 N_Y_c_788_n N_VGND_c_921_n 0.0143352f $X=7.85 $Y=0.39 $X2=0 $Y2=0
cc_518 N_Y_c_700_n N_VGND_c_921_n 0.00545596f $X=8.36 $Y=0.815 $X2=0 $Y2=0
cc_519 N_Y_c_709_n N_VGND_c_921_n 0.0065683f $X=8.495 $Y=0.905 $X2=0 $Y2=0
cc_520 N_Y_c_695_n N_VGND_c_923_n 0.00198695f $X=3.355 $Y=0.815 $X2=0 $Y2=0
cc_521 N_Y_c_743_n N_VGND_c_923_n 0.0231806f $X=3.57 $Y=0.39 $X2=0 $Y2=0
cc_522 N_Y_c_696_n N_VGND_c_923_n 0.00254521f $X=4.815 $Y=0.815 $X2=0 $Y2=0
cc_523 N_Y_c_696_n N_VGND_c_924_n 0.0528344f $X=4.815 $Y=0.815 $X2=0 $Y2=0
