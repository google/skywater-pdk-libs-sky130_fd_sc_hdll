# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__isobufsrc_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__isobufsrc_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.660000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.255000 0.315000 1.065000 ;
        RECT 0.085000 1.065000 0.505000 1.285000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  2.220000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.790000 1.075000 8.880000 1.275000 ;
    END
  END SLEEP
  PIN VGND
    ANTENNADIFFAREA  2.249000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.660000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.760000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.660000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  2.889000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.125000 0.255000 2.505000 0.725000 ;
        RECT 2.125000 0.725000 9.565000 0.905000 ;
        RECT 3.065000 0.255000 3.445000 0.725000 ;
        RECT 4.005000 0.255000 4.385000 0.725000 ;
        RECT 4.945000 0.255000 5.325000 0.725000 ;
        RECT 5.885000 0.255000 6.265000 0.725000 ;
        RECT 5.975000 1.445000 9.565000 1.615000 ;
        RECT 5.975000 1.615000 6.225000 2.125000 ;
        RECT 6.825000 0.255000 7.205000 0.725000 ;
        RECT 6.915000 1.615000 7.165000 2.125000 ;
        RECT 7.765000 0.255000 8.145000 0.725000 ;
        RECT 7.855000 1.615000 8.105000 2.125000 ;
        RECT 8.705000 0.255000 9.085000 0.725000 ;
        RECT 8.795000 1.615000 9.045000 2.125000 ;
        RECT 9.050000 0.905000 9.565000 1.445000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.660000 0.085000 ;
      RECT 0.000000  2.635000 9.660000 2.805000 ;
      RECT 0.125000  1.455000 0.345000 2.635000 ;
      RECT 0.485000  0.085000 0.705000 0.895000 ;
      RECT 0.515000  1.455000 0.945000 2.465000 ;
      RECT 0.725000  1.065000 1.235000 1.075000 ;
      RECT 0.725000  1.075000 5.520000 1.285000 ;
      RECT 0.725000  1.285000 0.945000 1.455000 ;
      RECT 0.875000  0.255000 1.235000 1.065000 ;
      RECT 1.165000  1.455000 1.460000 2.635000 ;
      RECT 1.445000  0.085000 1.955000 0.905000 ;
      RECT 1.675000  1.455000 5.755000 1.665000 ;
      RECT 1.675000  1.665000 1.995000 2.465000 ;
      RECT 2.215000  1.835000 2.465000 2.635000 ;
      RECT 2.685000  1.665000 2.935000 2.465000 ;
      RECT 2.725000  0.085000 2.895000 0.555000 ;
      RECT 3.155000  1.835000 3.405000 2.635000 ;
      RECT 3.625000  1.665000 3.875000 2.465000 ;
      RECT 3.665000  0.085000 3.835000 0.555000 ;
      RECT 4.095000  1.835000 4.345000 2.635000 ;
      RECT 4.565000  1.665000 4.815000 2.465000 ;
      RECT 4.605000  0.085000 4.775000 0.555000 ;
      RECT 5.035000  1.835000 5.285000 2.635000 ;
      RECT 5.505000  1.665000 5.755000 2.295000 ;
      RECT 5.505000  2.295000 9.515000 2.465000 ;
      RECT 5.545000  0.085000 5.715000 0.555000 ;
      RECT 6.445000  1.785000 6.695000 2.295000 ;
      RECT 6.485000  0.085000 6.655000 0.555000 ;
      RECT 7.385000  1.785000 7.635000 2.295000 ;
      RECT 7.425000  0.085000 7.595000 0.555000 ;
      RECT 8.325000  1.785000 8.575000 2.295000 ;
      RECT 8.365000  0.085000 8.535000 0.555000 ;
      RECT 9.265000  1.785000 9.515000 2.295000 ;
      RECT 9.305000  0.085000 9.575000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
      RECT 9.345000 -0.085000 9.515000 0.085000 ;
      RECT 9.345000  2.635000 9.515000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__isobufsrc_8
END LIBRARY
