* File: sky130_fd_sc_hdll__sdfxtp_2.pex.spice
* Created: Wed Sep  2 08:52:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%CLK 1 2 3 5 6 8 13
c38 1 0 2.71124e-20 $X=0.31 $Y=1.325
r39 13 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.25
+ $Y=1.16 $X2=0.25 $Y2=1.16
r40 6 9 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.5 $Y=1.665 $X2=0.31
+ $Y2=1.665
r41 6 8 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.5 $Y=1.74 $X2=0.5
+ $Y2=2.135
r42 3 16 89.156 $w=2.56e-07 $l=4.95076e-07 $layer=POLY_cond $X=0.47 $Y=0.73
+ $X2=0.33 $Y2=1.16
r43 3 5 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.47 $Y=0.73 $X2=0.47
+ $Y2=0.445
r44 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.31 $Y=1.59 $X2=0.31
+ $Y2=1.665
r45 1 16 39.2615 $w=2.56e-07 $l=1.74714e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.33 $Y2=1.16
r46 1 2 135.883 $w=1.5e-07 $l=2.65e-07 $layer=POLY_cond $X=0.31 $Y=1.325
+ $X2=0.31 $Y2=1.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_27_47# 1 2 9 12 13 15 18 20 21 23 24 26
+ 28 29 31 32 36 40 44 45 46 49 51 54 63 66 67 68 70 72 77 82 86
c238 66 0 1.55016e-19 $X=5.75 $Y=1.825
c239 46 0 1.76957e-19 $X=0.665 $Y=1.88
c240 36 0 7.21183e-20 $X=8.05 $Y=0.415
r241 85 87 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=7.275 $Y=1.41
+ $X2=7.275 $Y2=1.575
r242 85 86 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.25
+ $Y=1.41 $X2=7.25 $Y2=1.41
r243 82 85 16.2293 $w=3.2e-07 $l=9e-08 $layer=POLY_cond $X=7.275 $Y=1.32
+ $X2=7.275 $Y2=1.41
r244 80 81 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.55
+ $Y=1.74 $X2=5.55 $Y2=1.74
r245 76 77 6.66521 $w=2.7e-07 $l=3e-08 $layer=POLY_cond $X=0.94 $Y=1.235
+ $X2=0.97 $Y2=1.235
r246 71 86 19.9277 $w=2.38e-07 $l=4.15e-07 $layer=LI1_cond $X=7.285 $Y=1.825
+ $X2=7.285 $Y2=1.41
r247 70 72 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.31 $Y=1.825
+ $X2=7.115 $Y2=1.825
r248 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.31 $Y=1.825
+ $X2=7.31 $Y2=1.825
r249 68 72 1.5099 $w=1.4e-07 $l=1.22e-06 $layer=MET1_cond $X=5.895 $Y=1.87
+ $X2=7.115 $Y2=1.87
r250 66 81 6.49264 $w=3.53e-07 $l=2e-07 $layer=LI1_cond $X=5.75 $Y=1.832
+ $X2=5.55 $Y2=1.832
r251 65 68 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.895 $Y2=1.825
r252 65 67 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.75 $Y=1.825
+ $X2=5.555 $Y2=1.825
r253 65 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=1.825
+ $X2=5.75 $Y2=1.825
r254 63 67 5.76732 $w=1.4e-07 $l=4.66e-06 $layer=MET1_cond $X=0.895 $Y=1.87
+ $X2=5.555 $Y2=1.87
r255 60 63 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.75 $Y=1.825
+ $X2=0.895 $Y2=1.825
r256 60 61 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.75 $Y=1.825
+ $X2=0.75 $Y2=1.825
r257 52 76 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r258 51 52 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r259 49 61 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.88
r260 49 51 28.0595 $w=2.28e-07 $l=5.6e-07 $layer=LI1_cond $X=0.78 $Y=1.795
+ $X2=0.78 $Y2=1.235
r261 48 51 21.5457 $w=2.28e-07 $l=4.3e-07 $layer=LI1_cond $X=0.78 $Y=0.805
+ $X2=0.78 $Y2=1.235
r262 47 54 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.35 $Y=1.88
+ $X2=0.265 $Y2=1.88
r263 46 61 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.78 $Y2=1.88
r264 46 47 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.665 $Y=1.88
+ $X2=0.35 $Y2=1.88
r265 44 48 7.01789 $w=1.7e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.78 $Y2=0.805
r266 44 45 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=0.665 $Y=0.72
+ $X2=0.345 $Y2=0.72
r267 38 45 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.345 $Y2=0.72
r268 38 40 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.26 $Y=0.635
+ $X2=0.26 $Y2=0.51
r269 34 36 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=8.05 $Y=1.245
+ $X2=8.05 $Y2=0.415
r270 33 82 20.4921 $w=1.5e-07 $l=1.6e-07 $layer=POLY_cond $X=7.435 $Y=1.32
+ $X2=7.275 $Y2=1.32
r271 32 34 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=7.975 $Y=1.32
+ $X2=8.05 $Y2=1.245
r272 32 33 276.894 $w=1.5e-07 $l=5.4e-07 $layer=POLY_cond $X=7.975 $Y=1.32
+ $X2=7.435 $Y2=1.32
r273 29 31 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.28 $Y=1.99
+ $X2=7.28 $Y2=2.275
r274 28 29 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.28 $Y=1.89 $X2=7.28
+ $Y2=1.99
r275 28 87 104.447 $w=2e-07 $l=3.15e-07 $layer=POLY_cond $X=7.28 $Y=1.89
+ $X2=7.28 $Y2=1.575
r276 24 80 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.575 $Y2=1.74
r277 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.515 $Y=1.99
+ $X2=5.515 $Y2=2.275
r278 23 80 31.9848 $w=2.95e-07 $l=1.92678e-07 $layer=POLY_cond $X=5.515 $Y=1.575
+ $X2=5.575 $Y2=1.74
r279 22 23 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=5.515 $Y=1.395
+ $X2=5.515 $Y2=1.575
r280 20 22 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.515 $Y2=1.395
r281 20 21 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=5.415 $Y=1.32
+ $X2=5.055 $Y2=1.32
r282 16 21 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=5.055 $Y2=1.32
r283 16 18 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=4.98 $Y=1.245
+ $X2=4.98 $Y2=0.415
r284 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.97 $Y=1.74
+ $X2=0.97 $Y2=2.135
r285 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.97 $Y=1.64 $X2=0.97
+ $Y2=1.74
r286 11 77 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=0.97 $Y=1.37
+ $X2=0.97 $Y2=1.235
r287 11 12 89.5258 $w=2e-07 $l=2.7e-07 $layer=POLY_cond $X=0.97 $Y=1.37 $X2=0.97
+ $Y2=1.64
r288 7 76 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r289 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r290 2 54 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.14
+ $Y=1.815 $X2=0.265 $Y2=1.96
r291 1 40 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%SCE 1 3 6 8 10 13 15 19 22 28 33 35 37
c100 35 0 4.47538e-20 $X=2.047 $Y=0.785
c101 28 0 7.84804e-20 $X=1.965 $Y=1.52
c102 15 0 1.59107e-19 $X=3.335 $Y=0.7
c103 6 0 1.4868e-19 $X=1.95 $Y=0.445
r104 35 37 1.89207 $w=3.33e-07 $l=5.5e-08 $layer=LI1_cond $X=2.047 $Y=0.785
+ $X2=2.047 $Y2=0.84
r105 28 30 81.5018 $w=2.75e-07 $l=4.65e-07 $layer=POLY_cond $X=1.965 $Y=1.577
+ $X2=2.43 $Y2=1.577
r106 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.965
+ $Y=1.52 $X2=1.965 $Y2=1.52
r107 26 28 0.876364 $w=2.75e-07 $l=5e-09 $layer=POLY_cond $X=1.96 $Y=1.577
+ $X2=1.965 $Y2=1.577
r108 25 26 1.75273 $w=2.75e-07 $l=1e-08 $layer=POLY_cond $X=1.95 $Y=1.577
+ $X2=1.96 $Y2=1.577
r109 22 35 2.62343 $w=3.35e-07 $l=8.5e-08 $layer=LI1_cond $X=2.047 $Y=0.7
+ $X2=2.047 $Y2=0.785
r110 22 29 22.8081 $w=3.33e-07 $l=6.63e-07 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=1.52
r111 22 37 0.584822 $w=3.33e-07 $l=1.7e-08 $layer=LI1_cond $X=2.047 $Y=0.857
+ $X2=2.047 $Y2=0.84
r112 20 33 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=3.42 $Y=0.95
+ $X2=3.53 $Y2=0.95
r113 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.42
+ $Y=0.95 $X2=3.42 $Y2=0.95
r114 17 19 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.42 $Y=0.785
+ $X2=3.42 $Y2=0.95
r115 16 22 5.18513 $w=1.7e-07 $l=1.68e-07 $layer=LI1_cond $X=2.215 $Y=0.7
+ $X2=2.047 $Y2=0.7
r116 15 17 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=3.42 $Y2=0.785
r117 15 16 73.0695 $w=1.68e-07 $l=1.12e-06 $layer=LI1_cond $X=3.335 $Y=0.7
+ $X2=2.215 $Y2=0.7
r118 11 33 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.95
r119 11 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.53 $Y=0.785
+ $X2=3.53 $Y2=0.445
r120 8 30 12.7119 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=1.577
r121 8 10 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.43 $Y=1.77
+ $X2=2.43 $Y2=2.165
r122 4 25 16.9318 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.95 $Y=1.385
+ $X2=1.95 $Y2=1.577
r123 4 6 482 $w=1.5e-07 $l=9.4e-07 $layer=POLY_cond $X=1.95 $Y=1.385 $X2=1.95
+ $Y2=0.445
r124 1 26 12.7119 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=1.577
r125 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.96 $Y=1.77
+ $X2=1.96 $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_319_47# 1 2 9 11 13 15 18 20 23 24 28
+ 34 36 39 40 42
c118 39 0 2.2716e-19 $X=2.55 $Y=1.04
c119 28 0 1.61748e-19 $X=3.44 $Y=1.52
r120 40 44 45.2517 $w=3.8e-07 $l=1.65e-07 $layer=POLY_cond $X=2.525 $Y=1.04
+ $X2=2.525 $Y2=0.875
r121 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.55
+ $Y=1.04 $X2=2.55 $Y2=1.04
r122 31 34 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=1.62 $Y=0.36
+ $X2=1.74 $Y2=0.36
r123 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.44
+ $Y=1.52 $X2=3.44 $Y2=1.52
r124 26 28 19.338 $w=1.93e-07 $l=3.4e-07 $layer=LI1_cond $X=3.427 $Y=1.86
+ $X2=3.427 $Y2=1.52
r125 25 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.555 $Y=1.967
+ $X2=2.47 $Y2=1.967
r126 24 26 6.83761 $w=2.15e-07 $l=1.47743e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=3.427 $Y2=1.86
r127 24 25 41.5415 $w=2.13e-07 $l=7.75e-07 $layer=LI1_cond $X=3.33 $Y=1.967
+ $X2=2.555 $Y2=1.967
r128 23 42 2.20034 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=2.47 $Y=1.86
+ $X2=2.47 $Y2=1.967
r129 22 39 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.04
r130 22 23 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=2.47 $Y=1.125
+ $X2=2.47 $Y2=1.86
r131 21 36 1.46632 $w=2.15e-07 $l=1.38e-07 $layer=LI1_cond $X=1.81 $Y=1.967
+ $X2=1.672 $Y2=1.967
r132 20 42 4.23118 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=2.47 $Y2=1.967
r133 20 21 30.8211 $w=2.13e-07 $l=5.75e-07 $layer=LI1_cond $X=2.385 $Y=1.967
+ $X2=1.81 $Y2=1.967
r134 16 36 5.02022 $w=2.22e-07 $l=1.08e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=1.967
r135 16 18 4.1907 $w=2.73e-07 $l=1e-07 $layer=LI1_cond $X=1.672 $Y=2.075
+ $X2=1.672 $Y2=2.175
r136 15 36 5.02022 $w=2.22e-07 $l=1.30434e-07 $layer=LI1_cond $X=1.62 $Y=1.86
+ $X2=1.672 $Y2=1.967
r137 14 31 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=0.36
r138 14 15 92.3155 $w=1.68e-07 $l=1.415e-06 $layer=LI1_cond $X=1.62 $Y=0.445
+ $X2=1.62 $Y2=1.86
r139 11 29 48.1208 $w=2.95e-07 $l=2.7157e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.465 $Y2=1.52
r140 11 13 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.42 $Y=1.77
+ $X2=3.42 $Y2=2.165
r141 9 44 220.489 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.51 $Y=0.445
+ $X2=2.51 $Y2=0.875
r142 2 18 600 $w=1.7e-07 $l=3.87492e-07 $layer=licon1_PDIFF $count=1 $X=1.6
+ $Y=1.845 $X2=1.725 $Y2=2.175
r143 1 34 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.595
+ $Y=0.235 $X2=1.74 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%D 1 3 6 8 15
r39 11 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.91
+ $Y=1.52 $X2=2.91 $Y2=1.52
r40 8 15 2.7938 $w=3.28e-07 $l=8e-08 $layer=LI1_cond $X=2.99 $Y=1.52 $X2=2.91
+ $Y2=1.52
r41 4 11 38.535 $w=3.06e-07 $l=2.0106e-07 $layer=POLY_cond $X=3 $Y=1.355
+ $X2=2.92 $Y2=1.52
r42 4 6 466.617 $w=1.5e-07 $l=9.1e-07 $layer=POLY_cond $X=3 $Y=1.355 $X2=3
+ $Y2=0.445
r43 1 11 47.4839 $w=3.06e-07 $l=2.64575e-07 $layer=POLY_cond $X=2.95 $Y=1.77
+ $X2=2.92 $Y2=1.52
r44 1 3 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.95 $Y=1.77 $X2=2.95
+ $Y2=2.165
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%SCD 3 6 7 9 10 13
c53 6 0 1.61748e-19 $X=3.935 $Y=1.67
c54 3 0 1.59107e-19 $X=3.91 $Y=0.445
r55 13 16 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.52
r56 13 15 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=3.995 $Y=1.355
+ $X2=3.995 $Y2=1.19
r57 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.97
+ $Y=1.355 $X2=3.97 $Y2=1.355
r58 10 14 5.13927 $w=3.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.91 $Y=1.19
+ $X2=3.91 $Y2=1.355
r59 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.935 $Y=1.77
+ $X2=3.935 $Y2=2.165
r60 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.77
r61 6 16 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=3.935 $Y=1.67 $X2=3.935
+ $Y2=1.52
r62 3 15 382.011 $w=1.5e-07 $l=7.45e-07 $layer=POLY_cond $X=3.91 $Y=0.445
+ $X2=3.91 $Y2=1.19
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_203_47# 1 2 7 9 10 12 13 15 16 18 21 25
+ 26 30 41 45 46 48 50 55 57 62 67
c205 48 0 7.21183e-20 $X=7.31 $Y=0.805
c206 46 0 1.7664e-19 $X=5.385 $Y=0.805
r207 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.53
+ $Y=0.87 $X2=7.53 $Y2=0.87
r208 59 62 25.3549 $w=3.3e-07 $l=1.45e-07 $layer=POLY_cond $X=7.385 $Y=0.87
+ $X2=7.53 $Y2=0.87
r209 54 57 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=5.45 $Y=0.87
+ $X2=5.56 $Y2=0.87
r210 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.45
+ $Y=0.87 $X2=5.45 $Y2=0.87
r211 49 63 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=7.31 $Y=0.87
+ $X2=7.53 $Y2=0.87
r212 48 50 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.31 $Y=0.805
+ $X2=7.115 $Y2=0.805
r213 48 49 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.31 $Y=0.805
+ $X2=7.31 $Y2=0.805
r214 46 50 2.14109 $w=1.4e-07 $l=1.73e-06 $layer=MET1_cond $X=5.385 $Y=0.85
+ $X2=7.115 $Y2=0.85
r215 44 55 7.33373 $w=3.28e-07 $l=2.1e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.45 $Y2=0.87
r216 44 76 6.63528 $w=3.28e-07 $l=1.9e-07 $layer=LI1_cond $X=5.24 $Y=0.87
+ $X2=5.05 $Y2=0.87
r217 43 46 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.385 $Y2=0.805
r218 43 45 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.24 $Y=0.805
+ $X2=5.045 $Y2=0.805
r219 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.24 $Y=0.805
+ $X2=5.24 $Y2=0.805
r220 41 45 4.52969 $w=1.4e-07 $l=3.66e-06 $layer=MET1_cond $X=1.385 $Y=0.85
+ $X2=5.045 $Y2=0.85
r221 39 71 57.8727 $w=2.28e-07 $l=1.155e-06 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=1.96
r222 39 67 14.7813 $w=2.28e-07 $l=2.95e-07 $layer=LI1_cond $X=1.23 $Y=0.805
+ $X2=1.23 $Y2=0.51
r223 38 41 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.24 $Y=0.805
+ $X2=1.385 $Y2=0.805
r224 38 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.24 $Y=0.805
+ $X2=1.24 $Y2=0.805
r225 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.81
+ $Y=1.74 $X2=7.81 $Y2=1.74
r226 27 30 4.88915 $w=3.28e-07 $l=1.4e-07 $layer=LI1_cond $X=7.67 $Y=1.74
+ $X2=7.81 $Y2=1.74
r227 26 63 1.57151 $w=3.28e-07 $l=4.5e-08 $layer=LI1_cond $X=7.575 $Y=0.87
+ $X2=7.53 $Y2=0.87
r228 25 27 3.96751 $w=1.9e-07 $l=1.65e-07 $layer=LI1_cond $X=7.67 $Y=1.575
+ $X2=7.67 $Y2=1.74
r229 24 26 7.47963 $w=3.3e-07 $l=2.07123e-07 $layer=LI1_cond $X=7.67 $Y=1.035
+ $X2=7.575 $Y2=0.87
r230 24 25 31.5215 $w=1.88e-07 $l=5.4e-07 $layer=LI1_cond $X=7.67 $Y=1.035
+ $X2=7.67 $Y2=1.575
r231 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.99
+ $Y=1.74 $X2=4.99 $Y2=1.74
r232 19 76 1.49285 $w=2.9e-07 $l=1.65e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=0.87
r233 19 21 28.0163 $w=2.88e-07 $l=7.05e-07 $layer=LI1_cond $X=5.05 $Y=1.035
+ $X2=5.05 $Y2=1.74
r234 16 31 46.5577 $w=3.26e-07 $l=2.89396e-07 $layer=POLY_cond $X=7.75 $Y=1.99
+ $X2=7.835 $Y2=1.74
r235 16 18 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.75 $Y=1.99
+ $X2=7.75 $Y2=2.275
r236 13 59 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=7.385 $Y=0.705
+ $X2=7.385 $Y2=0.87
r237 13 15 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=7.385 $Y=0.705
+ $X2=7.385 $Y2=0.415
r238 10 57 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=5.56 $Y=0.705
+ $X2=5.56 $Y2=0.87
r239 10 12 93.1867 $w=1.5e-07 $l=2.9e-07 $layer=POLY_cond $X=5.56 $Y=0.705
+ $X2=5.56 $Y2=0.415
r240 7 22 46.5577 $w=3.26e-07 $l=2.57391e-07 $layer=POLY_cond $X=5 $Y=1.99
+ $X2=5.015 $Y2=1.74
r241 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5 $Y=1.99 $X2=5
+ $Y2=2.275
r242 2 71 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.06
+ $Y=1.815 $X2=1.205 $Y2=1.96
r243 1 67 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_1189_183# 1 2 8 9 11 14 16 22 25 27 29
+ 31 32 35
c98 9 0 1.55016e-19 $X=6.045 $Y=1.99
r99 34 35 10.6895 $w=2.48e-07 $l=5.5e-08 $layer=POLY_cond $X=6.045 $Y=0.93
+ $X2=6.1 $Y2=0.93
r100 31 32 7.18001 $w=2.98e-07 $l=1.65e-07 $layer=LI1_cond $X=6.925 $Y=2.3
+ $X2=6.925 $Y2=2.135
r101 25 27 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=6.995 $Y=0.45
+ $X2=7.12 $Y2=0.45
r102 23 29 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.885 $Y=1.065
+ $X2=6.885 $Y2=0.915
r103 23 32 56.0506 $w=2.18e-07 $l=1.07e-06 $layer=LI1_cond $X=6.885 $Y=1.065
+ $X2=6.885 $Y2=2.135
r104 22 29 6.6318 $w=2.2e-07 $l=1.5e-07 $layer=LI1_cond $X=6.885 $Y=0.765
+ $X2=6.885 $Y2=0.915
r105 21 25 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.885 $Y=0.535
+ $X2=6.995 $Y2=0.45
r106 21 22 12.0483 $w=2.18e-07 $l=2.3e-07 $layer=LI1_cond $X=6.885 $Y=0.535
+ $X2=6.885 $Y2=0.765
r107 19 35 25.2661 $w=2.48e-07 $l=1.3e-07 $layer=POLY_cond $X=6.23 $Y=0.93
+ $X2=6.1 $Y2=0.93
r108 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.23
+ $Y=0.93 $X2=6.23 $Y2=0.93
r109 16 29 0.253446 $w=3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.775 $Y=0.915
+ $X2=6.885 $Y2=0.915
r110 16 18 20.936 $w=2.98e-07 $l=5.45e-07 $layer=LI1_cond $X=6.775 $Y=0.915
+ $X2=6.23 $Y2=0.915
r111 12 35 14.534 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=6.1 $Y=0.795
+ $X2=6.1 $Y2=0.93
r112 12 14 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.1 $Y=0.795
+ $X2=6.1 $Y2=0.445
r113 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.045 $Y=1.99
+ $X2=6.045 $Y2=2.275
r114 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=6.045 $Y=1.89 $X2=6.045
+ $Y2=1.99
r115 7 34 7.89931 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=6.045 $Y=1.065
+ $X2=6.045 $Y2=0.93
r116 7 8 273.551 $w=2e-07 $l=8.25e-07 $layer=POLY_cond $X=6.045 $Y=1.065
+ $X2=6.045 $Y2=1.89
r117 2 31 600 $w=1.7e-07 $l=6.33364e-07 $layer=licon1_PDIFF $count=1 $X=6.845
+ $Y=1.735 $X2=6.99 $Y2=2.3
r118 1 27 182 $w=1.7e-07 $l=2.85832e-07 $layer=licon1_NDIFF $count=1 $X=6.955
+ $Y=0.235 $X2=7.12 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_1011_47# 1 2 8 9 11 14 15 16 17 18 19
+ 23 28 30 31 33
r117 36 37 15.25 $w=2.76e-07 $l=3.45e-07 $layer=LI1_cond $X=5.81 $Y=1.41
+ $X2=6.155 $Y2=1.41
r118 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.52
+ $Y=1.41 $X2=6.52 $Y2=1.41
r119 31 37 4.4292 $w=3.3e-07 $l=1.1e-07 $layer=LI1_cond $X=6.265 $Y=1.41
+ $X2=6.155 $Y2=1.41
r120 31 33 8.90524 $w=3.28e-07 $l=2.55e-07 $layer=LI1_cond $X=6.265 $Y=1.41
+ $X2=6.52 $Y2=1.41
r121 29 37 2.0678 $w=2.2e-07 $l=1.65e-07 $layer=LI1_cond $X=6.155 $Y=1.575
+ $X2=6.155 $Y2=1.41
r122 29 30 32.216 $w=2.18e-07 $l=6.15e-07 $layer=LI1_cond $X=6.155 $Y=1.575
+ $X2=6.155 $Y2=2.19
r123 28 36 3.57235 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.81 $Y=1.245
+ $X2=5.81 $Y2=1.41
r124 27 28 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=5.81 $Y=0.535
+ $X2=5.81 $Y2=1.245
r125 23 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.725 $Y=0.45
+ $X2=5.81 $Y2=0.535
r126 23 25 27.7273 $w=1.68e-07 $l=4.25e-07 $layer=LI1_cond $X=5.725 $Y=0.45
+ $X2=5.3 $Y2=0.45
r127 19 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=6.155 $Y2=2.19
r128 19 21 51.2139 $w=1.68e-07 $l=7.85e-07 $layer=LI1_cond $X=6.045 $Y=2.275
+ $X2=5.26 $Y2=2.275
r129 17 34 29.9935 $w=2.7e-07 $l=1.35e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.52 $Y2=1.41
r130 17 18 0.448535 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=6.655 $Y=1.41
+ $X2=6.755 $Y2=1.467
r131 15 16 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=6.805 $Y=0.95
+ $X2=6.805 $Y2=1.1
r132 14 15 126.927 $w=1.5e-07 $l=3.95e-07 $layer=POLY_cond $X=6.88 $Y=0.555
+ $X2=6.88 $Y2=0.95
r133 9 18 27.0491 $w=1.9e-07 $l=1.93e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=1.467
r134 9 11 120.5 $w=1.8e-07 $l=4.5e-07 $layer=POLY_cond $X=6.755 $Y=1.66
+ $X2=6.755 $Y2=2.11
r135 8 18 27.0491 $w=1.9e-07 $l=1.92e-07 $layer=POLY_cond $X=6.755 $Y=1.275
+ $X2=6.755 $Y2=1.467
r136 8 16 58.026 $w=2e-07 $l=1.75e-07 $layer=POLY_cond $X=6.755 $Y=1.275
+ $X2=6.755 $Y2=1.1
r137 2 21 600 $w=1.7e-07 $l=2.82489e-07 $layer=licon1_PDIFF $count=1 $X=5.09
+ $Y=2.065 $X2=5.26 $Y2=2.275
r138 1 25 182 $w=1.7e-07 $l=3.35708e-07 $layer=licon1_NDIFF $count=1 $X=5.055
+ $Y=0.235 $X2=5.3 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_1667_315# 1 2 7 9 12 14 16 17 19 20 22
+ 23 25 26 33 36 38 41 45 48 49 54
r94 54 55 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=10.48 $Y=1.202
+ $X2=10.505 $Y2=1.202
r95 51 52 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=9.985 $Y=1.202
+ $X2=10.01 $Y2=1.202
r96 45 47 16.9646 $w=3.58e-07 $l=4.4e-07 $layer=LI1_cond $X=9.32 $Y=0.385
+ $X2=9.32 $Y2=0.825
r97 42 54 55.1763 $w=3.8e-07 $l=4.35e-07 $layer=POLY_cond $X=10.045 $Y=1.202
+ $X2=10.48 $Y2=1.202
r98 42 52 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=10.045 $Y=1.202
+ $X2=10.01 $Y2=1.202
r99 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.045
+ $Y=1.16 $X2=10.045 $Y2=1.16
r100 39 49 0.674692 $w=3.3e-07 $l=9.3e-08 $layer=LI1_cond $X=9.505 $Y=1.16
+ $X2=9.412 $Y2=1.16
r101 39 41 18.8582 $w=3.28e-07 $l=5.4e-07 $layer=LI1_cond $X=9.505 $Y=1.16
+ $X2=10.045 $Y2=1.16
r102 38 48 6.7841 $w=2.35e-07 $l=1.88348e-07 $layer=LI1_cond $X=9.412 $Y=1.575
+ $X2=9.362 $Y2=1.74
r103 37 49 8.18839 $w=1.82e-07 $l=1.65e-07 $layer=LI1_cond $X=9.412 $Y=1.325
+ $X2=9.412 $Y2=1.16
r104 37 38 14.9877 $w=1.83e-07 $l=2.5e-07 $layer=LI1_cond $X=9.412 $Y=1.325
+ $X2=9.412 $Y2=1.575
r105 36 49 8.18839 $w=1.82e-07 $l=1.65997e-07 $layer=LI1_cond $X=9.41 $Y=0.995
+ $X2=9.412 $Y2=1.16
r106 36 47 10.4747 $w=1.78e-07 $l=1.7e-07 $layer=LI1_cond $X=9.41 $Y=0.995
+ $X2=9.41 $Y2=0.825
r107 31 48 6.7841 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=9.362 $Y=1.905
+ $X2=9.362 $Y2=1.74
r108 31 33 1.81965 $w=2.83e-07 $l=4.5e-08 $layer=LI1_cond $X=9.362 $Y=1.905
+ $X2=9.362 $Y2=1.95
r109 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.64
+ $Y=1.74 $X2=8.64 $Y2=1.74
r110 26 48 0.153733 $w=3.3e-07 $l=1.42e-07 $layer=LI1_cond $X=9.22 $Y=1.74
+ $X2=9.362 $Y2=1.74
r111 26 28 20.2551 $w=3.28e-07 $l=5.8e-07 $layer=LI1_cond $X=9.22 $Y=1.74
+ $X2=8.64 $Y2=1.74
r112 23 55 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=10.505 $Y=0.995
+ $X2=10.505 $Y2=1.202
r113 23 25 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=10.505 $Y=0.995
+ $X2=10.505 $Y2=0.56
r114 20 54 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.48 $Y=1.41
+ $X2=10.48 $Y2=1.202
r115 20 22 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.48 $Y=1.41
+ $X2=10.48 $Y2=1.985
r116 17 52 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.202
r117 17 19 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.01 $Y=1.41
+ $X2=10.01 $Y2=1.985
r118 14 51 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=9.985 $Y=0.995
+ $X2=9.985 $Y2=1.202
r119 14 16 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.985 $Y=0.995
+ $X2=9.985 $Y2=0.56
r120 10 29 39.3952 $w=3.9e-07 $l=1.79374e-07 $layer=POLY_cond $X=8.525 $Y=1.575
+ $X2=8.555 $Y2=1.74
r121 10 12 579.426 $w=1.5e-07 $l=1.13e-06 $layer=POLY_cond $X=8.525 $Y=1.575
+ $X2=8.525 $Y2=0.445
r122 7 29 44.9977 $w=3.9e-07 $l=3.04138e-07 $layer=POLY_cond $X=8.435 $Y=1.99
+ $X2=8.555 $Y2=1.74
r123 7 9 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=8.435 $Y=1.99
+ $X2=8.435 $Y2=2.275
r124 2 33 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=9.18
+ $Y=1.485 $X2=9.305 $Y2=1.95
r125 1 45 91 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_NDIFF $count=2 $X=9.18
+ $Y=0.235 $X2=9.305 $Y2=0.385
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_1474_413# 1 2 7 9 10 12 13 14 15 19 26
+ 29 32 33
c86 14 0 1.26472e-19 $X=9.54 $Y=1.202
r87 32 34 11.1226 $w=3.48e-07 $l=2.45e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=8.16 $Y2=1.405
r88 32 33 7.01492 $w=3.48e-07 $l=1.65e-07 $layer=LI1_cond $X=8.16 $Y=1.16
+ $X2=8.16 $Y2=0.995
r89 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.065
+ $Y=1.16 $X2=9.065 $Y2=1.16
r90 27 32 1.07274 $w=3.3e-07 $l=1.75e-07 $layer=LI1_cond $X=8.335 $Y=1.16
+ $X2=8.16 $Y2=1.16
r91 27 29 25.4934 $w=3.28e-07 $l=7.3e-07 $layer=LI1_cond $X=8.335 $Y=1.16
+ $X2=9.065 $Y2=1.16
r92 26 34 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=8.25 $Y=2.165
+ $X2=8.25 $Y2=1.405
r93 23 33 24.0965 $w=2.18e-07 $l=4.6e-07 $layer=LI1_cond $X=8.095 $Y=0.535
+ $X2=8.095 $Y2=0.995
r94 19 23 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=7.985 $Y=0.45
+ $X2=8.095 $Y2=0.535
r95 19 21 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=7.985 $Y=0.45
+ $X2=7.73 $Y2=0.45
r96 15 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=8.165 $Y=2.25
+ $X2=8.25 $Y2=2.165
r97 15 17 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=8.165 $Y=2.25
+ $X2=7.515 $Y2=2.25
r98 13 30 65.573 $w=3.3e-07 $l=3.75e-07 $layer=POLY_cond $X=9.44 $Y=1.16
+ $X2=9.065 $Y2=1.16
r99 13 14 3.90195 $w=3.3e-07 $l=1.19164e-07 $layer=POLY_cond $X=9.44 $Y=1.16
+ $X2=9.54 $Y2=1.202
r100 10 14 34.7346 $w=1.65e-07 $l=2.19144e-07 $layer=POLY_cond $X=9.565 $Y=0.995
+ $X2=9.54 $Y2=1.202
r101 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=9.565 $Y=0.995
+ $X2=9.565 $Y2=0.56
r102 7 14 34.7346 $w=1.65e-07 $l=2.08e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.202
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.54 $Y=1.41
+ $X2=9.54 $Y2=1.985
r104 2 17 600 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_PDIFF $count=1 $X=7.37
+ $Y=2.065 $X2=7.515 $Y2=2.25
r105 1 21 182 $w=1.7e-07 $l=3.6187e-07 $layer=licon1_NDIFF $count=1 $X=7.46
+ $Y=0.235 $X2=7.73 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%VPWR 1 2 3 4 5 6 7 24 28 32 36 40 44 46
+ 48 51 52 54 55 57 58 60 61 62 64 69 96 101 104 108
c156 1 0 1.76957e-19 $X=0.59 $Y=1.815
r157 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=2.72
+ $X2=10.81 $Y2=2.72
r158 104 105 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r159 101 102 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r160 99 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=10.81 $Y2=2.72
r161 98 99 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r162 96 107 3.40825 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=10.67 $Y=2.72
+ $X2=10.855 $Y2=2.72
r163 96 98 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.67 $Y=2.72
+ $X2=10.35 $Y2=2.72
r164 95 99 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r165 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r166 92 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r167 91 92 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r168 89 92 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r169 88 91 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=6.67 $Y=2.72
+ $X2=8.51 $Y2=2.72
r170 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r171 86 89 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r172 85 86 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r173 83 86 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r174 82 85 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r175 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r176 80 83 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r177 79 80 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r178 77 80 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r179 77 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r180 76 79 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r181 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r182 74 104 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.17 $Y2=2.72
r183 74 76 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.36 $Y=2.72
+ $X2=2.53 $Y2=2.72
r184 73 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r185 73 102 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r186 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r187 70 101 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.9 $Y=2.72
+ $X2=0.71 $Y2=2.72
r188 70 72 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=0.9 $Y=2.72
+ $X2=1.61 $Y2=2.72
r189 69 104 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=2.17 $Y2=2.72
r190 69 72 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=1.98 $Y=2.72
+ $X2=1.61 $Y2=2.72
r191 64 101 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.71 $Y2=2.72
r192 64 66 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=0.52 $Y=2.72
+ $X2=0.23 $Y2=2.72
r193 62 102 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r194 62 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r195 60 94 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.43 $Y2=2.72
r196 60 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=2.72
+ $X2=9.775 $Y2=2.72
r197 59 98 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=10.35 $Y2=2.72
r198 59 61 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=2.72
+ $X2=9.775 $Y2=2.72
r199 57 91 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.51 $Y2=2.72
r200 57 58 8.14251 $w=1.7e-07 $l=1.52e-07 $layer=LI1_cond $X=8.565 $Y=2.72
+ $X2=8.717 $Y2=2.72
r201 56 94 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=9.43 $Y2=2.72
r202 56 58 8.14251 $w=1.7e-07 $l=1.53e-07 $layer=LI1_cond $X=8.87 $Y=2.72
+ $X2=8.717 $Y2=2.72
r203 54 85 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=6.435 $Y=2.72
+ $X2=6.21 $Y2=2.72
r204 54 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.435 $Y=2.72
+ $X2=6.52 $Y2=2.72
r205 53 88 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.67 $Y2=2.72
r206 53 55 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.605 $Y=2.72
+ $X2=6.52 $Y2=2.72
r207 51 79 13.0481 $w=1.68e-07 $l=2e-07 $layer=LI1_cond $X=4.11 $Y=2.72 $X2=3.91
+ $Y2=2.72
r208 51 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.11 $Y=2.72
+ $X2=4.195 $Y2=2.72
r209 50 82 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4.28 $Y=2.72 $X2=4.37
+ $Y2=2.72
r210 50 52 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.28 $Y=2.72
+ $X2=4.195 $Y2=2.72
r211 46 107 3.40825 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=10.755 $Y=2.635
+ $X2=10.855 $Y2=2.72
r212 46 48 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=10.755 $Y=2.635
+ $X2=10.755 $Y2=2.01
r213 42 61 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=2.72
r214 42 44 55.1283 $w=1.68e-07 $l=8.45e-07 $layer=LI1_cond $X=9.775 $Y=2.635
+ $X2=9.775 $Y2=1.79
r215 38 58 0.649941 $w=3.05e-07 $l=8.5e-08 $layer=LI1_cond $X=8.717 $Y=2.635
+ $X2=8.717 $Y2=2.72
r216 38 40 12.658 $w=3.03e-07 $l=3.35e-07 $layer=LI1_cond $X=8.717 $Y=2.635
+ $X2=8.717 $Y2=2.3
r217 34 55 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=2.72
r218 34 36 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.52 $Y=2.635
+ $X2=6.52 $Y2=2
r219 30 52 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.72
r220 30 32 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.195 $Y=2.635
+ $X2=4.195 $Y2=2.33
r221 26 104 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.72
r222 26 28 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=2.17 $Y=2.635
+ $X2=2.17 $Y2=2.33
r223 22 101 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.72
r224 22 24 12.5859 $w=3.78e-07 $l=4.15e-07 $layer=LI1_cond $X=0.71 $Y=2.635
+ $X2=0.71 $Y2=2.22
r225 7 48 300 $w=1.7e-07 $l=6.10533e-07 $layer=licon1_PDIFF $count=2 $X=10.57
+ $Y=1.485 $X2=10.755 $Y2=2.01
r226 6 44 300 $w=1.7e-07 $l=3.70473e-07 $layer=licon1_PDIFF $count=2 $X=9.63
+ $Y=1.485 $X2=9.775 $Y2=1.79
r227 5 40 600 $w=1.7e-07 $l=3.53483e-07 $layer=licon1_PDIFF $count=1 $X=8.525
+ $Y=2.065 $X2=8.78 $Y2=2.3
r228 4 36 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=6.135
+ $Y=2.065 $X2=6.52 $Y2=2
r229 3 32 600 $w=1.7e-07 $l=5.63627e-07 $layer=licon1_PDIFF $count=1 $X=4.025
+ $Y=1.845 $X2=4.195 $Y2=2.33
r230 2 28 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=2.05
+ $Y=1.845 $X2=2.195 $Y2=2.33
r231 1 24 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=1.815 $X2=0.735 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%A_608_369# 1 2 3 4 13 17 22 24 25 26 27
+ 28 30 32 36 38 39
c113 30 0 1.7664e-19 $X=4.65 $Y=0.695
r114 39 41 21.3062 $w=2.09e-07 $l=3.65e-07 $layer=LI1_cond $X=4.682 $Y=1.91
+ $X2=4.682 $Y2=2.275
r115 33 36 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=4.65 $Y=0.45 $X2=4.75
+ $Y2=0.45
r116 32 39 5.42244 $w=2.09e-07 $l=9.97246e-08 $layer=LI1_cond $X=4.65 $Y=1.825
+ $X2=4.682 $Y2=1.91
r117 31 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=0.78
r118 31 32 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.65 $Y=0.865
+ $X2=4.65 $Y2=1.825
r119 30 38 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.695
+ $X2=4.65 $Y2=0.78
r120 29 33 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.45
r121 29 30 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=4.65 $Y=0.535
+ $X2=4.65 $Y2=0.695
r122 27 38 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=4.65 $Y2=0.78
r123 27 28 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=4.565 $Y=0.78
+ $X2=3.895 $Y2=0.78
r124 25 39 1.94907 $w=1.7e-07 $l=1.17e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=4.682 $Y2=1.91
r125 25 26 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.565 $Y=1.91
+ $X2=3.89 $Y2=1.91
r126 24 28 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.81 $Y=0.695
+ $X2=3.895 $Y2=0.78
r127 23 24 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.81 $Y=0.445
+ $X2=3.81 $Y2=0.695
r128 21 26 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.89 $Y2=1.91
r129 21 22 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=3.805 $Y=1.995
+ $X2=3.805 $Y2=2.245
r130 17 23 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.81 $Y2=0.445
r131 17 19 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=3.725 $Y=0.36
+ $X2=3.265 $Y2=0.36
r132 13 22 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.805 $Y2=2.245
r133 13 15 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=3.72 $Y=2.33
+ $X2=3.185 $Y2=2.33
r134 4 41 600 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_PDIFF $count=1 $X=4.59
+ $Y=2.065 $X2=4.715 $Y2=2.275
r135 3 15 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=1.845 $X2=3.185 $Y2=2.33
r136 2 36 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=4.625
+ $Y=0.235 $X2=4.75 $Y2=0.45
r137 1 19 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=3.075
+ $Y=0.235 $X2=3.265 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%Q 1 2 10 13 19 24 25
c32 25 0 1.26472e-19 $X=10.265 $Y=1.545
r33 24 25 7.30169 $w=4.68e-07 $l=8.5e-08 $layer=LI1_cond $X=10.265 $Y=1.63
+ $X2=10.265 $Y2=1.545
r34 19 21 11.3246 $w=4.68e-07 $l=4.45e-07 $layer=LI1_cond $X=10.265 $Y=1.865
+ $X2=10.265 $Y2=2.31
r35 13 16 0.203588 $w=4.68e-07 $l=8e-09 $layer=LI1_cond $X=10.265 $Y=1.772
+ $X2=10.265 $Y2=1.78
r36 13 24 3.61368 $w=4.68e-07 $l=1.42e-07 $layer=LI1_cond $X=10.265 $Y=1.772
+ $X2=10.265 $Y2=1.63
r37 13 19 0.203588 $w=4.68e-07 $l=8e-09 $layer=LI1_cond $X=10.265 $Y=1.857
+ $X2=10.265 $Y2=1.865
r38 13 16 1.95953 $w=4.68e-07 $l=7.7e-08 $layer=LI1_cond $X=10.265 $Y=1.857
+ $X2=10.265 $Y2=1.78
r39 12 25 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=10.415 $Y=0.82
+ $X2=10.415 $Y2=1.545
r40 10 12 15.9542 $w=4.68e-07 $l=4.25e-07 $layer=LI1_cond $X=10.265 $Y=0.395
+ $X2=10.265 $Y2=0.82
r41 2 24 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=1.63
r42 2 21 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=10.1
+ $Y=1.485 $X2=10.245 $Y2=2.31
r43 1 10 91 $w=1.7e-07 $l=2.52636e-07 $layer=licon1_NDIFF $count=2 $X=10.06
+ $Y=0.235 $X2=10.245 $Y2=0.395
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFXTP_2%VGND 1 2 3 4 5 6 7 24 28 32 36 40 42 44
+ 47 48 50 51 53 54 56 57 58 60 84 92 98 104 108
c157 108 0 2.71124e-20 $X=10.81 $Y=0
r158 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r159 104 105 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r160 98 101 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=0
+ $X2=0.705 $Y2=0.38
r161 98 99 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r162 95 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=10.81 $Y2=0
r163 94 95 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r164 92 107 3.40825 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=10.67 $Y=0
+ $X2=10.855 $Y2=0
r165 92 94 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=10.67 $Y=0 $X2=10.35
+ $Y2=0
r166 91 95 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r167 91 105 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=8.51 $Y2=0
r168 90 91 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0 $X2=9.43
+ $Y2=0
r169 88 104 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.87 $Y=0 $X2=8.66
+ $Y2=0
r170 88 90 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.87 $Y=0 $X2=9.43
+ $Y2=0
r171 87 105 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=8.51 $Y2=0
r172 86 87 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r173 84 104 10.1275 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=8.45 $Y=0 $X2=8.66
+ $Y2=0
r174 84 86 116.128 $w=1.68e-07 $l=1.78e-06 $layer=LI1_cond $X=8.45 $Y=0 $X2=6.67
+ $Y2=0
r175 83 87 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r176 82 83 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=0
+ $X2=6.21 $Y2=0
r177 80 83 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=6.21 $Y2=0
r178 79 82 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=6.21
+ $Y2=0
r179 79 80 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=0
+ $X2=4.37 $Y2=0
r180 77 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r181 76 77 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r182 74 77 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r183 73 76 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r184 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r185 71 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r186 70 71 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r187 68 71 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r188 68 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r189 67 70 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r190 67 68 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r191 65 98 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.705
+ $Y2=0
r192 65 67 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r193 60 98 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.705
+ $Y2=0
r194 60 62 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0
+ $X2=0.23 $Y2=0
r195 58 99 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r196 58 62 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r197 56 90 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=9.69 $Y=0 $X2=9.43
+ $Y2=0
r198 56 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.69 $Y=0 $X2=9.775
+ $Y2=0
r199 55 94 31.9679 $w=1.68e-07 $l=4.9e-07 $layer=LI1_cond $X=9.86 $Y=0 $X2=10.35
+ $Y2=0
r200 55 57 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.86 $Y=0 $X2=9.775
+ $Y2=0
r201 53 82 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.21
+ $Y2=0
r202 53 54 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.225 $Y=0 $X2=6.41
+ $Y2=0
r203 52 86 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.67
+ $Y2=0
r204 52 54 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=6.595 $Y=0 $X2=6.41
+ $Y2=0
r205 50 76 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=4.115 $Y=0
+ $X2=3.91 $Y2=0
r206 50 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.115 $Y=0 $X2=4.215
+ $Y2=0
r207 49 79 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.37
+ $Y2=0
r208 49 51 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=4.315 $Y=0 $X2=4.215
+ $Y2=0
r209 47 70 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.07
+ $Y2=0
r210 47 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r211 46 73 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.53
+ $Y2=0
r212 46 48 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r213 42 107 3.40825 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=10.755 $Y=0.085
+ $X2=10.855 $Y2=0
r214 42 44 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=10.755 $Y=0.085
+ $X2=10.755 $Y2=0.395
r215 38 57 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.775 $Y=0.085
+ $X2=9.775 $Y2=0
r216 38 40 29.0321 $w=1.68e-07 $l=4.45e-07 $layer=LI1_cond $X=9.775 $Y=0.085
+ $X2=9.775 $Y2=0.53
r217 34 104 1.60615 $w=4.2e-07 $l=8.5e-08 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0
r218 34 36 10.0153 $w=4.18e-07 $l=3.65e-07 $layer=LI1_cond $X=8.66 $Y=0.085
+ $X2=8.66 $Y2=0.45
r219 30 54 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0
r220 30 32 10.4343 $w=3.68e-07 $l=3.35e-07 $layer=LI1_cond $X=6.41 $Y=0.085
+ $X2=6.41 $Y2=0.42
r221 26 51 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0
r222 26 28 15.25 $w=1.98e-07 $l=2.75e-07 $layer=LI1_cond $X=4.215 $Y=0.085
+ $X2=4.215 $Y2=0.36
r223 22 48 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r224 22 24 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.36
r225 7 44 182 $w=1.7e-07 $l=2.42126e-07 $layer=licon1_NDIFF $count=1 $X=10.58
+ $Y=0.235 $X2=10.755 $Y2=0.395
r226 6 40 182 $w=1.7e-07 $l=3.5616e-07 $layer=licon1_NDIFF $count=1 $X=9.64
+ $Y=0.235 $X2=9.775 $Y2=0.53
r227 5 36 182 $w=1.7e-07 $l=2.93258e-07 $layer=licon1_NDIFF $count=1 $X=8.6
+ $Y=0.235 $X2=8.785 $Y2=0.45
r228 4 32 182 $w=1.7e-07 $l=3.86588e-07 $layer=licon1_NDIFF $count=1 $X=6.175
+ $Y=0.235 $X2=6.48 $Y2=0.42
r229 3 28 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=3.985
+ $Y=0.235 $X2=4.2 $Y2=0.36
r230 2 24 182 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=1 $X=2.025
+ $Y=0.235 $X2=2.29 $Y2=0.36
r231 1 101 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

