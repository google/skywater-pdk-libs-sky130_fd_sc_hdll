# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__or2b_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__or2b_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.730000 1.075000 2.470000 1.275000 ;
    END
  END A
  PIN B_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.425000 1.955000 ;
    END
  END B_N
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.475000 0.290000 2.855000 0.735000 ;
        RECT 2.475000 0.735000 4.490000 0.905000 ;
        RECT 2.565000 1.785000 3.755000 1.955000 ;
        RECT 2.565000 1.955000 2.815000 2.465000 ;
        RECT 3.080000 1.445000 4.490000 1.615000 ;
        RECT 3.080000 1.615000 3.755000 1.785000 ;
        RECT 3.415000 0.290000 3.795000 0.735000 ;
        RECT 3.505000 1.955000 3.755000 2.465000 ;
        RECT 4.105000 0.905000 4.490000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.640000  0.085000 1.295000 0.565000 ;
        RECT 2.130000  0.085000 2.305000 0.905000 ;
        RECT 3.075000  0.085000 3.245000 0.550000 ;
        RECT 4.015000  0.085000 4.185000 0.550000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.090000 2.125000 0.345000 2.635000 ;
        RECT 2.065000 1.835000 2.345000 2.635000 ;
        RECT 3.035000 2.135000 3.285000 2.635000 ;
        RECT 3.975000 1.795000 4.225000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.110000 0.265000 0.420000 0.735000 ;
      RECT 0.110000 0.735000 0.895000 0.905000 ;
      RECT 0.645000 0.905000 0.895000 0.995000 ;
      RECT 0.645000 0.995000 1.170000 1.325000 ;
      RECT 0.645000 1.325000 0.815000 2.465000 ;
      RECT 1.040000 1.495000 2.860000 1.615000 ;
      RECT 1.040000 1.615000 1.560000 2.465000 ;
      RECT 1.340000 0.735000 1.845000 0.905000 ;
      RECT 1.340000 0.905000 1.560000 1.445000 ;
      RECT 1.340000 1.445000 2.860000 1.495000 ;
      RECT 1.465000 0.305000 1.845000 0.735000 ;
      RECT 2.690000 1.075000 3.800000 1.245000 ;
      RECT 2.690000 1.245000 2.860000 1.445000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or2b_4
