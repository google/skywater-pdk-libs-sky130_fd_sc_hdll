* File: sky130_fd_sc_hdll__a211o_1.pex.spice
* Created: Wed Sep  2 08:15:42 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211O_1%A_80_21# 1 2 3 10 12 13 15 19 21 22 23 24
+ 27 29 33 37 39 41
r96 40 41 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=0.475 $Y=1.202
+ $X2=0.5 $Y2=1.202
r97 35 37 4.86587 $w=2.23e-07 $l=9.5e-08 $layer=LI1_cond $X=3.422 $Y=0.625
+ $X2=3.422 $Y2=0.53
r98 31 33 5.59274 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=3.375 $Y=1.685
+ $X2=3.375 $Y2=1.85
r99 30 39 7.86615 $w=1.9e-07 $l=1.63e-07 $layer=LI1_cond $X=2.52 $Y=0.72
+ $X2=2.357 $Y2=0.72
r100 29 35 6.87974 $w=1.9e-07 $l=1.52263e-07 $layer=LI1_cond $X=3.31 $Y=0.72
+ $X2=3.422 $Y2=0.625
r101 29 30 46.1148 $w=1.88e-07 $l=7.9e-07 $layer=LI1_cond $X=3.31 $Y=0.72
+ $X2=2.52 $Y2=0.72
r102 25 39 0.497779 $w=3.25e-07 $l=9.5e-08 $layer=LI1_cond $X=2.357 $Y=0.625
+ $X2=2.357 $Y2=0.72
r103 25 27 3.36868 $w=3.23e-07 $l=9.5e-08 $layer=LI1_cond $X=2.357 $Y=0.625
+ $X2=2.357 $Y2=0.53
r104 23 31 7.6914 $w=1.8e-07 $l=2.10238e-07 $layer=LI1_cond $X=3.205 $Y=1.595
+ $X2=3.375 $Y2=1.685
r105 23 24 145.414 $w=1.78e-07 $l=2.36e-06 $layer=LI1_cond $X=3.205 $Y=1.595
+ $X2=0.845 $Y2=1.595
r106 21 39 7.86615 $w=1.9e-07 $l=1.62e-07 $layer=LI1_cond $X=2.195 $Y=0.72
+ $X2=2.357 $Y2=0.72
r107 21 22 78.8038 $w=1.88e-07 $l=1.35e-06 $layer=LI1_cond $X=2.195 $Y=0.72
+ $X2=0.845 $Y2=0.72
r108 20 41 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=0.735 $Y=1.202
+ $X2=0.5 $Y2=1.202
r109 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.735
+ $Y=1.16 $X2=0.735 $Y2=1.16
r110 17 24 6.999 $w=1.8e-07 $l=1.58745e-07 $layer=LI1_cond $X=0.725 $Y=1.505
+ $X2=0.845 $Y2=1.595
r111 17 19 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.725 $Y=1.505
+ $X2=0.725 $Y2=1.16
r112 16 22 6.93705 $w=1.9e-07 $l=1.60624e-07 $layer=LI1_cond $X=0.725 $Y=0.815
+ $X2=0.845 $Y2=0.72
r113 16 19 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.725 $Y=0.815
+ $X2=0.725 $Y2=1.16
r114 13 41 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.5 $Y2=1.202
r115 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.5 $Y=1.41
+ $X2=0.5 $Y2=1.985
r116 10 40 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r117 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r118 3 33 300 $w=1.7e-07 $l=4.33561e-07 $layer=licon1_PDIFF $count=2 $X=3.26
+ $Y=1.485 $X2=3.41 $Y2=1.85
r119 2 37 182 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_NDIFF $count=1 $X=3.22
+ $Y=0.235 $X2=3.41 $Y2=0.53
r120 1 27 182 $w=1.7e-07 $l=3.60278e-07 $layer=licon1_NDIFF $count=1 $X=2.26
+ $Y=0.235 $X2=2.405 $Y2=0.53
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%A2 1 3 4 6 7 8 14 17
r33 14 15 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=1.5 $Y=1.202
+ $X2=1.525 $Y2=1.202
r34 12 14 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=1.265 $Y=1.202
+ $X2=1.5 $Y2=1.202
r35 7 8 11.8737 $w=3.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.21 $Y=1.16 $X2=1.55
+ $Y2=1.16
r36 7 17 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=1.21 $Y=1.16 $X2=1.16
+ $Y2=1.16
r37 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.265
+ $Y=1.16 $X2=1.265 $Y2=1.16
r38 4 15 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.525 $Y=0.995
+ $X2=1.525 $Y2=1.202
r39 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.525 $Y=0.995
+ $X2=1.525 $Y2=0.56
r40 1 14 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.5 $Y=1.41 $X2=1.5
+ $Y2=1.202
r41 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.5 $Y=1.41 $X2=1.5
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%A1 1 3 4 6 7 15
r30 10 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.125
+ $Y=1.16 $X2=2.125 $Y2=1.16
r31 7 15 0.523838 $w=3.28e-07 $l=1.5e-08 $layer=LI1_cond $X=2.09 $Y=1.16
+ $X2=2.105 $Y2=1.16
r32 4 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.185 $Y=0.995
+ $X2=2.1 $Y2=1.16
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.185 $Y=0.995
+ $X2=2.185 $Y2=0.56
r34 1 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.16 $Y=1.41
+ $X2=2.1 $Y2=1.16
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.16 $Y=1.41 $X2=2.16
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%B1 1 3 4 6 7 14
r30 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.675
+ $Y=1.16 $X2=2.675 $Y2=1.16
r31 7 14 9.25447 $w=3.28e-07 $l=2.65e-07 $layer=LI1_cond $X=2.94 $Y=1.16
+ $X2=2.675 $Y2=1.16
r32 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.64 $Y=1.41
+ $X2=2.7 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.64 $Y=1.41 $X2=2.64
+ $Y2=1.985
r34 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.615 $Y=0.995
+ $X2=2.7 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.615 $Y=0.995
+ $X2=2.615 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%C1 1 3 4 6 7 10 17
r27 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=3.17 $Y=1.202
+ $X2=3.405 $Y2=1.202
r28 9 10 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=3.145 $Y=1.202
+ $X2=3.17 $Y2=1.202
r29 7 17 1.74613 $w=3.28e-07 $l=5e-08 $layer=LI1_cond $X=3.405 $Y=1.16 $X2=3.455
+ $Y2=1.16
r30 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.405
+ $Y=1.16 $X2=3.405 $Y2=1.16
r31 4 10 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.17 $Y=1.41
+ $X2=3.17 $Y2=1.202
r32 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.17 $Y=1.41 $X2=3.17
+ $Y2=1.985
r33 1 9 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=1.202
r34 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.145 $Y=0.995
+ $X2=3.145 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%X 1 2 7 8 9 10 11 12 22 38
r16 20 38 0.412815 $w=3.33e-07 $l=1.2e-08 $layer=LI1_cond $X=0.257 $Y=1.518
+ $X2=0.257 $Y2=1.53
r17 11 12 14.7861 $w=2.63e-07 $l=3.4e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=2.21
r18 11 41 8.04536 $w=2.63e-07 $l=1.85e-07 $layer=LI1_cond $X=0.222 $Y=1.87
+ $X2=0.222 $Y2=1.685
r19 10 41 4.62931 $w=3.33e-07 $l=1.19e-07 $layer=LI1_cond $X=0.257 $Y=1.566
+ $X2=0.257 $Y2=1.685
r20 10 38 1.23845 $w=3.33e-07 $l=3.6e-08 $layer=LI1_cond $X=0.257 $Y=1.566
+ $X2=0.257 $Y2=1.53
r21 10 20 1.27285 $w=3.33e-07 $l=3.7e-08 $layer=LI1_cond $X=0.257 $Y=1.481
+ $X2=0.257 $Y2=1.518
r22 9 10 10.0108 $w=3.33e-07 $l=2.91e-07 $layer=LI1_cond $X=0.257 $Y=1.19
+ $X2=0.257 $Y2=1.481
r23 8 9 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=0.85
+ $X2=0.257 $Y2=1.19
r24 7 8 11.6964 $w=3.33e-07 $l=3.4e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.85
r25 7 22 3.78414 $w=3.33e-07 $l=1.1e-07 $layer=LI1_cond $X=0.257 $Y=0.51
+ $X2=0.257 $Y2=0.4
r26 2 10 300 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.65
r27 1 22 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%VPWR 1 2 9 11 13 25 26 29 34 40 44
r50 38 40 6.44552 $w=5.38e-07 $l=1.5e-08 $layer=LI1_cond $X=2.07 $Y=2.535
+ $X2=2.085 $Y2=2.535
r51 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r52 36 38 7.30937 $w=5.38e-07 $l=3.3e-07 $layer=LI1_cond $X=1.74 $Y=2.535
+ $X2=2.07 $Y2=2.535
r53 33 39 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r54 32 36 2.87945 $w=5.38e-07 $l=1.3e-07 $layer=LI1_cond $X=1.61 $Y=2.535
+ $X2=1.74 $Y2=2.535
r55 32 34 7.99599 $w=5.38e-07 $l=8.5e-08 $layer=LI1_cond $X=1.61 $Y=2.535
+ $X2=1.525 $Y2=2.535
r56 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r57 30 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=2.72
+ $X2=0.23 $Y2=2.72
r58 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 26 39 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.07 $Y2=2.72
r60 25 40 89.0535 $w=1.68e-07 $l=1.365e-06 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.085 $Y2=2.72
r61 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r62 22 33 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 22 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r64 21 34 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=1.525 $Y2=2.72
r65 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r66 19 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=0.715 $Y2=2.72
r67 19 21 15.984 $w=1.68e-07 $l=2.45e-07 $layer=LI1_cond $X=0.905 $Y=2.72
+ $X2=1.15 $Y2=2.72
r68 15 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r69 13 29 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.715 $Y2=2.72
r70 13 15 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r71 11 44 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=2.72
+ $X2=0.23 $Y2=2.72
r72 7 29 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2.72
r73 7 9 19.2579 $w=3.78e-07 $l=6.35e-07 $layer=LI1_cond $X=0.715 $Y=2.635
+ $X2=0.715 $Y2=2
r74 2 36 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.59
+ $Y=1.485 $X2=1.74 $Y2=2.36
r75 1 9 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=0.59
+ $Y=1.485 $X2=0.74 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%A_227_297# 1 2 7 9 11 13 15
r28 13 20 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=2.435 $Y=2.095
+ $X2=2.435 $Y2=1.98
r29 13 15 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=2.435 $Y=2.095
+ $X2=2.435 $Y2=2.29
r30 12 18 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=1.355 $Y=1.98
+ $X2=1.225 $Y2=1.98
r31 11 20 3.63458 $w=2.3e-07 $l=1.3e-07 $layer=LI1_cond $X=2.305 $Y=1.98
+ $X2=2.435 $Y2=1.98
r32 11 12 47.6009 $w=2.28e-07 $l=9.5e-07 $layer=LI1_cond $X=2.305 $Y=1.98
+ $X2=1.355 $Y2=1.98
r33 7 18 3.2152 $w=2.6e-07 $l=1.15e-07 $layer=LI1_cond $X=1.225 $Y=2.095
+ $X2=1.225 $Y2=1.98
r34 7 9 8.64332 $w=2.58e-07 $l=1.95e-07 $layer=LI1_cond $X=1.225 $Y=2.095
+ $X2=1.225 $Y2=2.29
r35 2 20 600 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.485 $X2=2.4 $Y2=1.95
r36 2 15 600 $w=1.7e-07 $l=8.76798e-07 $layer=licon1_PDIFF $count=1 $X=2.25
+ $Y=1.485 $X2=2.4 $Y2=2.29
r37 1 18 600 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.26 $Y2=1.95
r38 1 9 600 $w=1.7e-07 $l=8.65246e-07 $layer=licon1_PDIFF $count=1 $X=1.135
+ $Y=1.485 $X2=1.26 $Y2=2.29
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211O_1%VGND 1 2 9 11 21 22 25 33 36 44
r47 36 39 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=2.89 $Y=0 $X2=2.89
+ $Y2=0.36
r48 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r49 32 33 10.9862 $w=5.38e-07 $l=2.2e-07 $layer=LI1_cond $X=1.18 $Y=0.185
+ $X2=1.4 $Y2=0.185
r50 29 32 0.664488 $w=5.38e-07 $l=3e-08 $layer=LI1_cond $X=1.15 $Y=0.185
+ $X2=1.18 $Y2=0.185
r51 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r52 26 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r53 26 44 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r54 25 29 10.1888 $w=5.38e-07 $l=4.6e-07 $layer=LI1_cond $X=0.69 $Y=0.185
+ $X2=1.15 $Y2=0.185
r55 25 26 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r56 22 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.99
+ $Y2=0
r57 21 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r58 19 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=2.89
+ $Y2=0
r59 19 21 24.139 $w=1.68e-07 $l=3.7e-07 $layer=LI1_cond $X=3.08 $Y=0 $X2=3.45
+ $Y2=0
r60 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r61 17 18 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r62 15 18 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r63 15 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r64 14 17 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r65 14 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=1.4
+ $Y2=0
r66 14 15 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r67 11 36 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.89
+ $Y2=0
r68 11 17 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=2.7 $Y=0 $X2=2.53
+ $Y2=0
r69 9 44 0.00284542 $w=4.8e-07 $l=1e-08 $layer=MET1_cond $X=0.22 $Y=0 $X2=0.23
+ $Y2=0
r70 2 39 182 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_NDIFF $count=1 $X=2.69
+ $Y=0.235 $X2=2.915 $Y2=0.36
r71 1 32 91 $w=1.7e-07 $l=6.89674e-07 $layer=licon1_NDIFF $count=2 $X=0.55
+ $Y=0.235 $X2=1.18 $Y2=0.36
.ends

