* File: sky130_fd_sc_hdll__mux2_2.spice
* Created: Thu Aug 27 19:10:41 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__mux2_2.pex.spice"
.subckt sky130_fd_sc_hdll__mux2_2  VNB VPB A0 A1 S VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* S	S
* A1	A1
* A0	A0
* VPB	VPB
* VNB	VNB
MM1006 N_VGND_M1006_d N_A_79_21#_M1006_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.104 PD=1.82 PS=0.97 NRD=0 NRS=5.532 M=1 R=4.33333 SA=75000.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1012 N_VGND_M1012_d N_A_79_21#_M1012_g N_X_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.140145 AS=0.104 PD=1.25748 PS=0.97 NRD=8.304 NRS=1.836 M=1 R=4.33333
+ SA=75000.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1011 A_310_47# N_A_280_21#_M1011_g N_VGND_M1012_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0905551 PD=0.75 PS=0.812523 NRD=31.428 NRS=17.136 M=1 R=2.8
+ SA=75001.2 SB=75002.6 A=0.063 P=1.14 MULT=1
MM1004 N_A_79_21#_M1004_d N_A0_M1004_g A_310_47# VNB NSHORT L=0.15 W=0.42
+ AD=0.0693 AS=0.0693 PD=0.75 PS=0.75 NRD=0 NRS=31.428 M=1 R=2.8 SA=75001.7
+ SB=75002.1 A=0.063 P=1.14 MULT=1
MM1007 A_502_47# N_A1_M1007_g N_A_79_21#_M1004_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1554 AS=0.0693 PD=1.16 PS=0.75 NRD=90 NRS=15.708 M=1 R=2.8 SA=75002.1
+ SB=75001.6 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_S_M1005_g A_502_47# VNB NSHORT L=0.15 W=0.42 AD=0.0777
+ AS=0.1554 PD=0.79 PS=1.16 NRD=12.852 NRS=90 M=1 R=2.8 SA=75003 SB=75000.7
+ A=0.063 P=1.14 MULT=1
MM1013 N_A_280_21#_M1013_d N_S_M1013_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1155 AS=0.0777 PD=1.39 PS=0.79 NRD=2.856 NRS=12.852 M=1 R=2.8 SA=75003.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_79_21#_M1000_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.5 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1009_d N_A_79_21#_M1009_g N_X_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.19561 AS=0.145 PD=1.65244 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90002 A=0.18 P=2.36 MULT=1
MM1008 A_318_369# N_A_280_21#_M1008_g N_VPWR_M1009_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.2496 AS=0.12519 PD=1.42 PS=1.05756 NRD=103.11 NRS=21.5321 M=1 R=3.55556
+ SA=90001.2 SB=90002.5 A=0.1152 P=1.64 MULT=1
MM1010 N_A_79_21#_M1010_d N_A1_M1010_g A_318_369# VPB PHIGHVT L=0.18 W=0.64
+ AD=0.096 AS=0.2496 PD=0.94 PS=1.42 NRD=1.5366 NRS=103.11 M=1 R=3.55556
+ SA=90002.1 SB=90001.5 A=0.1152 P=1.64 MULT=1
MM1002 A_606_369# N_A0_M1002_g N_A_79_21#_M1010_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.0736 AS=0.096 PD=0.87 PS=0.94 NRD=18.4589 NRS=4.6098 M=1 R=3.55556
+ SA=90002.6 SB=90001.1 A=0.1152 P=1.64 MULT=1
MM1003 N_VPWR_M1003_d N_S_M1003_g A_606_369# VPB PHIGHVT L=0.18 W=0.64 AD=0.0928
+ AS=0.0736 PD=0.93 PS=0.87 NRD=1.5366 NRS=18.4589 M=1 R=3.55556 SA=90003
+ SB=90000.7 A=0.1152 P=1.64 MULT=1
MM1001 N_A_280_21#_M1001_d N_S_M1001_g N_VPWR_M1003_d VPB PHIGHVT L=0.18 W=0.64
+ AD=0.1792 AS=0.0928 PD=1.84 PS=0.93 NRD=4.6098 NRS=1.5366 M=1 R=3.55556
+ SA=90003.5 SB=90000.2 A=0.1152 P=1.64 MULT=1
DX14_noxref VNB VPB NWDIODE A=7.9929 P=13.17
c_76 VPB 0 1.25191e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__mux2_2.pxi.spice"
*
.ends
*
*
