* File: sky130_fd_sc_hdll__or2_1.pex.spice
* Created: Thu Aug 27 19:23:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__OR2_1%B 3 5 7 8 9 15
r26 15 16 10.0139 $w=3.61e-07 $l=7.5e-08 $layer=POLY_cond $X=0.475 $Y=1.202
+ $X2=0.55 $Y2=1.202
r27 13 15 28.0388 $w=3.61e-07 $l=2.1e-07 $layer=POLY_cond $X=0.265 $Y=1.202
+ $X2=0.475 $Y2=1.202
r28 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.265
+ $Y=1.16 $X2=0.265 $Y2=1.16
r29 8 9 10.0636 $w=3.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.262 $Y=0.85
+ $X2=0.262 $Y2=1.16
r30 5 16 19.0337 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.55 $Y=1.41
+ $X2=0.55 $Y2=1.202
r31 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.55 $Y=1.41 $X2=0.55
+ $Y2=1.695
r32 1 15 23.3725 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r33 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_1%A 3 5 7 8 9
r33 9 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.035
+ $Y=1.16 $X2=1.035 $Y2=1.16
r34 8 9 10.6644 $w=3.33e-07 $l=3.1e-07 $layer=LI1_cond $X=1.117 $Y=0.85
+ $X2=1.117 $Y2=1.16
r35 5 13 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=0.96 $Y=1.41
+ $X2=1.02 $Y2=1.16
r36 5 7 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.96 $Y=1.41 $X2=0.96
+ $Y2=1.695
r37 1 13 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=0.935 $Y=0.995
+ $X2=1.02 $Y2=1.16
r38 1 3 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.935 $Y=0.995
+ $X2=0.935 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_1%A_38_297# 1 2 7 9 10 12 14 15 16 19 26
c50 19 0 9.66706e-20 $X=1.61 $Y=1.16
c51 14 0 9.99956e-20 $X=0.695 $Y=1.495
r52 26 28 8.91885 $w=2.38e-07 $l=1.65e-07 $layer=LI1_cond $X=0.73 $Y=0.43
+ $X2=0.73 $Y2=0.595
r53 19 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.61
+ $Y=1.16 $X2=1.61 $Y2=1.16
r54 17 19 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.635 $Y=1.495
+ $X2=1.635 $Y2=1.16
r55 15 17 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=1.635 $Y2=1.495
r56 15 16 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=1.525 $Y=1.58
+ $X2=0.78 $Y2=1.58
r57 14 16 5.5252 $w=2.73e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.695 $Y=1.495
+ $X2=0.78 $Y2=1.58
r58 14 23 16.9817 $w=2.73e-07 $l=4.57996e-07 $layer=LI1_cond $X=0.695 $Y=1.495
+ $X2=0.315 $Y2=1.667
r59 14 28 58.7166 $w=1.68e-07 $l=9e-07 $layer=LI1_cond $X=0.695 $Y=1.495
+ $X2=0.695 $Y2=0.595
r60 10 20 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.61 $Y2=1.16
r61 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.495 $Y=1.41
+ $X2=1.495 $Y2=1.985
r62 7 20 39.2524 $w=3.82e-07 $l=2.24332e-07 $layer=POLY_cond $X=1.47 $Y=0.995
+ $X2=1.61 $Y2=1.16
r63 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.47 $Y=0.995 $X2=1.47
+ $Y2=0.56
r64 2 23 600 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.19
+ $Y=1.485 $X2=0.315 $Y2=1.66
r65 1 26 182 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.725 $Y2=0.43
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_1%VPWR 1 6 8 10 17 18 21
r21 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r22 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r23 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r24 15 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=1.26 $Y2=2.72
r25 15 17 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=1.425 $Y=2.72
+ $X2=2.07 $Y2=2.72
r26 10 21 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=1.26 $Y2=2.72
r27 10 12 56.4332 $w=1.68e-07 $l=8.65e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.23 $Y2=2.72
r28 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r29 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r30 4 21 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.26 $Y=2.635 $X2=1.26
+ $Y2=2.72
r31 4 6 24.9696 $w=3.28e-07 $l=7.15e-07 $layer=LI1_cond $X=1.26 $Y=2.635
+ $X2=1.26 $Y2=1.92
r32 1 6 300 $w=1.7e-07 $l=5.29693e-07 $layer=licon1_PDIFF $count=2 $X=1.05
+ $Y=1.485 $X2=1.26 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_1%X 1 2 10 13 19
c26 2 0 9.66706e-20 $X=1.585 $Y=1.485
r27 19 20 3.19486 $w=5.68e-07 $l=2.5e-08 $layer=LI1_cond $X=1.93 $Y=1.87
+ $X2=1.93 $Y2=1.845
r28 13 24 2.09838 $w=5.68e-07 $l=1e-07 $layer=LI1_cond $X=1.93 $Y=1.9 $X2=1.93
+ $Y2=2
r29 13 19 0.629515 $w=5.68e-07 $l=3e-08 $layer=LI1_cond $X=1.93 $Y=1.9 $X2=1.93
+ $Y2=1.87
r30 13 20 1.15244 $w=2.98e-07 $l=3e-08 $layer=LI1_cond $X=2.065 $Y=1.815
+ $X2=2.065 $Y2=1.845
r31 11 13 38.0306 $w=2.98e-07 $l=9.9e-07 $layer=LI1_cond $X=2.065 $Y=0.825
+ $X2=2.065 $Y2=1.815
r32 10 11 4.4967 $w=3e-07 $l=2.85e-07 $layer=LI1_cond $X=2.065 $Y=0.54 $X2=2.065
+ $Y2=0.825
r33 8 10 7.02958 $w=5.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.73 $Y=0.54
+ $X2=2.065 $Y2=0.54
r34 2 24 300 $w=1.7e-07 $l=6.17333e-07 $layer=licon1_PDIFF $count=2 $X=1.585
+ $Y=1.485 $X2=1.81 $Y2=2
r35 1 8 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=1.545
+ $Y=0.235 $X2=1.73 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__OR2_1%VGND 1 2 7 9 11 15 17 21 22 28
r30 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r31 22 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r32 21 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r33 19 28 6.25164 $w=1.7e-07 $l=1.08e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=1.237
+ $Y2=0
r34 19 21 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.345 $Y=0 $X2=2.07
+ $Y2=0
r35 17 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r36 17 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r37 13 28 0.512231 $w=2.15e-07 $l=8.5e-08 $layer=LI1_cond $X=1.237 $Y=0.085
+ $X2=1.237 $Y2=0
r38 13 15 18.4927 $w=2.13e-07 $l=3.45e-07 $layer=LI1_cond $X=1.237 $Y=0.085
+ $X2=1.237 $Y2=0.43
r39 12 25 3.9323 $w=1.7e-07 $l=1.75e-07 $layer=LI1_cond $X=0.35 $Y=0 $X2=0.175
+ $Y2=0
r40 11 28 6.25164 $w=1.7e-07 $l=1.07e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=1.237
+ $Y2=0
r41 11 12 50.8877 $w=1.68e-07 $l=7.8e-07 $layer=LI1_cond $X=1.13 $Y=0 $X2=0.35
+ $Y2=0
r42 7 25 3.14584 $w=2.4e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.175 $Y2=0
r43 7 9 16.5664 $w=2.38e-07 $l=3.45e-07 $layer=LI1_cond $X=0.23 $Y=0.085
+ $X2=0.23 $Y2=0.43
r44 2 15 182 $w=1.7e-07 $l=3.28329e-07 $layer=licon1_NDIFF $count=1 $X=1.01
+ $Y=0.235 $X2=1.255 $Y2=0.43
r45 1 9 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.14
+ $Y=0.235 $X2=0.265 $Y2=0.43
.ends

