* File: sky130_fd_sc_hdll__a21boi_1.pex.spice
* Created: Thu Aug 27 18:52:23 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%B1_N 1 2 3 5 6 8 11 13 14 18
r36 13 14 18.5393 $w=2.28e-07 $l=3.7e-07 $layer=LI1_cond $X=0.22 $Y=1.16
+ $X2=0.22 $Y2=1.53
r37 13 18 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r38 11 18 145.524 $w=2.7e-07 $l=6.55e-07 $layer=POLY_cond $X=0.24 $Y=1.815
+ $X2=0.24 $Y2=1.16
r39 9 18 56.6543 $w=2.7e-07 $l=2.55e-07 $layer=POLY_cond $X=0.24 $Y=0.905
+ $X2=0.24 $Y2=1.16
r40 6 8 99.6133 $w=1.5e-07 $l=3.1e-07 $layer=POLY_cond $X=0.865 $Y=0.755
+ $X2=0.865 $Y2=0.445
r41 3 11 78.325 $w=1.6e-07 $l=2.6e-07 $layer=POLY_cond $X=0.5 $Y=1.902 $X2=0.24
+ $Y2=1.902
r42 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.5 $Y=1.99 $X2=0.5
+ $Y2=2.275
r43 2 9 29.8935 $w=1.5e-07 $l=1.68375e-07 $layer=POLY_cond $X=0.375 $Y=0.83
+ $X2=0.24 $Y2=0.905
r44 1 6 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=0.79 $Y=0.83
+ $X2=0.865 $Y2=0.755
r45 1 2 212.798 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=0.79 $Y=0.83
+ $X2=0.375 $Y2=0.83
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%A_27_413# 1 2 7 11 13 15 16 20 23 25 32
+ 35
c66 16 0 1.57556e-19 $X=1.405 $Y=1.297
r67 32 34 7.60109 $w=4.88e-07 $l=2.65e-07 $layer=LI1_cond $X=0.61 $Y=0.45
+ $X2=0.61 $Y2=0.715
r68 26 35 27.9505 $w=3.2e-07 $l=1.55e-07 $layer=POLY_cond $X=0.795 $Y=1.44
+ $X2=0.795 $Y2=1.285
r69 25 34 24.5742 $w=3.38e-07 $l=7.25e-07 $layer=LI1_cond $X=0.685 $Y=1.44
+ $X2=0.685 $Y2=0.715
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.77
+ $Y=1.44 $X2=0.77 $Y2=1.44
r71 23 25 13.3887 $w=3.38e-07 $l=3.95e-07 $layer=LI1_cond $X=0.685 $Y=1.835
+ $X2=0.685 $Y2=1.44
r72 18 23 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=0.225 $Y=1.92
+ $X2=0.685 $Y2=1.92
r73 18 20 11.7461 $w=2.58e-07 $l=2.65e-07 $layer=LI1_cond $X=0.225 $Y=2.005
+ $X2=0.225 $Y2=2.27
r74 16 17 44.1268 $w=2.13e-07 $l=1.95e-07 $layer=POLY_cond $X=1.405 $Y=1.297
+ $X2=1.6 $Y2=1.297
r75 13 17 6.81225 $w=1.8e-07 $l=1.13e-07 $layer=POLY_cond $X=1.6 $Y=1.41 $X2=1.6
+ $Y2=1.297
r76 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.6 $Y=1.41 $X2=1.6
+ $Y2=1.985
r77 9 16 11.0275 $w=1.5e-07 $l=1.12e-07 $layer=POLY_cond $X=1.405 $Y=1.185
+ $X2=1.405 $Y2=1.297
r78 9 11 320.479 $w=1.5e-07 $l=6.25e-07 $layer=POLY_cond $X=1.405 $Y=1.185
+ $X2=1.405 $Y2=0.56
r79 8 35 13.7767 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=0.955 $Y=1.285
+ $X2=0.795 $Y2=1.285
r80 7 16 17.2128 $w=2.13e-07 $l=8.07775e-08 $layer=POLY_cond $X=1.33 $Y=1.285
+ $X2=1.405 $Y2=1.297
r81 7 8 124.341 $w=2e-07 $l=3.75e-07 $layer=POLY_cond $X=1.33 $Y=1.285 $X2=0.955
+ $Y2=1.285
r82 2 20 600 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.27
r83 1 32 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=0.425
+ $Y=0.235 $X2=0.55 $Y2=0.45
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%A1 1 3 4 6 7 8 9
c35 7 0 1.57556e-19 $X=2.07 $Y=0.51
r36 9 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.07
+ $Y=1.16 $X2=2.07 $Y2=1.16
r37 8 9 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=2.112 $Y=0.85
+ $X2=2.112 $Y2=1.16
r38 7 8 15.3659 $w=2.53e-07 $l=3.4e-07 $layer=LI1_cond $X=2.112 $Y=0.51
+ $X2=2.112 $Y2=0.85
r39 4 14 38.578 $w=2.95e-07 $l=1.72337e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.08 $Y2=1.16
r40 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.095 $Y=0.995
+ $X2=2.095 $Y2=0.56
r41 1 14 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=2.08 $Y=1.41
+ $X2=2.08 $Y2=1.16
r42 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.08 $Y=1.41 $X2=2.08
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%A2 1 3 4 6 7 14
r22 10 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.905
+ $Y=1.16 $X2=2.905 $Y2=1.16
r23 7 14 1.48171 $w=3.48e-07 $l=4.5e-08 $layer=LI1_cond $X=2.95 $Y=1.17
+ $X2=2.905 $Y2=1.17
r24 4 10 44.8379 $w=4.06e-07 $l=3.08221e-07 $layer=POLY_cond $X=2.68 $Y=1.41
+ $X2=2.81 $Y2=1.16
r25 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.68 $Y=1.41 $X2=2.68
+ $Y2=1.985
r26 1 10 39.7049 $w=4.06e-07 $l=2.29783e-07 $layer=POLY_cond $X=2.655 $Y=0.995
+ $X2=2.81 $Y2=1.16
r27 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.655 $Y=0.995
+ $X2=2.655 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%VPWR 1 2 9 13 16 17 18 20 33 34 37
r43 37 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r44 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r45 31 34 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r46 30 31 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r47 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r48 28 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r49 27 30 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 27 28 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r51 25 37 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.71 $Y2=2.72
r52 25 27 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r53 20 37 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.71 $Y2=2.72
r54 20 22 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.525 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 18 38 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r56 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r57 16 30 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 16 17 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.295 $Y2=2.72
r59 15 33 32.9465 $w=1.68e-07 $l=5.05e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.99 $Y2=2.72
r60 15 17 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.485 $Y=2.72
+ $X2=2.295 $Y2=2.72
r61 11 17 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.295 $Y=2.635
+ $X2=2.295 $Y2=2.72
r62 11 13 18.6514 $w=3.78e-07 $l=6.15e-07 $layer=LI1_cond $X=2.295 $Y=2.635
+ $X2=2.295 $Y2=2.02
r63 7 37 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.71 $Y=2.635 $X2=0.71
+ $Y2=2.72
r64 7 9 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.71 $Y=2.635 $X2=0.71
+ $Y2=2.34
r65 2 13 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=2.17
+ $Y=1.485 $X2=2.32 $Y2=2.02
r66 1 9 600 $w=1.7e-07 $l=3.4187e-07 $layer=licon1_PDIFF $count=1 $X=0.59
+ $Y=2.065 $X2=0.74 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%Y 1 2 7 8 9 10 11 29 37
r36 17 29 12.1007 $w=2.98e-07 $l=3.15e-07 $layer=LI1_cond $X=1.295 $Y=1.195
+ $X2=1.61 $Y2=1.195
r37 17 37 4.03355 $w=2.98e-07 $l=1.05e-07 $layer=LI1_cond $X=1.295 $Y=1.195
+ $X2=1.19 $Y2=1.195
r38 11 29 18.134 $w=3.38e-07 $l=5.35e-07 $layer=LI1_cond $X=1.61 $Y=0.51
+ $X2=1.61 $Y2=1.045
r39 10 21 6.24041 $w=4.58e-07 $l=2.4e-07 $layer=LI1_cond $X=1.295 $Y=1.87
+ $X2=1.295 $Y2=1.63
r40 9 21 2.60017 $w=4.58e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=1.53 $X2=1.295
+ $Y2=1.63
r41 9 17 4.81032 $w=4.58e-07 $l=1.85e-07 $layer=LI1_cond $X=1.295 $Y=1.53
+ $X2=1.295 $Y2=1.345
r42 8 27 2.60017 $w=4.58e-07 $l=1e-07 $layer=LI1_cond $X=1.295 $Y=2.21 $X2=1.295
+ $Y2=2.31
r43 8 10 8.84058 $w=4.58e-07 $l=3.4e-07 $layer=LI1_cond $X=1.295 $Y=2.21
+ $X2=1.295 $Y2=1.87
r44 7 37 0.576222 $w=2.98e-07 $l=1.5e-08 $layer=LI1_cond $X=1.175 $Y=1.195
+ $X2=1.19 $Y2=1.195
r45 2 27 400 $w=1.7e-07 $l=8.85297e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.485 $X2=1.31 $Y2=2.31
r46 2 21 400 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.185
+ $Y=1.485 $X2=1.31 $Y2=1.63
r47 1 11 182 $w=1.7e-07 $l=4.09115e-07 $layer=licon1_NDIFF $count=1 $X=1.48
+ $Y=0.235 $X2=1.67 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%A_338_297# 1 2 9 11 12 15
r16 13 15 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=2.92 $Y=1.725
+ $X2=2.92 $Y2=1.95
r17 11 13 6.87494 $w=2e-07 $l=1.36015e-07 $layer=LI1_cond $X=2.835 $Y=1.625
+ $X2=2.92 $Y2=1.725
r18 11 12 49.9091 $w=1.98e-07 $l=9e-07 $layer=LI1_cond $X=2.835 $Y=1.625
+ $X2=1.935 $Y2=1.625
r19 7 12 6.82232 $w=2e-07 $l=1.39642e-07 $layer=LI1_cond $X=1.84 $Y=1.725
+ $X2=1.935 $Y2=1.625
r20 7 9 13.134 $w=1.88e-07 $l=2.25e-07 $layer=LI1_cond $X=1.84 $Y=1.725 $X2=1.84
+ $Y2=1.95
r21 2 15 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=2.77
+ $Y=1.485 $X2=2.92 $Y2=1.95
r22 1 9 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.69
+ $Y=1.485 $X2=1.84 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BOI_1%VGND 1 2 9 11 13 15 17 22 31 35
r38 34 35 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r39 31 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r40 29 35 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.99
+ $Y2=0
r41 28 29 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r42 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r43 26 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=1.15
+ $Y2=0
r44 25 28 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r45 25 26 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r46 23 31 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.14
+ $Y2=0
r47 23 25 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=1.255 $Y=0 $X2=1.61
+ $Y2=0
r48 22 34 4.94333 $w=1.7e-07 $l=2.52e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.967
+ $Y2=0
r49 22 28 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.715 $Y=0 $X2=2.53
+ $Y2=0
r50 20 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r51 19 20 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r52 17 31 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=1.14
+ $Y2=0
r53 17 19 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.025 $Y=0 $X2=0.69
+ $Y2=0
r54 15 20 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r55 11 34 3.07978 $w=3.6e-07 $l=1.15521e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.967 $Y2=0
r56 11 13 9.44363 $w=3.58e-07 $l=2.95e-07 $layer=LI1_cond $X=2.895 $Y=0.085
+ $X2=2.895 $Y2=0.38
r57 7 31 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0
r58 7 9 13.7792 $w=2.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.14 $Y=0.085
+ $X2=1.14 $Y2=0.36
r59 2 13 91 $w=1.7e-07 $l=2.41868e-07 $layer=licon1_NDIFF $count=2 $X=2.73
+ $Y=0.235 $X2=2.91 $Y2=0.38
r60 1 9 91 $w=1.7e-07 $l=2.54951e-07 $layer=licon1_NDIFF $count=2 $X=0.94
+ $Y=0.235 $X2=1.14 $Y2=0.36
.ends

