* File: sky130_fd_sc_hdll__o21ba_4.pxi.spice
* Created: Wed Sep  2 08:44:00 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21BA_4%B1_N N_B1_N_c_103_n N_B1_N_M1004_g
+ N_B1_N_c_104_n N_B1_N_M1017_g B1_N B1_N N_B1_N_c_106_n
+ PM_SKY130_FD_SC_HDLL__O21BA_4%B1_N
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A_197_21# N_A_197_21#_M1003_s
+ N_A_197_21#_M1016_s N_A_197_21#_M1001_s N_A_197_21#_c_139_n
+ N_A_197_21#_M1007_g N_A_197_21#_c_148_n N_A_197_21#_M1000_g
+ N_A_197_21#_c_140_n N_A_197_21#_M1009_g N_A_197_21#_c_149_n
+ N_A_197_21#_M1006_g N_A_197_21#_c_141_n N_A_197_21#_M1013_g
+ N_A_197_21#_c_150_n N_A_197_21#_M1010_g N_A_197_21#_c_151_n
+ N_A_197_21#_M1014_g N_A_197_21#_c_142_n N_A_197_21#_M1021_g
+ N_A_197_21#_c_143_n N_A_197_21#_c_144_n N_A_197_21#_c_145_n
+ N_A_197_21#_c_256_p N_A_197_21#_c_164_p N_A_197_21#_c_169_p
+ N_A_197_21#_c_146_n N_A_197_21#_c_153_n N_A_197_21#_c_270_p
+ N_A_197_21#_c_154_n N_A_197_21#_c_176_p N_A_197_21#_c_155_n
+ N_A_197_21#_c_147_n PM_SKY130_FD_SC_HDLL__O21BA_4%A_197_21#
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A_27_297# N_A_27_297#_M1017_s
+ N_A_27_297#_M1004_s N_A_27_297#_c_306_n N_A_27_297#_M1016_g
+ N_A_27_297#_c_307_n N_A_27_297#_M1020_g N_A_27_297#_c_301_n
+ N_A_27_297#_M1003_g N_A_27_297#_c_302_n N_A_27_297#_M1011_g
+ N_A_27_297#_c_308_n N_A_27_297#_c_309_n N_A_27_297#_c_315_n
+ N_A_27_297#_c_342_n N_A_27_297#_c_310_n N_A_27_297#_c_303_n
+ N_A_27_297#_c_311_n N_A_27_297#_c_304_n N_A_27_297#_c_313_n
+ N_A_27_297#_c_351_n N_A_27_297#_c_305_n
+ PM_SKY130_FD_SC_HDLL__O21BA_4%A_27_297#
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A2 N_A2_c_409_n N_A2_M1002_g N_A2_c_413_n
+ N_A2_M1001_g N_A2_c_414_n N_A2_M1008_g N_A2_c_410_n N_A2_M1019_g A2
+ N_A2_c_412_n A2 PM_SKY130_FD_SC_HDLL__O21BA_4%A2
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A1 N_A1_c_463_n N_A1_M1005_g N_A1_c_467_n
+ N_A1_M1015_g N_A1_c_468_n N_A1_M1018_g N_A1_c_464_n N_A1_M1012_g A1
+ N_A1_c_466_n A1 PM_SKY130_FD_SC_HDLL__O21BA_4%A1
x_PM_SKY130_FD_SC_HDLL__O21BA_4%VPWR N_VPWR_M1004_d N_VPWR_M1006_d
+ N_VPWR_M1014_d N_VPWR_M1020_d N_VPWR_M1015_s N_VPWR_c_502_n N_VPWR_c_503_n
+ N_VPWR_c_504_n N_VPWR_c_505_n N_VPWR_c_506_n N_VPWR_c_507_n N_VPWR_c_508_n
+ N_VPWR_c_509_n N_VPWR_c_510_n N_VPWR_c_511_n N_VPWR_c_512_n VPWR
+ N_VPWR_c_513_n N_VPWR_c_501_n N_VPWR_c_515_n N_VPWR_c_516_n N_VPWR_c_517_n
+ PM_SKY130_FD_SC_HDLL__O21BA_4%VPWR
x_PM_SKY130_FD_SC_HDLL__O21BA_4%X N_X_M1007_d N_X_M1013_d N_X_M1000_s
+ N_X_M1010_s N_X_c_616_n N_X_c_609_n N_X_c_610_n N_X_c_612_n N_X_c_636_n X
+ N_X_c_638_n PM_SKY130_FD_SC_HDLL__O21BA_4%X
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A_823_297# N_A_823_297#_M1001_d
+ N_A_823_297#_M1008_d N_A_823_297#_M1018_d N_A_823_297#_c_672_n
+ N_A_823_297#_c_666_n N_A_823_297#_c_692_n N_A_823_297#_c_667_n
+ N_A_823_297#_c_668_n N_A_823_297#_c_669_n N_A_823_297#_c_670_n
+ PM_SKY130_FD_SC_HDLL__O21BA_4%A_823_297#
x_PM_SKY130_FD_SC_HDLL__O21BA_4%VGND N_VGND_M1017_d N_VGND_M1009_s
+ N_VGND_M1021_s N_VGND_M1002_d N_VGND_M1005_s N_VGND_c_705_n N_VGND_c_706_n
+ N_VGND_c_707_n N_VGND_c_708_n N_VGND_c_709_n N_VGND_c_710_n N_VGND_c_711_n
+ N_VGND_c_712_n N_VGND_c_713_n N_VGND_c_714_n N_VGND_c_715_n N_VGND_c_716_n
+ N_VGND_c_717_n N_VGND_c_718_n N_VGND_c_719_n VGND N_VGND_c_720_n
+ N_VGND_c_721_n PM_SKY130_FD_SC_HDLL__O21BA_4%VGND
x_PM_SKY130_FD_SC_HDLL__O21BA_4%A_635_47# N_A_635_47#_M1003_d
+ N_A_635_47#_M1011_d N_A_635_47#_M1019_s N_A_635_47#_M1012_d
+ N_A_635_47#_c_813_n N_A_635_47#_c_829_n N_A_635_47#_c_814_n
+ N_A_635_47#_c_815_n N_A_635_47#_c_837_n N_A_635_47#_c_816_n
+ N_A_635_47#_c_817_n N_A_635_47#_c_818_n
+ PM_SKY130_FD_SC_HDLL__O21BA_4%A_635_47#
cc_1 VNB N_B1_N_c_103_n 0.0287789f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.41
cc_2 VNB N_B1_N_c_104_n 0.0202057f $X=-0.19 $Y=-0.24 $X2=0.64 $Y2=0.995
cc_3 VNB B1_N 5.80836e-19 $X=-0.19 $Y=-0.24 $X2=0.605 $Y2=1.445
cc_4 VNB N_B1_N_c_106_n 0.00589029f $X=-0.19 $Y=-0.24 $X2=0.77 $Y2=1.285
cc_5 VNB N_A_197_21#_c_139_n 0.0166801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_197_21#_c_140_n 0.015981f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_197_21#_c_141_n 0.0171139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_197_21#_c_142_n 0.0191851f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_197_21#_c_143_n 0.00441285f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_197_21#_c_144_n 0.00402473f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_197_21#_c_145_n 0.0150708f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_197_21#_c_146_n 9.56934e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_197_21#_c_147_n 0.0747037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_297#_c_301_n 0.0204671f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_15 VNB N_A_27_297#_c_302_n 0.01669f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_297#_c_303_n 0.0265255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_297#_c_304_n 0.021664f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_297#_c_305_n 0.0692454f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A2_c_409_n 0.0173809f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.41
cc_20 VNB N_A2_c_410_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB A2 0.0124374f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_22 VNB N_A2_c_412_n 0.0365641f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A1_c_463_n 0.0169324f $X=-0.19 $Y=-0.24 $X2=0.615 $Y2=1.41
cc_24 VNB N_A1_c_464_n 0.0223965f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB A1 0.0186454f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_26 VNB N_A1_c_466_n 0.0430121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VPWR_c_501_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_609_n 0.00184153f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_610_n 0.00437891f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.18
cc_30 VNB N_VGND_c_705_n 0.00662136f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_706_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_707_n 0.00548869f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_708_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_709_n 0.00469739f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_710_n 0.0222618f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_711_n 0.00326991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_VGND_c_712_n 0.0203968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_713_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_VGND_c_714_n 0.0169949f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_715_n 0.00507229f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_716_n 0.0406466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_717_n 0.00323964f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_718_n 0.0191746f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_719_n 0.00324297f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_720_n 0.0202195f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_721_n 0.319382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_635_47#_c_813_n 0.00329212f $X=-0.19 $Y=-0.24 $X2=0.59 $Y2=1.16
cc_48 VNB N_A_635_47#_c_814_n 0.00299515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_635_47#_c_815_n 0.00276474f $X=-0.19 $Y=-0.24 $X2=0.69 $Y2=1.18
cc_50 VNB N_A_635_47#_c_816_n 0.0139603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_635_47#_c_817_n 0.0186133f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_635_47#_c_818_n 0.00253348f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VPB N_B1_N_c_103_n 0.0302064f $X=-0.19 $Y=1.305 $X2=0.615 $Y2=1.41
cc_54 VPB B1_N 0.00114226f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.445
cc_55 VPB N_A_197_21#_c_148_n 0.0158645f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_56 VPB N_A_197_21#_c_149_n 0.0151206f $X=-0.19 $Y=1.305 $X2=0.69 $Y2=1.18
cc_57 VPB N_A_197_21#_c_150_n 0.0156949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A_197_21#_c_151_n 0.0157354f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A_197_21#_c_146_n 0.00810112f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_A_197_21#_c_153_n 0.00681108f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_197_21#_c_154_n 0.0023495f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_197_21#_c_155_n 0.0029376f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_197_21#_c_147_n 0.045398f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_297#_c_306_n 0.0156315f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_65 VPB N_A_27_297#_c_307_n 0.0192331f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_297#_c_308_n 0.00956215f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_297#_c_309_n 0.0168446f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_297#_c_310_n 0.00495343f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_297#_c_311_n 0.00982421f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_A_27_297#_c_304_n 0.00715877f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_A_27_297#_c_313_n 0.00723806f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_A_27_297#_c_305_n 0.0380017f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_A2_c_413_n 0.0195777f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.995
cc_74 VPB N_A2_c_414_n 0.01642f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_75 VPB N_A2_c_412_n 0.0214781f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB N_A1_c_467_n 0.0156552f $X=-0.19 $Y=1.305 $X2=0.64 $Y2=0.995
cc_77 VPB N_A1_c_468_n 0.0201729f $X=-0.19 $Y=1.305 $X2=0.605 $Y2=1.105
cc_78 VPB N_A1_c_466_n 0.022695f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_502_n 4.04661e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_503_n 0.0133737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_504_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_505_n 0.0133737f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_506_n 3.34338e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_507_n 0.0077211f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_508_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_509_n 0.0172166f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_510_n 0.00478242f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_511_n 0.0382464f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_512_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_VPWR_c_513_n 0.0184169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_501_n 0.0497732f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_92 VPB N_VPWR_c_515_n 0.0222293f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_516_n 0.00502902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_VPWR_c_517_n 0.00502902f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_X_c_609_n 0.00137164f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_X_c_612_n 0.00347993f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_A_823_297#_c_666_n 0.00188899f $X=-0.19 $Y=1.305 $X2=0.59 $Y2=1.16
cc_98 VPB N_A_823_297#_c_667_n 0.00290609f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.285
cc_99 VPB N_A_823_297#_c_668_n 0.0116576f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_A_823_297#_c_669_n 0.0307403f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_A_823_297#_c_670_n 0.00493435f $X=-0.19 $Y=1.305 $X2=0.77 $Y2=1.18
cc_102 N_B1_N_c_104_n N_A_197_21#_c_139_n 0.0117969f $X=0.64 $Y=0.995 $X2=0
+ $Y2=0
cc_103 N_B1_N_c_103_n N_A_197_21#_c_148_n 0.0350274f $X=0.615 $Y=1.41 $X2=0
+ $Y2=0
cc_104 B1_N N_A_197_21#_c_148_n 0.00250598f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_105 N_B1_N_c_103_n N_A_197_21#_c_147_n 0.0259311f $X=0.615 $Y=1.41 $X2=0
+ $Y2=0
cc_106 B1_N N_A_197_21#_c_147_n 0.0010783f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_107 N_B1_N_c_106_n N_A_197_21#_c_147_n 0.00192841f $X=0.77 $Y=1.285 $X2=0
+ $Y2=0
cc_108 N_B1_N_c_103_n N_A_27_297#_c_315_n 0.0129228f $X=0.615 $Y=1.41 $X2=0
+ $Y2=0
cc_109 B1_N N_A_27_297#_c_315_n 0.0207078f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_110 N_B1_N_c_106_n N_A_27_297#_c_315_n 0.0036792f $X=0.77 $Y=1.285 $X2=0
+ $Y2=0
cc_111 N_B1_N_c_103_n N_A_27_297#_c_303_n 0.002158f $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B1_N_c_106_n N_A_27_297#_c_303_n 0.00653291f $X=0.77 $Y=1.285 $X2=0
+ $Y2=0
cc_113 N_B1_N_c_103_n N_A_27_297#_c_311_n 0.00511003f $X=0.615 $Y=1.41 $X2=0
+ $Y2=0
cc_114 B1_N N_A_27_297#_c_311_n 0.0194999f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_115 N_B1_N_c_106_n N_A_27_297#_c_311_n 7.71248e-19 $X=0.77 $Y=1.285 $X2=0
+ $Y2=0
cc_116 N_B1_N_c_103_n N_A_27_297#_c_304_n 0.00684842f $X=0.615 $Y=1.41 $X2=0
+ $Y2=0
cc_117 N_B1_N_c_104_n N_A_27_297#_c_304_n 0.00263902f $X=0.64 $Y=0.995 $X2=0
+ $Y2=0
cc_118 B1_N N_A_27_297#_c_304_n 0.00525983f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_119 N_B1_N_c_106_n N_A_27_297#_c_304_n 0.0171543f $X=0.77 $Y=1.285 $X2=0
+ $Y2=0
cc_120 B1_N N_VPWR_M1004_d 0.00436854f $X=0.605 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_121 N_B1_N_c_103_n N_VPWR_c_502_n 0.0117742f $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B1_N_c_103_n N_VPWR_c_501_n 0.00478793f $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B1_N_c_103_n N_VPWR_c_515_n 0.00315243f $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B1_N_c_103_n N_X_c_609_n 8.54878e-19 $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_125 B1_N N_X_c_609_n 0.0283819f $X=0.605 $Y=1.445 $X2=0 $Y2=0
cc_126 N_B1_N_c_106_n N_X_c_609_n 0.0146334f $X=0.77 $Y=1.285 $X2=0 $Y2=0
cc_127 N_B1_N_c_103_n N_VGND_c_705_n 2.31083e-19 $X=0.615 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B1_N_c_104_n N_VGND_c_705_n 0.00314514f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_129 N_B1_N_c_106_n N_VGND_c_705_n 0.0143616f $X=0.77 $Y=1.285 $X2=0 $Y2=0
cc_130 N_B1_N_c_104_n N_VGND_c_710_n 0.00585385f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_131 N_B1_N_c_104_n N_VGND_c_721_n 0.0116464f $X=0.64 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_197_21#_c_151_n N_A_27_297#_c_306_n 0.0319688f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_133 N_A_197_21#_c_164_p N_A_27_297#_c_307_n 0.0178703f $X=3.745 $Y=1.88 $X2=0
+ $Y2=0
cc_134 N_A_197_21#_c_146_n N_A_27_297#_c_307_n 0.0106027f $X=3.84 $Y=1.795 $X2=0
+ $Y2=0
cc_135 N_A_197_21#_c_144_n N_A_27_297#_c_301_n 0.00212658f $X=2.73 $Y=1.08 $X2=0
+ $Y2=0
cc_136 N_A_197_21#_c_145_n N_A_27_297#_c_301_n 0.0183654f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_137 N_A_197_21#_c_146_n N_A_27_297#_c_301_n 0.0021599f $X=3.84 $Y=1.795 $X2=0
+ $Y2=0
cc_138 N_A_197_21#_c_169_p N_A_27_297#_c_302_n 0.0034635f $X=3.84 $Y=0.895 $X2=0
+ $Y2=0
cc_139 N_A_197_21#_c_146_n N_A_27_297#_c_302_n 0.00256948f $X=3.84 $Y=1.795
+ $X2=0 $Y2=0
cc_140 N_A_197_21#_c_148_n N_A_27_297#_c_315_n 0.0183756f $X=1.085 $Y=1.41 $X2=0
+ $Y2=0
cc_141 N_A_197_21#_c_149_n N_A_27_297#_c_315_n 0.0130144f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_142 N_A_197_21#_c_150_n N_A_27_297#_c_315_n 0.0135034f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_143 N_A_197_21#_c_151_n N_A_27_297#_c_315_n 0.0148045f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_144 N_A_197_21#_c_143_n N_A_27_297#_c_315_n 0.0045399f $X=2.645 $Y=1.165
+ $X2=0 $Y2=0
cc_145 N_A_197_21#_c_176_p N_A_27_297#_c_315_n 0.0095715f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_146 N_A_197_21#_c_147_n N_A_27_297#_c_315_n 0.00105876f $X=2.495 $Y=1.202
+ $X2=0 $Y2=0
cc_147 N_A_197_21#_c_151_n N_A_27_297#_c_342_n 0.00479556f $X=2.495 $Y=1.41
+ $X2=0 $Y2=0
cc_148 N_A_197_21#_c_176_p N_A_27_297#_c_342_n 0.00425155f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_149 N_A_197_21#_M1016_s N_A_27_297#_c_310_n 0.00278173f $X=3.055 $Y=1.485
+ $X2=0 $Y2=0
cc_150 N_A_197_21#_c_151_n N_A_27_297#_c_310_n 0.00151723f $X=2.495 $Y=1.41
+ $X2=0 $Y2=0
cc_151 N_A_197_21#_c_143_n N_A_27_297#_c_310_n 0.0133161f $X=2.645 $Y=1.165
+ $X2=0 $Y2=0
cc_152 N_A_197_21#_c_145_n N_A_27_297#_c_310_n 0.00538384f $X=3.745 $Y=0.77
+ $X2=0 $Y2=0
cc_153 N_A_197_21#_c_146_n N_A_27_297#_c_310_n 0.0121236f $X=3.84 $Y=1.795 $X2=0
+ $Y2=0
cc_154 N_A_197_21#_c_176_p N_A_27_297#_c_310_n 0.00700741f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_155 N_A_197_21#_c_147_n N_A_27_297#_c_310_n 8.80522e-19 $X=2.495 $Y=1.202
+ $X2=0 $Y2=0
cc_156 N_A_197_21#_c_143_n N_A_27_297#_c_351_n 0.0141966f $X=2.645 $Y=1.165
+ $X2=0 $Y2=0
cc_157 N_A_197_21#_c_145_n N_A_27_297#_c_351_n 0.0318105f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_158 N_A_197_21#_c_164_p N_A_27_297#_c_351_n 0.00308902f $X=3.745 $Y=1.88
+ $X2=0 $Y2=0
cc_159 N_A_197_21#_c_146_n N_A_27_297#_c_351_n 0.00769191f $X=3.84 $Y=1.795
+ $X2=0 $Y2=0
cc_160 N_A_197_21#_c_176_p N_A_27_297#_c_351_n 0.00252632f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_161 N_A_197_21#_c_143_n N_A_27_297#_c_305_n 0.00168678f $X=2.645 $Y=1.165
+ $X2=0 $Y2=0
cc_162 N_A_197_21#_c_144_n N_A_27_297#_c_305_n 0.00216092f $X=2.73 $Y=1.08 $X2=0
+ $Y2=0
cc_163 N_A_197_21#_c_145_n N_A_27_297#_c_305_n 0.0187869f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_164 N_A_197_21#_c_164_p N_A_27_297#_c_305_n 0.00554968f $X=3.745 $Y=1.88
+ $X2=0 $Y2=0
cc_165 N_A_197_21#_c_146_n N_A_27_297#_c_305_n 0.0265093f $X=3.84 $Y=1.795 $X2=0
+ $Y2=0
cc_166 N_A_197_21#_c_153_n N_A_27_297#_c_305_n 0.00362047f $X=4.585 $Y=1.88
+ $X2=0 $Y2=0
cc_167 N_A_197_21#_c_176_p N_A_27_297#_c_305_n 0.00159385f $X=3.2 $Y=1.96 $X2=0
+ $Y2=0
cc_168 N_A_197_21#_c_147_n N_A_27_297#_c_305_n 0.0207f $X=2.495 $Y=1.202 $X2=0
+ $Y2=0
cc_169 N_A_197_21#_c_146_n N_A2_c_409_n 9.11308e-19 $X=3.84 $Y=1.795 $X2=-0.19
+ $Y2=-0.24
cc_170 N_A_197_21#_c_146_n N_A2_c_413_n 0.00703154f $X=3.84 $Y=1.795 $X2=0 $Y2=0
cc_171 N_A_197_21#_c_153_n N_A2_c_413_n 0.0149035f $X=4.585 $Y=1.88 $X2=0 $Y2=0
cc_172 N_A_197_21#_c_154_n N_A2_c_413_n 5.86193e-19 $X=4.71 $Y=1.62 $X2=0 $Y2=0
cc_173 N_A_197_21#_c_154_n N_A2_c_414_n 5.52341e-19 $X=4.71 $Y=1.62 $X2=0 $Y2=0
cc_174 N_A_197_21#_c_146_n A2 0.012255f $X=3.84 $Y=1.795 $X2=0 $Y2=0
cc_175 N_A_197_21#_c_153_n A2 0.0111726f $X=4.585 $Y=1.88 $X2=0 $Y2=0
cc_176 N_A_197_21#_c_154_n A2 0.0198142f $X=4.71 $Y=1.62 $X2=0 $Y2=0
cc_177 N_A_197_21#_c_146_n N_A2_c_412_n 0.00274868f $X=3.84 $Y=1.795 $X2=0 $Y2=0
cc_178 N_A_197_21#_c_154_n N_A2_c_412_n 0.00622399f $X=4.71 $Y=1.62 $X2=0 $Y2=0
cc_179 N_A_197_21#_c_164_p N_VPWR_M1020_d 0.00447905f $X=3.745 $Y=1.88 $X2=0
+ $Y2=0
cc_180 N_A_197_21#_c_146_n N_VPWR_M1020_d 0.00477104f $X=3.84 $Y=1.795 $X2=0
+ $Y2=0
cc_181 N_A_197_21#_c_155_n N_VPWR_M1020_d 0.00100143f $X=3.84 $Y=1.88 $X2=0
+ $Y2=0
cc_182 N_A_197_21#_c_148_n N_VPWR_c_502_n 0.00891164f $X=1.085 $Y=1.41 $X2=0
+ $Y2=0
cc_183 N_A_197_21#_c_149_n N_VPWR_c_502_n 0.0011802f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_197_21#_c_148_n N_VPWR_c_503_n 0.00458874f $X=1.085 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_197_21#_c_149_n N_VPWR_c_503_n 0.00315243f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_197_21#_c_148_n N_VPWR_c_504_n 0.001313f $X=1.085 $Y=1.41 $X2=0 $Y2=0
cc_187 N_A_197_21#_c_149_n N_VPWR_c_504_n 0.0119578f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_197_21#_c_150_n N_VPWR_c_504_n 0.00894471f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_197_21#_c_151_n N_VPWR_c_504_n 0.0011802f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_190 N_A_197_21#_c_150_n N_VPWR_c_505_n 0.00458874f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A_197_21#_c_151_n N_VPWR_c_505_n 0.00315243f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_192 N_A_197_21#_c_150_n N_VPWR_c_506_n 0.001313f $X=2.025 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_197_21#_c_151_n N_VPWR_c_506_n 0.0119247f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_194 N_A_197_21#_c_176_p N_VPWR_c_506_n 0.0153021f $X=3.2 $Y=1.96 $X2=0 $Y2=0
cc_195 N_A_197_21#_c_164_p N_VPWR_c_507_n 0.0128191f $X=3.745 $Y=1.88 $X2=0
+ $Y2=0
cc_196 N_A_197_21#_c_155_n N_VPWR_c_507_n 0.00467627f $X=3.84 $Y=1.88 $X2=0
+ $Y2=0
cc_197 N_A_197_21#_c_164_p N_VPWR_c_509_n 0.00285991f $X=3.745 $Y=1.88 $X2=0
+ $Y2=0
cc_198 N_A_197_21#_c_176_p N_VPWR_c_509_n 0.011801f $X=3.2 $Y=1.96 $X2=0 $Y2=0
cc_199 N_A_197_21#_c_153_n N_VPWR_c_511_n 0.00146078f $X=4.585 $Y=1.88 $X2=0
+ $Y2=0
cc_200 N_A_197_21#_c_155_n N_VPWR_c_511_n 0.00216841f $X=3.84 $Y=1.88 $X2=0
+ $Y2=0
cc_201 N_A_197_21#_M1016_s N_VPWR_c_501_n 0.00470726f $X=3.055 $Y=1.485 $X2=0
+ $Y2=0
cc_202 N_A_197_21#_M1001_s N_VPWR_c_501_n 0.00232895f $X=4.565 $Y=1.485 $X2=0
+ $Y2=0
cc_203 N_A_197_21#_c_148_n N_VPWR_c_501_n 0.00528719f $X=1.085 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_197_21#_c_149_n N_VPWR_c_501_n 0.00382819f $X=1.555 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_197_21#_c_150_n N_VPWR_c_501_n 0.00528719f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_197_21#_c_151_n N_VPWR_c_501_n 0.00382819f $X=2.495 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_197_21#_c_164_p N_VPWR_c_501_n 0.00654537f $X=3.745 $Y=1.88 $X2=0
+ $Y2=0
cc_208 N_A_197_21#_c_153_n N_VPWR_c_501_n 0.00373458f $X=4.585 $Y=1.88 $X2=0
+ $Y2=0
cc_209 N_A_197_21#_c_176_p N_VPWR_c_501_n 0.00646745f $X=3.2 $Y=1.96 $X2=0 $Y2=0
cc_210 N_A_197_21#_c_155_n N_VPWR_c_501_n 0.00397985f $X=3.84 $Y=1.88 $X2=0
+ $Y2=0
cc_211 N_A_197_21#_c_140_n N_X_c_616_n 0.00686626f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_197_21#_c_141_n N_X_c_616_n 5.46296e-19 $X=2 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_197_21#_c_139_n N_X_c_609_n 0.00267459f $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_197_21#_c_148_n N_X_c_609_n 0.00457989f $X=1.085 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_197_21#_c_140_n N_X_c_609_n 0.00268808f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_216 N_A_197_21#_c_149_n N_X_c_609_n 0.011794f $X=1.555 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_197_21#_c_141_n N_X_c_609_n 0.00209447f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A_197_21#_c_150_n N_X_c_609_n 8.32659e-19 $X=2.025 $Y=1.41 $X2=0 $Y2=0
cc_219 N_A_197_21#_c_143_n N_X_c_609_n 0.0139251f $X=2.645 $Y=1.165 $X2=0 $Y2=0
cc_220 N_A_197_21#_c_147_n N_X_c_609_n 0.0496141f $X=2.495 $Y=1.202 $X2=0 $Y2=0
cc_221 N_A_197_21#_c_141_n N_X_c_610_n 0.0103655f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_222 N_A_197_21#_c_142_n N_X_c_610_n 0.001178f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_197_21#_c_143_n N_X_c_610_n 0.0381594f $X=2.645 $Y=1.165 $X2=0 $Y2=0
cc_224 N_A_197_21#_c_144_n N_X_c_610_n 8.87833e-19 $X=2.73 $Y=1.08 $X2=0 $Y2=0
cc_225 N_A_197_21#_c_256_p N_X_c_610_n 0.00575362f $X=2.815 $Y=0.77 $X2=0 $Y2=0
cc_226 N_A_197_21#_c_147_n N_X_c_610_n 0.00870159f $X=2.495 $Y=1.202 $X2=0 $Y2=0
cc_227 N_A_197_21#_c_150_n N_X_c_612_n 0.0131867f $X=2.025 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_197_21#_c_151_n N_X_c_612_n 0.00404756f $X=2.495 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_197_21#_c_143_n N_X_c_612_n 0.0359366f $X=2.645 $Y=1.165 $X2=0 $Y2=0
cc_230 N_A_197_21#_c_147_n N_X_c_612_n 0.014314f $X=2.495 $Y=1.202 $X2=0 $Y2=0
cc_231 N_A_197_21#_c_139_n N_X_c_636_n 3.6982e-19 $X=1.06 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_197_21#_c_140_n N_X_c_636_n 0.00837496f $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_197_21#_c_140_n N_X_c_638_n 5.25321e-19 $X=1.53 $Y=0.995 $X2=0 $Y2=0
cc_234 N_A_197_21#_c_141_n N_X_c_638_n 0.00651696f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_235 N_A_197_21#_c_142_n N_X_c_638_n 0.00642131f $X=2.52 $Y=0.995 $X2=0 $Y2=0
cc_236 N_A_197_21#_c_153_n N_A_823_297#_M1001_d 0.00822237f $X=4.585 $Y=1.88
+ $X2=-0.19 $Y2=-0.24
cc_237 N_A_197_21#_M1001_s N_A_823_297#_c_672_n 0.00352392f $X=4.565 $Y=1.485
+ $X2=0 $Y2=0
cc_238 N_A_197_21#_c_153_n N_A_823_297#_c_672_n 0.00637037f $X=4.585 $Y=1.88
+ $X2=0 $Y2=0
cc_239 N_A_197_21#_c_270_p N_A_823_297#_c_672_n 0.0134104f $X=4.707 $Y=1.795
+ $X2=0 $Y2=0
cc_240 N_A_197_21#_c_154_n N_A_823_297#_c_666_n 0.00768652f $X=4.71 $Y=1.62
+ $X2=0 $Y2=0
cc_241 N_A_197_21#_c_153_n N_A_823_297#_c_670_n 0.0216429f $X=4.585 $Y=1.88
+ $X2=0 $Y2=0
cc_242 N_A_197_21#_c_145_n N_VGND_M1021_s 9.20278e-19 $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_243 N_A_197_21#_c_256_p N_VGND_M1021_s 0.00383f $X=2.815 $Y=0.77 $X2=0 $Y2=0
cc_244 N_A_197_21#_c_139_n N_VGND_c_705_n 0.00283672f $X=1.06 $Y=0.995 $X2=0
+ $Y2=0
cc_245 N_A_197_21#_c_140_n N_VGND_c_706_n 0.00379224f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_246 N_A_197_21#_c_141_n N_VGND_c_706_n 0.00276126f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_247 N_A_197_21#_c_141_n N_VGND_c_707_n 9.58281e-19 $X=2 $Y=0.995 $X2=0 $Y2=0
cc_248 N_A_197_21#_c_142_n N_VGND_c_707_n 0.00962528f $X=2.52 $Y=0.995 $X2=0
+ $Y2=0
cc_249 N_A_197_21#_c_143_n N_VGND_c_707_n 0.00150739f $X=2.645 $Y=1.165 $X2=0
+ $Y2=0
cc_250 N_A_197_21#_c_145_n N_VGND_c_707_n 0.00628317f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_251 N_A_197_21#_c_256_p N_VGND_c_707_n 0.0136659f $X=2.815 $Y=0.77 $X2=0
+ $Y2=0
cc_252 N_A_197_21#_c_139_n N_VGND_c_712_n 0.00585385f $X=1.06 $Y=0.995 $X2=0
+ $Y2=0
cc_253 N_A_197_21#_c_140_n N_VGND_c_712_n 0.00423225f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_254 N_A_197_21#_c_141_n N_VGND_c_714_n 0.00423334f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_255 N_A_197_21#_c_142_n N_VGND_c_714_n 0.0046653f $X=2.52 $Y=0.995 $X2=0
+ $Y2=0
cc_256 N_A_197_21#_c_145_n N_VGND_c_716_n 0.00385412f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_257 N_A_197_21#_M1003_s N_VGND_c_721_n 0.00256987f $X=3.585 $Y=0.235 $X2=0
+ $Y2=0
cc_258 N_A_197_21#_c_139_n N_VGND_c_721_n 0.0106913f $X=1.06 $Y=0.995 $X2=0
+ $Y2=0
cc_259 N_A_197_21#_c_140_n N_VGND_c_721_n 0.00609103f $X=1.53 $Y=0.995 $X2=0
+ $Y2=0
cc_260 N_A_197_21#_c_141_n N_VGND_c_721_n 0.00608558f $X=2 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_197_21#_c_142_n N_VGND_c_721_n 0.00821929f $X=2.52 $Y=0.995 $X2=0
+ $Y2=0
cc_262 N_A_197_21#_c_145_n N_VGND_c_721_n 0.00765093f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_263 N_A_197_21#_c_256_p N_VGND_c_721_n 8.32259e-19 $X=2.815 $Y=0.77 $X2=0
+ $Y2=0
cc_264 N_A_197_21#_c_145_n N_A_635_47#_M1003_d 0.00316796f $X=3.745 $Y=0.77
+ $X2=-0.19 $Y2=-0.24
cc_265 N_A_197_21#_M1003_s N_A_635_47#_c_813_n 0.0039919f $X=3.585 $Y=0.235
+ $X2=0 $Y2=0
cc_266 N_A_197_21#_c_145_n N_A_635_47#_c_813_n 0.0374711f $X=3.745 $Y=0.77 $X2=0
+ $Y2=0
cc_267 N_A_197_21#_c_169_p N_A_635_47#_c_813_n 0.0102417f $X=3.84 $Y=0.895 $X2=0
+ $Y2=0
cc_268 N_A_197_21#_c_169_p N_A_635_47#_c_814_n 0.0174391f $X=3.84 $Y=0.895 $X2=0
+ $Y2=0
cc_269 N_A_197_21#_c_146_n N_A_635_47#_c_814_n 6.42107e-19 $X=3.84 $Y=1.795
+ $X2=0 $Y2=0
cc_270 N_A_27_297#_c_302_n N_A2_c_409_n 0.0119754f $X=3.98 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_271 N_A_27_297#_c_305_n A2 0.00208754f $X=3.51 $Y=1.202 $X2=0 $Y2=0
cc_272 N_A_27_297#_c_305_n N_A2_c_412_n 0.0119754f $X=3.51 $Y=1.202 $X2=0 $Y2=0
cc_273 N_A_27_297#_c_315_n N_VPWR_M1004_d 0.00358615f $X=2.645 $Y=1.96 $X2=-0.19
+ $Y2=-0.24
cc_274 N_A_27_297#_c_315_n N_VPWR_M1006_d 0.00344677f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_275 N_A_27_297#_c_315_n N_VPWR_M1014_d 0.00402346f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_276 N_A_27_297#_c_342_n N_VPWR_M1014_d 0.00638008f $X=2.73 $Y=1.875 $X2=0
+ $Y2=0
cc_277 N_A_27_297#_c_310_n N_VPWR_M1014_d 0.00205406f $X=3.095 $Y=1.445 $X2=0
+ $Y2=0
cc_278 N_A_27_297#_c_309_n N_VPWR_c_502_n 0.017382f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_279 N_A_27_297#_c_315_n N_VPWR_c_502_n 0.0198692f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_280 N_A_27_297#_c_315_n N_VPWR_c_503_n 0.00784602f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_281 N_A_27_297#_c_315_n N_VPWR_c_504_n 0.0198692f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_282 N_A_27_297#_c_315_n N_VPWR_c_505_n 0.00784602f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_283 N_A_27_297#_c_306_n N_VPWR_c_506_n 0.00768171f $X=2.965 $Y=1.41 $X2=0
+ $Y2=0
cc_284 N_A_27_297#_c_307_n N_VPWR_c_506_n 5.34214e-19 $X=3.435 $Y=1.41 $X2=0
+ $Y2=0
cc_285 N_A_27_297#_c_315_n N_VPWR_c_506_n 0.0191257f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_286 N_A_27_297#_c_310_n N_VPWR_c_506_n 6.09944e-19 $X=3.095 $Y=1.445 $X2=0
+ $Y2=0
cc_287 N_A_27_297#_c_307_n N_VPWR_c_507_n 0.00341296f $X=3.435 $Y=1.41 $X2=0
+ $Y2=0
cc_288 N_A_27_297#_c_306_n N_VPWR_c_509_n 0.00622633f $X=2.965 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_27_297#_c_307_n N_VPWR_c_509_n 0.0053025f $X=3.435 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_27_297#_M1004_s N_VPWR_c_501_n 0.00352744f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_291 N_A_27_297#_c_306_n N_VPWR_c_501_n 0.0104011f $X=2.965 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_27_297#_c_307_n N_VPWR_c_501_n 0.00819982f $X=3.435 $Y=1.41 $X2=0
+ $Y2=0
cc_293 N_A_27_297#_c_309_n N_VPWR_c_501_n 0.0134021f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_294 N_A_27_297#_c_315_n N_VPWR_c_501_n 0.037451f $X=2.645 $Y=1.96 $X2=0 $Y2=0
cc_295 N_A_27_297#_c_309_n N_VPWR_c_515_n 0.0245389f $X=0.35 $Y=2.3 $X2=0 $Y2=0
cc_296 N_A_27_297#_c_315_n N_VPWR_c_515_n 0.00265325f $X=2.645 $Y=1.96 $X2=0
+ $Y2=0
cc_297 N_A_27_297#_c_315_n N_X_M1000_s 0.00489785f $X=2.645 $Y=1.96 $X2=0 $Y2=0
cc_298 N_A_27_297#_c_315_n N_X_M1010_s 0.00490173f $X=2.645 $Y=1.96 $X2=0 $Y2=0
cc_299 N_A_27_297#_c_315_n N_X_c_609_n 0.0296719f $X=2.645 $Y=1.96 $X2=0 $Y2=0
cc_300 N_A_27_297#_c_315_n N_X_c_612_n 0.0400839f $X=2.645 $Y=1.96 $X2=0 $Y2=0
cc_301 N_A_27_297#_c_342_n N_X_c_612_n 0.0057271f $X=2.73 $Y=1.875 $X2=0 $Y2=0
cc_302 N_A_27_297#_c_310_n N_X_c_612_n 0.0119093f $X=3.095 $Y=1.445 $X2=0 $Y2=0
cc_303 N_A_27_297#_c_301_n N_VGND_c_707_n 0.00217307f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_304 N_A_27_297#_c_303_n N_VGND_c_710_n 0.0290883f $X=0.38 $Y=0.39 $X2=0 $Y2=0
cc_305 N_A_27_297#_c_301_n N_VGND_c_716_n 0.00357877f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_306 N_A_27_297#_c_302_n N_VGND_c_716_n 0.00357877f $X=3.98 $Y=0.995 $X2=0
+ $Y2=0
cc_307 N_A_27_297#_M1017_s N_VGND_c_721_n 0.00357047f $X=0.21 $Y=0.235 $X2=0
+ $Y2=0
cc_308 N_A_27_297#_c_301_n N_VGND_c_721_n 0.00668309f $X=3.51 $Y=0.995 $X2=0
+ $Y2=0
cc_309 N_A_27_297#_c_302_n N_VGND_c_721_n 0.00550244f $X=3.98 $Y=0.995 $X2=0
+ $Y2=0
cc_310 N_A_27_297#_c_303_n N_VGND_c_721_n 0.0175126f $X=0.38 $Y=0.39 $X2=0 $Y2=0
cc_311 N_A_27_297#_c_301_n N_A_635_47#_c_813_n 0.00931157f $X=3.51 $Y=0.995
+ $X2=0 $Y2=0
cc_312 N_A_27_297#_c_302_n N_A_635_47#_c_813_n 0.0130858f $X=3.98 $Y=0.995 $X2=0
+ $Y2=0
cc_313 N_A_27_297#_c_305_n N_A_635_47#_c_813_n 3.367e-19 $X=3.51 $Y=1.202 $X2=0
+ $Y2=0
cc_314 N_A_27_297#_c_302_n N_A_635_47#_c_814_n 8.83927e-19 $X=3.98 $Y=0.995
+ $X2=0 $Y2=0
cc_315 N_A2_c_410_n N_A1_c_463_n 0.0176256f $X=4.97 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_316 N_A2_c_414_n N_A1_c_467_n 0.00966765f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_317 A2 A1 0.0136085f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_318 A2 N_A1_c_466_n 0.00578274f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_319 N_A2_c_412_n N_A1_c_466_n 0.0176256f $X=4.945 $Y=1.202 $X2=0 $Y2=0
cc_320 N_A2_c_413_n N_VPWR_c_507_n 0.00197731f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_321 N_A2_c_414_n N_VPWR_c_508_n 0.00110692f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_322 N_A2_c_413_n N_VPWR_c_511_n 0.00429453f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_323 N_A2_c_414_n N_VPWR_c_511_n 0.00429453f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_324 N_A2_c_413_n N_VPWR_c_501_n 0.00734734f $X=4.475 $Y=1.41 $X2=0 $Y2=0
cc_325 N_A2_c_414_n N_VPWR_c_501_n 0.00609021f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_326 N_A2_c_413_n N_A_823_297#_c_672_n 0.00991367f $X=4.475 $Y=1.41 $X2=0
+ $Y2=0
cc_327 N_A2_c_414_n N_A_823_297#_c_672_n 0.0143148f $X=4.945 $Y=1.41 $X2=0 $Y2=0
cc_328 N_A2_c_414_n N_A_823_297#_c_666_n 0.00133266f $X=4.945 $Y=1.41 $X2=0
+ $Y2=0
cc_329 A2 N_A_823_297#_c_666_n 0.0139423f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_330 A2 N_A_823_297#_c_667_n 0.0040358f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_331 N_A2_c_409_n N_VGND_c_708_n 0.00385178f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_332 N_A2_c_410_n N_VGND_c_708_n 0.00365402f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_333 N_A2_c_409_n N_VGND_c_716_n 0.00421816f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_334 N_A2_c_410_n N_VGND_c_718_n 0.00396605f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_335 N_A2_c_409_n N_VGND_c_721_n 0.00623587f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_336 N_A2_c_410_n N_VGND_c_721_n 0.00583042f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_337 N_A2_c_409_n N_A_635_47#_c_829_n 0.00284788f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_338 N_A2_c_409_n N_A_635_47#_c_814_n 0.0052094f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_339 N_A2_c_410_n N_A_635_47#_c_814_n 4.72003e-19 $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_340 A2 N_A_635_47#_c_814_n 0.0188951f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_341 N_A2_c_409_n N_A_635_47#_c_815_n 0.00929182f $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_342 N_A2_c_410_n N_A_635_47#_c_815_n 0.00650032f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_343 A2 N_A_635_47#_c_815_n 0.0399344f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_344 N_A2_c_412_n N_A_635_47#_c_815_n 0.00468948f $X=4.945 $Y=1.202 $X2=0
+ $Y2=0
cc_345 N_A2_c_409_n N_A_635_47#_c_837_n 5.69266e-19 $X=4.45 $Y=0.995 $X2=0 $Y2=0
cc_346 N_A2_c_410_n N_A_635_47#_c_837_n 0.00857123f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_347 N_A2_c_410_n N_A_635_47#_c_818_n 0.00269873f $X=4.97 $Y=0.995 $X2=0 $Y2=0
cc_348 A2 N_A_635_47#_c_818_n 0.0294984f $X=4.735 $Y=1.105 $X2=0 $Y2=0
cc_349 N_A1_c_467_n N_VPWR_c_508_n 0.0163934f $X=5.415 $Y=1.41 $X2=0 $Y2=0
cc_350 N_A1_c_468_n N_VPWR_c_508_n 0.0135516f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_351 N_A1_c_467_n N_VPWR_c_511_n 0.00427505f $X=5.415 $Y=1.41 $X2=0 $Y2=0
cc_352 N_A1_c_468_n N_VPWR_c_513_n 0.00622633f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_353 N_A1_c_467_n N_VPWR_c_501_n 0.00735499f $X=5.415 $Y=1.41 $X2=0 $Y2=0
cc_354 N_A1_c_468_n N_VPWR_c_501_n 0.0113638f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_355 N_A1_c_467_n N_A_823_297#_c_667_n 0.0170057f $X=5.415 $Y=1.41 $X2=0 $Y2=0
cc_356 N_A1_c_468_n N_A_823_297#_c_667_n 0.0166678f $X=5.885 $Y=1.41 $X2=0 $Y2=0
cc_357 A1 N_A_823_297#_c_667_n 0.0343628f $X=5.755 $Y=1.105 $X2=0 $Y2=0
cc_358 N_A1_c_466_n N_A_823_297#_c_667_n 0.00815835f $X=5.885 $Y=1.202 $X2=0
+ $Y2=0
cc_359 A1 N_A_823_297#_c_668_n 0.0225537f $X=5.755 $Y=1.105 $X2=0 $Y2=0
cc_360 N_A1_c_463_n N_VGND_c_709_n 0.00385467f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_361 N_A1_c_464_n N_VGND_c_709_n 0.00381583f $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_362 N_A1_c_463_n N_VGND_c_718_n 0.00423334f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_363 N_A1_c_464_n N_VGND_c_720_n 0.00397706f $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_364 N_A1_c_463_n N_VGND_c_721_n 0.00610858f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_365 N_A1_c_464_n N_VGND_c_721_n 0.00681132f $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_366 N_A1_c_463_n N_A_635_47#_c_837_n 0.00693563f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_367 N_A1_c_464_n N_A_635_47#_c_837_n 5.34196e-19 $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_368 N_A1_c_463_n N_A_635_47#_c_816_n 0.0107693f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_369 N_A1_c_464_n N_A_635_47#_c_816_n 0.00937294f $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_370 A1 N_A_635_47#_c_816_n 0.0599937f $X=5.755 $Y=1.105 $X2=0 $Y2=0
cc_371 N_A1_c_466_n N_A_635_47#_c_816_n 0.00468948f $X=5.885 $Y=1.202 $X2=0
+ $Y2=0
cc_372 N_A1_c_463_n N_A_635_47#_c_817_n 5.66376e-19 $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_373 N_A1_c_464_n N_A_635_47#_c_817_n 0.0084675f $X=5.91 $Y=0.995 $X2=0 $Y2=0
cc_374 N_A1_c_463_n N_A_635_47#_c_818_n 0.00142536f $X=5.39 $Y=0.995 $X2=0 $Y2=0
cc_375 N_VPWR_c_501_n N_X_M1000_s 0.0035556f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_376 N_VPWR_c_501_n N_X_M1010_s 0.0035556f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_377 N_VPWR_M1006_d N_X_c_612_n 0.00185701f $X=1.645 $Y=1.485 $X2=0 $Y2=0
cc_378 N_VPWR_c_501_n N_A_823_297#_M1001_d 0.0021672f $X=6.21 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_379 N_VPWR_c_501_n N_A_823_297#_M1008_d 0.00436089f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_380 N_VPWR_c_501_n N_A_823_297#_M1018_d 0.00442207f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_381 N_VPWR_c_511_n N_A_823_297#_c_672_n 0.0415876f $X=5.435 $Y=2.72 $X2=0
+ $Y2=0
cc_382 N_VPWR_c_501_n N_A_823_297#_c_672_n 0.0268901f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_383 N_VPWR_c_508_n N_A_823_297#_c_692_n 0.0484833f $X=5.65 $Y=2 $X2=0 $Y2=0
cc_384 N_VPWR_c_511_n N_A_823_297#_c_692_n 0.0119545f $X=5.435 $Y=2.72 $X2=0
+ $Y2=0
cc_385 N_VPWR_c_501_n N_A_823_297#_c_692_n 0.006547f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_386 N_VPWR_M1015_s N_A_823_297#_c_667_n 0.00188315f $X=5.505 $Y=1.485 $X2=0
+ $Y2=0
cc_387 N_VPWR_c_508_n N_A_823_297#_c_667_n 0.0212439f $X=5.65 $Y=2 $X2=0 $Y2=0
cc_388 N_VPWR_c_508_n N_A_823_297#_c_669_n 0.0399729f $X=5.65 $Y=2 $X2=0 $Y2=0
cc_389 N_VPWR_c_513_n N_A_823_297#_c_669_n 0.019258f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_390 N_VPWR_c_501_n N_A_823_297#_c_669_n 0.0105137f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_391 N_VPWR_c_507_n N_A_823_297#_c_670_n 0.0212565f $X=3.67 $Y=2.3 $X2=0 $Y2=0
cc_392 N_VPWR_c_511_n N_A_823_297#_c_670_n 0.0193258f $X=5.435 $Y=2.72 $X2=0
+ $Y2=0
cc_393 N_VPWR_c_501_n N_A_823_297#_c_670_n 0.0108939f $X=6.21 $Y=2.72 $X2=0
+ $Y2=0
cc_394 N_X_c_610_n N_VGND_M1009_s 0.00168466f $X=2.045 $Y=0.817 $X2=0 $Y2=0
cc_395 N_X_c_636_n N_VGND_M1009_s 8.66594e-19 $X=1.43 $Y=0.817 $X2=0 $Y2=0
cc_396 N_X_c_636_n N_VGND_c_705_n 0.00133683f $X=1.43 $Y=0.817 $X2=0 $Y2=0
cc_397 N_X_c_616_n N_VGND_c_706_n 0.0181628f $X=1.32 $Y=0.39 $X2=0 $Y2=0
cc_398 N_X_c_610_n N_VGND_c_706_n 0.01275f $X=2.045 $Y=0.817 $X2=0 $Y2=0
cc_399 N_X_c_638_n N_VGND_c_707_n 0.0156743f $X=2.21 $Y=0.39 $X2=0 $Y2=0
cc_400 N_X_c_616_n N_VGND_c_712_n 0.0197303f $X=1.32 $Y=0.39 $X2=0 $Y2=0
cc_401 N_X_c_636_n N_VGND_c_712_n 0.00289665f $X=1.43 $Y=0.817 $X2=0 $Y2=0
cc_402 N_X_c_610_n N_VGND_c_714_n 0.00198981f $X=2.045 $Y=0.817 $X2=0 $Y2=0
cc_403 N_X_c_638_n N_VGND_c_714_n 0.0209326f $X=2.21 $Y=0.39 $X2=0 $Y2=0
cc_404 N_X_M1007_d N_VGND_c_721_n 0.00324782f $X=1.135 $Y=0.235 $X2=0 $Y2=0
cc_405 N_X_M1013_d N_VGND_c_721_n 0.00542784f $X=2.075 $Y=0.235 $X2=0 $Y2=0
cc_406 N_X_c_616_n N_VGND_c_721_n 0.0124268f $X=1.32 $Y=0.39 $X2=0 $Y2=0
cc_407 N_X_c_610_n N_VGND_c_721_n 0.00450655f $X=2.045 $Y=0.817 $X2=0 $Y2=0
cc_408 N_X_c_636_n N_VGND_c_721_n 0.00553889f $X=1.43 $Y=0.817 $X2=0 $Y2=0
cc_409 N_X_c_638_n N_VGND_c_721_n 0.0124144f $X=2.21 $Y=0.39 $X2=0 $Y2=0
cc_410 N_A_823_297#_c_667_n N_A_635_47#_c_816_n 0.00554576f $X=6.035 $Y=1.56
+ $X2=0 $Y2=0
cc_411 N_A_823_297#_c_667_n N_A_635_47#_c_818_n 7.50318e-19 $X=6.035 $Y=1.56
+ $X2=0 $Y2=0
cc_412 N_VGND_c_721_n N_A_635_47#_M1003_d 0.00209344f $X=6.21 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_413 N_VGND_c_721_n N_A_635_47#_M1011_d 0.0025536f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_414 N_VGND_c_721_n N_A_635_47#_M1019_s 0.00215201f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_415 N_VGND_c_721_n N_A_635_47#_M1012_d 0.00226063f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_416 N_VGND_c_707_n N_A_635_47#_c_813_n 0.0166161f $X=2.73 $Y=0.39 $X2=0 $Y2=0
cc_417 N_VGND_c_716_n N_A_635_47#_c_813_n 0.0604763f $X=4.625 $Y=0 $X2=0 $Y2=0
cc_418 N_VGND_c_721_n N_A_635_47#_c_813_n 0.0378144f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_419 N_VGND_c_708_n N_A_635_47#_c_829_n 0.0141571f $X=4.71 $Y=0.39 $X2=0 $Y2=0
cc_420 N_VGND_c_716_n N_A_635_47#_c_829_n 0.015453f $X=4.625 $Y=0 $X2=0 $Y2=0
cc_421 N_VGND_c_721_n N_A_635_47#_c_829_n 0.00940698f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_422 N_VGND_c_708_n N_A_635_47#_c_814_n 0.00471242f $X=4.71 $Y=0.39 $X2=0
+ $Y2=0
cc_423 N_VGND_M1002_d N_A_635_47#_c_815_n 0.00348805f $X=4.525 $Y=0.235 $X2=0
+ $Y2=0
cc_424 N_VGND_c_708_n N_A_635_47#_c_815_n 0.0131987f $X=4.71 $Y=0.39 $X2=0 $Y2=0
cc_425 N_VGND_c_716_n N_A_635_47#_c_815_n 0.00266636f $X=4.625 $Y=0 $X2=0 $Y2=0
cc_426 N_VGND_c_718_n N_A_635_47#_c_815_n 0.00199443f $X=5.565 $Y=0 $X2=0 $Y2=0
cc_427 N_VGND_c_721_n N_A_635_47#_c_815_n 0.0100158f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_428 N_VGND_c_708_n N_A_635_47#_c_837_n 0.0223967f $X=4.71 $Y=0.39 $X2=0 $Y2=0
cc_429 N_VGND_c_709_n N_A_635_47#_c_837_n 0.0183628f $X=5.65 $Y=0.39 $X2=0 $Y2=0
cc_430 N_VGND_c_718_n N_A_635_47#_c_837_n 0.0222529f $X=5.565 $Y=0 $X2=0 $Y2=0
cc_431 N_VGND_c_721_n N_A_635_47#_c_837_n 0.0139016f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_432 N_VGND_M1005_s N_A_635_47#_c_816_n 0.00348805f $X=5.465 $Y=0.235 $X2=0
+ $Y2=0
cc_433 N_VGND_c_709_n N_A_635_47#_c_816_n 0.0131987f $X=5.65 $Y=0.39 $X2=0 $Y2=0
cc_434 N_VGND_c_718_n N_A_635_47#_c_816_n 0.00266636f $X=5.565 $Y=0 $X2=0 $Y2=0
cc_435 N_VGND_c_720_n N_A_635_47#_c_816_n 0.00199443f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_436 N_VGND_c_721_n N_A_635_47#_c_816_n 0.0100158f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_437 N_VGND_c_709_n N_A_635_47#_c_817_n 0.021759f $X=5.65 $Y=0.39 $X2=0 $Y2=0
cc_438 N_VGND_c_720_n N_A_635_47#_c_817_n 0.0245357f $X=6.21 $Y=0 $X2=0 $Y2=0
cc_439 N_VGND_c_721_n N_A_635_47#_c_817_n 0.0149859f $X=6.21 $Y=0 $X2=0 $Y2=0
