* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
M1000 a_27_297# B1 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=5.4e+11p pd=5.08e+06u as=6.4e+11p ps=5.28e+06u
M1001 X a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.9e+11p pd=2.58e+06u as=1.01e+12p ps=8.02e+06u
M1002 VGND a_27_297# X VNB nshort w=650000u l=150000u
+  ad=6.955e+11p pd=6.04e+06u as=2.08e+11p ps=1.94e+06u
M1003 VPWR A2 a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_27_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_117_297# B2 a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_411_47# A1 a_27_297# VNB nshort w=650000u l=150000u
+  ad=2.47e+11p pd=2.06e+06u as=4.03e+11p ps=3.84e+06u
M1007 VGND A2 a_411_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_117_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_119_47# B2 VGND VNB nshort w=650000u l=150000u
+  ad=1.495e+11p pd=1.76e+06u as=0p ps=0u
M1010 a_27_297# B1 a_119_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VPWR a_27_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends
