* File: sky130_fd_sc_hdll__nor4_1.pxi.spice
* Created: Wed Sep  2 08:40:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__NOR4_1%D N_D_c_41_n N_D_M1004_g N_D_c_38_n N_D_M1006_g D
+ D N_D_c_40_n PM_SKY130_FD_SC_HDLL__NOR4_1%D
x_PM_SKY130_FD_SC_HDLL__NOR4_1%C N_C_c_66_n N_C_M1001_g N_C_c_67_n N_C_M1000_g C
+ N_C_c_68_n PM_SKY130_FD_SC_HDLL__NOR4_1%C
x_PM_SKY130_FD_SC_HDLL__NOR4_1%B N_B_c_97_n N_B_M1003_g N_B_c_98_n N_B_M1005_g B
+ N_B_c_99_n PM_SKY130_FD_SC_HDLL__NOR4_1%B
x_PM_SKY130_FD_SC_HDLL__NOR4_1%A N_A_c_127_n N_A_M1007_g N_A_c_128_n N_A_M1002_g
+ A PM_SKY130_FD_SC_HDLL__NOR4_1%A
x_PM_SKY130_FD_SC_HDLL__NOR4_1%Y N_Y_M1006_d N_Y_M1003_d N_Y_M1004_s N_Y_c_153_n
+ N_Y_c_166_n N_Y_c_160_n N_Y_c_173_n Y PM_SKY130_FD_SC_HDLL__NOR4_1%Y
x_PM_SKY130_FD_SC_HDLL__NOR4_1%VPWR N_VPWR_M1002_d N_VPWR_c_202_n N_VPWR_c_203_n
+ VPWR N_VPWR_c_204_n N_VPWR_c_201_n PM_SKY130_FD_SC_HDLL__NOR4_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NOR4_1%VGND N_VGND_M1006_s N_VGND_M1001_d N_VGND_M1007_d
+ N_VGND_c_228_n N_VGND_c_229_n N_VGND_c_230_n N_VGND_c_231_n VGND
+ N_VGND_c_232_n N_VGND_c_233_n N_VGND_c_234_n N_VGND_c_235_n
+ PM_SKY130_FD_SC_HDLL__NOR4_1%VGND
cc_1 VNB N_D_c_38_n 0.01926f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB D 0.0213864f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.765
cc_3 VNB N_D_c_40_n 0.0417582f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_C_c_66_n 0.0171826f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_C_c_67_n 0.0218625f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_C_c_68_n 0.00389583f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_7 VNB N_B_c_97_n 0.0176471f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_B_c_98_n 0.0211587f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB N_B_c_99_n 0.00377655f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_10 VNB N_A_c_127_n 0.0199384f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_A_c_128_n 0.0262827f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB A 0.0152725f $X=-0.19 $Y=-0.24 $X2=0.14 $Y2=1.105
cc_13 VNB N_Y_c_153_n 0.00300781f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.202
cc_14 VNB N_VPWR_c_201_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_228_n 0.00988671f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_229_n 0.0184357f $X=-0.19 $Y=-0.24 $X2=0.25 $Y2=1.16
cc_17 VNB N_VGND_c_230_n 0.00224107f $X=-0.19 $Y=-0.24 $X2=0.21 $Y2=0.85
cc_18 VNB N_VGND_c_231_n 0.016743f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_232_n 0.0177254f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_233_n 0.00507288f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_234_n 0.0416087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_235_n 0.166414f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VPB N_D_c_41_n 0.0211914f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_24 VPB D 0.00299612f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.765
cc_25 VPB N_D_c_40_n 0.0176465f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_26 VPB N_C_c_67_n 0.0252944f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_27 VPB N_C_c_68_n 0.00106949f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.202
cc_28 VPB N_B_c_98_n 0.0252138f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_29 VPB N_B_c_99_n 0.00111671f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.202
cc_30 VPB N_A_c_128_n 0.0301237f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_31 VPB A 0.00654538f $X=-0.19 $Y=1.305 $X2=0.14 $Y2=1.105
cc_32 VPB N_Y_c_153_n 0.00867061f $X=-0.19 $Y=1.305 $X2=0.25 $Y2=1.202
cc_33 VPB Y 0.0310196f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_VPWR_c_202_n 0.0170461f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_35 VPB N_VPWR_c_203_n 0.042952f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_36 VPB N_VPWR_c_204_n 0.0615046f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_201_n 0.048765f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 N_D_c_38_n N_C_c_66_n 0.0166177f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_39 N_D_c_41_n N_C_c_67_n 0.0403886f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_40 N_D_c_40_n N_C_c_67_n 0.0166177f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_41 N_D_c_41_n N_C_c_68_n 0.0031054f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_42 N_D_c_40_n N_C_c_68_n 3.71802e-19 $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_43 N_D_c_41_n N_Y_c_153_n 0.0215417f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_D_c_38_n N_Y_c_153_n 0.003979f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_45 D N_Y_c_153_n 0.0190584f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_46 N_D_c_40_n N_Y_c_153_n 0.0182104f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_47 N_D_c_38_n N_Y_c_160_n 0.0138251f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_48 D N_Y_c_160_n 0.0407467f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_49 N_D_c_41_n Y 0.0146709f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_50 N_D_c_41_n N_VPWR_c_204_n 0.00674013f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_D_c_41_n N_VPWR_c_201_n 0.0130761f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 D N_VGND_M1006_s 0.00410474f $X=0.145 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_53 N_D_c_38_n N_VGND_c_229_n 0.00769729f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 D N_VGND_c_229_n 0.021476f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_55 N_D_c_40_n N_VGND_c_229_n 0.00136792f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_56 N_D_c_38_n N_VGND_c_230_n 0.00162892f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_57 N_D_c_38_n N_VGND_c_232_n 0.00478994f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 N_D_c_38_n N_VGND_c_235_n 0.0090185f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_59 D N_VGND_c_235_n 0.00102136f $X=0.145 $Y=0.765 $X2=0 $Y2=0
cc_60 N_C_c_66_n N_B_c_97_n 0.020459f $X=0.99 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_61 N_C_c_67_n N_B_c_98_n 0.0701222f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_62 N_C_c_68_n N_B_c_98_n 0.00979907f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_63 N_C_c_67_n N_B_c_99_n 0.00131025f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_64 N_C_c_68_n N_B_c_99_n 0.112305f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_65 N_C_c_66_n N_Y_c_153_n 0.00705937f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_66 N_C_c_67_n N_Y_c_153_n 0.00190512f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_67 N_C_c_68_n N_Y_c_153_n 0.0482985f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_68 N_C_c_66_n N_Y_c_166_n 0.0119268f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_69 N_C_c_67_n N_Y_c_166_n 7.17521e-19 $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_70 N_C_c_68_n N_Y_c_166_n 0.023124f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_71 N_C_c_67_n Y 0.00228373f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_72 N_C_c_68_n Y 0.0228026f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_73 N_C_c_68_n A_221_297# 0.00934502f $X=1.05 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_74 N_C_c_67_n N_VPWR_c_204_n 0.00494341f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_75 N_C_c_68_n N_VPWR_c_204_n 0.0183088f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_76 N_C_c_67_n N_VPWR_c_201_n 0.00782099f $X=1.015 $Y=1.41 $X2=0 $Y2=0
cc_77 N_C_c_68_n N_VPWR_c_201_n 0.0115173f $X=1.05 $Y=1.16 $X2=0 $Y2=0
cc_78 N_C_c_66_n N_VGND_c_230_n 0.00933018f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_79 N_C_c_66_n N_VGND_c_232_n 0.00341689f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_80 N_C_c_66_n N_VGND_c_235_n 0.00417721f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_81 N_B_c_97_n N_A_c_127_n 0.0231983f $X=1.47 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_82 N_B_c_98_n N_A_c_128_n 0.0680868f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_99_n N_A_c_128_n 0.0141513f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_84 N_B_c_97_n A 9.24895e-19 $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_85 N_B_c_98_n A 6.55017e-19 $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B_c_99_n A 0.0472753f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_87 N_B_c_97_n N_Y_c_166_n 0.0124573f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_88 N_B_c_99_n N_Y_c_166_n 0.00888581f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_89 N_B_c_98_n N_Y_c_173_n 5.83574e-19 $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B_c_99_n N_Y_c_173_n 0.0125774f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_91 N_B_c_99_n A_317_297# 0.0120367f $X=1.54 $Y=1.16 $X2=-0.19 $Y2=-0.24
cc_92 N_B_c_99_n N_VPWR_c_203_n 0.0268678f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_93 N_B_c_98_n N_VPWR_c_204_n 0.00509313f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_99_n N_VPWR_c_204_n 0.0164055f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_95 N_B_c_98_n N_VPWR_c_201_n 0.0081207f $X=1.495 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_99_n N_VPWR_c_201_n 0.0104164f $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_97 N_B_c_97_n N_VGND_c_230_n 0.00168834f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_98 N_B_c_97_n N_VGND_c_231_n 0.00428022f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_99 N_B_c_97_n N_VGND_c_234_n 8.82544e-19 $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_100 N_B_c_97_n N_VGND_c_235_n 0.00607415f $X=1.47 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_c_127_n N_Y_c_173_n 0.00577904f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_102 A N_Y_c_173_n 0.0123591f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_103 A N_VPWR_M1002_d 0.00801559f $X=1.97 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_104 N_A_c_128_n N_VPWR_c_203_n 0.0097201f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_105 A N_VPWR_c_203_n 0.006131f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_106 N_A_c_128_n N_VPWR_c_204_n 0.00702461f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_107 N_A_c_128_n N_VPWR_c_201_n 0.0137498f $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_108 A N_VGND_M1007_d 0.0104772f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_109 N_A_c_127_n N_VGND_c_231_n 0.00395127f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_110 A N_VGND_c_231_n 0.00117536f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_111 N_A_c_127_n N_VGND_c_234_n 0.0099956f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_112 N_A_c_128_n N_VGND_c_234_n 3.64048e-19 $X=1.985 $Y=1.41 $X2=0 $Y2=0
cc_113 A N_VGND_c_234_n 0.0118441f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_114 N_A_c_127_n N_VGND_c_235_n 0.00586748f $X=1.96 $Y=0.995 $X2=0 $Y2=0
cc_115 A N_VGND_c_235_n 0.00264706f $X=1.97 $Y=0.765 $X2=0 $Y2=0
cc_116 N_Y_c_153_n A_117_297# 0.00746405f $X=0.645 $Y=1.495 $X2=-0.19 $Y2=-0.24
cc_117 Y N_VPWR_c_204_n 0.0195512f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_118 N_Y_M1004_s N_VPWR_c_201_n 0.00218082f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_119 Y N_VPWR_c_201_n 0.0125731f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_120 N_Y_c_166_n N_VGND_M1001_d 0.00585587f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_121 N_Y_c_160_n N_VGND_c_229_n 0.0143789f $X=0.73 $Y=0.55 $X2=0 $Y2=0
cc_122 N_Y_c_166_n N_VGND_c_230_n 0.0186246f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_123 N_Y_c_160_n N_VGND_c_230_n 0.00632053f $X=0.73 $Y=0.55 $X2=0 $Y2=0
cc_124 N_Y_c_166_n N_VGND_c_231_n 0.00307136f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_125 N_Y_c_173_n N_VGND_c_231_n 0.00610094f $X=1.68 $Y=0.55 $X2=0 $Y2=0
cc_126 N_Y_c_166_n N_VGND_c_232_n 0.00310943f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_127 N_Y_c_160_n N_VGND_c_232_n 0.0101235f $X=0.73 $Y=0.55 $X2=0 $Y2=0
cc_128 N_Y_c_173_n N_VGND_c_234_n 0.0058852f $X=1.68 $Y=0.55 $X2=0 $Y2=0
cc_129 N_Y_M1006_d N_VGND_c_235_n 0.00309031f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_130 N_Y_M1003_d N_VGND_c_235_n 0.00722317f $X=1.545 $Y=0.235 $X2=0 $Y2=0
cc_131 N_Y_c_166_n N_VGND_c_235_n 0.0125677f $X=1.595 $Y=0.74 $X2=0 $Y2=0
cc_132 N_Y_c_160_n N_VGND_c_235_n 0.0102528f $X=0.73 $Y=0.55 $X2=0 $Y2=0
cc_133 N_Y_c_173_n N_VGND_c_235_n 0.00592513f $X=1.68 $Y=0.55 $X2=0 $Y2=0
cc_134 A_117_297# N_VPWR_c_201_n 0.0145335f $X=0.585 $Y=1.485 $X2=0.665 $Y2=0.55
cc_135 A_221_297# N_VPWR_c_201_n 0.00661333f $X=1.105 $Y=1.485 $X2=0 $Y2=0
cc_136 A_317_297# N_VPWR_c_201_n 0.00773468f $X=1.585 $Y=1.485 $X2=0 $Y2=0
