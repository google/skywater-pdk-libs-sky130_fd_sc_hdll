* File: sky130_fd_sc_hdll__a31o_1.pxi.spice
* Created: Wed Sep  2 08:19:53 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31O_1%A_80_21# N_A_80_21#_M1007_d N_A_80_21#_M1009_d
+ N_A_80_21#_c_53_n N_A_80_21#_M1004_g N_A_80_21#_c_54_n N_A_80_21#_M1003_g
+ N_A_80_21#_c_55_n N_A_80_21#_c_65_p N_A_80_21#_c_91_p N_A_80_21#_c_56_n
+ N_A_80_21#_c_57_n N_A_80_21#_c_74_p N_A_80_21#_c_61_n N_A_80_21#_c_58_n
+ PM_SKY130_FD_SC_HDLL__A31O_1%A_80_21#
x_PM_SKY130_FD_SC_HDLL__A31O_1%A3 N_A3_c_131_n N_A3_M1008_g N_A3_c_132_n
+ N_A3_M1005_g A3 A3 PM_SKY130_FD_SC_HDLL__A31O_1%A3
x_PM_SKY130_FD_SC_HDLL__A31O_1%A2 N_A2_c_163_n N_A2_M1006_g N_A2_c_164_n
+ N_A2_M1001_g A2 A2 PM_SKY130_FD_SC_HDLL__A31O_1%A2
x_PM_SKY130_FD_SC_HDLL__A31O_1%A1 N_A1_c_191_n N_A1_M1007_g N_A1_c_192_n
+ N_A1_M1002_g A1 A1 PM_SKY130_FD_SC_HDLL__A31O_1%A1
x_PM_SKY130_FD_SC_HDLL__A31O_1%B1 N_B1_c_220_n N_B1_M1000_g N_B1_c_221_n
+ N_B1_M1009_g B1 B1 N_B1_c_222_n PM_SKY130_FD_SC_HDLL__A31O_1%B1
x_PM_SKY130_FD_SC_HDLL__A31O_1%X N_X_M1004_s N_X_M1003_s N_X_c_245_n N_X_c_248_n
+ N_X_c_246_n X X X N_X_c_247_n PM_SKY130_FD_SC_HDLL__A31O_1%X
x_PM_SKY130_FD_SC_HDLL__A31O_1%VPWR N_VPWR_M1003_d N_VPWR_M1001_d N_VPWR_c_268_n
+ N_VPWR_c_269_n N_VPWR_c_270_n N_VPWR_c_271_n VPWR N_VPWR_c_272_n
+ N_VPWR_c_267_n N_VPWR_c_274_n VPWR PM_SKY130_FD_SC_HDLL__A31O_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A31O_1%A_225_297# N_A_225_297#_M1005_d
+ N_A_225_297#_M1002_d N_A_225_297#_c_310_n N_A_225_297#_c_312_n
+ N_A_225_297#_c_313_n N_A_225_297#_c_318_n N_A_225_297#_c_330_n
+ PM_SKY130_FD_SC_HDLL__A31O_1%A_225_297#
x_PM_SKY130_FD_SC_HDLL__A31O_1%VGND N_VGND_M1004_d N_VGND_M1000_d N_VGND_c_332_n
+ N_VGND_c_333_n N_VGND_c_334_n VGND N_VGND_c_335_n N_VGND_c_336_n
+ N_VGND_c_337_n N_VGND_c_338_n PM_SKY130_FD_SC_HDLL__A31O_1%VGND
cc_1 VNB N_A_80_21#_c_53_n 0.0203866f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_2 VNB N_A_80_21#_c_54_n 0.0276437f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_3 VNB N_A_80_21#_c_55_n 0.00210988f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.995
cc_4 VNB N_A_80_21#_c_56_n 0.00744674f $X=-0.19 $Y=-0.24 $X2=2.915 $Y2=0.74
cc_5 VNB N_A_80_21#_c_57_n 0.00209372f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=1.16
cc_6 VNB N_A_80_21#_c_58_n 0.0219389f $X=-0.19 $Y=-0.24 $X2=2.92 $Y2=1.825
cc_7 VNB N_A3_c_131_n 0.0183649f $X=-0.19 $Y=-0.24 $X2=2.145 $Y2=0.235
cc_8 VNB N_A3_c_132_n 0.0236497f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB A3 0.00425215f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.995
cc_10 VNB N_A2_c_163_n 0.0184029f $X=-0.19 $Y=-0.24 $X2=2.145 $Y2=0.235
cc_11 VNB N_A2_c_164_n 0.0236506f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB A2 0.00375716f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_13 VNB N_A1_c_191_n 0.0184068f $X=-0.19 $Y=-0.24 $X2=2.145 $Y2=0.235
cc_14 VNB N_A1_c_192_n 0.0234861f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB A1 0.00319932f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_16 VNB N_B1_c_220_n 0.0205907f $X=-0.19 $Y=-0.24 $X2=2.145 $Y2=0.235
cc_17 VNB N_B1_c_221_n 0.0252174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_B1_c_222_n 0.00322872f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.825
cc_19 VNB N_X_c_245_n 0.00638732f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.41
cc_20 VNB N_X_c_246_n 0.0228266f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.995
cc_21 VNB N_X_c_247_n 0.013624f $X=-0.19 $Y=-0.24 $X2=3 $Y2=1.825
cc_22 VNB N_VPWR_c_267_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_332_n 0.00561571f $X=-0.19 $Y=-0.24 $X2=0.475 $Y2=0.56
cc_24 VNB N_VGND_c_333_n 0.0136512f $X=-0.19 $Y=-0.24 $X2=0.5 $Y2=1.985
cc_25 VNB N_VGND_c_334_n 0.0149929f $X=-0.19 $Y=-0.24 $X2=0.73 $Y2=0.825
cc_26 VNB N_VGND_c_335_n 0.0185697f $X=-0.19 $Y=-0.24 $X2=2.915 $Y2=0.74
cc_27 VNB N_VGND_c_336_n 0.047698f $X=-0.19 $Y=-0.24 $X2=3 $Y2=1.825
cc_28 VNB N_VGND_c_337_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_VGND_c_338_n 0.182564f $X=-0.19 $Y=-0.24 $X2=2.92 $Y2=1.91
cc_30 VPB N_A_80_21#_c_54_n 0.0317461f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.41
cc_31 VPB N_A_80_21#_c_57_n 9.47786e-19 $X=-0.19 $Y=1.305 $X2=0.73 $Y2=1.16
cc_32 VPB N_A_80_21#_c_61_n 0.0234927f $X=-0.19 $Y=1.305 $X2=2.92 $Y2=1.91
cc_33 VPB N_A_80_21#_c_58_n 0.0204723f $X=-0.19 $Y=1.305 $X2=2.92 $Y2=1.825
cc_34 VPB N_A3_c_132_n 0.0274738f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB A3 9.55033e-19 $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_36 VPB N_A2_c_164_n 0.0271213f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB A2 0.00109924f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_38 VPB N_A1_c_192_n 0.0262759f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB A1 0.00218187f $X=-0.19 $Y=1.305 $X2=0.475 $Y2=0.56
cc_40 VPB N_B1_c_221_n 0.0311188f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_B1_c_222_n 0.00260753f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.825
cc_42 VPB N_X_c_248_n 0.00638732f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.825
cc_43 VPB N_X_c_246_n 0.0124631f $X=-0.19 $Y=1.305 $X2=0.73 $Y2=0.995
cc_44 VPB X 0.0267831f $X=-0.19 $Y=1.305 $X2=0.815 $Y2=0.74
cc_45 VPB N_VPWR_c_268_n 0.00516823f $X=-0.19 $Y=1.305 $X2=0.5 $Y2=1.985
cc_46 VPB N_VPWR_c_269_n 0.00561441f $X=-0.19 $Y=1.305 $X2=2.915 $Y2=0.74
cc_47 VPB N_VPWR_c_270_n 0.0208481f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_VPWR_c_271_n 0.00631953f $X=-0.19 $Y=1.305 $X2=3 $Y2=0.825
cc_49 VPB N_VPWR_c_272_n 0.035107f $X=-0.19 $Y=1.305 $X2=2.315 $Y2=0.74
cc_50 VPB N_VPWR_c_267_n 0.0459529f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_VPWR_c_274_n 0.0245976f $X=-0.19 $Y=1.305 $X2=2.92 $Y2=1.825
cc_52 N_A_80_21#_c_53_n N_A3_c_131_n 0.0194707f $X=0.475 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_53 N_A_80_21#_c_55_n N_A3_c_131_n 0.00391574f $X=0.73 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_80_21#_c_65_p N_A3_c_131_n 0.0140552f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A_80_21#_c_54_n N_A3_c_132_n 0.0309814f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_56 N_A_80_21#_c_65_p N_A3_c_132_n 0.00107f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_57 N_A_80_21#_c_57_n N_A3_c_132_n 0.00205493f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A_80_21#_c_54_n A3 3.15237e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A_80_21#_c_65_p A3 0.0253647f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_60 N_A_80_21#_c_57_n A3 0.0264036f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A_80_21#_c_54_n A3 8.22415e-19 $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_62 N_A_80_21#_c_65_p N_A2_c_163_n 0.0144433f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_63 N_A_80_21#_c_74_p N_A2_c_163_n 0.00164934f $X=2.34 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_64 N_A_80_21#_c_65_p N_A2_c_164_n 0.00107f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_65 N_A_80_21#_c_65_p A2 0.0211775f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_66 N_A_80_21#_c_65_p N_A1_c_191_n 0.00986875f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_80_21#_c_74_p N_A1_c_191_n 0.00797065f $X=2.34 $Y=0.4 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_80_21#_c_74_p N_A1_c_192_n 0.00257476f $X=2.34 $Y=0.4 $X2=0 $Y2=0
cc_69 N_A_80_21#_c_65_p A1 0.010296f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_70 N_A_80_21#_c_74_p A1 0.0100751f $X=2.34 $Y=0.4 $X2=0 $Y2=0
cc_71 N_A_80_21#_c_56_n N_B1_c_220_n 0.0115164f $X=2.915 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_80_21#_c_58_n N_B1_c_220_n 0.00536692f $X=2.92 $Y=1.825 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_80_21#_c_56_n N_B1_c_221_n 0.00415219f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_74 N_A_80_21#_c_61_n N_B1_c_221_n 0.00247342f $X=2.92 $Y=1.91 $X2=0 $Y2=0
cc_75 N_A_80_21#_c_58_n N_B1_c_221_n 0.0161882f $X=2.92 $Y=1.825 $X2=0 $Y2=0
cc_76 N_A_80_21#_c_56_n N_B1_c_222_n 0.0156236f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_77 N_A_80_21#_c_74_p N_B1_c_222_n 0.00365541f $X=2.34 $Y=0.4 $X2=0 $Y2=0
cc_78 N_A_80_21#_c_58_n N_B1_c_222_n 0.0433399f $X=2.92 $Y=1.825 $X2=0 $Y2=0
cc_79 N_A_80_21#_c_53_n N_X_c_245_n 0.00309617f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_80 N_A_80_21#_c_91_p N_X_c_245_n 0.0104924f $X=0.815 $Y=0.74 $X2=0 $Y2=0
cc_81 N_A_80_21#_c_54_n N_X_c_248_n 0.0025655f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_80_21#_c_53_n N_X_c_246_n 0.0137699f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_83 N_A_80_21#_c_54_n N_X_c_246_n 0.00310081f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_84 N_A_80_21#_c_55_n N_X_c_246_n 0.00600714f $X=0.73 $Y=0.995 $X2=0 $Y2=0
cc_85 N_A_80_21#_c_57_n N_X_c_246_n 0.0251475f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_80_21#_c_54_n X 0.00797211f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_80_21#_c_53_n N_X_c_247_n 0.00533946f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_88 N_A_80_21#_c_54_n N_VPWR_c_268_n 0.00474234f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A_80_21#_c_65_p N_VPWR_c_268_n 0.00196487f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_90 N_A_80_21#_c_57_n N_VPWR_c_268_n 0.0142812f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_80_21#_c_61_n N_VPWR_c_272_n 0.0178803f $X=2.92 $Y=1.91 $X2=0 $Y2=0
cc_92 N_A_80_21#_M1009_d N_VPWR_c_267_n 0.00412347f $X=2.715 $Y=1.485 $X2=0
+ $Y2=0
cc_93 N_A_80_21#_c_54_n N_VPWR_c_267_n 0.0131053f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A_80_21#_c_61_n N_VPWR_c_267_n 0.0123599f $X=2.92 $Y=1.91 $X2=0 $Y2=0
cc_95 N_A_80_21#_c_54_n N_VPWR_c_274_n 0.00681977f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A_80_21#_c_55_n N_VGND_M1004_d 0.00132169f $X=0.73 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_97 N_A_80_21#_c_65_p N_VGND_M1004_d 0.00194381f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_98 N_A_80_21#_c_91_p N_VGND_M1004_d 0.00439798f $X=0.815 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_99 N_A_80_21#_c_56_n N_VGND_M1000_d 0.00889881f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_100 N_A_80_21#_c_58_n N_VGND_M1000_d 0.00111605f $X=2.92 $Y=1.825 $X2=0 $Y2=0
cc_101 N_A_80_21#_c_53_n N_VGND_c_332_n 0.0043941f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_102 N_A_80_21#_c_54_n N_VGND_c_332_n 0.0010263f $X=0.5 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A_80_21#_c_65_p N_VGND_c_332_n 0.0048033f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_104 N_A_80_21#_c_91_p N_VGND_c_332_n 0.013745f $X=0.815 $Y=0.74 $X2=0 $Y2=0
cc_105 N_A_80_21#_c_57_n N_VGND_c_332_n 0.00136623f $X=0.73 $Y=1.16 $X2=0 $Y2=0
cc_106 N_A_80_21#_c_56_n N_VGND_c_333_n 5.86325e-19 $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_107 N_A_80_21#_c_56_n N_VGND_c_334_n 0.0258324f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_108 N_A_80_21#_c_53_n N_VGND_c_335_n 0.0055043f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_80_21#_c_65_p N_VGND_c_336_n 0.0177415f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_110 N_A_80_21#_c_56_n N_VGND_c_336_n 0.0029785f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_111 N_A_80_21#_c_74_p N_VGND_c_336_n 0.0165402f $X=2.34 $Y=0.4 $X2=0 $Y2=0
cc_112 N_A_80_21#_M1007_d N_VGND_c_338_n 0.00316154f $X=2.145 $Y=0.235 $X2=0
+ $Y2=0
cc_113 N_A_80_21#_c_53_n N_VGND_c_338_n 0.0110311f $X=0.475 $Y=0.995 $X2=0 $Y2=0
cc_114 N_A_80_21#_c_65_p N_VGND_c_338_n 0.0315558f $X=2.125 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_80_21#_c_91_p N_VGND_c_338_n 7.75073e-19 $X=0.815 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_80_21#_c_56_n N_VGND_c_338_n 0.00775267f $X=2.915 $Y=0.74 $X2=0 $Y2=0
cc_117 N_A_80_21#_c_74_p N_VGND_c_338_n 0.013831f $X=2.34 $Y=0.4 $X2=0 $Y2=0
cc_118 N_A_80_21#_c_65_p A_217_47# 0.00939126f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_80_21#_c_65_p A_323_47# 0.0109052f $X=2.125 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A3_c_131_n N_A2_c_163_n 0.0304877f $X=1.01 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_121 N_A3_c_132_n N_A2_c_164_n 0.0393549f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_122 A3 N_A2_c_164_n 0.00268102f $X=1.08 $Y=1.105 $X2=0 $Y2=0
cc_123 A3 N_A2_c_164_n 0.00176313f $X=1.09 $Y=1.445 $X2=0 $Y2=0
cc_124 N_A3_c_132_n A2 6.13446e-19 $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_125 A3 A2 0.050139f $X=1.08 $Y=1.105 $X2=0 $Y2=0
cc_126 N_A3_c_131_n N_X_c_247_n 5.67792e-19 $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A3_c_132_n N_VPWR_c_268_n 0.00293354f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A3_c_132_n N_VPWR_c_270_n 0.00645921f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A3_c_132_n N_VPWR_c_267_n 0.0114644f $X=1.035 $Y=1.41 $X2=0 $Y2=0
cc_130 A3 N_A_225_297#_M1005_d 0.00337293f $X=1.09 $Y=1.445 $X2=-0.19 $Y2=-0.24
cc_131 N_A3_c_132_n N_A_225_297#_c_310_n 0.00306579f $X=1.035 $Y=1.41 $X2=0
+ $Y2=0
cc_132 A3 N_A_225_297#_c_310_n 0.0172783f $X=1.09 $Y=1.445 $X2=0 $Y2=0
cc_133 N_A3_c_132_n N_A_225_297#_c_312_n 0.00564404f $X=1.035 $Y=1.41 $X2=0
+ $Y2=0
cc_134 N_A3_c_131_n N_VGND_c_332_n 0.00331705f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_135 N_A3_c_131_n N_VGND_c_336_n 0.00427293f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_136 N_A3_c_131_n N_VGND_c_338_n 0.00619412f $X=1.01 $Y=0.995 $X2=0 $Y2=0
cc_137 N_A2_c_163_n N_A1_c_191_n 0.0306517f $X=1.54 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_138 N_A2_c_164_n N_A1_c_192_n 0.0539674f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_139 A2 N_A1_c_192_n 0.00219945f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_140 N_A2_c_164_n A1 0.00150387f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_141 A2 A1 0.0467821f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_142 A2 N_VPWR_M1001_d 0.00258844f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_143 N_A2_c_164_n N_VPWR_c_269_n 0.00348239f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_164_n N_VPWR_c_270_n 0.00525423f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A2_c_164_n N_VPWR_c_267_n 0.00721835f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A2_c_164_n N_A_225_297#_c_313_n 0.0137409f $X=1.565 $Y=1.41 $X2=0 $Y2=0
cc_147 A2 N_A_225_297#_c_313_n 0.0188402f $X=1.55 $Y=1.105 $X2=0 $Y2=0
cc_148 N_A2_c_163_n N_VGND_c_336_n 0.00428022f $X=1.54 $Y=0.995 $X2=0 $Y2=0
cc_149 N_A2_c_163_n N_VGND_c_338_n 0.00649419f $X=1.54 $Y=0.995 $X2=0 $Y2=0
cc_150 N_A1_c_191_n N_B1_c_220_n 0.0088298f $X=2.07 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_151 N_A1_c_192_n N_B1_c_221_n 0.0409709f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_152 A1 N_B1_c_221_n 0.001298f $X=2.025 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A1_c_192_n N_B1_c_222_n 0.00296094f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_154 A1 N_B1_c_222_n 0.05218f $X=2.025 $Y=1.105 $X2=0 $Y2=0
cc_155 N_A1_c_192_n N_VPWR_c_269_n 0.00348239f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_156 N_A1_c_192_n N_VPWR_c_272_n 0.00525423f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_157 N_A1_c_192_n N_VPWR_c_267_n 0.00721835f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_158 A1 N_A_225_297#_M1002_d 0.00185056f $X=2.025 $Y=1.105 $X2=0 $Y2=0
cc_159 N_A1_c_192_n N_A_225_297#_c_313_n 0.0123755f $X=2.095 $Y=1.41 $X2=0 $Y2=0
cc_160 A1 N_A_225_297#_c_313_n 0.0162403f $X=2.025 $Y=1.105 $X2=0 $Y2=0
cc_161 N_A1_c_192_n N_A_225_297#_c_318_n 0.00122796f $X=2.095 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_A1_c_191_n N_VGND_c_336_n 0.00421711f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A1_c_191_n N_VGND_c_338_n 0.00635084f $X=2.07 $Y=0.995 $X2=0 $Y2=0
cc_164 N_B1_c_221_n N_VPWR_c_272_n 0.00702461f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B1_c_221_n N_VPWR_c_267_n 0.0139604f $X=2.625 $Y=1.41 $X2=0 $Y2=0
cc_166 N_B1_c_222_n N_A_225_297#_M1002_d 0.00185125f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_167 N_B1_c_222_n N_A_225_297#_c_318_n 0.00284875f $X=2.66 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B1_c_220_n N_VGND_c_334_n 0.00937902f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_169 N_B1_c_220_n N_VGND_c_336_n 0.00428022f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B1_c_220_n N_VGND_c_338_n 0.00714441f $X=2.6 $Y=0.995 $X2=0 $Y2=0
cc_171 N_X_M1003_s N_VPWR_c_267_n 0.00223991f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_172 X N_VPWR_c_267_n 0.0122458f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_173 X N_VPWR_c_274_n 0.0167868f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_174 N_X_c_247_n N_VGND_c_335_n 0.0162614f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_175 N_X_M1004_s N_VGND_c_338_n 0.00216172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_176 N_X_c_247_n N_VGND_c_338_n 0.012122f $X=0.26 $Y=0.385 $X2=0 $Y2=0
cc_177 N_VPWR_c_267_n N_A_225_297#_M1005_d 0.00328183f $X=2.99 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_178 N_VPWR_c_267_n N_A_225_297#_M1002_d 0.00366235f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_179 N_VPWR_c_270_n N_A_225_297#_c_312_n 0.0141504f $X=1.665 $Y=2.72 $X2=0
+ $Y2=0
cc_180 N_VPWR_c_267_n N_A_225_297#_c_312_n 0.0109465f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_181 N_VPWR_M1001_d N_A_225_297#_c_313_n 0.00855869f $X=1.655 $Y=1.485 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_269_n N_A_225_297#_c_313_n 0.0184724f $X=1.83 $Y=2.25 $X2=0
+ $Y2=0
cc_183 N_VPWR_c_270_n N_A_225_297#_c_313_n 0.0033873f $X=1.665 $Y=2.72 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_272_n N_A_225_297#_c_313_n 0.0033873f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_267_n N_A_225_297#_c_313_n 0.0142139f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_272_n N_A_225_297#_c_330_n 0.0118939f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_267_n N_A_225_297#_c_330_n 0.00927173f $X=2.99 $Y=2.72 $X2=0
+ $Y2=0
cc_188 N_VGND_c_338_n A_217_47# 0.00454783f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
cc_189 N_VGND_c_338_n A_323_47# 0.00454783f $X=2.99 $Y=0 $X2=-0.19 $Y2=-0.24
