* File: sky130_fd_sc_hdll__sdfstp_4.pex.spice
* Created: Thu Aug 27 19:27:27 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCD 1 2 3 5 6 8 13 14
c33 3 0 3.49297e-20 $X=0.495 $Y=1.77
r34 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.255
+ $Y=1.16 $X2=0.255 $Y2=1.16
r35 14 19 16.7217 $w=2.53e-07 $l=3.7e-07 $layer=LI1_cond $X=0.212 $Y=1.53
+ $X2=0.212 $Y2=1.16
r36 13 19 14.0101 $w=2.53e-07 $l=3.1e-07 $layer=LI1_cond $X=0.212 $Y=0.85
+ $X2=0.212 $Y2=1.16
r37 6 18 85.0704 $w=2.76e-07 $l=5.07937e-07 $layer=POLY_cond $X=0.52 $Y=0.73
+ $X2=0.35 $Y2=1.16
r38 6 8 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r39 3 9 92.2979 $w=1.5e-07 $l=1.8e-07 $layer=POLY_cond $X=0.495 $Y=1.695
+ $X2=0.315 $Y2=1.695
r40 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.77
+ $X2=0.495 $Y2=2.165
r41 2 9 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.315 $Y=1.62
+ $X2=0.315 $Y2=1.695
r42 1 18 38.7914 $w=2.76e-07 $l=1.81659e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.35 $Y2=1.16
r43 1 2 151.266 $w=1.5e-07 $l=2.95e-07 $layer=POLY_cond $X=0.315 $Y=1.325
+ $X2=0.315 $Y2=1.62
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%SCE 3 6 7 9 11 12 14 17 19 20 22 25 30 33
+ 34 38 46
c110 30 0 4.39648e-20 $X=0.93 $Y=1.25
c111 22 0 1.07953e-19 $X=2.73 $Y=1.19
c112 7 0 1.40323e-19 $X=0.965 $Y=1.77
r113 33 36 37.7919 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=1.325
r114 33 35 46.6671 $w=3.65e-07 $l=1.65e-07 $layer=POLY_cond $X=2.782 $Y=1.16
+ $X2=2.782 $Y2=0.995
r115 33 34 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.735
+ $Y=1.16 $X2=2.735 $Y2=1.16
r116 30 31 5.56766 $w=3.03e-07 $l=3.5e-08 $layer=POLY_cond $X=0.93 $Y=1.25
+ $X2=0.965 $Y2=1.25
r117 28 30 23.066 $w=3.03e-07 $l=1.45e-07 $layer=POLY_cond $X=0.785 $Y=1.25
+ $X2=0.93 $Y2=1.25
r118 28 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.785
+ $Y=1.25 $X2=0.785 $Y2=1.25
r119 25 46 0.0320802 $w=2.3e-07 $l=5e-08 $layer=MET1_cond $X=0.69 $Y=1.19
+ $X2=0.64 $Y2=1.19
r120 25 38 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.725 $Y=1.19
+ $X2=0.725 $Y2=1.19
r121 22 34 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.73 $Y=1.19
+ $X2=2.73 $Y2=1.19
r122 20 25 0.137923 $w=2.3e-07 $l=1.8e-07 $layer=MET1_cond $X=0.87 $Y=1.19
+ $X2=0.69 $Y2=1.19
r123 19 22 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=2.73 $Y2=1.19
r124 19 20 2.12252 $w=1.4e-07 $l=1.715e-06 $layer=MET1_cond $X=2.585 $Y=1.19
+ $X2=0.87 $Y2=1.19
r125 17 35 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=2.89 $Y=0.445
+ $X2=2.89 $Y2=0.995
r126 12 14 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.835 $Y=1.77
+ $X2=2.835 $Y2=2.165
r127 11 12 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.835 $Y=1.67 $X2=2.835
+ $Y2=1.77
r128 11 36 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=2.835 $Y=1.67
+ $X2=2.835 $Y2=1.325
r129 7 9 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.77
+ $X2=0.965 $Y2=2.165
r130 6 7 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.965 $Y=1.67 $X2=0.965
+ $Y2=1.77
r131 5 31 12.5184 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=0.965 $Y=1.415
+ $X2=0.965 $Y2=1.25
r132 5 6 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=0.965 $Y=1.415
+ $X2=0.965 $Y2=1.67
r133 1 30 19.2026 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.93 $Y=1.085
+ $X2=0.93 $Y2=1.25
r134 1 3 328.17 $w=1.5e-07 $l=6.4e-07 $layer=POLY_cond $X=0.93 $Y=1.085 $X2=0.93
+ $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%D 2 3 5 8 9 10 14 16
c49 9 0 3.49297e-20 $X=1.15 $Y=0.85
r50 14 16 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=0.93
+ $X2=1.375 $Y2=0.765
r51 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.35
+ $Y=0.93 $X2=1.35 $Y2=0.93
r52 10 15 15.5386 $w=4.43e-07 $l=6e-07 $layer=LI1_cond $X=1.262 $Y=1.53
+ $X2=1.262 $Y2=0.93
r53 9 15 2.07181 $w=4.43e-07 $l=8e-08 $layer=LI1_cond $X=1.262 $Y=0.85 $X2=1.262
+ $Y2=0.93
r54 8 16 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.4 $Y=0.445 $X2=1.4
+ $Y2=0.765
r55 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.375 $Y=1.77
+ $X2=1.375 $Y2=2.165
r56 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.375 $Y=1.67 $X2=1.375
+ $Y2=1.77
r57 1 14 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.375 $Y=1.095
+ $X2=1.375 $Y2=0.93
r58 1 2 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=1.375 $Y=1.095
+ $X2=1.375 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_349_21# 1 2 9 12 13 15 17 21 22 23 25
+ 35 37
c79 22 0 1.4475e-19 $X=2.15 $Y=1.16
r80 35 37 0.182927 $w=3.13e-07 $l=5e-09 $layer=LI1_cond $X=2.595 $Y=1.927
+ $X2=2.6 $Y2=1.927
r81 23 25 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=2.59 $Y=0.715
+ $X2=2.59 $Y2=0.44
r82 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.15
+ $Y=1.16 $X2=2.15 $Y2=1.16
r83 19 35 13.2805 $w=3.13e-07 $l=3.63e-07 $layer=LI1_cond $X=2.232 $Y=1.927
+ $X2=2.595 $Y2=1.927
r84 19 21 20.9848 $w=3.33e-07 $l=6.1e-07 $layer=LI1_cond $X=2.232 $Y=1.77
+ $X2=2.232 $Y2=1.16
r85 18 23 20.8976 $w=1.88e-07 $l=3.58e-07 $layer=LI1_cond $X=2.232 $Y=0.81
+ $X2=2.59 $Y2=0.81
r86 18 21 8.77233 $w=3.33e-07 $l=2.55e-07 $layer=LI1_cond $X=2.232 $Y=0.905
+ $X2=2.232 $Y2=1.16
r87 16 22 35.8466 $w=3.3e-07 $l=2.05e-07 $layer=POLY_cond $X=1.945 $Y=1.16
+ $X2=2.15 $Y2=1.16
r88 16 17 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.945 $Y=1.16
+ $X2=1.845 $Y2=1.16
r89 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.845 $Y=1.77
+ $X2=1.845 $Y2=2.165
r90 12 13 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.845 $Y=1.67 $X2=1.845
+ $Y2=1.77
r91 11 17 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.16
r92 11 12 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.845 $Y=1.325
+ $X2=1.845 $Y2=1.67
r93 7 17 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.82 $Y=0.995
+ $X2=1.845 $Y2=1.16
r94 7 9 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.82 $Y=0.995 $X2=1.82
+ $Y2=0.445
r95 2 37 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=2.475
+ $Y=1.845 $X2=2.6 $Y2=1.99
r96 1 25 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=2.505
+ $Y=0.235 $X2=2.63 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%CLK 7 8 10 13 15 16 17 20 21 22
c58 21 0 3.28604e-20 $X=3.68 $Y=1.255
c59 13 0 1.06712e-19 $X=3.88 $Y=0.805
r60 20 23 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.42
r61 20 22 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=3.68 $Y=1.255
+ $X2=3.68 $Y2=1.09
r62 20 21 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.68
+ $Y=1.255 $X2=3.68 $Y2=1.255
r63 17 21 4.6235 $w=5.93e-07 $l=2.3e-07 $layer=LI1_cond $X=3.45 $Y=1.352
+ $X2=3.68 $Y2=1.352
r64 15 16 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=3.795 $Y=1.62
+ $X2=3.795 $Y2=1.77
r65 15 23 102.553 $w=1.5e-07 $l=2e-07 $layer=POLY_cond $X=3.74 $Y=1.62 $X2=3.74
+ $Y2=1.42
r66 11 13 71.7872 $w=1.5e-07 $l=1.4e-07 $layer=POLY_cond $X=3.74 $Y=0.805
+ $X2=3.88 $Y2=0.805
r67 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.805
r68 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=3.88 $Y=0.73 $X2=3.88
+ $Y2=0.445
r69 7 16 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=3.825 $Y=2.165
+ $X2=3.825 $Y2=1.77
r70 1 11 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=0.805
r71 1 22 107.681 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=3.74 $Y=0.88 $X2=3.74
+ $Y2=1.09
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_693_369# 1 2 8 9 11 14 16 17 19 21 22
+ 24 26 27 29 32 34 37 41 43 44 45 46 48 50 51 55 56 57 58 61 64 65 66 67 68 77
+ 81 85 91
c285 91 0 6.70306e-20 $X=9.9 $Y=1.09
c286 85 0 1.8066e-19 $X=5.73 $Y=1.74
c287 81 0 3.28604e-20 $X=4.235 $Y=1.09
c288 77 0 2.08915e-19 $X=8.295 $Y=1.87
c289 67 0 1.36329e-19 $X=8.15 $Y=1.87
c290 61 0 1.97973e-19 $X=9.79 $Y=1.09
c291 34 0 6.74919e-20 $X=4.317 $Y=0.805
r292 84 85 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.74 $X2=5.73 $Y2=1.74
r293 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=8.295 $Y=1.87
+ $X2=8.295 $Y2=1.87
r294 74 85 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.69 $Y=1.87
+ $X2=5.69 $Y2=1.87
r295 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.21 $Y=1.87
+ $X2=4.21 $Y2=1.87
r296 68 74 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=5.885 $Y=1.87
+ $X2=5.69 $Y2=1.87
r297 67 77 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=8.15 $Y=1.87
+ $X2=8.295 $Y2=1.87
r298 67 68 2.80321 $w=1.4e-07 $l=2.265e-06 $layer=MET1_cond $X=8.15 $Y=1.87
+ $X2=5.885 $Y2=1.87
r299 66 70 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=4.405 $Y=1.87
+ $X2=4.21 $Y2=1.87
r300 65 74 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=5.69 $Y2=1.87
r301 65 66 1.41089 $w=1.4e-07 $l=1.14e-06 $layer=MET1_cond $X=5.545 $Y=1.87
+ $X2=4.405 $Y2=1.87
r302 64 78 11.7266 $w=2.83e-07 $l=2.9e-07 $layer=LI1_cond $X=8.585 $Y=1.812
+ $X2=8.295 $Y2=1.812
r303 62 91 19.2347 $w=3.3e-07 $l=1.1e-07 $layer=POLY_cond $X=9.79 $Y=1.09
+ $X2=9.9 $Y2=1.09
r304 61 62 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.79
+ $Y=1.09 $X2=9.79 $Y2=1.09
r305 59 61 6.36424 $w=3.33e-07 $l=1.85e-07 $layer=LI1_cond $X=9.837 $Y=0.905
+ $X2=9.837 $Y2=1.09
r306 57 59 7.58144 $w=1.85e-07 $l=2.08375e-07 $layer=LI1_cond $X=9.67 $Y=0.812
+ $X2=9.837 $Y2=0.905
r307 57 58 47.0614 $w=1.83e-07 $l=7.85e-07 $layer=LI1_cond $X=9.67 $Y=0.812
+ $X2=8.885 $Y2=0.812
r308 56 88 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=8.695 $Y=1.16
+ $X2=8.695 $Y2=1.325
r309 55 56 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.67
+ $Y=1.16 $X2=8.67 $Y2=1.16
r310 53 64 6.82232 $w=2.85e-07 $l=2.09285e-07 $layer=LI1_cond $X=8.735 $Y=1.67
+ $X2=8.585 $Y2=1.812
r311 53 55 19.5915 $w=2.98e-07 $l=5.1e-07 $layer=LI1_cond $X=8.735 $Y=1.67
+ $X2=8.735 $Y2=1.16
r312 52 58 7.32714 $w=1.85e-07 $l=1.90919e-07 $layer=LI1_cond $X=8.735 $Y=0.905
+ $X2=8.885 $Y2=0.812
r313 52 55 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=8.735 $Y=0.905
+ $X2=8.735 $Y2=1.16
r314 51 82 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.42
r315 51 81 39.9376 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=4.235 $Y=1.255
+ $X2=4.235 $Y2=1.09
r316 50 51 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.21
+ $Y=1.255 $X2=4.21 $Y2=1.255
r317 48 71 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=4.165 $Y=1.83
+ $X2=4.165 $Y2=1.915
r318 48 50 25.4867 $w=2.58e-07 $l=5.75e-07 $layer=LI1_cond $X=4.165 $Y=1.83
+ $X2=4.165 $Y2=1.255
r319 47 50 16.4002 $w=2.58e-07 $l=3.7e-07 $layer=LI1_cond $X=4.165 $Y=0.885
+ $X2=4.165 $Y2=1.255
r320 45 47 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=4.165 $Y2=0.885
r321 45 46 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=4.035 $Y=0.8
+ $X2=3.705 $Y2=0.8
r322 43 71 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=4.035 $Y=1.915
+ $X2=4.165 $Y2=1.915
r323 43 44 23.4866 $w=1.68e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=1.915
+ $X2=3.675 $Y2=1.915
r324 39 46 6.83233 $w=1.7e-07 $l=1.28662e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.705 $Y2=0.8
r325 39 41 16.4865 $w=1.83e-07 $l=2.75e-07 $layer=LI1_cond $X=3.612 $Y=0.715
+ $X2=3.612 $Y2=0.44
r326 35 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=3.59 $Y=2
+ $X2=3.675 $Y2=1.915
r327 35 37 10.4385 $w=1.68e-07 $l=1.6e-07 $layer=LI1_cond $X=3.59 $Y=2 $X2=3.59
+ $Y2=2.16
r328 30 91 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=9.9 $Y=0.925
+ $X2=9.9 $Y2=1.09
r329 30 32 246.128 $w=1.5e-07 $l=4.8e-07 $layer=POLY_cond $X=9.9 $Y=0.925
+ $X2=9.9 $Y2=0.445
r330 27 29 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.635 $Y=1.57
+ $X2=8.635 $Y2=2.065
r331 26 27 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.635 $Y=1.47 $X2=8.635
+ $Y2=1.57
r332 26 88 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.635 $Y=1.47
+ $X2=8.635 $Y2=1.325
r333 22 84 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=1.74
r334 22 24 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.755 $Y=1.99
+ $X2=5.755 $Y2=2.275
r335 19 21 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=5.34 $Y=0.73
+ $X2=5.34 $Y2=0.445
r336 18 34 6.88539 $w=1.5e-07 $l=1.08e-07 $layer=POLY_cond $X=4.425 $Y=0.805
+ $X2=4.317 $Y2=0.805
r337 17 19 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=5.34 $Y2=0.73
r338 17 18 430.723 $w=1.5e-07 $l=8.4e-07 $layer=POLY_cond $X=5.265 $Y=0.805
+ $X2=4.425 $Y2=0.805
r339 14 34 18.6014 $w=1.67e-07 $l=9e-08 $layer=POLY_cond $X=4.35 $Y=0.73
+ $X2=4.317 $Y2=0.805
r340 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=4.35 $Y=0.73
+ $X2=4.35 $Y2=0.445
r341 12 34 18.6014 $w=1.67e-07 $l=8.21584e-08 $layer=POLY_cond $X=4.302 $Y=0.88
+ $X2=4.317 $Y2=0.805
r342 12 81 77.5789 $w=1.85e-07 $l=2.1e-07 $layer=POLY_cond $X=4.302 $Y=0.88
+ $X2=4.302 $Y2=1.09
r343 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=4.295 $Y=1.77
+ $X2=4.295 $Y2=2.165
r344 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=4.295 $Y=1.67 $X2=4.295
+ $Y2=1.77
r345 8 82 82.8943 $w=2e-07 $l=2.5e-07 $layer=POLY_cond $X=4.295 $Y=1.67
+ $X2=4.295 $Y2=1.42
r346 2 37 600 $w=1.7e-07 $l=3.7229e-07 $layer=licon1_PDIFF $count=1 $X=3.465
+ $Y=1.845 $X2=3.59 $Y2=2.16
r347 1 41 182 $w=1.7e-07 $l=2.60096e-07 $layer=licon1_NDIFF $count=1 $X=3.495
+ $Y=0.235 $X2=3.62 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_877_369# 1 2 8 9 11 12 13 15 18 22 24
+ 26 29 34 35 37 39 41 42 46 48 54
c183 46 0 1.33492e-19 $X=4.72 $Y=1.185
c184 42 0 9.8756e-21 $X=9.365 $Y=1.19
c185 29 0 7.95993e-20 $X=4.56 $Y=0.42
c186 18 0 1.00357e-19 $X=5.81 $Y=0.445
c187 11 0 2.89743e-19 $X=5.195 $Y=1.915
c188 9 0 1.70908e-19 $X=5.735 $Y=1.165
c189 8 0 1.8066e-19 $X=4.965 $Y=1.84
r190 56 57 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=9.36
+ $Y=1.74 $X2=9.36 $Y2=1.74
r191 53 54 30.474 $w=3.3e-07 $l=7.5e-08 $layer=POLY_cond $X=4.965 $Y=1.255
+ $X2=5.04 $Y2=1.255
r192 50 53 36.7209 $w=3.3e-07 $l=2.1e-07 $layer=POLY_cond $X=4.755 $Y=1.255
+ $X2=4.965 $Y2=1.255
r193 46 64 7.6678 $w=3.63e-07 $l=2.35e-07 $layer=LI1_cond $X=4.657 $Y=1.185
+ $X2=4.657 $Y2=1.42
r194 46 63 5.21818 $w=3.63e-07 $l=1e-07 $layer=LI1_cond $X=4.657 $Y=1.185
+ $X2=4.657 $Y2=1.085
r195 46 50 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.755
+ $Y=1.255 $X2=4.755 $Y2=1.255
r196 45 48 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.72 $Y=1.185
+ $X2=4.865 $Y2=1.185
r197 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.72 $Y=1.185
+ $X2=4.72 $Y2=1.185
r198 42 57 19.5029 $w=3.23e-07 $l=5.5e-07 $layer=LI1_cond $X=9.337 $Y=1.19
+ $X2=9.337 $Y2=1.74
r199 41 42 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.365 $Y=1.19
+ $X2=9.365 $Y2=1.19
r200 39 41 0.0513283 $w=2.3e-07 $l=8e-08 $layer=MET1_cond $X=9.285 $Y=1.19
+ $X2=9.365 $Y2=1.19
r201 37 39 0.0850015 $w=2.3e-07 $l=1.15e-07 $layer=MET1_cond $X=9.17 $Y=1.19
+ $X2=9.285 $Y2=1.19
r202 37 48 5.32796 $w=1.4e-07 $l=4.305e-06 $layer=MET1_cond $X=9.17 $Y=1.19
+ $X2=4.865 $Y2=1.19
r203 35 64 26.1586 $w=3.13e-07 $l=7.15e-07 $layer=LI1_cond $X=4.632 $Y=2.135
+ $X2=4.632 $Y2=1.42
r204 34 35 5.62076 $w=3.43e-07 $l=1.65e-07 $layer=LI1_cond $X=4.617 $Y=2.3
+ $X2=4.617 $Y2=2.135
r205 29 63 35.1212 $w=2.08e-07 $l=6.65e-07 $layer=LI1_cond $X=4.58 $Y=0.42
+ $X2=4.58 $Y2=1.085
r206 24 56 45.2339 $w=3.74e-07 $l=2.78388e-07 $layer=POLY_cond $X=9.365 $Y=1.99
+ $X2=9.305 $Y2=1.74
r207 24 26 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.365 $Y=1.99
+ $X2=9.365 $Y2=2.275
r208 20 56 39.1188 $w=3.74e-07 $l=2.33345e-07 $layer=POLY_cond $X=9.14 $Y=1.575
+ $X2=9.305 $Y2=1.74
r209 20 22 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=9.14 $Y=1.575
+ $X2=9.14 $Y2=0.555
r210 16 18 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=5.81 $Y=1.09
+ $X2=5.81 $Y2=0.445
r211 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=5.285 $Y=1.99
+ $X2=5.285 $Y2=2.275
r212 11 13 27.2212 $w=1.5e-07 $l=1.21861e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.285 $Y2=1.99
r213 11 12 79.4787 $w=1.5e-07 $l=1.55e-07 $layer=POLY_cond $X=5.195 $Y=1.915
+ $X2=5.04 $Y2=1.915
r214 9 16 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.81 $Y2=1.09
r215 9 54 356.372 $w=1.5e-07 $l=6.95e-07 $layer=POLY_cond $X=5.735 $Y=1.165
+ $X2=5.04 $Y2=1.165
r216 8 12 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=4.965 $Y=1.84
+ $X2=5.04 $Y2=1.915
r217 7 53 21.2229 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.255
r218 7 8 215.362 $w=1.5e-07 $l=4.2e-07 $layer=POLY_cond $X=4.965 $Y=1.42
+ $X2=4.965 $Y2=1.84
r219 2 34 600 $w=1.7e-07 $l=5.22494e-07 $layer=licon1_PDIFF $count=1 $X=4.385
+ $Y=1.845 $X2=4.53 $Y2=2.3
r220 1 29 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=4.425
+ $Y=0.235 $X2=4.56 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1229_21# 1 2 9 12 13 15 18 21 23 24 27
+ 31 33 37
c95 33 0 4.30126e-20 $X=6.285 $Y=0.72
c96 23 0 3.13156e-20 $X=7.155 $Y=2.02
c97 21 0 3.91586e-20 $X=6.785 $Y=0.72
r98 37 41 32.4954 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.31 $Y=0.93
+ $X2=6.31 $Y2=1.065
r99 37 40 40.9657 $w=3.3e-07 $l=1.35e-07 $layer=POLY_cond $X=6.31 $Y=0.93
+ $X2=6.31 $Y2=0.795
r100 36 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.31
+ $Y=0.93 $X2=6.31 $Y2=0.93
r101 33 36 6.36876 $w=3.78e-07 $l=2.1e-07 $layer=LI1_cond $X=6.285 $Y=0.72
+ $X2=6.285 $Y2=0.93
r102 29 31 7.82791 $w=2.63e-07 $l=1.8e-07 $layer=LI1_cond $X=7.287 $Y=2.105
+ $X2=7.287 $Y2=2.285
r103 25 27 5.76222 $w=2.48e-07 $l=1.25e-07 $layer=LI1_cond $X=6.91 $Y=0.635
+ $X2=6.91 $Y2=0.51
r104 23 29 7.24806 $w=1.7e-07 $l=1.69245e-07 $layer=LI1_cond $X=7.155 $Y=2.02
+ $X2=7.287 $Y2=2.105
r105 23 24 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.155 $Y=2.02
+ $X2=6.595 $Y2=2.02
r106 22 33 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.475 $Y=0.72
+ $X2=6.285 $Y2=0.72
r107 21 25 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=6.785 $Y=0.72
+ $X2=6.91 $Y2=0.635
r108 21 22 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.785 $Y=0.72
+ $X2=6.475 $Y2=0.72
r109 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.51
+ $Y=1.74 $X2=6.51 $Y2=1.74
r110 16 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.595 $Y2=2.02
r111 16 18 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=6.51 $Y=1.935
+ $X2=6.51 $Y2=1.74
r112 13 19 45.1054 $w=3.82e-07 $l=3.02076e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.43 $Y2=1.74
r113 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=6.315 $Y=1.99
+ $X2=6.315 $Y2=2.275
r114 12 19 31.7097 $w=3.82e-07 $l=2.14942e-07 $layer=POLY_cond $X=6.315 $Y=1.575
+ $X2=6.43 $Y2=1.74
r115 12 41 169.104 $w=2e-07 $l=5.1e-07 $layer=POLY_cond $X=6.315 $Y=1.575
+ $X2=6.315 $Y2=1.065
r116 9 40 179.468 $w=1.5e-07 $l=3.5e-07 $layer=POLY_cond $X=6.22 $Y=0.445
+ $X2=6.22 $Y2=0.795
r117 2 31 600 $w=1.7e-07 $l=2.92916e-07 $layer=licon1_PDIFF $count=1 $X=7.095
+ $Y=2.065 $X2=7.265 $Y2=2.285
r118 1 27 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=6.825
+ $Y=0.235 $X2=6.95 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1075_413# 1 2 8 10 11 13 14 16 19 21 22
+ 24 27 29 35 38 40 41 49 50 53 56 59
c154 8 0 4.30126e-20 $X=7.005 $Y=1.095
r155 53 60 37.8338 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.14 $Y=1.16
+ $X2=8.14 $Y2=1.325
r156 53 59 46.7569 $w=3.7e-07 $l=1.65e-07 $layer=POLY_cond $X=8.14 $Y=1.16
+ $X2=8.14 $Y2=0.995
r157 52 53 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=8.09
+ $Y=1.16 $X2=8.09 $Y2=1.16
r158 48 56 25.55 $w=2.7e-07 $l=1.15e-07 $layer=POLY_cond $X=6.89 $Y=1.23
+ $X2=7.005 $Y2=1.23
r159 47 50 3.29018 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.185
+ $X2=6.975 $Y2=1.185
r160 47 49 6.54147 $w=4.18e-07 $l=8.5e-08 $layer=LI1_cond $X=6.89 $Y=1.185
+ $X2=6.805 $Y2=1.185
r161 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.89
+ $Y=1.23 $X2=6.89 $Y2=1.23
r162 41 52 3.24611 $w=3.5e-07 $l=8.5e-08 $layer=LI1_cond $X=8.005 $Y=1.125
+ $X2=8.09 $Y2=1.125
r163 41 50 39.5672 $w=2.98e-07 $l=1.03e-06 $layer=LI1_cond $X=8.005 $Y=1.125
+ $X2=6.975 $Y2=1.125
r164 40 45 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=6.12 $Y2=1.31
r165 40 49 39.1444 $w=1.68e-07 $l=6e-07 $layer=LI1_cond $X=6.205 $Y=1.31
+ $X2=6.805 $Y2=1.31
r166 37 45 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=6.12 $Y2=1.31
r167 37 38 48.2781 $w=1.68e-07 $l=7.4e-07 $layer=LI1_cond $X=6.12 $Y=1.395
+ $X2=6.12 $Y2=2.135
r168 33 45 28.9016 $w=1.68e-07 $l=4.43e-07 $layer=LI1_cond $X=5.677 $Y=1.31
+ $X2=6.12 $Y2=1.31
r169 33 35 21.8286 $w=4.23e-07 $l=8.05e-07 $layer=LI1_cond $X=5.677 $Y=1.225
+ $X2=5.677 $Y2=0.42
r170 29 38 7.76618 $w=3.3e-07 $l=2.03101e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=6.12 $Y2=2.135
r171 29 31 17.9851 $w=3.28e-07 $l=5.15e-07 $layer=LI1_cond $X=6.035 $Y=2.3
+ $X2=5.52 $Y2=2.3
r172 22 24 132.55 $w=1.8e-07 $l=4.95e-07 $layer=POLY_cond $X=8.225 $Y=1.57
+ $X2=8.225 $Y2=2.065
r173 21 22 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=8.225 $Y=1.47 $X2=8.225
+ $Y2=1.57
r174 21 60 48.0787 $w=2e-07 $l=1.45e-07 $layer=POLY_cond $X=8.225 $Y=1.47
+ $X2=8.225 $Y2=1.325
r175 19 59 141.387 $w=1.5e-07 $l=4.4e-07 $layer=POLY_cond $X=8.195 $Y=0.555
+ $X2=8.195 $Y2=0.995
r176 14 27 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.805
r177 14 16 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=7.26 $Y=0.73
+ $X2=7.26 $Y2=0.445
r178 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.005 $Y=1.99
+ $X2=7.005 $Y2=2.275
r179 10 11 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=7.005 $Y=1.89 $X2=7.005
+ $Y2=1.99
r180 9 56 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=7.005 $Y=1.365
+ $X2=7.005 $Y2=1.23
r181 9 10 174.078 $w=2e-07 $l=5.25e-07 $layer=POLY_cond $X=7.005 $Y=1.365
+ $X2=7.005 $Y2=1.89
r182 8 56 9.86319 $w=2e-07 $l=1.35e-07 $layer=POLY_cond $X=7.005 $Y=1.095
+ $X2=7.005 $Y2=1.23
r183 7 27 130.755 $w=1.5e-07 $l=2.55e-07 $layer=POLY_cond $X=7.005 $Y=0.805
+ $X2=7.26 $Y2=0.805
r184 7 8 71.2891 $w=2e-07 $l=2.15e-07 $layer=POLY_cond $X=7.005 $Y=0.88
+ $X2=7.005 $Y2=1.095
r185 2 31 600 $w=1.7e-07 $l=2.98831e-07 $layer=licon1_PDIFF $count=1 $X=5.375
+ $Y=2.065 $X2=5.52 $Y2=2.3
r186 1 35 182 $w=1.7e-07 $l=2.43311e-07 $layer=licon1_NDIFF $count=1 $X=5.415
+ $Y=0.235 $X2=5.55 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%SET_B 2 3 5 8 10 12 15 18 21 24 25 27 28
+ 30 37
c129 37 0 4.64199e-20 $X=7.52 $Y=1.53
c130 25 0 3.13156e-20 $X=7.715 $Y=1.53
c131 8 0 3.91586e-20 $X=7.67 $Y=0.445
c132 3 0 1.62495e-19 $X=7.595 $Y=1.99
r133 33 37 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=7.5
+ $Y=1.68 $X2=7.5 $Y2=1.68
r134 30 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.52 $Y=1.53
+ $X2=7.52 $Y2=1.53
r135 28 43 3.96743 $w=3.03e-07 $l=1.05e-07 $layer=LI1_cond $X=9.882 $Y=1.53
+ $X2=9.882 $Y2=1.635
r136 27 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=9.875 $Y=1.53
+ $X2=9.875 $Y2=1.53
r137 25 30 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=7.715 $Y=1.53
+ $X2=7.52 $Y2=1.53
r138 24 27 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=9.73 $Y=1.53
+ $X2=9.875 $Y2=1.53
r139 24 25 2.49381 $w=1.4e-07 $l=2.015e-06 $layer=MET1_cond $X=9.73 $Y=1.53
+ $X2=7.715 $Y2=1.53
r140 21 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.78
+ $Y=1.63 $X2=10.78 $Y2=1.63
r141 19 43 3.82255 $w=1.8e-07 $l=1.53e-07 $layer=LI1_cond $X=10.035 $Y=1.635
+ $X2=9.882 $Y2=1.635
r142 19 21 45.904 $w=1.78e-07 $l=7.45e-07 $layer=LI1_cond $X=10.035 $Y=1.635
+ $X2=10.78 $Y2=1.635
r143 17 18 54.0301 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.62 $Y=1.215
+ $X2=7.62 $Y2=1.365
r144 13 22 39.6847 $w=4.05e-07 $l=2.43926e-07 $layer=POLY_cond $X=10.89 $Y=1.465
+ $X2=10.715 $Y2=1.63
r145 13 15 523.021 $w=1.5e-07 $l=1.02e-06 $layer=POLY_cond $X=10.89 $Y=1.465
+ $X2=10.89 $Y2=0.445
r146 10 22 57.9372 $w=4.05e-07 $l=4.28486e-07 $layer=POLY_cond $X=10.565 $Y=1.99
+ $X2=10.715 $Y2=1.63
r147 10 12 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=10.565 $Y=1.99
+ $X2=10.565 $Y2=2.275
r148 8 17 394.83 $w=1.5e-07 $l=7.7e-07 $layer=POLY_cond $X=7.67 $Y=0.445
+ $X2=7.67 $Y2=1.215
r149 3 33 58.4175 $w=2.9e-07 $l=3.40955e-07 $layer=POLY_cond $X=7.595 $Y=1.99
+ $X2=7.53 $Y2=1.68
r150 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=7.595 $Y=1.99
+ $X2=7.595 $Y2=2.275
r151 2 33 32.1081 $w=2.9e-07 $l=1.94808e-07 $layer=POLY_cond $X=7.595 $Y=1.515
+ $X2=7.53 $Y2=1.68
r152 2 18 49.7366 $w=2e-07 $l=1.5e-07 $layer=POLY_cond $X=7.595 $Y=1.515
+ $X2=7.595 $Y2=1.365
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1951_295# 1 2 8 9 11 12 13 16 19 22 23
+ 25 26 29 32 34 37
c102 37 0 1.08045e-19 $X=11.885 $Y=1.28
c103 26 0 6.70306e-20 $X=10.48 $Y=1.28
c104 12 0 1.97973e-19 $X=10.185 $Y=1.55
c105 9 0 9.8756e-21 $X=9.855 $Y=1.99
r106 34 36 6.80499 $w=3.38e-07 $l=1.65e-07 $layer=LI1_cond $X=11.845 $Y=0.42
+ $X2=11.845 $Y2=0.585
r107 32 37 3.77418 $w=2.45e-07 $l=9.21954e-08 $layer=LI1_cond $X=11.9 $Y=1.195
+ $X2=11.885 $Y2=1.28
r108 32 36 30.5648 $w=2.28e-07 $l=6.1e-07 $layer=LI1_cond $X=11.9 $Y=1.195
+ $X2=11.9 $Y2=0.585
r109 27 37 3.77418 $w=2.45e-07 $l=8.5e-08 $layer=LI1_cond $X=11.885 $Y=1.365
+ $X2=11.885 $Y2=1.28
r110 27 29 40.7788 $w=2.58e-07 $l=9.2e-07 $layer=LI1_cond $X=11.885 $Y=1.365
+ $X2=11.885 $Y2=2.285
r111 25 37 2.68609 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=11.755 $Y=1.28
+ $X2=11.885 $Y2=1.28
r112 25 26 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=11.755 $Y=1.28
+ $X2=10.48 $Y2=1.28
r113 23 40 37.8241 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.345 $Y=1.02
+ $X2=10.345 $Y2=1.185
r114 23 39 46.1509 $w=3.2e-07 $l=1.65e-07 $layer=POLY_cond $X=10.345 $Y=1.02
+ $X2=10.345 $Y2=0.855
r115 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=10.32
+ $Y=1.02 $X2=10.32 $Y2=1.02
r116 20 26 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=10.35 $Y=1.195
+ $X2=10.48 $Y2=1.28
r117 20 22 7.75683 $w=2.58e-07 $l=1.75e-07 $layer=LI1_cond $X=10.35 $Y=1.195
+ $X2=10.35 $Y2=1.02
r118 19 40 96.1574 $w=2e-07 $l=2.9e-07 $layer=POLY_cond $X=10.285 $Y=1.475
+ $X2=10.285 $Y2=1.185
r119 16 39 210.234 $w=1.5e-07 $l=4.1e-07 $layer=POLY_cond $X=10.26 $Y=0.445
+ $X2=10.26 $Y2=0.855
r120 12 19 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=10.185 $Y=1.55
+ $X2=10.285 $Y2=1.475
r121 12 13 117.936 $w=1.5e-07 $l=2.3e-07 $layer=POLY_cond $X=10.185 $Y=1.55
+ $X2=9.955 $Y2=1.55
r122 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=9.855 $Y=1.99
+ $X2=9.855 $Y2=2.275
r123 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=9.855 $Y=1.89 $X2=9.855
+ $Y2=1.99
r124 7 13 27.6518 $w=1.5e-07 $l=1.32288e-07 $layer=POLY_cond $X=9.855 $Y=1.625
+ $X2=9.955 $Y2=1.55
r125 7 8 87.868 $w=2e-07 $l=2.65e-07 $layer=POLY_cond $X=9.855 $Y=1.625
+ $X2=9.855 $Y2=1.89
r126 2 29 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=11.695
+ $Y=2.065 $X2=11.84 $Y2=2.285
r127 1 34 182 $w=1.7e-07 $l=3.34963e-07 $layer=licon1_NDIFF $count=1 $X=11.585
+ $Y=0.235 $X2=11.84 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_1745_329# 1 2 3 12 13 15 16 18 20 23 25
+ 26 27 28 32 36 39 40 42 43 45 47 57
c140 23 0 1.61945e-19 $X=12.62 $Y=0.56
r141 62 64 11.2698 $w=4.1e-07 $l=8.87412e-08 $layer=POLY_cond $X=11.425 $Y=1.205
+ $X2=11.455 $Y2=1.28
r142 58 64 48.2 $w=4.1e-07 $l=4.1e-07 $layer=POLY_cond $X=11.455 $Y=1.69
+ $X2=11.455 $Y2=1.28
r143 57 60 8.79496 $w=3.78e-07 $l=2.9e-07 $layer=LI1_cond $X=11.395 $Y=1.69
+ $X2=11.395 $Y2=1.98
r144 57 58 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.37
+ $Y=1.69 $X2=11.37 $Y2=1.69
r145 45 60 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.205 $Y=1.98
+ $X2=11.395 $Y2=1.98
r146 45 46 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=11.205 $Y=1.98
+ $X2=11.015 $Y2=1.98
r147 43 62 49.5896 $w=3.2e-07 $l=2.75e-07 $layer=POLY_cond $X=11.425 $Y=0.93
+ $X2=11.425 $Y2=1.205
r148 42 43 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=11.4
+ $Y=0.93 $X2=11.4 $Y2=0.93
r149 40 42 24.552 $w=2.28e-07 $l=4.9e-07 $layer=LI1_cond $X=10.91 $Y=0.9
+ $X2=11.4 $Y2=0.9
r150 39 40 6.85974 $w=2.3e-07 $l=1.57242e-07 $layer=LI1_cond $X=10.81 $Y=0.785
+ $X2=10.91 $Y2=0.9
r151 38 39 13.3091 $w=1.98e-07 $l=2.4e-07 $layer=LI1_cond $X=10.81 $Y=0.545
+ $X2=10.81 $Y2=0.785
r152 37 47 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.84 $Y=1.98
+ $X2=9.755 $Y2=1.98
r153 36 54 8.67889 $w=4.03e-07 $l=3.05e-07 $layer=LI1_cond $X=10.812 $Y=1.98
+ $X2=10.812 $Y2=2.285
r154 36 46 5.85399 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=10.812 $Y=1.98
+ $X2=11.015 $Y2=1.98
r155 36 37 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=10.61 $Y=1.98
+ $X2=9.84 $Y2=1.98
r156 32 38 7.01501 $w=2.7e-07 $l=1.78115e-07 $layer=LI1_cond $X=10.71 $Y=0.41
+ $X2=10.81 $Y2=0.545
r157 32 34 54.6343 $w=2.68e-07 $l=1.28e-06 $layer=LI1_cond $X=10.71 $Y=0.41
+ $X2=9.43 $Y2=0.41
r158 28 47 20.3551 $w=1.68e-07 $l=3.12e-07 $layer=LI1_cond $X=9.755 $Y=2.292
+ $X2=9.755 $Y2=1.98
r159 28 30 22.3608 $w=3.33e-07 $l=6.5e-07 $layer=LI1_cond $X=9.67 $Y=2.292
+ $X2=9.02 $Y2=2.292
r160 25 43 0.901628 $w=3.2e-07 $l=5e-09 $layer=POLY_cond $X=11.425 $Y=0.925
+ $X2=11.425 $Y2=0.93
r161 25 26 45.2492 $w=3.2e-07 $l=1.6e-07 $layer=POLY_cond $X=11.425 $Y=0.925
+ $X2=11.425 $Y2=0.765
r162 21 27 18.8402 $w=1.65e-07 $l=1.13816e-07 $layer=POLY_cond $X=12.62 $Y=1.205
+ $X2=12.595 $Y2=1.307
r163 21 23 330.734 $w=1.5e-07 $l=6.45e-07 $layer=POLY_cond $X=12.62 $Y=1.205
+ $X2=12.62 $Y2=0.56
r164 18 27 18.8402 $w=1.65e-07 $l=1.03e-07 $layer=POLY_cond $X=12.595 $Y=1.41
+ $X2=12.595 $Y2=1.307
r165 18 20 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=12.595 $Y=1.41
+ $X2=12.595 $Y2=1.985
r166 17 64 26.4667 $w=1.5e-07 $l=2.5e-07 $layer=POLY_cond $X=11.705 $Y=1.28
+ $X2=11.455 $Y2=1.28
r167 16 27 6.66866 $w=1.5e-07 $l=1.12694e-07 $layer=POLY_cond $X=12.495 $Y=1.28
+ $X2=12.595 $Y2=1.307
r168 16 17 405.085 $w=1.5e-07 $l=7.9e-07 $layer=POLY_cond $X=12.495 $Y=1.28
+ $X2=11.705 $Y2=1.28
r169 13 58 50.6865 $w=4.1e-07 $l=3.67423e-07 $layer=POLY_cond $X=11.605 $Y=1.99
+ $X2=11.455 $Y2=1.69
r170 13 15 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=11.605 $Y=1.99
+ $X2=11.605 $Y2=2.275
r171 12 26 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=11.51 $Y=0.445
+ $X2=11.51 $Y2=0.765
r172 3 54 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=10.655
+ $Y=2.065 $X2=10.8 $Y2=2.285
r173 2 30 600 $w=1.7e-07 $l=7.78653e-07 $layer=licon1_PDIFF $count=1 $X=8.725
+ $Y=1.645 $X2=9.02 $Y2=2.29
r174 1 34 182 $w=1.7e-07 $l=2.7037e-07 $layer=licon1_NDIFF $count=1 $X=9.215
+ $Y=0.235 $X2=9.43 $Y2=0.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_2447_47# 1 2 7 9 10 12 13 15 16 18 19
+ 21 22 24 25 27 28 30 33 37 41 44 52
r99 52 53 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=14.58 $Y=1.202
+ $X2=14.605 $Y2=1.202
r100 51 52 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=14.135 $Y=1.202
+ $X2=14.58 $Y2=1.202
r101 50 51 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=14.11 $Y=1.202
+ $X2=14.135 $Y2=1.202
r102 49 50 64.8342 $w=3.68e-07 $l=4.95e-07 $layer=POLY_cond $X=13.615 $Y=1.202
+ $X2=14.11 $Y2=1.202
r103 48 49 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=13.59 $Y=1.202
+ $X2=13.615 $Y2=1.202
r104 47 48 58.2853 $w=3.68e-07 $l=4.45e-07 $layer=POLY_cond $X=13.145 $Y=1.202
+ $X2=13.59 $Y2=1.202
r105 46 47 3.27446 $w=3.68e-07 $l=2.5e-08 $layer=POLY_cond $X=13.12 $Y=1.202
+ $X2=13.145 $Y2=1.202
r106 42 46 10.4783 $w=3.68e-07 $l=8e-08 $layer=POLY_cond $X=13.04 $Y=1.202
+ $X2=13.12 $Y2=1.202
r107 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=13.04
+ $Y=1.16 $X2=13.04 $Y2=1.16
r108 39 44 0.499868 $w=3.3e-07 $l=1.3e-07 $layer=LI1_cond $X=12.445 $Y=1.16
+ $X2=12.315 $Y2=1.16
r109 39 41 20.7789 $w=3.28e-07 $l=5.95e-07 $layer=LI1_cond $X=12.445 $Y=1.16
+ $X2=13.04 $Y2=1.16
r110 35 44 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=12.315 $Y=1.325
+ $X2=12.315 $Y2=1.16
r111 35 37 27.9246 $w=2.58e-07 $l=6.3e-07 $layer=LI1_cond $X=12.315 $Y=1.325
+ $X2=12.315 $Y2=1.955
r112 31 44 6.26932 $w=2.6e-07 $l=1.65e-07 $layer=LI1_cond $X=12.315 $Y=0.995
+ $X2=12.315 $Y2=1.16
r113 31 33 25.2651 $w=2.58e-07 $l=5.7e-07 $layer=LI1_cond $X=12.315 $Y=0.995
+ $X2=12.315 $Y2=0.425
r114 28 53 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.605 $Y=0.995
+ $X2=14.605 $Y2=1.202
r115 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.605 $Y=0.995
+ $X2=14.605 $Y2=0.56
r116 25 52 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.58 $Y=1.41
+ $X2=14.58 $Y2=1.202
r117 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.58 $Y=1.41
+ $X2=14.58 $Y2=1.985
r118 22 51 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=14.135 $Y=0.995
+ $X2=14.135 $Y2=1.202
r119 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=14.135 $Y=0.995
+ $X2=14.135 $Y2=0.56
r120 19 50 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=14.11 $Y=1.41
+ $X2=14.11 $Y2=1.202
r121 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=14.11 $Y=1.41
+ $X2=14.11 $Y2=1.985
r122 16 49 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.615 $Y=0.995
+ $X2=13.615 $Y2=1.202
r123 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.615 $Y=0.995
+ $X2=13.615 $Y2=0.56
r124 13 48 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.59 $Y=1.41
+ $X2=13.59 $Y2=1.202
r125 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.59 $Y=1.41
+ $X2=13.59 $Y2=1.985
r126 10 47 23.8357 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=13.145 $Y=0.995
+ $X2=13.145 $Y2=1.202
r127 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=13.145 $Y=0.995
+ $X2=13.145 $Y2=0.56
r128 7 46 19.486 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=13.12 $Y=1.41
+ $X2=13.12 $Y2=1.202
r129 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=13.12 $Y=1.41
+ $X2=13.12 $Y2=1.985
r130 2 37 300 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_PDIFF $count=2 $X=12.235
+ $Y=1.485 $X2=12.36 $Y2=1.955
r131 1 33 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=12.235
+ $Y=0.235 $X2=12.36 $Y2=0.425
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_27_369# 1 2 7 10 11 13 14 16
r46 14 16 45.1558 $w=2.08e-07 $l=8.55e-07 $layer=LI1_cond $X=1.225 $Y=2.36
+ $X2=2.08 $Y2=2.36
r47 13 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.14 $Y=2.255
+ $X2=1.225 $Y2=2.36
r48 12 13 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.14 $Y=2.025
+ $X2=1.14 $Y2=2.255
r49 10 12 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.055 $Y=1.935
+ $X2=1.14 $Y2=2.025
r50 10 11 43.7475 $w=1.78e-07 $l=7.1e-07 $layer=LI1_cond $X=1.055 $Y=1.935
+ $X2=0.345 $Y2=1.935
r51 7 11 7.11373 $w=1.8e-07 $l=1.69115e-07 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.345 $Y2=1.935
r52 7 9 2.11154 $w=2.6e-07 $l=4.5e-08 $layer=LI1_cond $X=0.215 $Y=2.025
+ $X2=0.215 $Y2=2.07
r53 2 16 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=1.935
+ $Y=1.845 $X2=2.08 $Y2=2.34
r54 1 9 600 $w=1.7e-07 $l=2.80624e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.845 $X2=0.26 $Y2=2.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%VPWR 1 2 3 4 5 6 7 8 9 10 33 37 39 41 42
+ 45 47 51 55 61 65 67 74 76 77 78 80 85 90 102 110 119 124 127 130 137 146 148
+ 151 154 158
c211 158 0 1.2037e-19 $X=14.95 $Y=2.72
c212 5 0 1.36329e-19 $X=7.685 $Y=2.065
r213 157 158 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=2.72
+ $X2=14.95 $Y2=2.72
r214 154 155 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.65 $Y=2.72
+ $X2=12.65 $Y2=2.72
r215 151 152 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r216 149 152 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r217 148 149 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r218 144 146 12.2594 $w=6.78e-07 $l=2.55e-07 $layer=LI1_cond $X=8.51 $Y=2.465
+ $X2=8.765 $Y2=2.465
r219 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r220 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r221 130 133 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=2.36
+ $X2=4.035 $Y2=2.72
r222 128 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r223 127 128 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r224 124 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r225 122 158 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=2.72
+ $X2=14.95 $Y2=2.72
r226 121 122 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=2.72
+ $X2=14.49 $Y2=2.72
r227 119 157 4.31409 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=14.78 $Y=2.72
+ $X2=14.98 $Y2=2.72
r228 119 121 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=14.78 $Y=2.72
+ $X2=14.49 $Y2=2.72
r229 118 122 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=14.49 $Y2=2.72
r230 118 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=2.72
+ $X2=12.65 $Y2=2.72
r231 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=2.72
+ $X2=13.57 $Y2=2.72
r232 115 154 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=13.02 $Y=2.72
+ $X2=12.817 $Y2=2.72
r233 115 117 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=13.02 $Y=2.72
+ $X2=13.57 $Y2=2.72
r234 114 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=12.65 $Y2=2.72
r235 114 152 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=2.72
+ $X2=11.27 $Y2=2.72
r236 113 114 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.73 $Y=2.72
+ $X2=11.73 $Y2=2.72
r237 111 151 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.585 $Y=2.72
+ $X2=11.395 $Y2=2.72
r238 111 113 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=11.585 $Y=2.72
+ $X2=11.73 $Y2=2.72
r239 110 154 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=12.615 $Y=2.72
+ $X2=12.817 $Y2=2.72
r240 110 113 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=12.615 $Y=2.72
+ $X2=11.73 $Y2=2.72
r241 109 149 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=9.89 $Y=2.72
+ $X2=10.35 $Y2=2.72
r242 108 109 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=9.89 $Y=2.72
+ $X2=9.89 $Y2=2.72
r243 106 109 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r244 106 145 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.97 $Y=2.72
+ $X2=8.51 $Y2=2.72
r245 105 108 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=9.89 $Y2=2.72
r246 105 146 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=8.97 $Y=2.72
+ $X2=8.765 $Y2=2.72
r247 105 106 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=8.97 $Y=2.72
+ $X2=8.97 $Y2=2.72
r248 102 148 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.06 $Y=2.72
+ $X2=10.25 $Y2=2.72
r249 102 108 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=10.06 $Y=2.72
+ $X2=9.89 $Y2=2.72
r250 101 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r251 101 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=6.67 $Y2=2.72
r252 100 101 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r253 98 100 49.5829 $w=1.68e-07 $l=7.6e-07 $layer=LI1_cond $X=6.83 $Y=2.72
+ $X2=7.59 $Y2=2.72
r254 97 141 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r255 96 97 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r256 94 97 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r257 94 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=3.91 $Y2=2.72
r258 93 96 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=4.37 $Y=2.72
+ $X2=6.21 $Y2=2.72
r259 93 94 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r260 91 133 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.035 $Y2=2.72
r261 91 93 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.225 $Y=2.72
+ $X2=4.37 $Y2=2.72
r262 90 98 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=6.637 $Y=2.72
+ $X2=6.83 $Y2=2.72
r263 90 141 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r264 90 137 10.7761 $w=3.83e-07 $l=3.6e-07 $layer=LI1_cond $X=6.637 $Y=2.72
+ $X2=6.637 $Y2=2.36
r265 90 96 15.3316 $w=1.68e-07 $l=2.35e-07 $layer=LI1_cond $X=6.445 $Y=2.72
+ $X2=6.21 $Y2=2.72
r266 89 128 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.99 $Y2=2.72
r267 89 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r268 88 89 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r269 86 124 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=0.675 $Y2=2.72
r270 86 88 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.835 $Y=2.72
+ $X2=1.15 $Y2=2.72
r271 85 127 7.94884 $w=1.7e-07 $l=1.47e-07 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=3.087 $Y2=2.72
r272 85 88 116.781 $w=1.68e-07 $l=1.79e-06 $layer=LI1_cond $X=2.94 $Y=2.72
+ $X2=1.15 $Y2=2.72
r273 80 124 8.42608 $w=1.7e-07 $l=1.6e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.675 $Y2=2.72
r274 80 82 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r275 78 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r276 78 82 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r277 76 117 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.79 $Y=2.72
+ $X2=13.57 $Y2=2.72
r278 76 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=2.72
+ $X2=13.875 $Y2=2.72
r279 75 121 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.96 $Y=2.72
+ $X2=14.49 $Y2=2.72
r280 75 77 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.96 $Y=2.72
+ $X2=13.875 $Y2=2.72
r281 74 100 7.82888 $w=1.68e-07 $l=1.2e-07 $layer=LI1_cond $X=7.71 $Y=2.72
+ $X2=7.59 $Y2=2.72
r282 73 74 10.6764 $w=6.78e-07 $l=1.65e-07 $layer=LI1_cond $X=7.875 $Y=2.465
+ $X2=7.71 $Y2=2.465
r283 67 70 27.4969 $w=2.83e-07 $l=6.8e-07 $layer=LI1_cond $X=14.922 $Y=1.66
+ $X2=14.922 $Y2=2.34
r284 65 157 3.08458 $w=2.85e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.922 $Y=2.635
+ $X2=14.98 $Y2=2.72
r285 65 70 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=14.922 $Y=2.635
+ $X2=14.922 $Y2=2.34
r286 61 64 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=13.875 $Y=1.66
+ $X2=13.875 $Y2=2.34
r287 59 77 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.875 $Y=2.635
+ $X2=13.875 $Y2=2.72
r288 59 64 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.875 $Y=2.635
+ $X2=13.875 $Y2=2.34
r289 55 58 19.3497 $w=4.03e-07 $l=6.8e-07 $layer=LI1_cond $X=12.817 $Y=1.68
+ $X2=12.817 $Y2=2.36
r290 53 154 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=12.817 $Y=2.635
+ $X2=12.817 $Y2=2.72
r291 53 58 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=12.817 $Y=2.635
+ $X2=12.817 $Y2=2.36
r292 49 151 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=11.395 $Y=2.635
+ $X2=11.395 $Y2=2.72
r293 49 51 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=11.395 $Y=2.635
+ $X2=11.395 $Y2=2.34
r294 48 148 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.44 $Y=2.72
+ $X2=10.25 $Y2=2.72
r295 47 151 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=11.395 $Y2=2.72
r296 47 48 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=11.205 $Y=2.72
+ $X2=10.44 $Y2=2.72
r297 43 148 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.25 $Y=2.635
+ $X2=10.25 $Y2=2.72
r298 43 45 8.34005 $w=3.78e-07 $l=2.75e-07 $layer=LI1_cond $X=10.25 $Y=2.635
+ $X2=10.25 $Y2=2.36
r299 42 73 3.07814 $w=6.78e-07 $l=1.75e-07 $layer=LI1_cond $X=8.05 $Y=2.465
+ $X2=7.875 $Y2=2.465
r300 41 144 1.4951 $w=6.78e-07 $l=8.5e-08 $layer=LI1_cond $X=8.425 $Y=2.465
+ $X2=8.51 $Y2=2.465
r301 41 42 6.59602 $w=6.78e-07 $l=3.75e-07 $layer=LI1_cond $X=8.425 $Y=2.465
+ $X2=8.05 $Y2=2.465
r302 40 127 7.94884 $w=1.7e-07 $l=1.48e-07 $layer=LI1_cond $X=3.235 $Y=2.72
+ $X2=3.087 $Y2=2.72
r303 39 133 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=4.035 $Y2=2.72
r304 39 40 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=3.235 $Y2=2.72
r305 35 127 0.543863 $w=2.95e-07 $l=8.5e-08 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=2.72
r306 35 37 11.5244 $w=2.93e-07 $l=2.95e-07 $layer=LI1_cond $X=3.087 $Y=2.635
+ $X2=3.087 $Y2=2.34
r307 31 124 0.800721 $w=3.2e-07 $l=8.5e-08 $layer=LI1_cond $X=0.675 $Y=2.635
+ $X2=0.675 $Y2=2.72
r308 31 33 9.90381 $w=3.18e-07 $l=2.75e-07 $layer=LI1_cond $X=0.675 $Y=2.635
+ $X2=0.675 $Y2=2.36
r309 10 70 400 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=14.67
+ $Y=1.485 $X2=14.865 $Y2=2.34
r310 10 67 400 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=14.67
+ $Y=1.485 $X2=14.865 $Y2=1.66
r311 9 64 400 $w=1.7e-07 $l=9.47497e-07 $layer=licon1_PDIFF $count=1 $X=13.68
+ $Y=1.485 $X2=13.875 $Y2=2.34
r312 9 61 400 $w=1.7e-07 $l=2.68608e-07 $layer=licon1_PDIFF $count=1 $X=13.68
+ $Y=1.485 $X2=13.875 $Y2=1.66
r313 8 58 400 $w=1.7e-07 $l=9.5623e-07 $layer=licon1_PDIFF $count=1 $X=12.685
+ $Y=1.485 $X2=12.855 $Y2=2.36
r314 8 55 400 $w=1.7e-07 $l=2.66786e-07 $layer=licon1_PDIFF $count=1 $X=12.685
+ $Y=1.485 $X2=12.855 $Y2=1.68
r315 7 51 600 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_PDIFF $count=1 $X=11.245
+ $Y=2.065 $X2=11.37 $Y2=2.34
r316 6 45 600 $w=1.7e-07 $l=4.11856e-07 $layer=licon1_PDIFF $count=1 $X=9.945
+ $Y=2.065 $X2=10.225 $Y2=2.36
r317 5 73 600 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_PDIFF $count=1 $X=7.685
+ $Y=2.065 $X2=7.875 $Y2=2.36
r318 4 137 600 $w=1.7e-07 $l=3.84057e-07 $layer=licon1_PDIFF $count=1 $X=6.405
+ $Y=2.065 $X2=6.61 $Y2=2.36
r319 3 130 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=3.915
+ $Y=1.845 $X2=4.06 $Y2=2.36
r320 2 37 600 $w=1.7e-07 $l=5.6285e-07 $layer=licon1_PDIFF $count=1 $X=2.925
+ $Y=1.845 $X2=3.07 $Y2=2.34
r321 1 33 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.845 $X2=0.73 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%A_201_47# 1 2 3 4 13 19 21 23 28 33 36 37
+ 40 43 44
c126 43 0 4.73773e-19 $X=5.095 $Y=1.53
c127 37 0 1.4475e-19 $X=1.955 $Y=1.53
c128 33 0 1.00357e-19 $X=5.017 $Y=0.78
c129 28 0 1.40323e-19 $X=1.75 $Y=1.965
c130 13 0 4.39648e-20 $X=1.655 $Y=0.425
r131 43 44 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.095 $Y=1.53
+ $X2=5.095 $Y2=1.53
r132 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.76 $Y=1.53
+ $X2=1.76 $Y2=1.53
r133 37 39 0.147547 $w=2.3e-07 $l=1.95e-07 $layer=MET1_cond $X=1.955 $Y=1.53
+ $X2=1.76 $Y2=1.53
r134 36 43 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=5.095 $Y2=1.53
r135 36 37 3.70668 $w=1.4e-07 $l=2.995e-06 $layer=MET1_cond $X=4.95 $Y=1.53
+ $X2=1.955 $Y2=1.53
r136 35 44 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=5.095 $Y=1.59
+ $X2=5.095 $Y2=1.53
r137 33 44 48.9305 $w=1.68e-07 $l=7.5e-07 $layer=LI1_cond $X=5.095 $Y=0.78
+ $X2=5.095 $Y2=1.53
r138 31 40 54.5789 $w=1.88e-07 $l=9.35e-07 $layer=LI1_cond $X=1.75 $Y=0.595
+ $X2=1.75 $Y2=1.53
r139 29 40 18.3876 $w=1.88e-07 $l=3.15e-07 $layer=LI1_cond $X=1.75 $Y=1.845
+ $X2=1.75 $Y2=1.53
r140 28 29 2.10789 $w=1.9e-07 $l=1.2e-07 $layer=LI1_cond $X=1.75 $Y=1.965
+ $X2=1.75 $Y2=1.845
r141 26 28 6.72258 $w=2.38e-07 $l=1.4e-07 $layer=LI1_cond $X=1.61 $Y=1.965
+ $X2=1.75 $Y2=1.965
r142 21 35 6.27261 $w=2.13e-07 $l=1.07e-07 $layer=LI1_cond $X=5.072 $Y=1.697
+ $X2=5.072 $Y2=1.59
r143 21 23 32.322 $w=2.13e-07 $l=6.03e-07 $layer=LI1_cond $X=5.072 $Y=1.697
+ $X2=5.072 $Y2=2.3
r144 17 33 8.35379 $w=3.23e-07 $l=1.62e-07 $layer=LI1_cond $X=5.017 $Y=0.618
+ $X2=5.017 $Y2=0.78
r145 17 19 7.02104 $w=3.23e-07 $l=1.98e-07 $layer=LI1_cond $X=5.017 $Y=0.618
+ $X2=5.017 $Y2=0.42
r146 13 31 7.55181 $w=3.4e-07 $l=2.1225e-07 $layer=LI1_cond $X=1.655 $Y=0.425
+ $X2=1.75 $Y2=0.595
r147 13 15 17.4561 $w=3.38e-07 $l=5.15e-07 $layer=LI1_cond $X=1.655 $Y=0.425
+ $X2=1.14 $Y2=0.425
r148 4 23 600 $w=1.7e-07 $l=2.90861e-07 $layer=licon1_PDIFF $count=1 $X=4.925
+ $Y=2.065 $X2=5.05 $Y2=2.3
r149 3 26 600 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=1 $X=1.465
+ $Y=1.845 $X2=1.61 $Y2=1.97
r150 2 19 182 $w=1.7e-07 $l=2.39479e-07 $layer=licon1_NDIFF $count=1 $X=4.955
+ $Y=0.235 $X2=5.08 $Y2=0.42
r151 1 15 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.005
+ $Y=0.235 $X2=1.14 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%Q 1 2 3 4 15 17 19 22 25 26 28 29 30 31
+ 32 33 34 35 43 45 49
c49 28 0 1.03354e-19 $X=13.457 $Y=1.19
c50 22 0 2.30468e-20 $X=13.457 $Y=1.055
r51 35 65 3.61315 $w=4.78e-07 $l=1.45e-07 $layer=LI1_cond $X=14.37 $Y=2.21
+ $X2=14.37 $Y2=2.355
r52 34 35 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=14.37 $Y=1.87
+ $X2=14.37 $Y2=2.21
r53 34 59 4.85907 $w=4.78e-07 $l=1.95e-07 $layer=LI1_cond $X=14.37 $Y=1.87
+ $X2=14.37 $Y2=1.675
r54 33 59 3.61315 $w=4.78e-07 $l=1.45e-07 $layer=LI1_cond $X=14.37 $Y=1.53
+ $X2=14.37 $Y2=1.675
r55 33 55 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=14.37 $Y=1.53
+ $X2=14.37 $Y2=1.325
r56 32 43 3.47601 $w=2.7e-07 $l=2.4e-07 $layer=LI1_cond $X=14.37 $Y=1.19
+ $X2=14.13 $Y2=1.19
r57 32 47 3.128 $w=4.8e-07 $l=1.35e-07 $layer=LI1_cond $X=14.37 $Y=1.19
+ $X2=14.37 $Y2=1.055
r58 32 55 3.128 $w=4.8e-07 $l=1.35e-07 $layer=LI1_cond $X=14.37 $Y=1.19
+ $X2=14.37 $Y2=1.325
r59 31 47 5.10825 $w=4.78e-07 $l=2.05e-07 $layer=LI1_cond $X=14.37 $Y=0.85
+ $X2=14.37 $Y2=1.055
r60 30 31 8.47222 $w=4.78e-07 $l=3.4e-07 $layer=LI1_cond $X=14.37 $Y=0.51
+ $X2=14.37 $Y2=0.85
r61 30 49 3.73775 $w=4.78e-07 $l=1.5e-07 $layer=LI1_cond $X=14.37 $Y=0.51
+ $X2=14.37 $Y2=0.36
r62 29 43 5.76222 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=13.995 $Y=1.19
+ $X2=14.13 $Y2=1.19
r63 29 45 0.213415 $w=2.68e-07 $l=5e-09 $layer=LI1_cond $X=13.995 $Y=1.19
+ $X2=13.99 $Y2=1.19
r64 27 45 17.9269 $w=2.68e-07 $l=4.2e-07 $layer=LI1_cond $X=13.57 $Y=1.19
+ $X2=13.99 $Y2=1.19
r65 27 28 0.695019 $w=2.7e-07 $l=1.13e-07 $layer=LI1_cond $X=13.57 $Y=1.19
+ $X2=13.457 $Y2=1.19
r66 23 28 5.99569 $w=2.25e-07 $l=1.35e-07 $layer=LI1_cond $X=13.457 $Y=1.325
+ $X2=13.457 $Y2=1.19
r67 23 26 8.70735 $w=2.23e-07 $l=1.7e-07 $layer=LI1_cond $X=13.457 $Y=1.325
+ $X2=13.457 $Y2=1.495
r68 22 28 5.99569 $w=2.25e-07 $l=1.35e-07 $layer=LI1_cond $X=13.457 $Y=1.055
+ $X2=13.457 $Y2=1.19
r69 22 25 11.7805 $w=2.23e-07 $l=2.3e-07 $layer=LI1_cond $X=13.457 $Y=1.055
+ $X2=13.457 $Y2=0.825
r70 17 26 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=1.66
+ $X2=13.405 $Y2=1.495
r71 17 19 21.8266 $w=3.28e-07 $l=6.25e-07 $layer=LI1_cond $X=13.405 $Y=1.66
+ $X2=13.405 $Y2=2.285
r72 13 25 6.93655 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=13.405 $Y=0.66
+ $X2=13.405 $Y2=0.825
r73 13 15 7.68295 $w=3.28e-07 $l=2.2e-07 $layer=LI1_cond $X=13.405 $Y=0.66
+ $X2=13.405 $Y2=0.44
r74 4 65 400 $w=1.7e-07 $l=9.39707e-07 $layer=licon1_PDIFF $count=1 $X=14.2
+ $Y=1.485 $X2=14.345 $Y2=2.355
r75 4 59 400 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_PDIFF $count=1 $X=14.2
+ $Y=1.485 $X2=14.345 $Y2=1.675
r76 3 19 600 $w=1.7e-07 $l=8.69483e-07 $layer=licon1_PDIFF $count=1 $X=13.21
+ $Y=1.485 $X2=13.355 $Y2=2.285
r77 2 49 91 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=2 $X=14.21
+ $Y=0.235 $X2=14.345 $Y2=0.36
r78 1 15 182 $w=1.7e-07 $l=2.64008e-07 $layer=licon1_NDIFF $count=1 $X=13.22
+ $Y=0.235 $X2=13.355 $Y2=0.44
.ends

.subckt PM_SKY130_FD_SC_HDLL__SDFSTP_4%VGND 1 2 3 4 5 6 7 8 9 10 31 32 35 37 41
+ 45 49 53 57 59 61 64 65 67 68 69 75 87 95 104 117 120 131 135 137 140 144
c197 144 0 2.71124e-20 $X=14.95 $Y=0
c198 75 0 6.74919e-20 $X=6.06 $Y=0
r199 143 144 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=14.95 $Y=0
+ $X2=14.95 $Y2=0
r200 140 141 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=12.65 $Y=0
+ $X2=12.65 $Y2=0
r201 137 138 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r202 133 135 14.9552 $w=8.88e-07 $l=3.65e-07 $layer=LI1_cond $X=8.05 $Y=0.36
+ $X2=8.415 $Y2=0.36
r203 133 134 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.05 $Y=0
+ $X2=8.05 $Y2=0
r204 130 133 2.19326 $w=8.88e-07 $l=1.6e-07 $layer=LI1_cond $X=7.89 $Y=0.36
+ $X2=8.05 $Y2=0.36
r205 130 131 18.6563 $w=8.88e-07 $l=6.35e-07 $layer=LI1_cond $X=7.89 $Y=0.36
+ $X2=7.255 $Y2=0.36
r206 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r207 118 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0
+ $X2=2.99 $Y2=0
r208 117 118 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r209 115 118 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0
+ $X2=2.07 $Y2=0
r210 114 115 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0
+ $X2=0.69 $Y2=0
r211 112 114 8.43408 $w=6.22e-07 $l=4.3e-07 $layer=LI1_cond $X=0.26 $Y=0.255
+ $X2=0.69 $Y2=0.255
r212 109 112 0.588424 $w=6.22e-07 $l=3e-08 $layer=LI1_cond $X=0.23 $Y=0.255
+ $X2=0.26 $Y2=0.255
r213 107 144 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=14.49 $Y=0
+ $X2=14.95 $Y2=0
r214 106 107 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=14.49 $Y=0
+ $X2=14.49 $Y2=0
r215 104 143 4.31409 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=14.78 $Y=0 $X2=14.98
+ $Y2=0
r216 104 106 18.9198 $w=1.68e-07 $l=2.9e-07 $layer=LI1_cond $X=14.78 $Y=0
+ $X2=14.49 $Y2=0
r217 103 107 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=14.49 $Y2=0
r218 103 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=13.57 $Y=0
+ $X2=12.65 $Y2=0
r219 102 103 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=13.57 $Y=0
+ $X2=13.57 $Y2=0
r220 100 140 9.89127 $w=1.7e-07 $l=2.03e-07 $layer=LI1_cond $X=13.02 $Y=0
+ $X2=12.817 $Y2=0
r221 100 102 35.8824 $w=1.68e-07 $l=5.5e-07 $layer=LI1_cond $X=13.02 $Y=0
+ $X2=13.57 $Y2=0
r222 99 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=12.65 $Y2=0
r223 99 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=11.73 $Y=0
+ $X2=11.27 $Y2=0
r224 98 99 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=11.73 $Y=0
+ $X2=11.73 $Y2=0
r225 96 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.415 $Y=0
+ $X2=11.29 $Y2=0
r226 96 98 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=11.415 $Y=0
+ $X2=11.73 $Y2=0
r227 95 140 9.89127 $w=1.7e-07 $l=2.02e-07 $layer=LI1_cond $X=12.615 $Y=0
+ $X2=12.817 $Y2=0
r228 95 98 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=12.615 $Y=0
+ $X2=11.73 $Y2=0
r229 94 138 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=10.81 $Y=0
+ $X2=11.27 $Y2=0
r230 93 94 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=10.81 $Y=0
+ $X2=10.81 $Y2=0
r231 91 94 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=10.81 $Y2=0
r232 91 134 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=8.05 $Y2=0
r233 90 93 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=8.51 $Y=0 $X2=10.81
+ $Y2=0
r234 90 135 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=8.51 $Y=0
+ $X2=8.415 $Y2=0
r235 90 91 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=8.51 $Y=0 $X2=8.51
+ $Y2=0
r236 87 137 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=11.165 $Y=0
+ $X2=11.29 $Y2=0
r237 87 93 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=11.165 $Y=0
+ $X2=10.81 $Y2=0
r238 86 134 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=8.05 $Y2=0
r239 86 125 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.13 $Y=0
+ $X2=6.21 $Y2=0
r240 85 131 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=7.13 $Y=0
+ $X2=7.255 $Y2=0
r241 85 86 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r242 83 85 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=6.595 $Y=0
+ $X2=7.13 $Y2=0
r243 81 125 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.21 $Y2=0
r244 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r245 78 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=4.37 $Y=0
+ $X2=5.75 $Y2=0
r246 77 80 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.75
+ $Y2=0
r247 77 78 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r248 75 127 8.49551 $w=5.33e-07 $l=3.8e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.327 $Y2=0.38
r249 75 83 7.58357 $w=1.7e-07 $l=2.68e-07 $layer=LI1_cond $X=6.327 $Y=0
+ $X2=6.595 $Y2=0
r250 75 125 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r251 75 80 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=6.06 $Y=0 $X2=5.75
+ $Y2=0
r252 74 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.37
+ $Y2=0
r253 74 121 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=2.99 $Y2=0
r254 73 74 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r255 71 120 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=3.35 $Y=0
+ $X2=3.145 $Y2=0
r256 71 73 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=3.35 $Y=0 $X2=3.91
+ $Y2=0
r257 69 115 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=0.69 $Y2=0
r258 69 109 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r259 67 102 14.3529 $w=1.68e-07 $l=2.2e-07 $layer=LI1_cond $X=13.79 $Y=0
+ $X2=13.57 $Y2=0
r260 67 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.79 $Y=0
+ $X2=13.875 $Y2=0
r261 66 106 34.5775 $w=1.68e-07 $l=5.3e-07 $layer=LI1_cond $X=13.96 $Y=0
+ $X2=14.49 $Y2=0
r262 66 68 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.96 $Y=0
+ $X2=13.875 $Y2=0
r263 64 73 0.97861 $w=1.68e-07 $l=1.5e-08 $layer=LI1_cond $X=3.925 $Y=0 $X2=3.91
+ $Y2=0
r264 64 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.925 $Y=0 $X2=4.09
+ $Y2=0
r265 63 77 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=4.255 $Y=0
+ $X2=4.37 $Y2=0
r266 63 65 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.255 $Y=0 $X2=4.09
+ $Y2=0
r267 59 143 3.08458 $w=2.85e-07 $l=1.1025e-07 $layer=LI1_cond $X=14.922 $Y=0.085
+ $X2=14.98 $Y2=0
r268 59 61 11.9288 $w=2.83e-07 $l=2.95e-07 $layer=LI1_cond $X=14.922 $Y=0.085
+ $X2=14.922 $Y2=0.38
r269 55 68 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=13.875 $Y=0.085
+ $X2=13.875 $Y2=0
r270 55 57 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=13.875 $Y=0.085
+ $X2=13.875 $Y2=0.38
r271 51 140 1.50354 $w=4.05e-07 $l=8.5e-08 $layer=LI1_cond $X=12.817 $Y=0.085
+ $X2=12.817 $Y2=0
r272 51 53 7.82523 $w=4.03e-07 $l=2.75e-07 $layer=LI1_cond $X=12.817 $Y=0.085
+ $X2=12.817 $Y2=0.36
r273 47 137 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=11.29 $Y=0.085
+ $X2=11.29 $Y2=0
r274 47 49 12.6769 $w=2.48e-07 $l=2.75e-07 $layer=LI1_cond $X=11.29 $Y=0.085
+ $X2=11.29 $Y2=0.36
r275 43 65 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0
r276 43 45 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=4.09 $Y=0.085
+ $X2=4.09 $Y2=0.36
r277 39 120 1.53834 $w=4.1e-07 $l=8.5e-08 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0
r278 39 41 8.29197 $w=4.08e-07 $l=2.95e-07 $layer=LI1_cond $X=3.145 $Y=0.085
+ $X2=3.145 $Y2=0.38
r279 38 117 7.34436 $w=1.7e-07 $l=1.33e-07 $layer=LI1_cond $X=2.29 $Y=0
+ $X2=2.157 $Y2=0
r280 37 120 9.97069 $w=1.7e-07 $l=2.05e-07 $layer=LI1_cond $X=2.94 $Y=0
+ $X2=3.145 $Y2=0
r281 37 38 42.4064 $w=1.68e-07 $l=6.5e-07 $layer=LI1_cond $X=2.94 $Y=0 $X2=2.29
+ $Y2=0
r282 33 117 0.195364 $w=2.65e-07 $l=8.5e-08 $layer=LI1_cond $X=2.157 $Y=0.085
+ $X2=2.157 $Y2=0
r283 33 35 12.8291 $w=2.63e-07 $l=2.95e-07 $layer=LI1_cond $X=2.157 $Y=0.085
+ $X2=2.157 $Y2=0.38
r284 32 114 8.44605 $w=6.22e-07 $l=2.83417e-07 $layer=LI1_cond $X=0.75 $Y=0
+ $X2=0.69 $Y2=0.255
r285 31 117 7.34436 $w=1.7e-07 $l=1.32e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=2.157 $Y2=0
r286 31 32 83.1818 $w=1.68e-07 $l=1.275e-06 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=0.75 $Y2=0
r287 10 61 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=14.68
+ $Y=0.235 $X2=14.865 $Y2=0.38
r288 9 57 91 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=2 $X=13.69
+ $Y=0.235 $X2=13.875 $Y2=0.38
r289 8 53 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=12.695
+ $Y=0.235 $X2=12.855 $Y2=0.36
r290 7 49 182 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_NDIFF $count=1 $X=10.965
+ $Y=0.235 $X2=11.25 $Y2=0.36
r291 6 130 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=7.745
+ $Y=0.235 $X2=7.89 $Y2=0.36
r292 5 127 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.295
+ $Y=0.235 $X2=6.43 $Y2=0.38
r293 4 45 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=3.955
+ $Y=0.235 $X2=4.09 $Y2=0.36
r294 3 41 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.965
+ $Y=0.235 $X2=3.1 $Y2=0.38
r295 2 35 182 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=1 $X=1.895
+ $Y=0.235 $X2=2.11 $Y2=0.38
r296 1 112 182 $w=1.7e-07 $l=2.498e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.43
.ends

