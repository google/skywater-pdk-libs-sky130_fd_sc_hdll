* File: sky130_fd_sc_hdll__buf_16.pex.spice
* Created: Thu Aug 27 19:00:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__BUF_16%A 3 5 7 10 12 14 17 19 21 24 26 28 31 33 35
+ 36 38 41 43 44 62 63 68 71
c124 62 0 1.34672e-19 $X=2.5 $Y=1.16
c125 41 0 1.25206e-19 $X=2.87 $Y=0.56
c126 36 0 1.26528e-19 $X=2.845 $Y=1.41
r127 63 64 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.845 $Y=1.217
+ $X2=2.87 $Y2=1.217
r128 61 63 51.3241 $w=3.24e-07 $l=3.45e-07 $layer=POLY_cond $X=2.5 $Y=1.217
+ $X2=2.845 $Y2=1.217
r129 61 62 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=2.5
+ $Y=1.16 $X2=2.5 $Y2=1.16
r130 59 61 18.5957 $w=3.24e-07 $l=1.25e-07 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.5 $Y2=1.217
r131 58 59 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=2.35 $Y=1.217
+ $X2=2.375 $Y2=1.217
r132 57 58 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=2.35 $Y2=1.217
r133 56 57 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.88 $Y=1.217
+ $X2=1.905 $Y2=1.217
r134 55 56 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=1.435 $Y=1.217
+ $X2=1.88 $Y2=1.217
r135 54 55 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.217
+ $X2=1.435 $Y2=1.217
r136 53 54 66.2006 $w=3.24e-07 $l=4.45e-07 $layer=POLY_cond $X=0.965 $Y=1.217
+ $X2=1.41 $Y2=1.217
r137 52 53 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.94 $Y=1.217
+ $X2=0.965 $Y2=1.217
r138 51 68 56.2864 $w=1.98e-07 $l=1.015e-06 $layer=LI1_cond $X=0.6 $Y=1.175
+ $X2=1.615 $Y2=1.175
r139 50 52 50.5802 $w=3.24e-07 $l=3.4e-07 $layer=POLY_cond $X=0.6 $Y=1.217
+ $X2=0.94 $Y2=1.217
r140 50 51 48.4267 $w=1.7e-07 $l=5.1e-07 $layer=licon1_POLY $count=3 $X=0.6
+ $Y=1.16 $X2=0.6 $Y2=1.16
r141 48 50 15.6204 $w=3.24e-07 $l=1.05e-07 $layer=POLY_cond $X=0.495 $Y=1.217
+ $X2=0.6 $Y2=1.217
r142 47 48 3.71914 $w=3.24e-07 $l=2.5e-08 $layer=POLY_cond $X=0.47 $Y=1.217
+ $X2=0.495 $Y2=1.217
r143 44 62 23.2909 $w=1.98e-07 $l=4.2e-07 $layer=LI1_cond $X=2.08 $Y=1.175
+ $X2=2.5 $Y2=1.175
r144 44 71 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=2.08 $Y=1.175
+ $X2=2.075 $Y2=1.175
r145 43 71 25.2318 $w=1.98e-07 $l=4.55e-07 $layer=LI1_cond $X=1.62 $Y=1.175
+ $X2=2.075 $Y2=1.175
r146 43 68 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=1.62 $Y=1.175
+ $X2=1.615 $Y2=1.175
r147 39 64 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r148 39 41 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r149 36 63 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.217
r150 36 38 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.845 $Y=1.41
+ $X2=2.845 $Y2=1.985
r151 33 59 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r152 33 35 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r153 29 58 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=1.217
r154 29 31 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.35 $Y=1.025
+ $X2=2.35 $Y2=0.56
r155 26 57 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r156 26 28 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r157 22 56 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=1.217
r158 22 24 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.88 $Y=1.025
+ $X2=1.88 $Y2=0.56
r159 19 55 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.217
r160 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r161 15 54 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=1.217
r162 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.41 $Y=1.025
+ $X2=1.41 $Y2=0.56
r163 12 53 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.217
r164 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r165 8 52 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=1.217
r166 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.94 $Y=1.025
+ $X2=0.94 $Y2=0.56
r167 5 48 16.5046 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r168 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r169 1 47 20.7868 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=1.217
r170 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_16%A_109_47# 1 2 3 4 5 6 21 23 25 28 30 32 35
+ 37 39 42 44 46 49 51 53 56 58 60 63 65 67 70 72 74 77 79 81 84 86 88 91 93 95
+ 98 100 102 105 107 109 112 114 116 119 121 123 124 126 129 133 137 141 142 143
+ 144 147 151 155 157 161 165 169 171 174 176 182 185 186 187 188 189 222
c459 222 0 1.34672e-19 $X=10.365 $Y=1.217
r460 222 223 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=10.365 $Y=1.217
+ $X2=10.39 $Y2=1.217
r461 221 222 70.7937 $w=3.2e-07 $l=4.7e-07 $layer=POLY_cond $X=9.895 $Y=1.217
+ $X2=10.365 $Y2=1.217
r462 218 219 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=9.425 $Y=1.217
+ $X2=9.87 $Y2=1.217
r463 217 218 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=9.4 $Y=1.217
+ $X2=9.425 $Y2=1.217
r464 216 217 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.955 $Y=1.217
+ $X2=9.4 $Y2=1.217
r465 215 216 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.93 $Y=1.217
+ $X2=8.955 $Y2=1.217
r466 214 215 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.485 $Y=1.217
+ $X2=8.93 $Y2=1.217
r467 213 214 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=8.46 $Y=1.217
+ $X2=8.485 $Y2=1.217
r468 212 213 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=8.015 $Y=1.217
+ $X2=8.46 $Y2=1.217
r469 211 212 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.99 $Y=1.217
+ $X2=8.015 $Y2=1.217
r470 210 211 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.545 $Y=1.217
+ $X2=7.99 $Y2=1.217
r471 209 210 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.52 $Y=1.217
+ $X2=7.545 $Y2=1.217
r472 208 209 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=7.075 $Y=1.217
+ $X2=7.52 $Y2=1.217
r473 207 208 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=7.05 $Y=1.217
+ $X2=7.075 $Y2=1.217
r474 206 207 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.605 $Y=1.217
+ $X2=7.05 $Y2=1.217
r475 205 206 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.58 $Y=1.217
+ $X2=6.605 $Y2=1.217
r476 204 205 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=6.135 $Y=1.217
+ $X2=6.58 $Y2=1.217
r477 203 204 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=6.11 $Y=1.217
+ $X2=6.135 $Y2=1.217
r478 202 203 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=5.665 $Y=1.217
+ $X2=6.11 $Y2=1.217
r479 201 202 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=5.64 $Y=1.217
+ $X2=5.665 $Y2=1.217
r480 200 201 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=5.195 $Y=1.217
+ $X2=5.64 $Y2=1.217
r481 199 200 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=5.17 $Y=1.217
+ $X2=5.195 $Y2=1.217
r482 198 199 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=4.725 $Y=1.217
+ $X2=5.17 $Y2=1.217
r483 197 198 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=4.7 $Y=1.217
+ $X2=4.725 $Y2=1.217
r484 196 197 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=4.255 $Y=1.217
+ $X2=4.7 $Y2=1.217
r485 195 196 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=4.23 $Y=1.217
+ $X2=4.255 $Y2=1.217
r486 194 195 67.0281 $w=3.2e-07 $l=4.45e-07 $layer=POLY_cond $X=3.785 $Y=1.217
+ $X2=4.23 $Y2=1.217
r487 193 194 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=3.76 $Y=1.217
+ $X2=3.785 $Y2=1.217
r488 190 191 3.76562 $w=3.2e-07 $l=2.5e-08 $layer=POLY_cond $X=3.29 $Y=1.217
+ $X2=3.315 $Y2=1.217
r489 183 221 2.25938 $w=3.2e-07 $l=1.5e-08 $layer=POLY_cond $X=9.88 $Y=1.217
+ $X2=9.895 $Y2=1.217
r490 183 219 1.50625 $w=3.2e-07 $l=1e-08 $layer=POLY_cond $X=9.88 $Y=1.217
+ $X2=9.87 $Y2=1.217
r491 182 183 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=9.88
+ $Y=1.16 $X2=9.88 $Y2=1.16
r492 180 193 54.225 $w=3.2e-07 $l=3.6e-07 $layer=POLY_cond $X=3.4 $Y=1.217
+ $X2=3.76 $Y2=1.217
r493 180 191 12.8031 $w=3.2e-07 $l=8.5e-08 $layer=POLY_cond $X=3.4 $Y=1.217
+ $X2=3.315 $Y2=1.217
r494 179 182 359.345 $w=1.98e-07 $l=6.48e-06 $layer=LI1_cond $X=3.4 $Y=1.175
+ $X2=9.88 $Y2=1.175
r495 179 180 16.1422 $w=1.7e-07 $l=1.53e-06 $layer=licon1_POLY $count=9 $X=3.4
+ $Y=1.16 $X2=3.4 $Y2=1.16
r496 177 189 0.866423 $w=2e-07 $l=8.8e-08 $layer=LI1_cond $X=3.165 $Y=1.175
+ $X2=3.077 $Y2=1.175
r497 177 179 13.0318 $w=1.98e-07 $l=2.35e-07 $layer=LI1_cond $X=3.165 $Y=1.175
+ $X2=3.4 $Y2=1.175
r498 175 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=3.077 $Y=1.275
+ $X2=3.077 $Y2=1.175
r499 175 176 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=3.077 $Y=1.275
+ $X2=3.077 $Y2=1.445
r500 174 189 5.7647 $w=1.75e-07 $l=1e-07 $layer=LI1_cond $X=3.077 $Y=1.075
+ $X2=3.077 $Y2=1.175
r501 173 174 10.774 $w=1.73e-07 $l=1.7e-07 $layer=LI1_cond $X=3.077 $Y=0.905
+ $X2=3.077 $Y2=1.075
r502 172 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=1.53
+ $X2=2.585 $Y2=1.53
r503 171 176 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.99 $Y=1.53
+ $X2=3.077 $Y2=1.445
r504 171 172 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.99 $Y=1.53
+ $X2=2.775 $Y2=1.53
r505 170 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.775 $Y=0.82
+ $X2=2.585 $Y2=0.82
r506 169 173 6.81835 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=2.99 $Y=0.82
+ $X2=3.077 $Y2=0.905
r507 169 170 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.99 $Y=0.82
+ $X2=2.775 $Y2=0.82
r508 165 167 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=2.585 $Y=1.63
+ $X2=2.585 $Y2=2.31
r509 163 188 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=1.615
+ $X2=2.585 $Y2=1.53
r510 163 165 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=2.585 $Y=1.615
+ $X2=2.585 $Y2=1.63
r511 159 187 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.585 $Y=0.735
+ $X2=2.585 $Y2=0.82
r512 159 161 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.585 $Y=0.735
+ $X2=2.585 $Y2=0.4
r513 158 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=1.53
+ $X2=1.645 $Y2=1.53
r514 157 188 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=1.53
+ $X2=2.585 $Y2=1.53
r515 157 158 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=1.53
+ $X2=1.835 $Y2=1.53
r516 156 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=0.82
+ $X2=1.645 $Y2=0.82
r517 155 187 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0.82
+ $X2=2.585 $Y2=0.82
r518 155 156 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=2.395 $Y=0.82
+ $X2=1.835 $Y2=0.82
r519 151 153 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.645 $Y=1.63
+ $X2=1.645 $Y2=2.31
r520 149 186 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=1.615
+ $X2=1.645 $Y2=1.53
r521 149 151 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=1.645 $Y=1.615
+ $X2=1.645 $Y2=1.63
r522 145 185 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.645 $Y=0.735
+ $X2=1.645 $Y2=0.82
r523 145 147 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=1.645 $Y=0.735
+ $X2=1.645 $Y2=0.4
r524 143 186 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=1.53
+ $X2=1.645 $Y2=1.53
r525 143 144 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=1.53
+ $X2=0.895 $Y2=1.53
r526 141 185 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=0.82
+ $X2=1.645 $Y2=0.82
r527 141 142 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=1.455 $Y=0.82
+ $X2=0.895 $Y2=0.82
r528 137 139 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.705 $Y=1.63
+ $X2=0.705 $Y2=2.31
r529 135 144 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.705 $Y=1.615
+ $X2=0.895 $Y2=1.53
r530 135 137 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=0.705 $Y=1.615
+ $X2=0.705 $Y2=1.63
r531 131 142 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.895 $Y2=0.82
r532 131 133 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=0.705 $Y=0.735
+ $X2=0.705 $Y2=0.4
r533 127 223 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=10.39 $Y=1.025
+ $X2=10.39 $Y2=1.217
r534 127 129 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=10.39 $Y=1.025
+ $X2=10.39 $Y2=0.56
r535 124 222 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.217
r536 124 126 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=10.365 $Y=1.41
+ $X2=10.365 $Y2=1.985
r537 121 221 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.217
r538 121 123 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.895 $Y=1.41
+ $X2=9.895 $Y2=1.985
r539 117 219 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.87 $Y=1.025
+ $X2=9.87 $Y2=1.217
r540 117 119 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.87 $Y=1.025
+ $X2=9.87 $Y2=0.56
r541 114 218 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.217
r542 114 116 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=9.425 $Y=1.41
+ $X2=9.425 $Y2=1.985
r543 110 217 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=9.4 $Y=1.025
+ $X2=9.4 $Y2=1.217
r544 110 112 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=9.4 $Y=1.025
+ $X2=9.4 $Y2=0.56
r545 107 216 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.217
r546 107 109 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.955 $Y=1.41
+ $X2=8.955 $Y2=1.985
r547 103 215 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.93 $Y=1.025
+ $X2=8.93 $Y2=1.217
r548 103 105 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.93 $Y=1.025
+ $X2=8.93 $Y2=0.56
r549 100 214 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.217
r550 100 102 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.485 $Y=1.41
+ $X2=8.485 $Y2=1.985
r551 96 213 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=8.46 $Y=1.025
+ $X2=8.46 $Y2=1.217
r552 96 98 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=8.46 $Y=1.025
+ $X2=8.46 $Y2=0.56
r553 93 212 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.217
r554 93 95 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=8.015 $Y=1.41
+ $X2=8.015 $Y2=1.985
r555 89 211 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.99 $Y=1.025
+ $X2=7.99 $Y2=1.217
r556 89 91 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.99 $Y=1.025
+ $X2=7.99 $Y2=0.56
r557 86 210 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.217
r558 86 88 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.545 $Y=1.41
+ $X2=7.545 $Y2=1.985
r559 82 209 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=1.217
r560 82 84 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.52 $Y=1.025
+ $X2=7.52 $Y2=0.56
r561 79 208 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.217
r562 79 81 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.075 $Y=1.41
+ $X2=7.075 $Y2=1.985
r563 75 207 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=1.217
r564 75 77 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.05 $Y=1.025
+ $X2=7.05 $Y2=0.56
r565 72 206 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.217
r566 72 74 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.605 $Y=1.41
+ $X2=6.605 $Y2=1.985
r567 68 205 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=1.217
r568 68 70 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.58 $Y=1.025
+ $X2=6.58 $Y2=0.56
r569 65 204 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.217
r570 65 67 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.135 $Y=1.41
+ $X2=6.135 $Y2=1.985
r571 61 203 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=1.217
r572 61 63 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.11 $Y=1.025
+ $X2=6.11 $Y2=0.56
r573 58 202 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.217
r574 58 60 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.665 $Y=1.41
+ $X2=5.665 $Y2=1.985
r575 54 201 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=1.217
r576 54 56 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.64 $Y=1.025
+ $X2=5.64 $Y2=0.56
r577 51 200 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.217
r578 51 53 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.195 $Y=1.41
+ $X2=5.195 $Y2=1.985
r579 47 199 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=1.217
r580 47 49 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.17 $Y=1.025
+ $X2=5.17 $Y2=0.56
r581 44 198 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.217
r582 44 46 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.725 $Y=1.41
+ $X2=4.725 $Y2=1.985
r583 40 197 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=1.217
r584 40 42 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.7 $Y=1.025
+ $X2=4.7 $Y2=0.56
r585 37 196 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.217
r586 37 39 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.255 $Y=1.41
+ $X2=4.255 $Y2=1.985
r587 33 195 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=1.217
r588 33 35 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.23 $Y=1.025
+ $X2=4.23 $Y2=0.56
r589 30 194 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.217
r590 30 32 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.785 $Y=1.41
+ $X2=3.785 $Y2=1.985
r591 26 193 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=1.217
r592 26 28 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.76 $Y=1.025
+ $X2=3.76 $Y2=0.56
r593 23 191 16.2157 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.217
r594 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.315 $Y=1.41
+ $X2=3.315 $Y2=1.985
r595 19 190 20.4921 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r596 19 21 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r597 6 167 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.31
r598 6 165 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=1.63
r599 5 153 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.31
r600 5 151 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.63
r601 4 139 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.31
r602 4 137 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.63
r603 3 161 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=2.425
+ $Y=0.235 $X2=2.61 $Y2=0.4
r604 2 147 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.4
r605 1 133 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_16%VPWR 1 2 3 4 5 6 7 8 9 10 11 12 37 39 43 47
+ 49 53 57 61 65 69 73 77 81 85 89 92 93 95 96 98 99 101 102 104 105 107 108 110
+ 111 113 114 116 117 118 149 150 156 159
r187 159 160 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r188 157 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r189 156 157 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r190 149 150 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=2.72
+ $X2=11.27 $Y2=2.72
r191 147 150 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=2.72
+ $X2=11.27 $Y2=2.72
r192 146 147 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=2.72
+ $X2=10.35 $Y2=2.72
r193 144 147 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=2.72
+ $X2=10.35 $Y2=2.72
r194 143 144 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=2.72
+ $X2=9.43 $Y2=2.72
r195 141 144 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=2.72
+ $X2=9.43 $Y2=2.72
r196 140 141 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=2.72
+ $X2=8.51 $Y2=2.72
r197 138 141 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=2.72
+ $X2=8.51 $Y2=2.72
r198 137 138 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r199 135 138 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=2.72
+ $X2=7.59 $Y2=2.72
r200 134 135 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r201 132 135 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=2.72
+ $X2=6.67 $Y2=2.72
r202 131 132 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r203 129 132 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r204 128 129 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r205 126 129 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r206 125 126 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r207 123 126 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r208 123 160 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r209 122 123 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r210 120 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.14 $Y2=2.72
r211 120 122 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=2.72
+ $X2=2.99 $Y2=2.72
r212 118 157 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r213 118 153 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r214 116 146 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.515 $Y=2.72
+ $X2=10.35 $Y2=2.72
r215 116 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=2.72
+ $X2=10.6 $Y2=2.72
r216 115 149 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=10.685 $Y=2.72
+ $X2=11.27 $Y2=2.72
r217 115 117 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.685 $Y=2.72
+ $X2=10.6 $Y2=2.72
r218 113 143 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=9.575 $Y=2.72
+ $X2=9.43 $Y2=2.72
r219 113 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=2.72
+ $X2=9.66 $Y2=2.72
r220 112 146 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.745 $Y=2.72
+ $X2=10.35 $Y2=2.72
r221 112 114 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.745 $Y=2.72
+ $X2=9.66 $Y2=2.72
r222 110 140 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.635 $Y=2.72
+ $X2=8.51 $Y2=2.72
r223 110 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.635 $Y=2.72
+ $X2=8.72 $Y2=2.72
r224 109 143 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.805 $Y=2.72
+ $X2=9.43 $Y2=2.72
r225 109 111 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.805 $Y=2.72
+ $X2=8.72 $Y2=2.72
r226 107 137 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.695 $Y=2.72
+ $X2=7.59 $Y2=2.72
r227 107 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.695 $Y=2.72
+ $X2=7.78 $Y2=2.72
r228 106 140 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=7.865 $Y=2.72
+ $X2=8.51 $Y2=2.72
r229 106 108 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=2.72
+ $X2=7.78 $Y2=2.72
r230 104 134 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.67 $Y2=2.72
r231 104 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=2.72
+ $X2=6.84 $Y2=2.72
r232 103 137 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.925 $Y=2.72
+ $X2=7.59 $Y2=2.72
r233 103 105 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=2.72
+ $X2=6.84 $Y2=2.72
r234 101 131 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=5.75 $Y2=2.72
r235 101 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.815 $Y=2.72
+ $X2=5.9 $Y2=2.72
r236 100 134 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=6.67 $Y2=2.72
r237 100 102 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=2.72
+ $X2=5.9 $Y2=2.72
r238 98 128 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.83 $Y2=2.72
r239 98 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=2.72
+ $X2=4.96 $Y2=2.72
r240 97 131 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=5.75 $Y2=2.72
r241 97 99 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=2.72
+ $X2=4.96 $Y2=2.72
r242 95 125 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=3.91 $Y2=2.72
r243 95 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=2.72
+ $X2=4.02 $Y2=2.72
r244 94 128 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.83 $Y2=2.72
r245 94 96 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=2.72
+ $X2=4.02 $Y2=2.72
r246 92 122 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=2.99 $Y2=2.72
r247 92 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=2.72
+ $X2=3.08 $Y2=2.72
r248 91 125 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.91 $Y2=2.72
r249 91 93 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=2.72
+ $X2=3.08 $Y2=2.72
r250 87 117 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2.72
r251 87 89 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=10.6 $Y=2.635
+ $X2=10.6 $Y2=2
r252 83 114 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2.72
r253 83 85 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=9.66 $Y=2.635
+ $X2=9.66 $Y2=2
r254 79 111 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2.72
r255 79 81 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=8.72 $Y=2.635
+ $X2=8.72 $Y2=2
r256 75 108 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2.72
r257 75 77 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=7.78 $Y=2.635
+ $X2=7.78 $Y2=2
r258 71 105 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2.72
r259 71 73 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.84 $Y=2.635
+ $X2=6.84 $Y2=2
r260 67 102 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2.72
r261 67 69 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=5.9 $Y=2.635
+ $X2=5.9 $Y2=2
r262 63 99 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2.72
r263 63 65 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.96 $Y=2.635
+ $X2=4.96 $Y2=2
r264 59 96 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2.72
r265 59 61 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.02 $Y=2.635
+ $X2=4.02 $Y2=2
r266 55 93 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2.72
r267 55 57 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=3.08 $Y=2.635
+ $X2=3.08 $Y2=2
r268 51 159 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2.72
r269 51 53 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.14 $Y=2.635
+ $X2=2.14 $Y2=2
r270 50 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.72
+ $X2=1.2 $Y2=2.72
r271 49 159 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.14 $Y2=2.72
r272 49 50 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.285 $Y2=2.72
r273 45 156 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2.72
r274 45 47 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.2 $Y=2.635
+ $X2=1.2 $Y2=2
r275 44 153 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=2.72
+ $X2=0.172 $Y2=2.72
r276 43 156 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=1.2 $Y2=2.72
r277 43 44 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.72
+ $X2=0.345 $Y2=2.72
r278 39 42 44.3636 $w=1.68e-07 $l=6.8e-07 $layer=LI1_cond $X=0.26 $Y=1.66
+ $X2=0.26 $Y2=2.34
r279 37 153 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.172 $Y2=2.72
r280 37 42 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=2.635
+ $X2=0.26 $Y2=2.34
r281 12 89 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=10.455
+ $Y=1.485 $X2=10.6 $Y2=2
r282 11 85 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=9.515
+ $Y=1.485 $X2=9.66 $Y2=2
r283 10 81 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=8.575
+ $Y=1.485 $X2=8.72 $Y2=2
r284 9 77 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=7.635
+ $Y=1.485 $X2=7.78 $Y2=2
r285 8 73 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.695
+ $Y=1.485 $X2=6.84 $Y2=2
r286 7 69 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=5.755
+ $Y=1.485 $X2=5.9 $Y2=2
r287 6 65 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.815
+ $Y=1.485 $X2=4.96 $Y2=2
r288 5 61 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.875
+ $Y=1.485 $X2=4.02 $Y2=2
r289 4 57 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.935
+ $Y=1.485 $X2=3.08 $Y2=2
r290 3 53 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2
r291 2 47 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=2
r292 1 42 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r293 1 39 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_16%X 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 49
+ 50 53 57 58 59 60 61 62 65 69 71 73 74 77 81 83 87 91 95 97 101 105 109 111
+ 115 119 123 125 129 133 137 139 143 145 155 156 159 160 161 162 163 164 165
+ 166 167 168 169 171 173 174 175 176 184 191
c370 60 0 1.26528e-19 $X=3.715 $Y=1.53
c371 58 0 1.25206e-19 $X=3.715 $Y=0.82
r372 191 194 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=10.105 $Y=1.63
+ $X2=10.105 $Y2=2.31
r373 175 181 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.105 $Y=1.53
+ $X2=10.295 $Y2=1.53
r374 175 191 0.501524 $w=4.08e-07 $l=1.5e-08 $layer=LI1_cond $X=10.105 $Y=1.615
+ $X2=10.105 $Y2=1.63
r375 175 184 10.1123 $w=1.68e-07 $l=1.55e-07 $layer=LI1_cond $X=10.365 $Y=1.53
+ $X2=10.52 $Y2=1.53
r376 175 181 4.56684 $w=1.68e-07 $l=7e-08 $layer=LI1_cond $X=10.365 $Y=1.53
+ $X2=10.295 $Y2=1.53
r377 173 184 7.50267 $w=1.68e-07 $l=1.15e-07 $layer=LI1_cond $X=10.635 $Y=1.53
+ $X2=10.52 $Y2=1.53
r378 173 174 4.42191 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=10.635 $Y=1.53
+ $X2=10.885 $Y2=1.53
r379 172 176 6.1 $w=4.98e-07 $l=2.55e-07 $layer=LI1_cond $X=10.885 $Y=1.445
+ $X2=10.885 $Y2=1.19
r380 172 174 2.49074 $w=3.87e-07 $l=8.5e-08 $layer=LI1_cond $X=10.885 $Y=1.445
+ $X2=10.885 $Y2=1.53
r381 170 176 6.81765 $w=4.98e-07 $l=2.85e-07 $layer=LI1_cond $X=10.885 $Y=0.905
+ $X2=10.885 $Y2=1.19
r382 170 171 2.49074 $w=3.87e-07 $l=8.5e-08 $layer=LI1_cond $X=10.885 $Y=0.905
+ $X2=10.885 $Y2=0.82
r383 146 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=10.295 $Y=0.82
+ $X2=10.105 $Y2=0.82
r384 145 171 4.42191 $w=1.7e-07 $l=2.5e-07 $layer=LI1_cond $X=10.635 $Y=0.82
+ $X2=10.885 $Y2=0.82
r385 145 146 22.1818 $w=1.68e-07 $l=3.4e-07 $layer=LI1_cond $X=10.635 $Y=0.82
+ $X2=10.295 $Y2=0.82
r386 141 169 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=10.105 $Y=0.735
+ $X2=10.105 $Y2=0.82
r387 141 143 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=10.105 $Y=0.735
+ $X2=10.105 $Y2=0.4
r388 140 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.355 $Y=1.53
+ $X2=9.165 $Y2=1.53
r389 139 175 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.915 $Y=1.53
+ $X2=10.105 $Y2=1.53
r390 139 140 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.915 $Y=1.53
+ $X2=9.355 $Y2=1.53
r391 138 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.355 $Y=0.82
+ $X2=9.165 $Y2=0.82
r392 137 169 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=9.915 $Y=0.82
+ $X2=10.105 $Y2=0.82
r393 137 138 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=9.915 $Y=0.82
+ $X2=9.355 $Y2=0.82
r394 133 135 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=9.165 $Y=1.63
+ $X2=9.165 $Y2=2.31
r395 131 168 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=1.615
+ $X2=9.165 $Y2=1.53
r396 131 133 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=9.165 $Y=1.615
+ $X2=9.165 $Y2=1.63
r397 127 167 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=9.165 $Y=0.735
+ $X2=9.165 $Y2=0.82
r398 127 129 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=9.165 $Y=0.735
+ $X2=9.165 $Y2=0.4
r399 126 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.415 $Y=1.53
+ $X2=8.225 $Y2=1.53
r400 125 168 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.975 $Y=1.53
+ $X2=9.165 $Y2=1.53
r401 125 126 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.975 $Y=1.53
+ $X2=8.415 $Y2=1.53
r402 124 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.415 $Y=0.82
+ $X2=8.225 $Y2=0.82
r403 123 167 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.975 $Y=0.82
+ $X2=9.165 $Y2=0.82
r404 123 124 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.975 $Y=0.82
+ $X2=8.415 $Y2=0.82
r405 119 121 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=8.225 $Y=1.63
+ $X2=8.225 $Y2=2.31
r406 117 166 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.225 $Y=1.615
+ $X2=8.225 $Y2=1.53
r407 117 119 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=8.225 $Y=1.615
+ $X2=8.225 $Y2=1.63
r408 113 165 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=8.225 $Y=0.735
+ $X2=8.225 $Y2=0.82
r409 113 115 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=8.225 $Y=0.735
+ $X2=8.225 $Y2=0.4
r410 112 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.475 $Y=1.53
+ $X2=7.285 $Y2=1.53
r411 111 166 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.035 $Y=1.53
+ $X2=8.225 $Y2=1.53
r412 111 112 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.035 $Y=1.53
+ $X2=7.475 $Y2=1.53
r413 110 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.475 $Y=0.82
+ $X2=7.285 $Y2=0.82
r414 109 165 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=8.035 $Y=0.82
+ $X2=8.225 $Y2=0.82
r415 109 110 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=8.035 $Y=0.82
+ $X2=7.475 $Y2=0.82
r416 105 107 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=7.285 $Y=1.63
+ $X2=7.285 $Y2=2.31
r417 103 164 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.285 $Y=1.615
+ $X2=7.285 $Y2=1.53
r418 103 105 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=7.285 $Y=1.615
+ $X2=7.285 $Y2=1.63
r419 99 163 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=7.285 $Y=0.735
+ $X2=7.285 $Y2=0.82
r420 99 101 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=7.285 $Y=0.735
+ $X2=7.285 $Y2=0.4
r421 98 162 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.535 $Y=1.53
+ $X2=6.345 $Y2=1.53
r422 97 164 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.095 $Y=1.53
+ $X2=7.285 $Y2=1.53
r423 97 98 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.095 $Y=1.53
+ $X2=6.535 $Y2=1.53
r424 96 161 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.535 $Y=0.82
+ $X2=6.345 $Y2=0.82
r425 95 163 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=7.095 $Y=0.82
+ $X2=7.285 $Y2=0.82
r426 95 96 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=7.095 $Y=0.82
+ $X2=6.535 $Y2=0.82
r427 91 93 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=6.345 $Y=1.63
+ $X2=6.345 $Y2=2.31
r428 89 162 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=1.615
+ $X2=6.345 $Y2=1.53
r429 89 91 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=6.345 $Y=1.615
+ $X2=6.345 $Y2=1.63
r430 85 161 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=6.345 $Y=0.735
+ $X2=6.345 $Y2=0.82
r431 85 87 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.345 $Y=0.735
+ $X2=6.345 $Y2=0.4
r432 84 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.595 $Y=1.53
+ $X2=5.405 $Y2=1.53
r433 83 162 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.155 $Y=1.53
+ $X2=6.345 $Y2=1.53
r434 83 84 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.155 $Y=1.53
+ $X2=5.595 $Y2=1.53
r435 82 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.595 $Y=0.82
+ $X2=5.405 $Y2=0.82
r436 81 161 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=6.155 $Y=0.82
+ $X2=6.345 $Y2=0.82
r437 81 82 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=6.155 $Y=0.82
+ $X2=5.595 $Y2=0.82
r438 77 79 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=5.405 $Y=1.63
+ $X2=5.405 $Y2=2.31
r439 75 160 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=1.615
+ $X2=5.405 $Y2=1.53
r440 75 77 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=5.405 $Y=1.615
+ $X2=5.405 $Y2=1.63
r441 74 159 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=5.405 $Y=0.735
+ $X2=5.405 $Y2=0.82
r442 73 158 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=5.405 $Y=0.45
+ $X2=5.405 $Y2=0.4
r443 73 74 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=5.405 $Y=0.45
+ $X2=5.405 $Y2=0.735
r444 72 156 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=1.53
+ $X2=4.465 $Y2=1.53
r445 71 160 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.215 $Y=1.53
+ $X2=5.405 $Y2=1.53
r446 71 72 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=1.53
+ $X2=4.655 $Y2=1.53
r447 70 155 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.655 $Y=0.82
+ $X2=4.465 $Y2=0.82
r448 69 159 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.215 $Y=0.82
+ $X2=5.405 $Y2=0.82
r449 69 70 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=5.215 $Y=0.82
+ $X2=4.655 $Y2=0.82
r450 65 67 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=4.465 $Y=1.63
+ $X2=4.465 $Y2=2.31
r451 63 156 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=1.615
+ $X2=4.465 $Y2=1.53
r452 63 65 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=4.465 $Y=1.615
+ $X2=4.465 $Y2=1.63
r453 62 155 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=4.465 $Y=0.735
+ $X2=4.465 $Y2=0.82
r454 61 154 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=4.465 $Y=0.45
+ $X2=4.465 $Y2=0.4
r455 61 62 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=4.465 $Y=0.45
+ $X2=4.465 $Y2=0.735
r456 59 156 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=1.53
+ $X2=4.465 $Y2=1.53
r457 59 60 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.275 $Y=1.53
+ $X2=3.715 $Y2=1.53
r458 57 155 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.275 $Y=0.82
+ $X2=4.465 $Y2=0.82
r459 57 58 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.275 $Y=0.82
+ $X2=3.715 $Y2=0.82
r460 53 55 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=3.525 $Y=1.63
+ $X2=3.525 $Y2=2.31
r461 51 60 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.525 $Y=1.615
+ $X2=3.715 $Y2=1.53
r462 51 53 0.454912 $w=3.78e-07 $l=1.5e-08 $layer=LI1_cond $X=3.525 $Y=1.615
+ $X2=3.525 $Y2=1.63
r463 50 58 8.19669 $w=1.7e-07 $l=2.28583e-07 $layer=LI1_cond $X=3.525 $Y=0.735
+ $X2=3.715 $Y2=0.82
r464 49 152 1.60526 $w=3.8e-07 $l=5e-08 $layer=LI1_cond $X=3.525 $Y=0.45
+ $X2=3.525 $Y2=0.4
r465 49 50 8.64332 $w=3.78e-07 $l=2.85e-07 $layer=LI1_cond $X=3.525 $Y=0.45
+ $X2=3.525 $Y2=0.735
r466 16 194 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=2.31
r467 16 191 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.985
+ $Y=1.485 $X2=10.13 $Y2=1.63
r468 15 135 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=2.31
r469 15 133 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=9.045
+ $Y=1.485 $X2=9.19 $Y2=1.63
r470 14 121 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=2.31
r471 14 119 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=8.105
+ $Y=1.485 $X2=8.25 $Y2=1.63
r472 13 107 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=2.31
r473 13 105 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=7.165
+ $Y=1.485 $X2=7.31 $Y2=1.63
r474 12 93 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=2.31
r475 12 91 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=6.225
+ $Y=1.485 $X2=6.37 $Y2=1.63
r476 11 79 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=2.31
r477 11 77 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=5.285
+ $Y=1.485 $X2=5.43 $Y2=1.63
r478 10 67 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=2.31
r479 10 65 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=4.345
+ $Y=1.485 $X2=4.49 $Y2=1.63
r480 9 55 400 $w=1.7e-07 $l=8.94567e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=2.31
r481 9 53 400 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.405
+ $Y=1.485 $X2=3.55 $Y2=1.63
r482 8 143 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.945
+ $Y=0.235 $X2=10.13 $Y2=0.4
r483 7 129 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=9.005
+ $Y=0.235 $X2=9.19 $Y2=0.4
r484 6 115 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=8.065
+ $Y=0.235 $X2=8.25 $Y2=0.4
r485 5 101 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=7.125
+ $Y=0.235 $X2=7.31 $Y2=0.4
r486 4 87 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=6.185
+ $Y=0.235 $X2=6.37 $Y2=0.4
r487 3 158 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=5.245
+ $Y=0.235 $X2=5.43 $Y2=0.4
r488 2 154 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=4.305
+ $Y=0.235 $X2=4.49 $Y2=0.4
r489 1 152 91 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=2 $X=3.365
+ $Y=0.235 $X2=3.55 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__BUF_16%VGND 1 2 3 4 5 6 7 8 9 10 11 12 37 39 41 45
+ 47 51 55 59 63 67 71 75 79 83 87 90 91 93 94 96 97 99 100 102 103 105 106 108
+ 109 111 112 114 115 116 147 148 154 157
r207 157 158 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0
+ $X2=2.07 $Y2=0
r208 155 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0
+ $X2=2.07 $Y2=0
r209 154 155 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r210 147 148 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=11.27 $Y=0
+ $X2=11.27 $Y2=0
r211 145 148 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=10.35 $Y=0
+ $X2=11.27 $Y2=0
r212 144 145 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=10.35 $Y=0
+ $X2=10.35 $Y2=0
r213 142 145 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=9.43 $Y=0
+ $X2=10.35 $Y2=0
r214 141 142 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=9.43 $Y=0
+ $X2=9.43 $Y2=0
r215 139 142 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=8.51 $Y=0
+ $X2=9.43 $Y2=0
r216 138 139 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=8.51 $Y=0
+ $X2=8.51 $Y2=0
r217 136 139 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=7.59 $Y=0
+ $X2=8.51 $Y2=0
r218 135 136 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.59 $Y=0
+ $X2=7.59 $Y2=0
r219 133 136 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.67 $Y=0
+ $X2=7.59 $Y2=0
r220 132 133 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.67 $Y=0
+ $X2=6.67 $Y2=0
r221 130 133 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.75 $Y=0
+ $X2=6.67 $Y2=0
r222 129 130 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0
+ $X2=5.75 $Y2=0
r223 127 130 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0
+ $X2=5.75 $Y2=0
r224 126 127 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r225 124 127 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0
+ $X2=4.83 $Y2=0
r226 123 124 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0
+ $X2=3.91 $Y2=0
r227 121 124 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=3.91 $Y2=0
r228 121 158 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=0
+ $X2=2.07 $Y2=0
r229 120 121 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0
+ $X2=2.99 $Y2=0
r230 118 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.14 $Y2=0
r231 118 120 49.9091 $w=1.68e-07 $l=7.65e-07 $layer=LI1_cond $X=2.225 $Y=0
+ $X2=2.99 $Y2=0
r232 116 155 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0
+ $X2=1.15 $Y2=0
r233 116 151 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0
+ $X2=0.23 $Y2=0
r234 114 144 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.35 $Y2=0
r235 114 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.515 $Y=0
+ $X2=10.6 $Y2=0
r236 113 147 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=10.685 $Y=0
+ $X2=11.27 $Y2=0
r237 113 115 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.685 $Y=0
+ $X2=10.6 $Y2=0
r238 111 141 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=9.575 $Y=0
+ $X2=9.43 $Y2=0
r239 111 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.575 $Y=0
+ $X2=9.66 $Y2=0
r240 110 144 39.4706 $w=1.68e-07 $l=6.05e-07 $layer=LI1_cond $X=9.745 $Y=0
+ $X2=10.35 $Y2=0
r241 110 112 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.745 $Y=0
+ $X2=9.66 $Y2=0
r242 108 138 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.51 $Y2=0
r243 108 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.635 $Y=0
+ $X2=8.72 $Y2=0
r244 107 141 40.7754 $w=1.68e-07 $l=6.25e-07 $layer=LI1_cond $X=8.805 $Y=0
+ $X2=9.43 $Y2=0
r245 107 109 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.805 $Y=0
+ $X2=8.72 $Y2=0
r246 105 135 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=7.695 $Y=0
+ $X2=7.59 $Y2=0
r247 105 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.695 $Y=0
+ $X2=7.78 $Y2=0
r248 104 138 42.0802 $w=1.68e-07 $l=6.45e-07 $layer=LI1_cond $X=7.865 $Y=0
+ $X2=8.51 $Y2=0
r249 104 106 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.865 $Y=0
+ $X2=7.78 $Y2=0
r250 102 132 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.67 $Y2=0
r251 102 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.755 $Y=0
+ $X2=6.84 $Y2=0
r252 101 135 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=6.925 $Y=0
+ $X2=7.59 $Y2=0
r253 101 103 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.925 $Y=0
+ $X2=6.84 $Y2=0
r254 99 129 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=5.815 $Y=0
+ $X2=5.75 $Y2=0
r255 99 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.815 $Y=0 $X2=5.9
+ $Y2=0
r256 98 132 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=5.985 $Y=0
+ $X2=6.67 $Y2=0
r257 98 100 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.985 $Y=0 $X2=5.9
+ $Y2=0
r258 96 126 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=4.875 $Y=0
+ $X2=4.83 $Y2=0
r259 96 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.875 $Y=0 $X2=4.96
+ $Y2=0
r260 95 129 45.9947 $w=1.68e-07 $l=7.05e-07 $layer=LI1_cond $X=5.045 $Y=0
+ $X2=5.75 $Y2=0
r261 95 97 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.045 $Y=0 $X2=4.96
+ $Y2=0
r262 93 123 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=3.935 $Y=0
+ $X2=3.91 $Y2=0
r263 93 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.935 $Y=0 $X2=4.02
+ $Y2=0
r264 92 126 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=4.105 $Y=0
+ $X2=4.83 $Y2=0
r265 92 94 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.105 $Y=0 $X2=4.02
+ $Y2=0
r266 90 120 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=2.995 $Y=0 $X2=2.99
+ $Y2=0
r267 90 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.995 $Y=0 $X2=3.08
+ $Y2=0
r268 89 123 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=3.165 $Y=0
+ $X2=3.91 $Y2=0
r269 89 91 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.165 $Y=0 $X2=3.08
+ $Y2=0
r270 85 115 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=10.6 $Y=0.085
+ $X2=10.6 $Y2=0
r271 85 87 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=10.6 $Y=0.085
+ $X2=10.6 $Y2=0.4
r272 81 112 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0
r273 81 83 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=9.66 $Y=0.085
+ $X2=9.66 $Y2=0.4
r274 77 109 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=8.72 $Y=0.085
+ $X2=8.72 $Y2=0
r275 77 79 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=8.72 $Y=0.085
+ $X2=8.72 $Y2=0.4
r276 73 106 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=7.78 $Y=0.085
+ $X2=7.78 $Y2=0
r277 73 75 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=7.78 $Y=0.085
+ $X2=7.78 $Y2=0.4
r278 69 103 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0
r279 69 71 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=6.84 $Y=0.085
+ $X2=6.84 $Y2=0.4
r280 65 100 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0
r281 65 67 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=5.9 $Y=0.085
+ $X2=5.9 $Y2=0.4
r282 61 97 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0
r283 61 63 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.96 $Y=0.085
+ $X2=4.96 $Y2=0.4
r284 57 94 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0
r285 57 59 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=4.02 $Y=0.085
+ $X2=4.02 $Y2=0.4
r286 53 91 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0
r287 53 55 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=3.08 $Y=0.085
+ $X2=3.08 $Y2=0.4
r288 49 157 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0
r289 49 51 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.14 $Y=0.085
+ $X2=2.14 $Y2=0.4
r290 48 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=0 $X2=1.2
+ $Y2=0
r291 47 157 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.055 $Y=0 $X2=2.14
+ $Y2=0
r292 47 48 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=0
+ $X2=1.285 $Y2=0
r293 43 154 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0
r294 43 45 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.2 $Y=0.085
+ $X2=1.2 $Y2=0.4
r295 42 151 3.40825 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0
+ $X2=0.172 $Y2=0
r296 41 154 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=0 $X2=1.2
+ $Y2=0
r297 41 42 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=0
+ $X2=0.345 $Y2=0
r298 37 151 3.40825 $w=1.7e-07 $l=1.23386e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.172 $Y2=0
r299 37 39 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.4
r300 12 87 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=10.465
+ $Y=0.235 $X2=10.6 $Y2=0.4
r301 11 83 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=9.475
+ $Y=0.235 $X2=9.66 $Y2=0.4
r302 10 79 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=8.535
+ $Y=0.235 $X2=8.72 $Y2=0.4
r303 9 75 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=7.595
+ $Y=0.235 $X2=7.78 $Y2=0.4
r304 8 71 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=6.655
+ $Y=0.235 $X2=6.84 $Y2=0.4
r305 7 67 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=5.715
+ $Y=0.235 $X2=5.9 $Y2=0.4
r306 6 63 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=4.775
+ $Y=0.235 $X2=4.96 $Y2=0.4
r307 5 59 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=3.835
+ $Y=0.235 $X2=4.02 $Y2=0.4
r308 4 55 182 $w=1.7e-07 $l=2.22486e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.4
r309 3 51 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.955
+ $Y=0.235 $X2=2.14 $Y2=0.4
r310 2 45 182 $w=1.7e-07 $l=2.5446e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.2 $Y2=0.4
r311 1 39 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

