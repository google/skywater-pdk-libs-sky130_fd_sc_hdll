* File: sky130_fd_sc_hdll__o21a_2.pxi.spice
* Created: Thu Aug 27 19:18:59 2020
* 
x_PM_SKY130_FD_SC_HDLL__O21A_2%A_79_21# N_A_79_21#_M1002_s N_A_79_21#_M1000_d
+ N_A_79_21#_c_51_n N_A_79_21#_M1005_g N_A_79_21#_c_59_n N_A_79_21#_M1001_g
+ N_A_79_21#_c_52_n N_A_79_21#_M1009_g N_A_79_21#_c_60_n N_A_79_21#_M1006_g
+ N_A_79_21#_c_53_n N_A_79_21#_c_61_n N_A_79_21#_c_54_n N_A_79_21#_c_55_n
+ N_A_79_21#_c_67_p N_A_79_21#_c_83_p N_A_79_21#_c_56_n N_A_79_21#_c_75_p
+ N_A_79_21#_c_76_p N_A_79_21#_c_57_n N_A_79_21#_c_58_n
+ PM_SKY130_FD_SC_HDLL__O21A_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__O21A_2%B1 N_B1_c_124_n N_B1_M1000_g N_B1_c_125_n
+ N_B1_M1002_g B1 N_B1_c_126_n PM_SKY130_FD_SC_HDLL__O21A_2%B1
x_PM_SKY130_FD_SC_HDLL__O21A_2%A2 N_A2_c_153_n N_A2_M1004_g N_A2_c_154_n
+ N_A2_M1007_g N_A2_c_155_n A2 PM_SKY130_FD_SC_HDLL__O21A_2%A2
x_PM_SKY130_FD_SC_HDLL__O21A_2%A1 N_A1_c_189_n N_A1_M1003_g N_A1_c_192_n
+ N_A1_M1008_g A1 N_A1_c_191_n PM_SKY130_FD_SC_HDLL__O21A_2%A1
x_PM_SKY130_FD_SC_HDLL__O21A_2%VPWR N_VPWR_M1001_s N_VPWR_M1006_s N_VPWR_M1008_d
+ N_VPWR_c_219_n N_VPWR_c_220_n N_VPWR_c_221_n N_VPWR_c_222_n VPWR
+ N_VPWR_c_223_n N_VPWR_c_224_n N_VPWR_c_225_n N_VPWR_c_218_n
+ PM_SKY130_FD_SC_HDLL__O21A_2%VPWR
x_PM_SKY130_FD_SC_HDLL__O21A_2%X N_X_M1005_d N_X_M1001_d X N_X_c_264_n
+ PM_SKY130_FD_SC_HDLL__O21A_2%X
x_PM_SKY130_FD_SC_HDLL__O21A_2%VGND N_VGND_M1005_s N_VGND_M1009_s N_VGND_M1004_d
+ N_VGND_c_282_n N_VGND_c_283_n VGND N_VGND_c_284_n N_VGND_c_285_n
+ N_VGND_c_286_n N_VGND_c_287_n N_VGND_c_288_n N_VGND_c_289_n
+ PM_SKY130_FD_SC_HDLL__O21A_2%VGND
x_PM_SKY130_FD_SC_HDLL__O21A_2%A_414_47# N_A_414_47#_M1002_d N_A_414_47#_M1003_d
+ N_A_414_47#_c_333_n N_A_414_47#_c_347_n N_A_414_47#_c_332_n
+ PM_SKY130_FD_SC_HDLL__O21A_2%A_414_47#
cc_1 VNB N_A_79_21#_c_51_n 0.0220353f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_52_n 0.0195555f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.995
cc_3 VNB N_A_79_21#_c_53_n 0.00335532f $X=-0.19 $Y=-0.24 $X2=1.175 $Y2=1.15
cc_4 VNB N_A_79_21#_c_54_n 0.0110603f $X=-0.19 $Y=-0.24 $X2=1.565 $Y2=0.737
cc_5 VNB N_A_79_21#_c_55_n 3.01577e-19 $X=-0.19 $Y=-0.24 $X2=1.355 $Y2=0.737
cc_6 VNB N_A_79_21#_c_56_n 0.00488867f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.385
cc_7 VNB N_A_79_21#_c_57_n 9.92848e-19 $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.16
cc_8 VNB N_A_79_21#_c_58_n 0.0593356f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.202
cc_9 VNB N_B1_c_124_n 0.0342249f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=0.235
cc_10 VNB N_B1_c_125_n 0.0204042f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_B1_c_126_n 0.0028651f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_12 VNB N_A2_c_153_n 0.0182976f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=0.235
cc_13 VNB N_A2_c_154_n 0.0238236f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A2_c_155_n 0.00653127f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_15 VNB N_A1_c_189_n 0.0239352f $X=-0.19 $Y=-0.24 $X2=1.605 $Y2=0.235
cc_16 VNB A1 0.0137693f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_17 VNB N_A1_c_191_n 0.0396619f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_18 VNB N_VPWR_c_218_n 0.155873f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.202
cc_19 VNB N_X_c_264_n 6.35937e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_20 VNB N_VGND_c_282_n 0.0101667f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_21 VNB N_VGND_c_283_n 0.0379064f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_22 VNB N_VGND_c_284_n 0.0167192f $X=-0.19 $Y=-0.24 $X2=0.97 $Y2=1.41
cc_23 VNB N_VGND_c_285_n 0.0285809f $X=-0.19 $Y=-0.24 $X2=1.27 $Y2=1.33
cc_24 VNB N_VGND_c_286_n 0.0190528f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.385
cc_25 VNB N_VGND_c_287_n 0.204886f $X=-0.19 $Y=-0.24 $X2=1.73 $Y2=0.385
cc_26 VNB N_VGND_c_288_n 0.0117459f $X=-0.19 $Y=-0.24 $X2=1.08 $Y2=1.16
cc_27 VNB N_VGND_c_289_n 0.00964473f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=1.202
cc_28 VNB N_A_414_47#_c_332_n 0.0130293f $X=-0.19 $Y=-0.24 $X2=0.945 $Y2=0.56
cc_29 VPB N_A_79_21#_c_59_n 0.0208002f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_A_79_21#_c_60_n 0.0181297f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_31 VPB N_A_79_21#_c_61_n 0.00225704f $X=-0.19 $Y=1.305 $X2=1.27 $Y2=1.785
cc_32 VPB N_A_79_21#_c_57_n 0.00486079f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.16
cc_33 VPB N_A_79_21#_c_58_n 0.0306287f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.202
cc_34 VPB N_B1_c_124_n 0.0342434f $X=-0.19 $Y=1.305 $X2=1.605 $Y2=0.235
cc_35 VPB N_B1_c_126_n 0.00127301f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_36 VPB N_A2_c_154_n 0.0279872f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_A2_c_155_n 0.0106372f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_38 VPB A2 9.47552e-19 $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.995
cc_39 VPB N_A1_c_192_n 0.0211382f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB A1 0.00869997f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.995
cc_41 VPB N_A1_c_191_n 0.0166505f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_VPWR_c_219_n 0.00995082f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_43 VPB N_VPWR_c_220_n 0.0384221f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_44 VPB N_VPWR_c_221_n 0.0123393f $X=-0.19 $Y=1.305 $X2=0.945 $Y2=0.56
cc_45 VPB N_VPWR_c_222_n 0.037138f $X=-0.19 $Y=1.305 $X2=0.97 $Y2=1.41
cc_46 VPB N_VPWR_c_223_n 0.0374541f $X=-0.19 $Y=1.305 $X2=2.115 $Y2=1.895
cc_47 VPB N_VPWR_c_224_n 0.0166741f $X=-0.19 $Y=1.305 $X2=2.245 $Y2=1.895
cc_48 VPB N_VPWR_c_225_n 0.0176591f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_49 VPB N_VPWR_c_218_n 0.0453595f $X=-0.19 $Y=1.305 $X2=1.08 $Y2=1.202
cc_50 VPB N_X_c_264_n 0.00112635f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 N_A_79_21#_c_53_n N_B1_c_124_n 0.00131615f $X=1.175 $Y=1.15 $X2=-0.19
+ $Y2=-0.24
cc_52 N_A_79_21#_c_61_n N_B1_c_124_n 0.0047735f $X=1.27 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_53 N_A_79_21#_c_54_n N_B1_c_124_n 0.0063366f $X=1.565 $Y=0.737 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A_79_21#_c_67_p N_B1_c_124_n 0.019857f $X=2.115 $Y=1.895 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A_79_21#_c_57_n N_B1_c_124_n 2.89858e-19 $X=1.08 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_56 N_A_79_21#_c_58_n N_B1_c_124_n 0.00890385f $X=0.97 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_57 N_A_79_21#_c_53_n N_B1_c_125_n 0.00332331f $X=1.175 $Y=1.15 $X2=0 $Y2=0
cc_58 N_A_79_21#_c_53_n N_B1_c_126_n 0.0499795f $X=1.175 $Y=1.15 $X2=0 $Y2=0
cc_59 N_A_79_21#_c_54_n N_B1_c_126_n 0.0304611f $X=1.565 $Y=0.737 $X2=0 $Y2=0
cc_60 N_A_79_21#_c_67_p N_B1_c_126_n 0.0300452f $X=2.115 $Y=1.895 $X2=0 $Y2=0
cc_61 N_A_79_21#_c_58_n N_B1_c_126_n 9.30587e-19 $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_62 N_A_79_21#_c_75_p N_A2_c_154_n 0.00404646f $X=2.245 $Y=2.005 $X2=0 $Y2=0
cc_63 N_A_79_21#_c_76_p N_A2_c_154_n 0.00971236f $X=2.21 $Y=2.3 $X2=0 $Y2=0
cc_64 N_A_79_21#_c_75_p N_A2_c_155_n 0.00152662f $X=2.245 $Y=2.005 $X2=0 $Y2=0
cc_65 N_A_79_21#_c_75_p A2 0.00798412f $X=2.245 $Y=2.005 $X2=0 $Y2=0
cc_66 N_A_79_21#_c_75_p N_A1_c_192_n 2.35169e-19 $X=2.245 $Y=2.005 $X2=0 $Y2=0
cc_67 N_A_79_21#_c_76_p N_A1_c_192_n 0.00193653f $X=2.21 $Y=2.3 $X2=0 $Y2=0
cc_68 N_A_79_21#_c_61_n N_VPWR_M1006_s 0.00983811f $X=1.27 $Y=1.785 $X2=0 $Y2=0
cc_69 N_A_79_21#_c_67_p N_VPWR_M1006_s 0.0187668f $X=2.115 $Y=1.895 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_83_p N_VPWR_M1006_s 0.00651216f $X=1.355 $Y=1.895 $X2=0 $Y2=0
cc_71 N_A_79_21#_c_59_n N_VPWR_c_220_n 0.00872587f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_67_p N_VPWR_c_223_n 0.00271905f $X=2.115 $Y=1.895 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_76_p N_VPWR_c_223_n 0.0160594f $X=2.21 $Y=2.3 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_59_n N_VPWR_c_224_n 0.00620483f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_60_n N_VPWR_c_224_n 0.00447018f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_59_n N_VPWR_c_225_n 5.20907e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_60_n N_VPWR_c_225_n 0.0142428f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_67_p N_VPWR_c_225_n 0.0361623f $X=2.115 $Y=1.895 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_83_p N_VPWR_c_225_n 0.0137948f $X=1.355 $Y=1.895 $X2=0 $Y2=0
cc_80 N_A_79_21#_M1000_d N_VPWR_c_218_n 0.00264529f $X=2.06 $Y=1.485 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_59_n N_VPWR_c_218_n 0.0114735f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_60_n N_VPWR_c_218_n 0.00760114f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_67_p N_VPWR_c_218_n 0.00722617f $X=2.115 $Y=1.895 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_83_p N_VPWR_c_218_n 7.64972e-19 $X=1.355 $Y=1.895 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_76_p N_VPWR_c_218_n 0.00979433f $X=2.21 $Y=2.3 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_51_n N_X_c_264_n 0.0154423f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_59_n N_X_c_264_n 0.0251587f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_52_n N_X_c_264_n 0.00220545f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_60_n N_X_c_264_n 0.00184943f $X=0.97 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_53_n N_X_c_264_n 0.0353331f $X=1.175 $Y=1.15 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_61_n N_X_c_264_n 0.0134026f $X=1.27 $Y=1.785 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_58_n N_X_c_264_n 0.0425185f $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_55_n N_VGND_M1009_s 0.00409231f $X=1.355 $Y=0.737 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_51_n N_VGND_c_283_n 0.00318444f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_51_n N_VGND_c_284_n 0.00564131f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_52_n N_VGND_c_284_n 0.00487821f $X=0.945 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_54_n N_VGND_c_285_n 0.00351026f $X=1.565 $Y=0.737 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_56_n N_VGND_c_285_n 0.0218088f $X=1.73 $Y=0.385 $X2=0 $Y2=0
cc_99 N_A_79_21#_M1002_s N_VGND_c_287_n 0.00341197f $X=1.605 $Y=0.235 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_51_n N_VGND_c_287_n 0.0111495f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_52_n N_VGND_c_287_n 0.00833798f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_54_n N_VGND_c_287_n 0.00554211f $X=1.565 $Y=0.737 $X2=0
+ $Y2=0
cc_103 N_A_79_21#_c_55_n N_VGND_c_287_n 0.0018018f $X=1.355 $Y=0.737 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_56_n N_VGND_c_287_n 0.0125824f $X=1.73 $Y=0.385 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_51_n N_VGND_c_288_n 4.68063e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_52_n N_VGND_c_288_n 0.00789681f $X=0.945 $Y=0.995 $X2=0
+ $Y2=0
cc_107 N_A_79_21#_c_54_n N_VGND_c_288_n 0.00148828f $X=1.565 $Y=0.737 $X2=0
+ $Y2=0
cc_108 N_A_79_21#_c_55_n N_VGND_c_288_n 0.0253682f $X=1.355 $Y=0.737 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_56_n N_VGND_c_288_n 0.016345f $X=1.73 $Y=0.385 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_58_n N_VGND_c_288_n 6.23957e-19 $X=0.97 $Y=1.202 $X2=0 $Y2=0
cc_111 N_B1_c_125_n N_A2_c_153_n 0.0209519f $X=1.995 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_112 N_B1_c_124_n N_A2_c_154_n 0.0413184f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B1_c_126_n N_A2_c_154_n 0.00156815f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_124_n N_A2_c_155_n 0.00326852f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B1_c_126_n N_A2_c_155_n 0.0181252f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_116 N_B1_c_126_n N_VPWR_M1006_s 0.00554778f $X=1.79 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B1_c_124_n N_VPWR_c_223_n 0.00479351f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_118 N_B1_c_124_n N_VPWR_c_225_n 0.00996638f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B1_c_124_n N_VPWR_c_218_n 0.0055283f $X=1.97 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_125_n N_VGND_c_285_n 0.00585385f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_121 N_B1_c_125_n N_VGND_c_287_n 0.0121155f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_122 N_B1_c_125_n N_VGND_c_288_n 0.00247598f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_123 N_B1_c_125_n N_VGND_c_289_n 0.00171866f $X=1.995 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A2_c_153_n N_A1_c_189_n 0.0191445f $X=2.425 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_125 N_A2_c_154_n N_A1_c_192_n 0.0266259f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_126 A2 N_A1_c_192_n 0.0219411f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_127 N_A2_c_154_n A1 2.91106e-19 $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A2_c_155_n A1 0.0261206f $X=2.8 $Y=1.212 $X2=0 $Y2=0
cc_129 A2 A1 0.00332746f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_130 N_A2_c_154_n N_A1_c_191_n 0.0123782f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A2_c_155_n N_A1_c_191_n 0.0134124f $X=2.8 $Y=1.212 $X2=0 $Y2=0
cc_132 A2 N_A1_c_191_n 4.75184e-19 $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_133 N_A2_c_154_n N_VPWR_c_223_n 0.00681208f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_134 A2 N_VPWR_c_223_n 0.00379002f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_135 N_A2_c_154_n N_VPWR_c_225_n 0.00103117f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_136 N_A2_c_154_n N_VPWR_c_218_n 0.0127129f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_137 A2 N_VPWR_c_218_n 0.00745471f $X=2.9 $Y=1.785 $X2=0 $Y2=0
cc_138 A2 A_508_297# 0.0117719f $X=2.9 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_139 N_A2_c_153_n N_VGND_c_285_n 0.00410924f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A2_c_153_n N_VGND_c_287_n 0.00475403f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_141 N_A2_c_153_n N_VGND_c_289_n 0.0131295f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_142 N_A2_c_153_n N_A_414_47#_c_333_n 0.0115145f $X=2.425 $Y=0.995 $X2=0 $Y2=0
cc_143 N_A2_c_154_n N_A_414_47#_c_333_n 0.00367389f $X=2.45 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A2_c_155_n N_A_414_47#_c_333_n 0.0473731f $X=2.8 $Y=1.212 $X2=0 $Y2=0
cc_145 N_A1_c_192_n N_VPWR_c_222_n 0.00705937f $X=3.13 $Y=1.41 $X2=0 $Y2=0
cc_146 A1 N_VPWR_c_222_n 0.0200607f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_147 N_A1_c_191_n N_VPWR_c_222_n 0.00142072f $X=3.13 $Y=1.202 $X2=0 $Y2=0
cc_148 N_A1_c_192_n N_VPWR_c_223_n 0.00669297f $X=3.13 $Y=1.41 $X2=0 $Y2=0
cc_149 N_A1_c_192_n N_VPWR_c_218_n 0.0128547f $X=3.13 $Y=1.41 $X2=0 $Y2=0
cc_150 N_A1_c_189_n N_VGND_c_286_n 0.00410924f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A1_c_189_n N_VGND_c_287_n 0.00578113f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_152 N_A1_c_189_n N_VGND_c_289_n 0.0191915f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_153 N_A1_c_189_n N_A_414_47#_c_333_n 0.0146153f $X=3.105 $Y=0.995 $X2=0 $Y2=0
cc_154 N_A1_c_191_n N_A_414_47#_c_333_n 0.00200568f $X=3.13 $Y=1.202 $X2=0 $Y2=0
cc_155 A1 N_A_414_47#_c_332_n 0.0204086f $X=3.31 $Y=1.105 $X2=0 $Y2=0
cc_156 N_A1_c_191_n N_A_414_47#_c_332_n 0.00262059f $X=3.13 $Y=1.202 $X2=0 $Y2=0
cc_157 N_VPWR_c_218_n N_X_M1001_d 0.00426212f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_158 N_VPWR_c_220_n N_X_c_264_n 0.0586842f $X=0.26 $Y=1.815 $X2=0 $Y2=0
cc_159 N_VPWR_c_224_n N_X_c_264_n 0.018435f $X=0.995 $Y=2.495 $X2=0 $Y2=0
cc_160 N_VPWR_c_218_n N_X_c_264_n 0.0109593f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_161 N_VPWR_c_218_n A_508_297# 0.0143195f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_162 N_X_c_264_n N_VGND_c_284_n 0.0181722f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_163 N_X_M1005_d N_VGND_c_287_n 0.00415586f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_164 N_X_c_264_n N_VGND_c_287_n 0.0111475f $X=0.73 $Y=0.42 $X2=0 $Y2=0
cc_165 N_VGND_c_287_n N_A_414_47#_M1002_d 0.00421987f $X=3.45 $Y=0 $X2=-0.19
+ $Y2=-0.24
cc_166 N_VGND_c_287_n N_A_414_47#_M1003_d 0.00323627f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_167 N_VGND_M1004_d N_A_414_47#_c_333_n 0.0105422f $X=2.5 $Y=0.235 $X2=0 $Y2=0
cc_168 N_VGND_c_285_n N_A_414_47#_c_333_n 0.00262712f $X=2.495 $Y=0 $X2=0 $Y2=0
cc_169 N_VGND_c_286_n N_A_414_47#_c_333_n 0.00325763f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_170 N_VGND_c_287_n N_A_414_47#_c_333_n 0.0121028f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_171 N_VGND_c_289_n N_A_414_47#_c_333_n 0.0325446f $X=2.53 $Y=0 $X2=0 $Y2=0
cc_172 N_VGND_c_285_n N_A_414_47#_c_347_n 0.00533689f $X=2.495 $Y=0 $X2=0 $Y2=0
cc_173 N_VGND_c_287_n N_A_414_47#_c_347_n 0.00689411f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_174 N_VGND_c_286_n N_A_414_47#_c_332_n 0.007063f $X=3.45 $Y=0 $X2=0 $Y2=0
cc_175 N_VGND_c_287_n N_A_414_47#_c_332_n 0.0088263f $X=3.45 $Y=0 $X2=0 $Y2=0
