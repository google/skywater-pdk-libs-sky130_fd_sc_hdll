* File: sky130_fd_sc_hdll__o22ai_4.spice
* Created: Wed Sep  2 08:45:51 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22ai_4.pex.spice"
.subckt sky130_fd_sc_hdll__o22ai_4  VNB VPB A1 A2 B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2	A2
* A1	A1
* VPB	VPB
* VNB	VNB
MM1005 N_A_33_47#_M1005_d N_A1_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75007.3 A=0.0975 P=1.6 MULT=1
MM1006 N_A_33_47#_M1006_d N_A1_M1006_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75006.8 A=0.0975 P=1.6 MULT=1
MM1019 N_A_33_47#_M1006_d N_A1_M1019_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.2
+ SB=75006.3 A=0.0975 P=1.6 MULT=1
MM1002 N_A_33_47#_M1002_d N_A2_M1002_g N_VGND_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1016 N_A_33_47#_M1002_d N_A2_M1016_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75005.5 A=0.0975 P=1.6 MULT=1
MM1024 N_A_33_47#_M1024_d N_A2_M1024_g N_VGND_M1016_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.5
+ SB=75005 A=0.0975 P=1.6 MULT=1
MM1026 N_A_33_47#_M1024_d N_A2_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75003.1
+ SB=75004.5 A=0.0975 P=1.6 MULT=1
MM1031 N_A_33_47#_M1031_d N_A1_M1031_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75003.5
+ SB=75004 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_B1_M1004_g N_A_33_47#_M1031_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=8.304 M=1 R=4.33333 SA=75004
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1014 N_Y_M1004_d N_B1_M1014_g N_A_33_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75004.5
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1020_d N_B1_M1020_g N_A_33_47#_M1014_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1009 N_A_33_47#_M1009_d N_B2_M1009_g N_Y_M1020_d VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.08775 PD=0.97 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75005.4
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1010 N_A_33_47#_M1009_d N_B2_M1010_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75005.9
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1017 N_A_33_47#_M1017_d N_B2_M1017_g N_Y_M1010_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.3
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1021 N_A_33_47#_M1017_d N_B2_M1021_g N_Y_M1021_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.104 PD=1.02 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75006.9
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1029 N_Y_M1021_s N_B1_M1029_g N_A_33_47#_M1029_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.169 PD=0.97 PS=1.82 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75007.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_123_297#_M1007_d N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.3 PD=1.29 PS=2.6 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90007.3 A=0.18 P=2.36 MULT=1
MM1011 N_A_123_297#_M1007_d N_A1_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90006.8 A=0.18 P=2.36 MULT=1
MM1012 N_A_123_297#_M1012_d N_A1_M1012_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90006.3 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_A2_M1000_g N_A_123_297#_M1012_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90005.9 A=0.18 P=2.36 MULT=1
MM1015 N_Y_M1000_d N_A2_M1015_g N_A_123_297#_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90005.4 A=0.18 P=2.36 MULT=1
MM1022 N_Y_M1022_d N_A2_M1022_g N_A_123_297#_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1025 N_Y_M1022_d N_A2_M1025_g N_A_123_297#_M1025_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90004.5 A=0.18 P=2.36 MULT=1
MM1027 N_A_123_297#_M1025_s N_A1_M1027_g N_VPWR_M1027_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.17 PD=1.29 PS=1.34 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90003.5 SB=90004 A=0.18 P=2.36 MULT=1
MM1003 N_A_885_297#_M1003_d N_B1_M1003_g N_VPWR_M1027_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.17 PD=1.29 PS=1.34 NRD=0.9653 NRS=2.9353 M=1 R=5.55556 SA=90004
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1018 N_A_885_297#_M1003_d N_B1_M1018_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.5 SB=90003 A=0.18 P=2.36 MULT=1
MM1023 N_A_885_297#_M1023_d N_B1_M1023_g N_VPWR_M1018_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1001 N_Y_M1001_d N_B2_M1001_g N_A_885_297#_M1023_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.4 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1008 N_Y_M1001_d N_B2_M1008_g N_A_885_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.9 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1013 N_Y_M1013_d N_B2_M1013_g N_A_885_297#_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.4 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1028 N_Y_M1013_d N_B2_M1028_g N_A_885_297#_M1028_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90006.8 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1030 N_A_885_297#_M1028_s N_B1_M1030_g N_VPWR_M1030_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90007.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX32_noxref VNB VPB NWDIODE A=13.8993 P=20.53
pX33_noxref noxref_13 A1 A1 PROBETYPE=1
pX34_noxref noxref_14 A2 A2 PROBETYPE=1
pX35_noxref noxref_15 B1 B1 PROBETYPE=1
pX36_noxref noxref_16 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o22ai_4.pxi.spice"
*
.ends
*
*
