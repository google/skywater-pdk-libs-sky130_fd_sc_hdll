* File: sky130_fd_sc_hdll__a32o_2.pxi.spice
* Created: Wed Sep  2 08:20:41 2020
* 
x_PM_SKY130_FD_SC_HDLL__A32O_2%A_21_199# N_A_21_199#_M1004_d N_A_21_199#_M1008_d
+ N_A_21_199#_c_69_n N_A_21_199#_M1000_g N_A_21_199#_c_64_n N_A_21_199#_M1001_g
+ N_A_21_199#_c_70_n N_A_21_199#_M1003_g N_A_21_199#_c_65_n N_A_21_199#_M1009_g
+ N_A_21_199#_c_66_n N_A_21_199#_c_72_n N_A_21_199#_c_118_p N_A_21_199#_c_67_n
+ N_A_21_199#_c_74_n N_A_21_199#_c_82_p N_A_21_199#_c_83_p N_A_21_199#_c_78_p
+ N_A_21_199#_c_79_p N_A_21_199#_c_84_p N_A_21_199#_c_68_n
+ PM_SKY130_FD_SC_HDLL__A32O_2%A_21_199#
x_PM_SKY130_FD_SC_HDLL__A32O_2%B2 N_B2_c_161_n N_B2_M1012_g N_B2_c_162_n
+ N_B2_M1008_g N_B2_c_163_n B2 B2 PM_SKY130_FD_SC_HDLL__A32O_2%B2
x_PM_SKY130_FD_SC_HDLL__A32O_2%B1 N_B1_c_198_n N_B1_M1004_g N_B1_c_199_n
+ N_B1_M1005_g N_B1_c_200_n B1 PM_SKY130_FD_SC_HDLL__A32O_2%B1
x_PM_SKY130_FD_SC_HDLL__A32O_2%A1 N_A1_c_238_n N_A1_M1007_g N_A1_c_239_n
+ N_A1_M1002_g A1 PM_SKY130_FD_SC_HDLL__A32O_2%A1
x_PM_SKY130_FD_SC_HDLL__A32O_2%A2 N_A2_c_272_n N_A2_M1011_g N_A2_c_273_n
+ N_A2_M1010_g A2 A2 A2 A2 PM_SKY130_FD_SC_HDLL__A32O_2%A2
x_PM_SKY130_FD_SC_HDLL__A32O_2%A3 N_A3_c_307_n N_A3_M1013_g N_A3_c_310_n
+ N_A3_M1006_g A3 A3 N_A3_c_309_n PM_SKY130_FD_SC_HDLL__A32O_2%A3
x_PM_SKY130_FD_SC_HDLL__A32O_2%X N_X_M1001_s N_X_M1000_d N_X_M1003_d N_X_c_337_n
+ N_X_c_341_n N_X_c_346_n X X X X X N_X_c_332_n X PM_SKY130_FD_SC_HDLL__A32O_2%X
x_PM_SKY130_FD_SC_HDLL__A32O_2%VPWR N_VPWR_M1000_s N_VPWR_M1002_d N_VPWR_M1006_d
+ N_VPWR_c_375_n N_VPWR_c_376_n N_VPWR_c_377_n N_VPWR_c_378_n VPWR
+ N_VPWR_c_379_n N_VPWR_c_380_n N_VPWR_c_381_n N_VPWR_c_382_n N_VPWR_c_383_n
+ N_VPWR_c_374_n PM_SKY130_FD_SC_HDLL__A32O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A32O_2%A_319_297# N_A_319_297#_M1008_s
+ N_A_319_297#_M1005_d N_A_319_297#_M1011_d N_A_319_297#_c_443_n
+ N_A_319_297#_c_445_n N_A_319_297#_c_460_n N_A_319_297#_c_447_n
+ N_A_319_297#_c_449_n N_A_319_297#_c_454_n N_A_319_297#_c_458_n
+ PM_SKY130_FD_SC_HDLL__A32O_2%A_319_297#
x_PM_SKY130_FD_SC_HDLL__A32O_2%VGND N_VGND_M1001_d N_VGND_M1009_d N_VGND_M1013_d
+ N_VGND_c_479_n N_VGND_c_480_n N_VGND_c_481_n N_VGND_c_482_n VGND
+ N_VGND_c_483_n N_VGND_c_484_n N_VGND_c_485_n N_VGND_c_486_n
+ PM_SKY130_FD_SC_HDLL__A32O_2%VGND
cc_1 VNB N_A_21_199#_c_64_n 0.0196754f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB N_A_21_199#_c_65_n 0.0187056f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_A_21_199#_c_66_n 6.46921e-19 $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.16
cc_4 VNB N_A_21_199#_c_67_n 0.00114743f $X=-0.19 $Y=-0.24 $X2=1.92 $Y2=1.445
cc_5 VNB N_A_21_199#_c_68_n 0.0677561f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_6 VNB N_B2_c_161_n 0.0192854f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.235
cc_7 VNB N_B2_c_162_n 0.0190177f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_B2_c_163_n 0.0312788f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_9 VNB B2 0.00746941f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_10 VNB N_B1_c_198_n 0.0181522f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.235
cc_11 VNB N_B1_c_199_n 0.0225267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_B1_c_200_n 0.0038461f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_13 VNB B1 6.1667e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_14 VNB N_A1_c_238_n 0.0187296f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.235
cc_15 VNB N_A1_c_239_n 0.0283838f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB A1 7.25193e-19 $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_17 VNB N_A2_c_272_n 0.0245135f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.235
cc_18 VNB N_A2_c_273_n 0.017115f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB A2 0.00381859f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_20 VNB N_A3_c_307_n 0.0213114f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=0.235
cc_21 VNB A3 0.0181035f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_22 VNB N_A3_c_309_n 0.0394908f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_23 VNB N_X_c_332_n 0.00692367f $X=-0.19 $Y=-0.24 $X2=2.04 $Y2=0.76
cc_24 VNB X 0.00492f $X=-0.19 $Y=-0.24 $X2=2.62 $Y2=0.51
cc_25 VNB N_VPWR_c_374_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0.62 $Y2=1.202
cc_26 VNB N_VGND_c_479_n 0.0114823f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_27 VNB N_VGND_c_480_n 0.0148471f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_28 VNB N_VGND_c_481_n 0.0147433f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_29 VNB N_VGND_c_482_n 0.0259025f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_30 VNB N_VGND_c_483_n 0.0621069f $X=-0.19 $Y=-0.24 $X2=0.755 $Y2=1.53
cc_31 VNB N_VGND_c_484_n 0.0147015f $X=-0.19 $Y=-0.24 $X2=2.15 $Y2=1.53
cc_32 VNB N_VGND_c_485_n 0.0177781f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_33 VNB N_VGND_c_486_n 0.241603f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_34 VPB N_A_21_199#_c_69_n 0.018351f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_35 VPB N_A_21_199#_c_70_n 0.0199096f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_36 VPB N_A_21_199#_c_66_n 0.00114011f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.16
cc_37 VPB N_A_21_199#_c_72_n 0.0179612f $X=-0.19 $Y=1.305 $X2=1.8 $Y2=1.53
cc_38 VPB N_A_21_199#_c_67_n 0.00448371f $X=-0.19 $Y=1.305 $X2=1.92 $Y2=1.445
cc_39 VPB N_A_21_199#_c_74_n 0.00339638f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.615
cc_40 VPB N_A_21_199#_c_68_n 0.0329382f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_41 VPB N_B2_c_162_n 0.0294298f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_B2_c_163_n 0.011407f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_43 VPB N_B1_c_199_n 0.0262074f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_44 VPB B1 0.00166918f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_45 VPB N_A1_c_239_n 0.0292201f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB A1 0.00215509f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_47 VPB N_A2_c_272_n 0.0265272f $X=-0.19 $Y=1.305 $X2=2.415 $Y2=0.235
cc_48 VPB A2 0.00336577f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_49 VPB N_A3_c_310_n 0.0181963f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A3 0.0189911f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_51 VPB N_A3_c_309_n 0.0166497f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_52 VPB X 0.00692367f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB X 0.00659625f $X=-0.19 $Y=1.305 $X2=2.62 $Y2=0.51
cc_54 VPB N_VPWR_c_375_n 4.89699e-19 $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.56
cc_55 VPB N_VPWR_c_376_n 0.00287591f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_56 VPB N_VPWR_c_377_n 0.0144807f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.56
cc_57 VPB N_VPWR_c_378_n 0.0257878f $X=-0.19 $Y=1.305 $X2=0.645 $Y2=1.16
cc_58 VPB N_VPWR_c_379_n 0.015528f $X=-0.19 $Y=1.305 $X2=1.8 $Y2=1.53
cc_59 VPB N_VPWR_c_380_n 0.0492252f $X=-0.19 $Y=1.305 $X2=2.15 $Y2=1.945
cc_60 VPB N_VPWR_c_381_n 0.0188829f $X=-0.19 $Y=1.305 $X2=2.555 $Y2=0.675
cc_61 VPB N_VPWR_c_382_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_VPWR_c_383_n 0.00580298f $X=-0.19 $Y=1.305 $X2=2.19 $Y2=1.945
cc_63 VPB N_VPWR_c_374_n 0.0608534f $X=-0.19 $Y=1.305 $X2=0.62 $Y2=1.202
cc_64 N_A_21_199#_c_65_n N_B2_c_161_n 0.00782949f $X=0.99 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_65 N_A_21_199#_c_67_n N_B2_c_161_n 0.00367864f $X=1.92 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_66 N_A_21_199#_c_78_p N_B2_c_161_n 0.0104442f $X=2.04 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_67 N_A_21_199#_c_79_p N_B2_c_161_n 0.00151464f $X=2.62 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_68 N_A_21_199#_c_67_n N_B2_c_162_n 0.0253675f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_69 N_A_21_199#_c_74_n N_B2_c_162_n 0.0228882f $X=2.15 $Y=1.615 $X2=0 $Y2=0
cc_70 N_A_21_199#_c_82_p N_B2_c_162_n 0.00926687f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_71 N_A_21_199#_c_83_p N_B2_c_162_n 4.36275e-19 $X=2.405 $Y=0.76 $X2=0 $Y2=0
cc_72 N_A_21_199#_c_84_p N_B2_c_162_n 0.00235935f $X=2.19 $Y=2.03 $X2=0 $Y2=0
cc_73 N_A_21_199#_c_66_n N_B2_c_163_n 3.79417e-19 $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_21_199#_c_72_n N_B2_c_163_n 0.00702957f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_75 N_A_21_199#_c_68_n N_B2_c_163_n 0.0167085f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_76 N_A_21_199#_c_65_n B2 0.00920453f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_77 N_A_21_199#_c_66_n B2 0.0144183f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_78 N_A_21_199#_c_72_n B2 0.0452692f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_79 N_A_21_199#_c_67_n B2 0.0334038f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_80 N_A_21_199#_c_78_p B2 0.00857643f $X=2.04 $Y=0.76 $X2=0 $Y2=0
cc_81 N_A_21_199#_c_67_n N_B1_c_198_n 0.00318895f $X=1.92 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_21_199#_c_83_p N_B1_c_198_n 0.0125489f $X=2.405 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_83 N_A_21_199#_c_79_p N_B1_c_198_n 0.0117833f $X=2.62 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_84 N_A_21_199#_c_67_n N_B1_c_199_n 0.00150261f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_85 N_A_21_199#_c_74_n N_B1_c_199_n 0.00109995f $X=2.15 $Y=1.615 $X2=0 $Y2=0
cc_86 N_A_21_199#_c_82_p N_B1_c_199_n 0.00463218f $X=2.19 $Y=1.63 $X2=0 $Y2=0
cc_87 N_A_21_199#_c_83_p N_B1_c_199_n 0.00437651f $X=2.405 $Y=0.76 $X2=0 $Y2=0
cc_88 N_A_21_199#_c_84_p N_B1_c_199_n 0.00381353f $X=2.19 $Y=2.03 $X2=0 $Y2=0
cc_89 N_A_21_199#_c_67_n N_B1_c_200_n 0.0120484f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_90 N_A_21_199#_c_74_n N_B1_c_200_n 0.00264867f $X=2.15 $Y=1.615 $X2=0 $Y2=0
cc_91 N_A_21_199#_c_83_p N_B1_c_200_n 0.0229481f $X=2.405 $Y=0.76 $X2=0 $Y2=0
cc_92 N_A_21_199#_c_67_n B1 0.007028f $X=1.92 $Y=1.445 $X2=0 $Y2=0
cc_93 N_A_21_199#_c_74_n B1 0.01358f $X=2.15 $Y=1.615 $X2=0 $Y2=0
cc_94 N_A_21_199#_c_83_p N_A1_c_238_n 0.00132568f $X=2.405 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_95 N_A_21_199#_c_79_p N_A1_c_238_n 0.00345111f $X=2.62 $Y=0.51 $X2=-0.19
+ $Y2=-0.24
cc_96 N_A_21_199#_c_83_p A1 0.0138445f $X=2.405 $Y=0.76 $X2=0 $Y2=0
cc_97 N_A_21_199#_c_79_p A1 0.0197003f $X=2.62 $Y=0.51 $X2=0 $Y2=0
cc_98 N_A_21_199#_c_72_n N_X_M1003_d 0.00397597f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_99 N_A_21_199#_c_64_n N_X_c_337_n 0.0140761f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_100 N_A_21_199#_c_66_n N_X_c_337_n 0.0147504f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A_21_199#_c_72_n N_X_c_337_n 0.00343508f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_102 N_A_21_199#_c_68_n N_X_c_337_n 0.00532881f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_103 N_A_21_199#_c_69_n N_X_c_341_n 0.0145782f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_A_21_199#_c_70_n N_X_c_341_n 0.0111137f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_105 N_A_21_199#_c_72_n N_X_c_341_n 0.0168151f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_106 N_A_21_199#_c_118_p N_X_c_341_n 0.0128629f $X=0.755 $Y=1.53 $X2=0 $Y2=0
cc_107 N_A_21_199#_c_68_n N_X_c_341_n 6.24009e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_108 N_A_21_199#_c_72_n N_X_c_346_n 0.013831f $X=1.8 $Y=1.53 $X2=0 $Y2=0
cc_109 N_A_21_199#_c_69_n X 0.0109525f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_21_199#_c_64_n X 0.0064012f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_21_199#_c_66_n X 0.029329f $X=0.62 $Y=1.16 $X2=0 $Y2=0
cc_112 N_A_21_199#_c_118_p X 0.0124935f $X=0.755 $Y=1.53 $X2=0 $Y2=0
cc_113 N_A_21_199#_c_68_n X 0.0352168f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_114 N_A_21_199#_c_72_n N_VPWR_M1000_s 6.60679e-19 $X=1.8 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_115 N_A_21_199#_c_118_p N_VPWR_M1000_s 0.00123897f $X=0.755 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_116 N_A_21_199#_c_69_n N_VPWR_c_375_n 0.0139134f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_21_199#_c_70_n N_VPWR_c_375_n 0.0109769f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_21_199#_c_69_n N_VPWR_c_379_n 0.00427505f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_21_199#_c_70_n N_VPWR_c_380_n 0.00622633f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_21_199#_M1008_d N_VPWR_c_374_n 0.00232895f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_121 N_A_21_199#_c_69_n N_VPWR_c_374_n 0.00485802f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_122 N_A_21_199#_c_70_n N_VPWR_c_374_n 0.0067625f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_21_199#_c_72_n N_A_319_297#_M1008_s 0.00382182f $X=1.8 $Y=1.53
+ $X2=-0.19 $Y2=-0.24
cc_124 N_A_21_199#_c_72_n N_A_319_297#_c_443_n 0.0136318f $X=1.8 $Y=1.53 $X2=0
+ $Y2=0
cc_125 N_A_21_199#_c_82_p N_A_319_297#_c_443_n 0.0197461f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_126 N_A_21_199#_M1008_d N_A_319_297#_c_445_n 0.00350851f $X=2.045 $Y=1.485
+ $X2=0 $Y2=0
cc_127 N_A_21_199#_c_84_p N_A_319_297#_c_445_n 0.0148109f $X=2.19 $Y=2.03 $X2=0
+ $Y2=0
cc_128 N_A_21_199#_c_82_p N_A_319_297#_c_447_n 0.00820492f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_129 N_A_21_199#_c_84_p N_A_319_297#_c_447_n 0.00135384f $X=2.19 $Y=2.03 $X2=0
+ $Y2=0
cc_130 N_A_21_199#_c_84_p N_A_319_297#_c_449_n 0.00905129f $X=2.19 $Y=2.03 $X2=0
+ $Y2=0
cc_131 N_A_21_199#_c_64_n N_VGND_c_480_n 0.00330856f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_132 N_A_21_199#_c_68_n N_VGND_c_480_n 0.00177805f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_133 N_A_21_199#_c_83_p N_VGND_c_483_n 0.00527747f $X=2.405 $Y=0.76 $X2=0
+ $Y2=0
cc_134 N_A_21_199#_c_78_p N_VGND_c_483_n 0.0036069f $X=2.04 $Y=0.76 $X2=0 $Y2=0
cc_135 N_A_21_199#_c_79_p N_VGND_c_483_n 0.0148919f $X=2.62 $Y=0.51 $X2=0 $Y2=0
cc_136 N_A_21_199#_c_64_n N_VGND_c_484_n 0.00428022f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_137 N_A_21_199#_c_65_n N_VGND_c_484_n 0.00271402f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_138 N_A_21_199#_c_64_n N_VGND_c_485_n 0.00119847f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_139 N_A_21_199#_c_65_n N_VGND_c_485_n 0.0148934f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_140 N_A_21_199#_M1004_d N_VGND_c_486_n 0.00623554f $X=2.415 $Y=0.235 $X2=0
+ $Y2=0
cc_141 N_A_21_199#_c_64_n N_VGND_c_486_n 0.00681489f $X=0.52 $Y=0.995 $X2=0
+ $Y2=0
cc_142 N_A_21_199#_c_65_n N_VGND_c_486_n 0.00505489f $X=0.99 $Y=0.995 $X2=0
+ $Y2=0
cc_143 N_A_21_199#_c_83_p N_VGND_c_486_n 0.00931653f $X=2.405 $Y=0.76 $X2=0
+ $Y2=0
cc_144 N_A_21_199#_c_78_p N_VGND_c_486_n 0.00644623f $X=2.04 $Y=0.76 $X2=0 $Y2=0
cc_145 N_A_21_199#_c_79_p N_VGND_c_486_n 0.0111373f $X=2.62 $Y=0.51 $X2=0 $Y2=0
cc_146 N_A_21_199#_c_67_n A_382_47# 4.90902e-19 $X=1.92 $Y=1.445 $X2=-0.19
+ $Y2=-0.24
cc_147 N_A_21_199#_c_83_p A_382_47# 0.00609277f $X=2.405 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_148 N_A_21_199#_c_78_p A_382_47# 0.00139636f $X=2.04 $Y=0.76 $X2=-0.19
+ $Y2=-0.24
cc_149 N_B2_c_161_n N_B1_c_198_n 0.0301168f $X=1.835 $Y=0.995 $X2=-0.19
+ $Y2=-0.24
cc_150 N_B2_c_162_n N_B1_c_199_n 0.0469587f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_151 N_B2_c_162_n N_B1_c_200_n 0.0011151f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_152 N_B2_c_162_n B1 6.70716e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_153 N_B2_c_162_n N_VPWR_c_380_n 0.00429453f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_154 N_B2_c_162_n N_VPWR_c_374_n 0.00737353f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_155 N_B2_c_162_n N_A_319_297#_c_445_n 0.0137415f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_156 B2 N_VGND_M1009_d 0.0102623f $X=1.105 $Y=0.765 $X2=0 $Y2=0
cc_157 N_B2_c_161_n N_VGND_c_483_n 0.00471988f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_158 N_B2_c_161_n N_VGND_c_485_n 0.00389079f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B2_c_163_n N_VGND_c_485_n 0.00397473f $X=1.76 $Y=1.16 $X2=0 $Y2=0
cc_160 B2 N_VGND_c_485_n 0.0256744f $X=1.105 $Y=0.765 $X2=0 $Y2=0
cc_161 N_B2_c_161_n N_VGND_c_486_n 0.00797598f $X=1.835 $Y=0.995 $X2=0 $Y2=0
cc_162 B2 N_VGND_c_486_n 0.00309731f $X=1.105 $Y=0.765 $X2=0 $Y2=0
cc_163 N_B1_c_198_n N_A1_c_238_n 0.0218401f $X=2.34 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_164 N_B1_c_199_n N_A1_c_239_n 0.0460562f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_165 N_B1_c_200_n N_A1_c_239_n 0.0011722f $X=2.557 $Y=1.245 $X2=0 $Y2=0
cc_166 B1 N_A1_c_239_n 0.0039184f $X=2.46 $Y=1.445 $X2=0 $Y2=0
cc_167 N_B1_c_198_n A1 0.00108273f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_168 N_B1_c_199_n A1 7.1502e-19 $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B1_c_200_n A1 0.0116995f $X=2.557 $Y=1.245 $X2=0 $Y2=0
cc_170 B1 A1 0.00525992f $X=2.46 $Y=1.445 $X2=0 $Y2=0
cc_171 B1 A2 0.00875757f $X=2.46 $Y=1.445 $X2=0 $Y2=0
cc_172 N_B1_c_199_n N_VPWR_c_376_n 0.00110692f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B1_c_199_n N_VPWR_c_380_n 0.00429453f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B1_c_199_n N_VPWR_c_374_n 0.00611639f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_175 B1 N_A_319_297#_M1005_d 0.00293265f $X=2.46 $Y=1.445 $X2=0 $Y2=0
cc_176 N_B1_c_199_n N_A_319_297#_c_445_n 0.0137415f $X=2.425 $Y=1.41 $X2=0 $Y2=0
cc_177 B1 N_A_319_297#_c_447_n 0.0077591f $X=2.46 $Y=1.445 $X2=0 $Y2=0
cc_178 N_B1_c_198_n N_VGND_c_483_n 0.00428026f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B1_c_198_n N_VGND_c_486_n 0.00643382f $X=2.34 $Y=0.995 $X2=0 $Y2=0
cc_180 N_A1_c_239_n N_A2_c_272_n 0.0473494f $X=2.895 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_181 A1 N_A2_c_272_n 3.67601e-19 $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_182 N_A1_c_238_n N_A2_c_273_n 0.0180892f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_183 A1 N_A2_c_273_n 0.0017862f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_184 N_A1_c_238_n A2 0.00149717f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_185 N_A1_c_239_n A2 0.00503701f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_186 A1 A2 0.0711977f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_187 N_A1_c_239_n N_VPWR_c_376_n 0.0132763f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A1_c_239_n N_VPWR_c_380_n 0.00323221f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A1_c_239_n N_VPWR_c_374_n 0.00395348f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A1_c_239_n N_A_319_297#_c_454_n 0.0160917f $X=2.895 $Y=1.41 $X2=0 $Y2=0
cc_191 A1 N_A_319_297#_c_454_n 0.00829823f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_192 N_A1_c_238_n N_VGND_c_483_n 0.00494995f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_193 A1 N_VGND_c_483_n 0.00816915f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_194 N_A1_c_238_n N_VGND_c_486_n 0.0091727f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_195 A1 N_VGND_c_486_n 0.0090742f $X=2.9 $Y=0.425 $X2=0 $Y2=0
cc_196 A1 A_589_47# 0.00660945f $X=2.9 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_197 N_A2_c_273_n N_A3_c_307_n 0.0404083f $X=3.55 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_198 A2 N_A3_c_307_n 0.00363067f $X=3.47 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_199 N_A2_c_272_n N_A3_c_310_n 0.0219414f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_200 A2 N_A3_c_310_n 0.00108197f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_201 N_A2_c_272_n A3 7.78486e-19 $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_202 A2 A3 0.0186433f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_203 N_A2_c_272_n N_A3_c_309_n 0.0255549f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_204 A2 N_A3_c_309_n 0.00212107f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_205 A2 N_VPWR_M1002_d 0.00292509f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_206 N_A2_c_272_n N_VPWR_c_376_n 0.00682201f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_272_n N_VPWR_c_378_n 0.00125077f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A2_c_272_n N_VPWR_c_381_n 0.0053025f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A2_c_272_n N_VPWR_c_374_n 0.00754605f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A2_c_272_n N_A_319_297#_c_454_n 0.0128873f $X=3.525 $Y=1.41 $X2=0 $Y2=0
cc_211 A2 N_A_319_297#_c_454_n 0.0187217f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_212 N_A2_c_272_n N_A_319_297#_c_458_n 3.21564e-19 $X=3.525 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A2_c_273_n N_VGND_c_482_n 0.00238769f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A2_c_273_n N_VGND_c_483_n 0.00390689f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_215 A2 N_VGND_c_483_n 0.00956464f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_216 N_A2_c_273_n N_VGND_c_486_n 0.00601726f $X=3.55 $Y=0.995 $X2=0 $Y2=0
cc_217 A2 N_VGND_c_486_n 0.0108789f $X=3.47 $Y=0.425 $X2=0 $Y2=0
cc_218 A2 A_589_47# 0.00563257f $X=3.47 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_219 A3 N_VPWR_M1006_d 0.00587217f $X=4.175 $Y=1.105 $X2=0 $Y2=0
cc_220 N_A3_c_310_n N_VPWR_c_378_n 0.0188674f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_221 A3 N_VPWR_c_378_n 0.0144066f $X=4.175 $Y=1.105 $X2=0 $Y2=0
cc_222 N_A3_c_309_n N_VPWR_c_378_n 0.0022376f $X=3.995 $Y=1.202 $X2=0 $Y2=0
cc_223 N_A3_c_310_n N_VPWR_c_381_n 0.00427505f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A3_c_310_n N_VPWR_c_374_n 0.00735499f $X=3.995 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A3_c_307_n N_VGND_c_482_n 0.0167063f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_226 A3 N_VGND_c_482_n 0.018723f $X=4.175 $Y=1.105 $X2=0 $Y2=0
cc_227 N_A3_c_309_n N_VGND_c_482_n 0.00578686f $X=3.995 $Y=1.202 $X2=0 $Y2=0
cc_228 N_A3_c_307_n N_VGND_c_483_n 0.0046653f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_229 N_A3_c_307_n N_VGND_c_486_n 0.00799591f $X=3.97 $Y=0.995 $X2=0 $Y2=0
cc_230 N_X_c_341_n N_VPWR_M1000_s 0.00346733f $X=1.115 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_231 N_X_c_341_n N_VPWR_c_375_n 0.0203395f $X=1.115 $Y=1.87 $X2=0 $Y2=0
cc_232 N_X_c_346_n N_VPWR_c_375_n 0.0208109f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_233 X N_VPWR_c_375_n 0.0257801f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_234 X N_VPWR_c_379_n 0.0146267f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_235 N_X_c_346_n N_VPWR_c_380_n 0.0118139f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_236 N_X_M1000_d N_VPWR_c_374_n 0.00248768f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_237 N_X_M1003_d N_VPWR_c_374_n 0.00391905f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_238 N_X_c_341_n N_VPWR_c_374_n 0.0134894f $X=1.115 $Y=1.87 $X2=0 $Y2=0
cc_239 N_X_c_346_n N_VPWR_c_374_n 0.00646998f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_240 X N_VPWR_c_374_n 0.00801045f $X=0.15 $Y=2.125 $X2=0 $Y2=0
cc_241 N_X_c_346_n N_A_319_297#_c_443_n 0.0225975f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_242 N_X_c_346_n N_A_319_297#_c_460_n 0.00811595f $X=1.2 $Y=1.95 $X2=0 $Y2=0
cc_243 N_X_c_337_n N_VGND_M1001_d 9.38157e-19 $X=0.73 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_244 N_X_c_332_n N_VGND_M1001_d 0.0111686f $X=0.24 $Y=0.825 $X2=-0.19
+ $Y2=-0.24
cc_245 X N_VGND_M1001_d 0.0029848f $X=0.235 $Y=0.85 $X2=-0.19 $Y2=-0.24
cc_246 N_X_c_337_n N_VGND_c_480_n 0.00296116f $X=0.73 $Y=0.74 $X2=0 $Y2=0
cc_247 N_X_c_332_n N_VGND_c_480_n 0.0161059f $X=0.24 $Y=0.825 $X2=0 $Y2=0
cc_248 N_X_c_337_n N_VGND_c_484_n 0.00683865f $X=0.73 $Y=0.74 $X2=0 $Y2=0
cc_249 N_X_M1001_s N_VGND_c_486_n 0.0044638f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_250 N_X_c_337_n N_VGND_c_486_n 0.0126594f $X=0.73 $Y=0.74 $X2=0 $Y2=0
cc_251 N_X_c_332_n N_VGND_c_486_n 0.00107851f $X=0.24 $Y=0.825 $X2=0 $Y2=0
cc_252 N_VPWR_c_374_n N_A_319_297#_M1008_s 0.00356385f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_253 N_VPWR_c_374_n N_A_319_297#_M1005_d 0.00263241f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_254 N_VPWR_c_374_n N_A_319_297#_M1011_d 0.00470726f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_255 N_VPWR_c_376_n N_A_319_297#_c_445_n 0.0141783f $X=3.13 $Y=2.225 $X2=0
+ $Y2=0
cc_256 N_VPWR_c_380_n N_A_319_297#_c_445_n 0.0534447f $X=2.915 $Y=2.72 $X2=0
+ $Y2=0
cc_257 N_VPWR_c_374_n N_A_319_297#_c_445_n 0.0334225f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_258 N_VPWR_c_380_n N_A_319_297#_c_460_n 0.0119545f $X=2.915 $Y=2.72 $X2=0
+ $Y2=0
cc_259 N_VPWR_c_374_n N_A_319_297#_c_460_n 0.006547f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_260 N_VPWR_c_376_n N_A_319_297#_c_449_n 0.0115352f $X=3.13 $Y=2.225 $X2=0
+ $Y2=0
cc_261 N_VPWR_M1002_d N_A_319_297#_c_454_n 0.0135729f $X=2.985 $Y=1.485 $X2=0
+ $Y2=0
cc_262 N_VPWR_c_376_n N_A_319_297#_c_454_n 0.0243049f $X=3.13 $Y=2.225 $X2=0
+ $Y2=0
cc_263 N_VPWR_c_380_n N_A_319_297#_c_454_n 0.00180073f $X=2.915 $Y=2.72 $X2=0
+ $Y2=0
cc_264 N_VPWR_c_381_n N_A_319_297#_c_454_n 0.00422212f $X=4.015 $Y=2.72 $X2=0
+ $Y2=0
cc_265 N_VPWR_c_374_n N_A_319_297#_c_454_n 0.0140634f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_266 N_VPWR_c_376_n N_A_319_297#_c_458_n 0.0138781f $X=3.13 $Y=2.225 $X2=0
+ $Y2=0
cc_267 N_VPWR_c_378_n N_A_319_297#_c_458_n 0.0415036f $X=4.23 $Y=2 $X2=0 $Y2=0
cc_268 N_VPWR_c_381_n N_A_319_297#_c_458_n 0.011801f $X=4.015 $Y=2.72 $X2=0
+ $Y2=0
cc_269 N_VPWR_c_374_n N_A_319_297#_c_458_n 0.00646745f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_270 N_VGND_c_486_n A_382_47# 0.00435064f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_271 N_VGND_c_486_n A_589_47# 0.0105864f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_272 N_VGND_c_486_n A_725_47# 0.0107316f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
