# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb4to1_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb4to1_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.740000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[0]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.335000 1.055000 0.730000 1.325000 ;
        RECT 0.560000 0.395000 0.835000 0.625000 ;
        RECT 0.560000 0.625000 0.730000 1.055000 ;
    END
  END D[0]
  PIN D[1]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.765000 0.395000 4.040000 0.625000 ;
        RECT 3.870000 0.625000 4.040000 1.055000 ;
        RECT 3.870000 1.055000 4.265000 1.325000 ;
    END
  END D[1]
  PIN D[2]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.475000 1.055000 4.870000 1.325000 ;
        RECT 4.700000 0.395000 4.975000 0.625000 ;
        RECT 4.700000 0.625000 4.870000 1.055000 ;
    END
  END D[2]
  PIN D[3]
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.905000 0.395000 8.180000 0.625000 ;
        RECT 8.010000 0.625000 8.180000 1.055000 ;
        RECT 8.010000 1.055000 8.405000 1.325000 ;
    END
  END D[3]
  PIN S[0]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.805000 0.945000 2.155000 1.295000 ;
    END
  END S[0]
  PIN S[1]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.945000 2.795000 1.295000 ;
    END
  END S[1]
  PIN S[2]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.945000 0.945000 6.295000 1.295000 ;
    END
  END S[2]
  PIN S[3]
    ANTENNAGATEAREA  0.336000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.585000 0.945000 6.935000 1.295000 ;
    END
  END S[3]
  PIN VGND
    ANTENNADIFFAREA  0.999700 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.740000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  1.690000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 8.740000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  1.426400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1.005000 1.755000 1.295000 1.800000 ;
        RECT 1.005000 1.800000 7.735000 1.940000 ;
        RECT 1.005000 1.940000 1.295000 1.985000 ;
        RECT 3.305000 1.755000 3.595000 1.800000 ;
        RECT 3.305000 1.940000 3.595000 1.985000 ;
        RECT 5.145000 1.755000 5.435000 1.800000 ;
        RECT 5.145000 1.940000 5.435000 1.985000 ;
        RECT 7.445000 1.755000 7.735000 1.800000 ;
        RECT 7.445000 1.940000 7.735000 1.985000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 8.740000 0.085000 ;
      RECT 0.000000  2.635000 8.740000 2.805000 ;
      RECT 0.095000  1.495000 0.425000 2.635000 ;
      RECT 0.130000  0.085000 0.390000 0.885000 ;
      RECT 0.900000  0.835000 1.290000 1.005000 ;
      RECT 0.900000  1.005000 1.070000 1.755000 ;
      RECT 0.900000  1.755000 1.295000 1.805000 ;
      RECT 0.900000  1.805000 1.420000 1.985000 ;
      RECT 1.045000  0.330000 1.290000 0.835000 ;
      RECT 1.090000  1.985000 1.420000 2.465000 ;
      RECT 1.240000  1.175000 1.630000 1.465000 ;
      RECT 1.240000  1.465000 1.940000 1.505000 ;
      RECT 1.460000  0.585000 1.900000 0.755000 ;
      RECT 1.460000  0.755000 1.630000 1.175000 ;
      RECT 1.460000  1.505000 1.940000 1.635000 ;
      RECT 1.610000  1.635000 1.940000 2.465000 ;
      RECT 1.650000  0.330000 1.900000 0.585000 ;
      RECT 2.135000  0.085000 2.465000 0.660000 ;
      RECT 2.165000  1.465000 2.465000 2.635000 ;
      RECT 2.660000  1.465000 3.360000 1.505000 ;
      RECT 2.660000  1.505000 3.140000 1.635000 ;
      RECT 2.660000  1.635000 2.990000 2.465000 ;
      RECT 2.700000  0.330000 2.950000 0.585000 ;
      RECT 2.700000  0.585000 3.140000 0.755000 ;
      RECT 2.970000  0.755000 3.140000 1.175000 ;
      RECT 2.970000  1.175000 3.360000 1.465000 ;
      RECT 3.180000  1.805000 3.700000 1.985000 ;
      RECT 3.180000  1.985000 3.510000 2.465000 ;
      RECT 3.305000  1.755000 3.700000 1.805000 ;
      RECT 3.310000  0.330000 3.555000 0.835000 ;
      RECT 3.310000  0.835000 3.700000 1.005000 ;
      RECT 3.530000  1.005000 3.700000 1.755000 ;
      RECT 4.175000  1.495000 4.565000 2.635000 ;
      RECT 4.210000  0.085000 4.530000 0.885000 ;
      RECT 5.040000  0.835000 5.430000 1.005000 ;
      RECT 5.040000  1.005000 5.210000 1.755000 ;
      RECT 5.040000  1.755000 5.435000 1.805000 ;
      RECT 5.040000  1.805000 5.560000 1.985000 ;
      RECT 5.185000  0.330000 5.430000 0.835000 ;
      RECT 5.230000  1.985000 5.560000 2.465000 ;
      RECT 5.380000  1.175000 5.770000 1.465000 ;
      RECT 5.380000  1.465000 6.080000 1.505000 ;
      RECT 5.600000  0.585000 6.040000 0.755000 ;
      RECT 5.600000  0.755000 5.770000 1.175000 ;
      RECT 5.600000  1.505000 6.080000 1.635000 ;
      RECT 5.750000  1.635000 6.080000 2.465000 ;
      RECT 5.790000  0.330000 6.040000 0.585000 ;
      RECT 6.275000  0.085000 6.605000 0.660000 ;
      RECT 6.275000  1.465000 6.575000 2.635000 ;
      RECT 6.800000  1.465000 7.500000 1.505000 ;
      RECT 6.800000  1.505000 7.280000 1.635000 ;
      RECT 6.800000  1.635000 7.130000 2.465000 ;
      RECT 6.840000  0.330000 7.090000 0.585000 ;
      RECT 6.840000  0.585000 7.280000 0.755000 ;
      RECT 7.110000  0.755000 7.280000 1.175000 ;
      RECT 7.110000  1.175000 7.500000 1.465000 ;
      RECT 7.320000  1.805000 7.840000 1.985000 ;
      RECT 7.320000  1.985000 7.650000 2.465000 ;
      RECT 7.445000  1.755000 7.840000 1.805000 ;
      RECT 7.450000  0.330000 7.695000 0.835000 ;
      RECT 7.450000  0.835000 7.840000 1.005000 ;
      RECT 7.670000  1.005000 7.840000 1.755000 ;
      RECT 8.315000  1.495000 8.645000 2.635000 ;
      RECT 8.350000  0.085000 8.610000 0.885000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  1.785000 1.235000 1.955000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  1.785000 3.535000 1.955000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  1.785000 5.375000 1.955000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  1.785000 7.675000 1.955000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb4to1_1
END LIBRARY
