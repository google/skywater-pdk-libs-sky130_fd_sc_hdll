* File: sky130_fd_sc_hdll__clkmux2_2.pxi.spice
* Created: Wed Sep  2 08:27:04 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_79_199# N_A_79_199#_M1013_d
+ N_A_79_199#_M1011_d N_A_79_199#_c_83_n N_A_79_199#_M1000_g N_A_79_199#_M1003_g
+ N_A_79_199#_M1010_g N_A_79_199#_c_84_n N_A_79_199#_M1005_g N_A_79_199#_c_79_n
+ N_A_79_199#_c_80_n N_A_79_199#_c_147_p N_A_79_199#_c_81_n N_A_79_199#_c_109_p
+ N_A_79_199#_c_92_p N_A_79_199#_c_103_p N_A_79_199#_c_98_p N_A_79_199#_c_82_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_79_199#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%S N_S_c_175_n N_S_M1002_g N_S_M1008_g
+ N_S_c_177_n N_S_M1009_g N_S_M1004_g N_S_c_183_n N_S_c_201_n N_S_c_249_p
+ N_S_c_184_n N_S_c_224_p N_S_c_241_p N_S_c_179_n N_S_c_180_n S S
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%S
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A1 N_A1_M1013_g N_A1_c_271_n N_A1_M1006_g
+ N_A1_c_272_n N_A1_c_273_n N_A1_c_288_n N_A1_c_290_n A1 A1
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A1
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A0 N_A0_c_343_n N_A0_M1011_g N_A0_c_344_n
+ N_A0_c_345_n N_A0_M1007_g N_A0_c_340_n A0 N_A0_c_341_n N_A0_c_342_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A0
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_741_21# N_A_741_21#_M1004_d
+ N_A_741_21#_M1009_d N_A_741_21#_M1001_g N_A_741_21#_c_390_n
+ N_A_741_21#_c_399_n N_A_741_21#_M1012_g N_A_741_21#_c_391_n
+ N_A_741_21#_c_392_n N_A_741_21#_c_393_n N_A_741_21#_c_394_n
+ N_A_741_21#_c_395_n N_A_741_21#_c_400_n N_A_741_21#_c_396_n
+ N_A_741_21#_c_397_n PM_SKY130_FD_SC_HDLL__CLKMUX2_2%A_741_21#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VPWR N_VPWR_M1000_d N_VPWR_M1005_d
+ N_VPWR_M1012_d N_VPWR_c_458_n N_VPWR_c_459_n N_VPWR_c_460_n N_VPWR_c_461_n
+ N_VPWR_c_462_n N_VPWR_c_463_n N_VPWR_c_464_n VPWR N_VPWR_c_465_n
+ N_VPWR_c_457_n N_VPWR_c_467_n PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%X N_X_M1003_d N_X_M1000_s N_X_c_511_n X X X
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%X
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VGND N_VGND_M1003_s N_VGND_M1010_s
+ N_VGND_M1001_d N_VGND_c_537_n N_VGND_c_538_n N_VGND_c_539_n VGND
+ N_VGND_c_540_n N_VGND_c_541_n N_VGND_c_542_n N_VGND_c_543_n N_VGND_c_544_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_2%VGND
cc_1 VNB N_A_79_199#_M1003_g 0.0313714f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_2 VNB N_A_79_199#_M1010_g 0.0241174f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_3 VNB N_A_79_199#_c_79_n 0.00195867f $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=1.16
cc_4 VNB N_A_79_199#_c_80_n 0.0184511f $X=-0.19 $Y=-0.24 $X2=1.895 $Y2=0.74
cc_5 VNB N_A_79_199#_c_81_n 0.0051489f $X=-0.19 $Y=-0.24 $X2=1.985 $Y2=1.955
cc_6 VNB N_A_79_199#_c_82_n 0.0586569f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.202
cc_7 VNB N_S_c_175_n 0.0252834f $X=-0.19 $Y=-0.24 $X2=2.195 $Y2=0.235
cc_8 VNB N_S_M1008_g 0.0320387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_S_c_177_n 0.0209544f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_10 VNB N_S_M1004_g 0.0335245f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_S_c_179_n 5.74134e-19 $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=1.16
cc_12 VNB N_S_c_180_n 0.0037048f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=0.74
cc_13 VNB N_A1_M1013_g 0.0228368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_271_n 0.0236121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_272_n 0.00497652f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_16 VNB N_A1_c_273_n 0.0366468f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_17 VNB A1 0.00997405f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_18 VNB N_A0_M1007_g 0.0254644f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_19 VNB N_A0_c_340_n 0.00955013f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_20 VNB N_A0_c_341_n 0.028761f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_21 VNB N_A0_c_342_n 0.00455985f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_22 VNB N_A_741_21#_M1001_g 0.02497f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_23 VNB N_A_741_21#_c_390_n 0.0070328f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_24 VNB N_A_741_21#_c_391_n 5.32232e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_25 VNB N_A_741_21#_c_392_n 0.0308747f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_26 VNB N_A_741_21#_c_393_n 0.00551271f $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=0.825
cc_27 VNB N_A_741_21#_c_394_n 8.46441e-19 $X=-0.19 $Y=-0.24 $X2=1.06 $Y2=1.16
cc_28 VNB N_A_741_21#_c_395_n 0.0158392f $X=-0.19 $Y=-0.24 $X2=1.145 $Y2=0.74
cc_29 VNB N_A_741_21#_c_396_n 0.0211382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_741_21#_c_397_n 0.0166335f $X=-0.19 $Y=-0.24 $X2=2.07 $Y2=2.04
cc_31 VNB N_VPWR_c_457_n 0.212805f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_32 VNB X 0.00145735f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_33 VNB N_VGND_c_537_n 0.0113126f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.995
cc_34 VNB N_VGND_c_538_n 0.00451978f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=0.495
cc_35 VNB N_VGND_c_539_n 0.00301626f $X=-0.19 $Y=-0.24 $X2=0.93 $Y2=0.495
cc_36 VNB N_VGND_c_540_n 0.0152053f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.985
cc_37 VNB N_VGND_c_541_n 0.0702689f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_VGND_c_542_n 0.0249556f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=2.04
cc_39 VNB N_VGND_c_543_n 0.265148f $X=-0.19 $Y=-0.24 $X2=2.415 $Y2=2.04
cc_40 VNB N_VGND_c_544_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.202
cc_41 VPB N_A_79_199#_c_83_n 0.0207617f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_42 VPB N_A_79_199#_c_84_n 0.0174347f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_43 VPB N_A_79_199#_c_79_n 0.00108432f $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.16
cc_44 VPB N_A_79_199#_c_81_n 0.00429564f $X=-0.19 $Y=1.305 $X2=1.985 $Y2=1.955
cc_45 VPB N_A_79_199#_c_82_n 0.0280519f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_46 VPB N_S_c_175_n 0.0328546f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=0.235
cc_47 VPB N_S_c_177_n 0.0330042f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_48 VPB N_S_c_183_n 0.0014488f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_49 VPB N_S_c_184_n 6.63611e-19 $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_50 VPB N_S_c_179_n 6.16925e-19 $X=-0.19 $Y=1.305 $X2=1.06 $Y2=1.16
cc_51 VPB N_S_c_180_n 0.00125389f $X=-0.19 $Y=1.305 $X2=1.145 $Y2=0.74
cc_52 VPB S 0.00455426f $X=-0.19 $Y=1.305 $X2=2.495 $Y2=0.455
cc_53 VPB N_A1_c_271_n 0.0304527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A1_c_272_n 0.00280866f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_55 VPB A1 0.00558813f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_56 VPB N_A0_c_343_n 0.020637f $X=-0.19 $Y=1.305 $X2=2.195 $Y2=0.235
cc_57 VPB N_A0_c_344_n 0.0406981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A0_c_345_n 0.00988826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_59 VPB N_A0_c_340_n 8.40892e-19 $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_60 VPB N_A0_c_342_n 0.0023903f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_61 VPB N_A_741_21#_c_390_n 0.00378234f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_62 VPB N_A_741_21#_c_399_n 0.0224682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_741_21#_c_400_n 0.0267191f $X=-0.19 $Y=1.305 $X2=2.495 $Y2=0.455
cc_64 VPB N_A_741_21#_c_396_n 0.0225129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_458_n 0.0111924f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.995
cc_66 VPB N_VPWR_c_459_n 0.00513559f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_67 VPB N_VPWR_c_460_n 0.0186422f $X=-0.19 $Y=1.305 $X2=0.93 $Y2=0.495
cc_68 VPB N_VPWR_c_461_n 0.00518f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_69 VPB N_VPWR_c_462_n 0.00497347f $X=-0.19 $Y=1.305 $X2=1.895 $Y2=0.74
cc_70 VPB N_VPWR_c_463_n 0.0638297f $X=-0.19 $Y=1.305 $X2=1.985 $Y2=1.955
cc_71 VPB N_VPWR_c_464_n 0.00439107f $X=-0.19 $Y=1.305 $X2=2.07 $Y2=0.437
cc_72 VPB N_VPWR_c_465_n 0.0232568f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_73 VPB N_VPWR_c_457_n 0.0518412f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.202
cc_74 VPB N_VPWR_c_467_n 0.0047828f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB X 0.0015278f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=0.495
cc_76 N_A_79_199#_c_84_n N_S_c_175_n 0.0152976f $X=0.965 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_79_199#_c_79_n N_S_c_175_n 0.00107569f $X=1.06 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_79_199#_c_80_n N_S_c_175_n 0.00246858f $X=1.895 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_79_199#_c_81_n N_S_c_175_n 0.00361956f $X=1.985 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_79_199#_c_92_p N_S_c_175_n 6.54365e-19 $X=2.07 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_81 N_A_79_199#_c_82_n N_S_c_175_n 0.0237573f $X=0.965 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_82 N_A_79_199#_M1010_g N_S_M1008_g 0.013677f $X=0.93 $Y=0.495 $X2=0 $Y2=0
cc_83 N_A_79_199#_c_79_n N_S_M1008_g 0.00297788f $X=1.06 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_79_199#_c_80_n N_S_M1008_g 0.0133748f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_85 N_A_79_199#_c_81_n N_S_M1008_g 0.00343808f $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_86 N_A_79_199#_c_98_p N_S_M1008_g 0.00699958f $X=1.982 $Y=0.54 $X2=0 $Y2=0
cc_87 N_A_79_199#_c_84_n N_S_c_183_n 6.47769e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A_79_199#_c_82_n N_S_c_183_n 4.6068e-19 $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_89 N_A_79_199#_M1011_d N_S_c_201_n 0.02385f $X=2.27 $Y=1.545 $X2=0 $Y2=0
cc_90 N_A_79_199#_c_92_p N_S_c_201_n 0.0100943f $X=2.07 $Y=2.04 $X2=0 $Y2=0
cc_91 N_A_79_199#_c_103_p N_S_c_201_n 0.0768599f $X=3.13 $Y=2.04 $X2=0 $Y2=0
cc_92 N_A_79_199#_c_79_n N_S_c_180_n 0.014361f $X=1.06 $Y=1.16 $X2=0 $Y2=0
cc_93 N_A_79_199#_c_80_n N_S_c_180_n 0.0211311f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_94 N_A_79_199#_c_81_n N_S_c_180_n 0.0573317f $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_95 N_A_79_199#_c_82_n N_S_c_180_n 0.00127031f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_96 N_A_79_199#_c_81_n N_A1_M1013_g 2.53446e-19 $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_97 N_A_79_199#_c_109_p N_A1_M1013_g 0.0166772f $X=2.495 $Y=0.455 $X2=0 $Y2=0
cc_98 N_A_79_199#_c_98_p N_A1_M1013_g 0.0116551f $X=1.982 $Y=0.54 $X2=0 $Y2=0
cc_99 N_A_79_199#_c_103_p N_A1_c_271_n 0.00495514f $X=3.13 $Y=2.04 $X2=0 $Y2=0
cc_100 N_A_79_199#_M1011_d N_A1_c_272_n 0.00263273f $X=2.27 $Y=1.545 $X2=0 $Y2=0
cc_101 N_A_79_199#_c_81_n N_A1_c_272_n 0.053476f $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_102 N_A_79_199#_c_109_p N_A1_c_272_n 0.0126222f $X=2.495 $Y=0.455 $X2=0 $Y2=0
cc_103 N_A_79_199#_c_98_p N_A1_c_272_n 0.00119858f $X=1.982 $Y=0.54 $X2=0 $Y2=0
cc_104 N_A_79_199#_c_81_n N_A1_c_273_n 0.0072307f $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_105 N_A_79_199#_c_109_p N_A1_c_273_n 0.00418341f $X=2.495 $Y=0.455 $X2=0
+ $Y2=0
cc_106 N_A_79_199#_M1011_d N_A1_c_288_n 0.0262928f $X=2.27 $Y=1.545 $X2=0 $Y2=0
cc_107 N_A_79_199#_c_103_p N_A1_c_288_n 0.0639496f $X=3.13 $Y=2.04 $X2=0 $Y2=0
cc_108 N_A_79_199#_M1011_d N_A1_c_290_n 9.09665e-19 $X=2.27 $Y=1.545 $X2=0 $Y2=0
cc_109 N_A_79_199#_c_103_p N_A1_c_290_n 0.00891696f $X=3.13 $Y=2.04 $X2=0 $Y2=0
cc_110 N_A_79_199#_c_81_n N_A0_c_343_n 0.00341414f $X=1.985 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_111 N_A_79_199#_c_103_p N_A0_c_343_n 0.0138951f $X=3.13 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_112 N_A_79_199#_c_103_p N_A0_c_344_n 0.00104228f $X=3.13 $Y=2.04 $X2=0 $Y2=0
cc_113 N_A_79_199#_c_81_n N_A0_c_345_n 0.00178945f $X=1.985 $Y=1.955 $X2=0 $Y2=0
cc_114 N_A_79_199#_c_109_p N_A0_M1007_g 0.00342458f $X=2.495 $Y=0.455 $X2=0
+ $Y2=0
cc_115 N_A_79_199#_c_98_p N_A0_M1007_g 8.26503e-19 $X=1.982 $Y=0.54 $X2=0 $Y2=0
cc_116 N_A_79_199#_c_109_p N_A0_c_342_n 0.0299622f $X=2.495 $Y=0.455 $X2=0 $Y2=0
cc_117 N_A_79_199#_c_83_n N_VPWR_c_459_n 0.00474293f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_118 N_A_79_199#_c_83_n N_VPWR_c_460_n 0.00658436f $X=0.495 $Y=1.41 $X2=0
+ $Y2=0
cc_119 N_A_79_199#_c_84_n N_VPWR_c_460_n 0.00673617f $X=0.965 $Y=1.41 $X2=0
+ $Y2=0
cc_120 N_A_79_199#_c_84_n N_VPWR_c_461_n 0.0032377f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A_79_199#_c_79_n N_VPWR_c_461_n 0.00431418f $X=1.06 $Y=1.16 $X2=0 $Y2=0
cc_122 N_A_79_199#_c_80_n N_VPWR_c_461_n 0.00540521f $X=1.895 $Y=0.74 $X2=0
+ $Y2=0
cc_123 N_A_79_199#_c_82_n N_VPWR_c_461_n 0.00198236f $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_124 N_A_79_199#_M1011_d N_VPWR_c_457_n 0.00817943f $X=2.27 $Y=1.545 $X2=0
+ $Y2=0
cc_125 N_A_79_199#_c_83_n N_VPWR_c_457_n 0.0122976f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_126 N_A_79_199#_c_84_n N_VPWR_c_457_n 0.0120826f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_79_199#_c_83_n N_X_c_511_n 0.00201828f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_79_199#_c_84_n N_X_c_511_n 0.00280049f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_79_199#_c_82_n N_X_c_511_n 0.00176607f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_130 N_A_79_199#_c_83_n X 0.00423085f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_79_199#_M1003_g X 0.0221059f $X=0.51 $Y=0.495 $X2=0 $Y2=0
cc_132 N_A_79_199#_M1010_g X 0.00216963f $X=0.93 $Y=0.495 $X2=0 $Y2=0
cc_133 N_A_79_199#_c_84_n X 0.00209972f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_79_199#_c_79_n X 0.0355257f $X=1.06 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_79_199#_c_147_p X 0.00992523f $X=1.145 $Y=0.74 $X2=0 $Y2=0
cc_136 N_A_79_199#_c_82_n X 0.0397638f $X=0.965 $Y=1.202 $X2=0 $Y2=0
cc_137 N_A_79_199#_c_83_n X 0.00972579f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_79_199#_c_84_n X 0.00892448f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_79_199#_c_81_n A_335_309# 0.00526835f $X=1.985 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_140 N_A_79_199#_c_92_p A_335_309# 0.00300196f $X=2.07 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_141 N_A_79_199#_c_80_n N_VGND_M1010_s 0.00244694f $X=1.895 $Y=0.74 $X2=0
+ $Y2=0
cc_142 N_A_79_199#_c_147_p N_VGND_M1010_s 8.75693e-19 $X=1.145 $Y=0.74 $X2=0
+ $Y2=0
cc_143 N_A_79_199#_M1003_g N_VGND_c_538_n 0.00426039f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_144 N_A_79_199#_M1003_g N_VGND_c_539_n 6.01892e-19 $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_145 N_A_79_199#_M1010_g N_VGND_c_539_n 0.00756751f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_146 N_A_79_199#_c_80_n N_VGND_c_539_n 0.0160584f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_147 N_A_79_199#_c_147_p N_VGND_c_539_n 0.00929542f $X=1.145 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_79_199#_c_98_p N_VGND_c_539_n 0.00832873f $X=1.982 $Y=0.54 $X2=0
+ $Y2=0
cc_149 N_A_79_199#_c_82_n N_VGND_c_539_n 5.28291e-19 $X=0.965 $Y=1.202 $X2=0
+ $Y2=0
cc_150 N_A_79_199#_M1003_g N_VGND_c_540_n 0.00541359f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_151 N_A_79_199#_M1010_g N_VGND_c_540_n 0.0046653f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_152 N_A_79_199#_c_80_n N_VGND_c_541_n 0.00916117f $X=1.895 $Y=0.74 $X2=0
+ $Y2=0
cc_153 N_A_79_199#_c_109_p N_VGND_c_541_n 0.0319877f $X=2.495 $Y=0.455 $X2=0
+ $Y2=0
cc_154 N_A_79_199#_c_98_p N_VGND_c_541_n 0.0102622f $X=1.982 $Y=0.54 $X2=0 $Y2=0
cc_155 N_A_79_199#_M1013_d N_VGND_c_543_n 0.00824573f $X=2.195 $Y=0.235 $X2=0
+ $Y2=0
cc_156 N_A_79_199#_M1003_g N_VGND_c_543_n 0.0106446f $X=0.51 $Y=0.495 $X2=0
+ $Y2=0
cc_157 N_A_79_199#_M1010_g N_VGND_c_543_n 0.00796766f $X=0.93 $Y=0.495 $X2=0
+ $Y2=0
cc_158 N_A_79_199#_c_80_n N_VGND_c_543_n 0.0152428f $X=1.895 $Y=0.74 $X2=0 $Y2=0
cc_159 N_A_79_199#_c_147_p N_VGND_c_543_n 8.0899e-19 $X=1.145 $Y=0.74 $X2=0
+ $Y2=0
cc_160 N_A_79_199#_c_109_p N_VGND_c_543_n 0.0187496f $X=2.495 $Y=0.455 $X2=0
+ $Y2=0
cc_161 N_A_79_199#_c_98_p N_VGND_c_543_n 0.00662435f $X=1.982 $Y=0.54 $X2=0
+ $Y2=0
cc_162 N_A_79_199#_c_98_p A_337_47# 0.00653116f $X=1.982 $Y=0.54 $X2=-0.19
+ $Y2=-0.24
cc_163 N_S_M1008_g N_A1_M1013_g 0.0156947f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_164 N_S_c_201_n N_A1_c_271_n 0.0140173f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_165 N_S_c_184_n N_A1_c_271_n 3.3557e-19 $X=3.79 $Y=1.63 $X2=0 $Y2=0
cc_166 N_S_c_175_n N_A1_c_273_n 0.0156947f $X=1.585 $Y=1.47 $X2=0 $Y2=0
cc_167 N_S_c_180_n N_A1_c_273_n 2.95407e-19 $X=1.54 $Y=1.16 $X2=0 $Y2=0
cc_168 N_S_c_201_n N_A1_c_288_n 0.00421347f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_169 N_S_c_184_n A1 0.0117446f $X=3.79 $Y=1.63 $X2=0 $Y2=0
cc_170 N_S_c_175_n N_A0_c_343_n 0.0291584f $X=1.585 $Y=1.47 $X2=-0.19 $Y2=-0.24
cc_171 N_S_c_201_n N_A0_c_343_n 0.0135571f $X=3.705 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_172 N_S_c_175_n N_A0_c_345_n 0.00409565f $X=1.585 $Y=1.47 $X2=0 $Y2=0
cc_173 N_S_M1004_g N_A_741_21#_M1001_g 0.0166525f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_174 N_S_c_177_n N_A_741_21#_c_390_n 0.00791167f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_175 N_S_c_179_n N_A_741_21#_c_390_n 0.00114571f $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_176 N_S_c_177_n N_A_741_21#_c_399_n 0.0253237f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_177 N_S_c_201_n N_A_741_21#_c_399_n 0.00665392f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_178 N_S_c_184_n N_A_741_21#_c_399_n 0.00936369f $X=3.79 $Y=1.63 $X2=0 $Y2=0
cc_179 N_S_c_224_p N_A_741_21#_c_399_n 0.0169742f $X=3.79 $Y=2.295 $X2=0 $Y2=0
cc_180 N_S_c_179_n N_A_741_21#_c_399_n 9.61528e-19 $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_181 S N_A_741_21#_c_399_n 0.00468862f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_182 N_S_c_177_n N_A_741_21#_c_391_n 4.2108e-19 $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_183 N_S_M1004_g N_A_741_21#_c_391_n 0.00105012f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_184 N_S_c_184_n N_A_741_21#_c_391_n 0.00529971f $X=3.79 $Y=1.63 $X2=0 $Y2=0
cc_185 N_S_c_179_n N_A_741_21#_c_391_n 0.00549551f $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_186 S N_A_741_21#_c_391_n 0.00442941f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_187 N_S_c_177_n N_A_741_21#_c_392_n 0.0078874f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_188 N_S_M1004_g N_A_741_21#_c_392_n 0.00773768f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_189 N_S_c_179_n N_A_741_21#_c_392_n 4.28614e-19 $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_190 S N_A_741_21#_c_392_n 0.00155646f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_191 N_S_c_177_n N_A_741_21#_c_393_n 0.00210123f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_192 N_S_M1004_g N_A_741_21#_c_393_n 0.0151946f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_193 N_S_c_179_n N_A_741_21#_c_393_n 0.0131349f $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_194 S N_A_741_21#_c_393_n 0.00986081f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_195 N_S_c_177_n N_A_741_21#_c_400_n 0.00747341f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_196 N_S_c_241_p N_A_741_21#_c_400_n 6.43652e-19 $X=4.36 $Y=1.44 $X2=0 $Y2=0
cc_197 N_S_c_177_n N_A_741_21#_c_396_n 0.0171101f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_198 N_S_M1004_g N_A_741_21#_c_396_n 0.00462428f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_199 N_S_c_241_p N_A_741_21#_c_396_n 0.0123401f $X=4.36 $Y=1.44 $X2=0 $Y2=0
cc_200 N_S_c_179_n N_A_741_21#_c_396_n 0.0228671f $X=4.35 $Y=1.22 $X2=0 $Y2=0
cc_201 S N_VPWR_M1012_d 0.00577639f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_202 N_S_c_175_n N_VPWR_c_461_n 0.010595f $X=1.585 $Y=1.47 $X2=0 $Y2=0
cc_203 N_S_c_183_n N_VPWR_c_461_n 0.0506953f $X=1.63 $Y=2.295 $X2=0 $Y2=0
cc_204 N_S_c_249_p N_VPWR_c_461_n 0.011874f $X=1.73 $Y=2.38 $X2=0 $Y2=0
cc_205 N_S_c_177_n N_VPWR_c_462_n 0.00324489f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_206 N_S_c_201_n N_VPWR_c_462_n 0.0136491f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_207 N_S_c_224_p N_VPWR_c_462_n 0.0330344f $X=3.79 $Y=2.295 $X2=0 $Y2=0
cc_208 S N_VPWR_c_462_n 0.0129774f $X=4.265 $Y=1.445 $X2=0 $Y2=0
cc_209 N_S_c_175_n N_VPWR_c_463_n 0.00482335f $X=1.585 $Y=1.47 $X2=0 $Y2=0
cc_210 N_S_c_201_n N_VPWR_c_463_n 0.127998f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_211 N_S_c_249_p N_VPWR_c_463_n 0.0118049f $X=1.73 $Y=2.38 $X2=0 $Y2=0
cc_212 N_S_c_177_n N_VPWR_c_465_n 0.00673617f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_213 N_S_c_175_n N_VPWR_c_457_n 0.00805617f $X=1.585 $Y=1.47 $X2=0 $Y2=0
cc_214 N_S_c_177_n N_VPWR_c_457_n 0.0130085f $X=4.375 $Y=1.47 $X2=0 $Y2=0
cc_215 N_S_c_201_n N_VPWR_c_457_n 0.077726f $X=3.705 $Y=2.38 $X2=0 $Y2=0
cc_216 N_S_c_249_p N_VPWR_c_457_n 0.00702939f $X=1.73 $Y=2.38 $X2=0 $Y2=0
cc_217 N_S_c_201_n A_335_309# 0.0111518f $X=3.705 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_218 N_S_c_201_n A_691_309# 0.00646556f $X=3.705 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_219 N_S_M1008_g N_VGND_c_539_n 0.00593008f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_220 N_S_M1008_g N_VGND_c_541_n 0.00428022f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_221 N_S_M1004_g N_VGND_c_541_n 0.00646436f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_222 N_S_M1004_g N_VGND_c_542_n 0.00433717f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_223 N_S_M1008_g N_VGND_c_543_n 0.00672742f $X=1.61 $Y=0.445 $X2=0 $Y2=0
cc_224 N_S_M1004_g N_VGND_c_543_n 0.00761805f $X=4.4 $Y=0.495 $X2=0 $Y2=0
cc_225 N_A1_c_272_n N_A0_c_343_n 0.00409325f $X=2.325 $Y=0.975 $X2=-0.19
+ $Y2=-0.24
cc_226 N_A1_c_290_n N_A0_c_343_n 0.00649866f $X=2.41 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_227 N_A1_c_271_n N_A0_c_344_n 0.00277644f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_228 N_A1_c_272_n N_A0_c_344_n 0.0101853f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_229 N_A1_c_288_n N_A0_c_344_n 0.016411f $X=3.245 $Y=1.7 $X2=0 $Y2=0
cc_230 A1 N_A0_c_344_n 0.00120799f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_231 N_A1_c_272_n N_A0_c_345_n 0.0020234f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_232 N_A1_c_273_n N_A0_c_345_n 0.0292599f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_233 N_A1_M1013_g N_A0_M1007_g 0.0140866f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_234 N_A1_c_272_n N_A0_M1007_g 2.42785e-19 $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_235 A1 N_A0_M1007_g 0.00248702f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A1_c_271_n N_A0_c_340_n 0.00936614f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_237 A1 N_A0_c_340_n 2.12428e-19 $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_238 N_A1_c_271_n N_A0_c_341_n 0.00503691f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_239 N_A1_c_272_n N_A0_c_341_n 0.00486025f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_240 N_A1_c_273_n N_A0_c_341_n 0.0169793f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_241 N_A1_c_288_n N_A0_c_341_n 2.70133e-19 $X=3.245 $Y=1.7 $X2=0 $Y2=0
cc_242 A1 N_A0_c_341_n 0.00144026f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_243 N_A1_M1013_g N_A0_c_342_n 0.00121146f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_244 N_A1_c_271_n N_A0_c_342_n 0.00240846f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_245 N_A1_c_272_n N_A0_c_342_n 0.0256133f $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_246 N_A1_c_273_n N_A0_c_342_n 9.69032e-19 $X=2.325 $Y=0.975 $X2=0 $Y2=0
cc_247 N_A1_c_288_n N_A0_c_342_n 0.0231818f $X=3.245 $Y=1.7 $X2=0 $Y2=0
cc_248 A1 N_A0_c_342_n 0.0929962f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_249 A1 N_A_741_21#_M1001_g 0.0260542f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_250 N_A1_c_271_n N_A_741_21#_c_399_n 0.0556404f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_251 N_A1_c_288_n N_A_741_21#_c_399_n 6.59428e-19 $X=3.245 $Y=1.7 $X2=0 $Y2=0
cc_252 A1 N_A_741_21#_c_399_n 5.7392e-19 $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_253 A1 N_A_741_21#_c_391_n 0.0179199f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_254 N_A1_c_271_n N_A_741_21#_c_392_n 0.0213383f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_255 A1 N_A_741_21#_c_394_n 0.0105375f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_256 N_A1_c_271_n N_VPWR_c_463_n 0.00429453f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_257 N_A1_c_271_n N_VPWR_c_457_n 0.0073872f $X=3.365 $Y=1.47 $X2=0 $Y2=0
cc_258 N_A1_c_288_n A_691_309# 0.0019065f $X=3.245 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_259 A1 A_691_309# 5.87758e-19 $X=3.365 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_260 N_A1_M1013_g N_VGND_c_541_n 0.00357842f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_261 A1 N_VGND_c_541_n 0.041242f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_262 N_A1_M1013_g N_VGND_c_543_n 0.006025f $X=2.12 $Y=0.445 $X2=0 $Y2=0
cc_263 A1 N_VGND_c_543_n 0.0110914f $X=3.365 $Y=0.765 $X2=0 $Y2=0
cc_264 A1 A_570_47# 0.0167608f $X=3.365 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_265 N_A0_c_343_n N_VPWR_c_463_n 0.00429453f $X=2.18 $Y=1.47 $X2=0 $Y2=0
cc_266 N_A0_c_343_n N_VPWR_c_457_n 0.00774138f $X=2.18 $Y=1.47 $X2=0 $Y2=0
cc_267 N_A0_M1007_g N_VGND_c_541_n 0.00435091f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_268 N_A0_c_342_n N_VGND_c_541_n 0.0205158f $X=2.835 $Y=0.98 $X2=0 $Y2=0
cc_269 N_A0_M1007_g N_VGND_c_543_n 0.00904666f $X=2.775 $Y=0.445 $X2=0 $Y2=0
cc_270 N_A0_c_342_n N_VGND_c_543_n 0.0119866f $X=2.835 $Y=0.98 $X2=0 $Y2=0
cc_271 N_A0_c_342_n A_570_47# 0.00656391f $X=2.835 $Y=0.98 $X2=-0.19 $Y2=-0.24
cc_272 N_A_741_21#_c_399_n N_VPWR_c_462_n 0.00744201f $X=3.805 $Y=1.47 $X2=0
+ $Y2=0
cc_273 N_A_741_21#_c_399_n N_VPWR_c_463_n 0.00459563f $X=3.805 $Y=1.47 $X2=0
+ $Y2=0
cc_274 N_A_741_21#_c_400_n N_VPWR_c_465_n 0.0259839f $X=4.61 $Y=2 $X2=0 $Y2=0
cc_275 N_A_741_21#_M1009_d N_VPWR_c_457_n 0.00233913f $X=4.465 $Y=1.545 $X2=0
+ $Y2=0
cc_276 N_A_741_21#_c_399_n N_VPWR_c_457_n 0.00704825f $X=3.805 $Y=1.47 $X2=0
+ $Y2=0
cc_277 N_A_741_21#_c_400_n N_VPWR_c_457_n 0.0151509f $X=4.61 $Y=2 $X2=0 $Y2=0
cc_278 N_A_741_21#_c_393_n N_VGND_M1001_d 0.00234003f $X=4.495 $Y=0.78 $X2=0
+ $Y2=0
cc_279 N_A_741_21#_M1001_g N_VGND_c_541_n 0.023697f $X=3.78 $Y=0.445 $X2=0 $Y2=0
cc_280 N_A_741_21#_c_392_n N_VGND_c_541_n 6.87788e-19 $X=3.87 $Y=1.02 $X2=0
+ $Y2=0
cc_281 N_A_741_21#_c_393_n N_VGND_c_541_n 0.0210008f $X=4.495 $Y=0.78 $X2=0
+ $Y2=0
cc_282 N_A_741_21#_c_394_n N_VGND_c_541_n 0.0115145f $X=3.955 $Y=0.78 $X2=0
+ $Y2=0
cc_283 N_A_741_21#_c_393_n N_VGND_c_542_n 0.00345018f $X=4.495 $Y=0.78 $X2=0
+ $Y2=0
cc_284 N_A_741_21#_c_395_n N_VGND_c_542_n 0.0157596f $X=4.61 $Y=0.455 $X2=0
+ $Y2=0
cc_285 N_A_741_21#_c_397_n N_VGND_c_542_n 0.00189167f $X=4.67 $Y=0.78 $X2=0
+ $Y2=0
cc_286 N_A_741_21#_M1004_d N_VGND_c_543_n 0.00218371f $X=4.475 $Y=0.235 $X2=0
+ $Y2=0
cc_287 N_A_741_21#_M1001_g N_VGND_c_543_n 0.00251647f $X=3.78 $Y=0.445 $X2=0
+ $Y2=0
cc_288 N_A_741_21#_c_393_n N_VGND_c_543_n 0.00766116f $X=4.495 $Y=0.78 $X2=0
+ $Y2=0
cc_289 N_A_741_21#_c_394_n N_VGND_c_543_n 7.21038e-19 $X=3.955 $Y=0.78 $X2=0
+ $Y2=0
cc_290 N_A_741_21#_c_395_n N_VGND_c_543_n 0.0093388f $X=4.61 $Y=0.455 $X2=0
+ $Y2=0
cc_291 N_A_741_21#_c_397_n N_VGND_c_543_n 0.00302259f $X=4.67 $Y=0.78 $X2=0
+ $Y2=0
cc_292 N_VPWR_c_457_n N_X_M1000_s 0.00231261f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_460_n X 0.0196285f $X=1.075 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_c_457_n X 0.0126526f $X=4.83 $Y=2.72 $X2=0 $Y2=0
cc_295 N_VPWR_c_457_n A_335_309# 0.003342f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_296 N_VPWR_c_457_n A_691_309# 0.00208801f $X=4.83 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_297 X N_VGND_c_540_n 0.0151826f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_298 N_X_M1003_d N_VGND_c_543_n 0.00393857f $X=0.585 $Y=0.235 $X2=0 $Y2=0
cc_299 X N_VGND_c_543_n 0.00941829f $X=0.61 $Y=0.425 $X2=0 $Y2=0
cc_300 N_VGND_c_543_n A_337_47# 0.00371776f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
cc_301 N_VGND_c_543_n A_570_47# 0.0188707f $X=4.83 $Y=0 $X2=-0.19 $Y2=-0.24
