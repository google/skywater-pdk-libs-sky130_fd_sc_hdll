* File: sky130_fd_sc_hdll__clkbuf_12.pxi.spice
* Created: Wed Sep  2 08:25:12 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKBUF_12%A N_A_c_137_n N_A_M1002_g N_A_M1009_g
+ N_A_M1022_g N_A_c_138_n N_A_M1013_g N_A_c_139_n N_A_M1019_g N_A_M1028_g
+ N_A_M1031_g N_A_c_140_n N_A_M1027_g A N_A_c_136_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_12%A
x_PM_SKY130_FD_SC_HDLL__CLKBUF_12%A_117_297# N_A_117_297#_M1009_s
+ N_A_117_297#_M1028_s N_A_117_297#_M1002_s N_A_117_297#_M1019_s
+ N_A_117_297#_c_224_n N_A_117_297#_M1000_g N_A_117_297#_M1001_g
+ N_A_117_297#_M1006_g N_A_117_297#_c_225_n N_A_117_297#_M1003_g
+ N_A_117_297#_c_226_n N_A_117_297#_M1004_g N_A_117_297#_M1010_g
+ N_A_117_297#_M1011_g N_A_117_297#_c_227_n N_A_117_297#_M1005_g
+ N_A_117_297#_c_228_n N_A_117_297#_M1007_g N_A_117_297#_M1012_g
+ N_A_117_297#_M1014_g N_A_117_297#_c_229_n N_A_117_297#_M1008_g
+ N_A_117_297#_c_230_n N_A_117_297#_M1015_g N_A_117_297#_M1017_g
+ N_A_117_297#_M1018_g N_A_117_297#_c_231_n N_A_117_297#_M1016_g
+ N_A_117_297#_c_232_n N_A_117_297#_M1021_g N_A_117_297#_M1020_g
+ N_A_117_297#_M1024_g N_A_117_297#_c_233_n N_A_117_297#_M1023_g
+ N_A_117_297#_c_234_n N_A_117_297#_M1026_g N_A_117_297#_M1025_g
+ N_A_117_297#_M1030_g N_A_117_297#_c_235_n N_A_117_297#_M1029_g
+ N_A_117_297#_c_236_n N_A_117_297#_c_247_n N_A_117_297#_c_219_n
+ N_A_117_297#_c_220_n N_A_117_297#_c_256_n N_A_117_297#_c_237_n
+ N_A_117_297#_c_221_n N_A_117_297#_c_266_n N_A_117_297#_c_238_n
+ N_A_117_297#_c_319_p N_A_117_297#_c_222_n N_A_117_297#_c_271_n
+ N_A_117_297#_c_274_n N_A_117_297#_c_281_p N_A_117_297#_c_223_n
+ PM_SKY130_FD_SC_HDLL__CLKBUF_12%A_117_297#
x_PM_SKY130_FD_SC_HDLL__CLKBUF_12%VPWR N_VPWR_M1002_d N_VPWR_M1013_d
+ N_VPWR_M1027_d N_VPWR_M1003_d N_VPWR_M1005_d N_VPWR_M1008_d N_VPWR_M1016_d
+ N_VPWR_M1023_d N_VPWR_M1029_d N_VPWR_c_479_n N_VPWR_c_480_n N_VPWR_c_481_n
+ N_VPWR_c_482_n N_VPWR_c_483_n N_VPWR_c_484_n N_VPWR_c_485_n N_VPWR_c_486_n
+ N_VPWR_c_487_n N_VPWR_c_488_n N_VPWR_c_489_n N_VPWR_c_490_n N_VPWR_c_491_n
+ N_VPWR_c_492_n N_VPWR_c_493_n N_VPWR_c_494_n N_VPWR_c_495_n N_VPWR_c_496_n
+ VPWR N_VPWR_c_497_n N_VPWR_c_498_n N_VPWR_c_499_n N_VPWR_c_478_n
+ N_VPWR_c_501_n N_VPWR_c_502_n N_VPWR_c_503_n N_VPWR_c_504_n N_VPWR_c_505_n
+ N_VPWR_c_506_n PM_SKY130_FD_SC_HDLL__CLKBUF_12%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKBUF_12%X N_X_M1001_d N_X_M1010_d N_X_M1012_d
+ N_X_M1017_d N_X_M1020_d N_X_M1025_d N_X_M1000_s N_X_M1004_s N_X_M1007_s
+ N_X_M1015_s N_X_M1021_s N_X_M1026_s N_X_c_630_n N_X_c_645_n N_X_c_612_n
+ N_X_c_613_n N_X_c_614_n N_X_c_631_n N_X_c_615_n N_X_c_748_n N_X_c_616_n
+ N_X_c_632_n N_X_c_617_n N_X_c_752_n N_X_c_618_n N_X_c_633_n N_X_c_619_n
+ N_X_c_756_n N_X_c_620_n N_X_c_634_n N_X_c_621_n N_X_c_760_n N_X_c_622_n
+ N_X_c_635_n N_X_c_623_n N_X_c_764_n N_X_c_624_n N_X_c_636_n N_X_c_625_n
+ N_X_c_637_n N_X_c_626_n N_X_c_638_n N_X_c_627_n N_X_c_639_n N_X_c_628_n
+ N_X_c_728_n X PM_SKY130_FD_SC_HDLL__CLKBUF_12%X
x_PM_SKY130_FD_SC_HDLL__CLKBUF_12%VGND N_VGND_M1009_d N_VGND_M1022_d
+ N_VGND_M1031_d N_VGND_M1006_s N_VGND_M1011_s N_VGND_M1014_s N_VGND_M1018_s
+ N_VGND_M1024_s N_VGND_M1030_s N_VGND_c_809_n N_VGND_c_810_n N_VGND_c_811_n
+ N_VGND_c_812_n N_VGND_c_813_n N_VGND_c_814_n N_VGND_c_815_n N_VGND_c_816_n
+ N_VGND_c_817_n N_VGND_c_818_n N_VGND_c_819_n N_VGND_c_820_n N_VGND_c_821_n
+ N_VGND_c_822_n N_VGND_c_823_n N_VGND_c_824_n N_VGND_c_825_n N_VGND_c_826_n
+ VGND N_VGND_c_827_n N_VGND_c_828_n N_VGND_c_829_n N_VGND_c_830_n
+ N_VGND_c_831_n N_VGND_c_832_n N_VGND_c_833_n N_VGND_c_834_n N_VGND_c_835_n
+ N_VGND_c_836_n PM_SKY130_FD_SC_HDLL__CLKBUF_12%VGND
cc_1 VNB N_A_M1009_g 0.0319831f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.445
cc_2 VNB N_A_M1022_g 0.0225773f $X=-0.19 $Y=-0.24 $X2=0.94 $Y2=0.445
cc_3 VNB N_A_M1028_g 0.0225773f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.445
cc_4 VNB N_A_M1031_g 0.0237781f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.445
cc_5 VNB N_A_c_136_n 0.112639f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.155
cc_6 VNB N_A_117_297#_M1001_g 0.0264336f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.9
cc_7 VNB N_A_117_297#_M1006_g 0.025215f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=0.9
cc_8 VNB N_A_117_297#_M1010_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.155
cc_9 VNB N_A_117_297#_M1011_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=1.155 $Y2=1.16
cc_10 VNB N_A_117_297#_M1012_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_M1014_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_117_297#_M1017_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_117_297#_M1018_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_117_297#_M1020_g 0.0252407f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_117_297#_M1024_g 0.0252085f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_117_297#_M1025_g 0.0248481f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_117_297#_M1030_g 0.0359475f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_117_297#_c_219_n 0.00124412f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_117_297#_c_220_n 0.00334909f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_117_297#_c_221_n 0.00124486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_117_297#_c_222_n 0.00653071f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_117_297#_c_223_n 0.266585f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_478_n 0.345644f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_612_n 0.00124486f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_X_c_613_n 0.00617255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_X_c_614_n 0.00280924f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_X_c_615_n 9.92465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_616_n 0.00617255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_617_n 9.92465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_X_c_618_n 0.00617255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_X_c_619_n 9.92465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_X_c_620_n 0.00617255f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_X_c_621_n 9.92465e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_X_c_622_n 0.00563362f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_X_c_623_n 0.00124194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_X_c_624_n 0.00220003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_X_c_625_n 0.00220003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_X_c_626_n 0.00220003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_X_c_627_n 0.00220003f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_X_c_628_n 8.55634e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB X 9.87143e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_809_n 0.0115537f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_43 VNB N_VGND_c_810_n 0.0210194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_811_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.155
cc_45 VNB N_VGND_c_812_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.155
cc_46 VNB N_VGND_c_813_n 0.0162809f $X=-0.19 $Y=-0.24 $X2=1.88 $Y2=1.155
cc_47 VNB N_VGND_c_814_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_815_n 0.0156408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_816_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_817_n 0.0156408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_VGND_c_818_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_VGND_c_819_n 0.0156408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_VGND_c_820_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_VGND_c_821_n 0.00442069f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_VGND_c_822_n 0.0210194f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_VGND_c_823_n 0.0156408f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VGND_c_824_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_VGND_c_825_n 0.0162797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_VGND_c_826_n 0.00632231f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_VGND_c_827_n 0.0162809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_VGND_c_828_n 0.0162809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_VGND_c_829_n 0.0128037f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_VGND_c_830_n 0.399295f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_VGND_c_831_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_VGND_c_832_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_VGND_c_833_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_VGND_c_834_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_VGND_c_835_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_VGND_c_836_n 0.006319f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VPB N_A_c_137_n 0.0210307f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_71 VPB N_A_c_138_n 0.0161166f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_72 VPB N_A_c_139_n 0.0161015f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_73 VPB N_A_c_140_n 0.0161299f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_74 VPB N_A_c_136_n 0.05028f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.155
cc_75 VPB N_A_117_297#_c_224_n 0.01638f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.985
cc_76 VPB N_A_117_297#_c_225_n 0.0159704f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=0.445
cc_77 VPB N_A_117_297#_c_226_n 0.0159704f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_78 VPB N_A_117_297#_c_227_n 0.0159704f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.155
cc_79 VPB N_A_117_297#_c_228_n 0.0159704f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.155
cc_80 VPB N_A_117_297#_c_229_n 0.0159704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_A_117_297#_c_230_n 0.0159704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_A_117_297#_c_231_n 0.0159704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_A_117_297#_c_232_n 0.0159704f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_A_117_297#_c_233_n 0.0159413f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_A_117_297#_c_234_n 0.0153999f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_A_117_297#_c_235_n 0.0198008f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_A_117_297#_c_236_n 0.00176214f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_A_117_297#_c_237_n 0.0018532f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_A_117_297#_c_238_n 0.00284451f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_A_117_297#_c_223_n 0.153289f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_91 VPB N_VPWR_c_479_n 0.0109725f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.985
cc_92 VPB N_VPWR_c_480_n 0.0442531f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_93 VPB N_VPWR_c_481_n 0.0041482f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_94 VPB N_VPWR_c_482_n 0.00464704f $X=-0.19 $Y=1.305 $X2=1.88 $Y2=1.155
cc_95 VPB N_VPWR_c_483_n 0.0163297f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB N_VPWR_c_484_n 3.40287e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB N_VPWR_c_485_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 VPB N_VPWR_c_486_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_99 VPB N_VPWR_c_487_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_100 VPB N_VPWR_c_488_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_101 VPB N_VPWR_c_489_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_102 VPB N_VPWR_c_490_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_103 VPB N_VPWR_c_491_n 3.35805e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_104 VPB N_VPWR_c_492_n 0.0545118f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_105 VPB N_VPWR_c_493_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_106 VPB N_VPWR_c_494_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_107 VPB N_VPWR_c_495_n 0.0147329f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_108 VPB N_VPWR_c_496_n 0.00513801f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_109 VPB N_VPWR_c_497_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_110 VPB N_VPWR_c_498_n 0.0167344f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_111 VPB N_VPWR_c_499_n 0.0128037f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_112 VPB N_VPWR_c_478_n 0.0536543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_113 VPB N_VPWR_c_501_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_114 VPB N_VPWR_c_502_n 0.00455763f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_115 VPB N_VPWR_c_503_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_116 VPB N_VPWR_c_504_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_117 VPB N_VPWR_c_505_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_118 VPB N_VPWR_c_506_n 0.00436868f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_119 VPB N_X_c_630_n 0.00170286f $X=-0.19 $Y=1.305 $X2=1.155 $Y2=1.16
cc_120 VPB N_X_c_631_n 0.00183209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_X_c_632_n 0.00183209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_X_c_633_n 0.00183209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_X_c_634_n 0.00183209f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_X_c_635_n 0.0022065f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_X_c_636_n 0.00164358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_X_c_637_n 0.00164358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_X_c_638_n 0.00164358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_X_c_639_n 0.00164358f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB X 0.00323163f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 N_A_c_140_n N_A_117_297#_c_224_n 0.00928797f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_M1031_g N_A_117_297#_M1001_g 0.012839f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_132 N_A_c_136_n N_A_117_297#_M1001_g 0.00227284f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_133 N_A_c_137_n N_A_117_297#_c_236_n 0.00322357f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_c_138_n N_A_117_297#_c_236_n 7.41548e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_135 A N_A_117_297#_c_236_n 0.0269456f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_c_136_n N_A_117_297#_c_236_n 0.00789737f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_137 N_A_c_137_n N_A_117_297#_c_247_n 0.00897418f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_138 N_A_c_138_n N_A_117_297#_c_247_n 0.0100971f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_139_n N_A_117_297#_c_247_n 5.97234e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_M1009_g N_A_117_297#_c_219_n 0.00169095f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_141 N_A_M1022_g N_A_117_297#_c_219_n 9.75885e-19 $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_142 N_A_M1022_g N_A_117_297#_c_220_n 0.00902836f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_143 N_A_M1028_g N_A_117_297#_c_220_n 0.00902836f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_144 A N_A_117_297#_c_220_n 0.0318053f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_145 N_A_c_136_n N_A_117_297#_c_220_n 0.0154003f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_146 N_A_M1009_g N_A_117_297#_c_256_n 0.00620653f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_147 N_A_M1022_g N_A_117_297#_c_256_n 0.00206962f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_148 A N_A_117_297#_c_256_n 0.0208607f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_149 N_A_c_136_n N_A_117_297#_c_256_n 0.00633209f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_150 N_A_c_138_n N_A_117_297#_c_237_n 0.014439f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_151 N_A_c_139_n N_A_117_297#_c_237_n 0.0182506f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_152 A N_A_117_297#_c_237_n 0.0307126f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_153 N_A_c_136_n N_A_117_297#_c_237_n 0.00782413f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_154 N_A_M1028_g N_A_117_297#_c_221_n 9.75885e-19 $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_155 N_A_M1031_g N_A_117_297#_c_221_n 9.75885e-19 $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_156 N_A_c_136_n N_A_117_297#_c_266_n 0.0149752f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_157 N_A_c_139_n N_A_117_297#_c_238_n 0.00178892f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_158 N_A_c_140_n N_A_117_297#_c_238_n 0.00178892f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_159 N_A_c_136_n N_A_117_297#_c_238_n 0.0131756f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_160 N_A_c_136_n N_A_117_297#_c_222_n 0.0231863f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_161 N_A_M1028_g N_A_117_297#_c_271_n 0.00206962f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_162 N_A_M1031_g N_A_117_297#_c_271_n 0.00335799f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_163 N_A_c_136_n N_A_117_297#_c_271_n 0.00232955f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_164 A N_A_117_297#_c_274_n 0.0159631f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_165 N_A_c_136_n N_A_117_297#_c_274_n 0.00958118f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_166 N_A_c_136_n N_A_117_297#_c_223_n 0.0241539f $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_167 N_A_c_137_n N_VPWR_c_480_n 0.00356412f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_168 N_A_c_138_n N_VPWR_c_481_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_c_139_n N_VPWR_c_481_n 0.00170062f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_c_139_n N_VPWR_c_482_n 6.96617e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_171 N_A_c_140_n N_VPWR_c_482_n 0.0147456f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_172 N_A_c_136_n N_VPWR_c_482_n 2.88532e-19 $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_173 N_A_c_137_n N_VPWR_c_497_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_c_138_n N_VPWR_c_497_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_175 N_A_c_139_n N_VPWR_c_498_n 0.00702461f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_176 N_A_c_140_n N_VPWR_c_498_n 0.00622633f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_c_137_n N_VPWR_c_478_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_c_138_n N_VPWR_c_478_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_179 N_A_c_139_n N_VPWR_c_478_n 0.0123841f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_180 N_A_c_140_n N_VPWR_c_478_n 0.0104011f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_181 N_A_M1031_g N_X_c_614_n 5.50882e-19 $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_182 N_A_M1009_g N_VGND_c_810_n 0.00366311f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_183 N_A_M1022_g N_VGND_c_811_n 0.00183908f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_184 N_A_M1028_g N_VGND_c_811_n 0.00183908f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_185 N_A_c_136_n N_VGND_c_811_n 9.63051e-19 $X=1.88 $Y=1.155 $X2=0 $Y2=0
cc_186 N_A_M1031_g N_VGND_c_812_n 0.00183908f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_187 N_A_M1009_g N_VGND_c_827_n 0.00585385f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A_M1022_g N_VGND_c_827_n 0.00436487f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A_M1028_g N_VGND_c_828_n 0.00436487f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A_M1031_g N_VGND_c_828_n 0.00585385f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_191 N_A_M1009_g N_VGND_c_830_n 0.0116506f $X=0.52 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A_M1022_g N_VGND_c_830_n 0.00612685f $X=0.94 $Y=0.445 $X2=0 $Y2=0
cc_193 N_A_M1028_g N_VGND_c_830_n 0.00612685f $X=1.46 $Y=0.445 $X2=0 $Y2=0
cc_194 N_A_M1031_g N_VGND_c_830_n 0.0108765f $X=1.88 $Y=0.445 $X2=0 $Y2=0
cc_195 N_A_117_297#_c_237_n N_VPWR_M1013_d 0.00187735f $X=1.535 $Y=1.57 $X2=0
+ $Y2=0
cc_196 N_A_117_297#_c_237_n N_VPWR_c_481_n 0.0144271f $X=1.535 $Y=1.57 $X2=0
+ $Y2=0
cc_197 N_A_117_297#_c_224_n N_VPWR_c_482_n 0.0017965f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A_117_297#_c_222_n N_VPWR_c_482_n 0.0254987f $X=6.52 $Y=1.16 $X2=0
+ $Y2=0
cc_199 N_A_117_297#_c_281_p N_VPWR_c_482_n 0.00747887f $X=1.67 $Y=1.62 $X2=0
+ $Y2=0
cc_200 N_A_117_297#_c_224_n N_VPWR_c_483_n 0.00673617f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_201 N_A_117_297#_c_225_n N_VPWR_c_483_n 0.00622633f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A_117_297#_c_224_n N_VPWR_c_484_n 4.46241e-19 $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_203 N_A_117_297#_c_225_n N_VPWR_c_484_n 0.0111329f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_204 N_A_117_297#_c_226_n N_VPWR_c_484_n 0.0110732f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_205 N_A_117_297#_c_227_n N_VPWR_c_484_n 5.94261e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_206 N_A_117_297#_c_226_n N_VPWR_c_485_n 0.00622633f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_207 N_A_117_297#_c_227_n N_VPWR_c_485_n 0.00622633f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_208 N_A_117_297#_c_226_n N_VPWR_c_486_n 5.94261e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_209 N_A_117_297#_c_227_n N_VPWR_c_486_n 0.0110732f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_210 N_A_117_297#_c_228_n N_VPWR_c_486_n 0.0110732f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_211 N_A_117_297#_c_229_n N_VPWR_c_486_n 5.94261e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A_117_297#_c_228_n N_VPWR_c_487_n 0.00622633f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_213 N_A_117_297#_c_229_n N_VPWR_c_487_n 0.00622633f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_214 N_A_117_297#_c_228_n N_VPWR_c_488_n 5.94261e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_215 N_A_117_297#_c_229_n N_VPWR_c_488_n 0.0110732f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_216 N_A_117_297#_c_230_n N_VPWR_c_488_n 0.0110732f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_217 N_A_117_297#_c_231_n N_VPWR_c_488_n 5.94261e-19 $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_218 N_A_117_297#_c_230_n N_VPWR_c_489_n 0.00622633f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_219 N_A_117_297#_c_231_n N_VPWR_c_489_n 0.00622633f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_220 N_A_117_297#_c_230_n N_VPWR_c_490_n 5.94261e-19 $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_221 N_A_117_297#_c_231_n N_VPWR_c_490_n 0.0110732f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_222 N_A_117_297#_c_232_n N_VPWR_c_490_n 0.0110732f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_223 N_A_117_297#_c_233_n N_VPWR_c_490_n 5.94261e-19 $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_224 N_A_117_297#_c_232_n N_VPWR_c_491_n 5.94261e-19 $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_225 N_A_117_297#_c_233_n N_VPWR_c_491_n 0.0110732f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_226 N_A_117_297#_c_234_n N_VPWR_c_491_n 0.0110724f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_227 N_A_117_297#_c_235_n N_VPWR_c_491_n 5.94261e-19 $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_228 N_A_117_297#_c_223_n N_VPWR_c_491_n 3.03461e-19 $X=7.52 $Y=1.18 $X2=0
+ $Y2=0
cc_229 N_A_117_297#_c_234_n N_VPWR_c_492_n 6.96996e-19 $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_230 N_A_117_297#_c_235_n N_VPWR_c_492_n 0.0170427f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_231 N_A_117_297#_c_223_n N_VPWR_c_492_n 5.21878e-19 $X=7.52 $Y=1.18 $X2=0
+ $Y2=0
cc_232 N_A_117_297#_c_232_n N_VPWR_c_493_n 0.00622633f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_233 N_A_117_297#_c_233_n N_VPWR_c_493_n 0.00622633f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_234 N_A_117_297#_c_234_n N_VPWR_c_495_n 0.00622633f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_235 N_A_117_297#_c_235_n N_VPWR_c_495_n 0.00622633f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_236 N_A_117_297#_c_247_n N_VPWR_c_497_n 0.0189467f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_237 N_A_117_297#_c_319_p N_VPWR_c_498_n 0.0156407f $X=1.67 $Y=2.3 $X2=0 $Y2=0
cc_238 N_A_117_297#_M1002_s N_VPWR_c_478_n 0.00231261f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_239 N_A_117_297#_M1019_s N_VPWR_c_478_n 0.00300692f $X=1.525 $Y=1.485 $X2=0
+ $Y2=0
cc_240 N_A_117_297#_c_224_n N_VPWR_c_478_n 0.0117436f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_241 N_A_117_297#_c_225_n N_VPWR_c_478_n 0.0104011f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_242 N_A_117_297#_c_226_n N_VPWR_c_478_n 0.0104011f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_243 N_A_117_297#_c_227_n N_VPWR_c_478_n 0.0104011f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_244 N_A_117_297#_c_228_n N_VPWR_c_478_n 0.0104011f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_245 N_A_117_297#_c_229_n N_VPWR_c_478_n 0.0104011f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_246 N_A_117_297#_c_230_n N_VPWR_c_478_n 0.0104011f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_247 N_A_117_297#_c_231_n N_VPWR_c_478_n 0.0104011f $X=5.665 $Y=1.41 $X2=0
+ $Y2=0
cc_248 N_A_117_297#_c_232_n N_VPWR_c_478_n 0.0104011f $X=6.135 $Y=1.41 $X2=0
+ $Y2=0
cc_249 N_A_117_297#_c_233_n N_VPWR_c_478_n 0.0104011f $X=6.605 $Y=1.41 $X2=0
+ $Y2=0
cc_250 N_A_117_297#_c_234_n N_VPWR_c_478_n 0.0104011f $X=7.075 $Y=1.41 $X2=0
+ $Y2=0
cc_251 N_A_117_297#_c_235_n N_VPWR_c_478_n 0.0104011f $X=7.545 $Y=1.41 $X2=0
+ $Y2=0
cc_252 N_A_117_297#_c_247_n N_VPWR_c_478_n 0.0123132f $X=0.73 $Y=2.3 $X2=0 $Y2=0
cc_253 N_A_117_297#_c_319_p N_VPWR_c_478_n 0.0103212f $X=1.67 $Y=2.3 $X2=0 $Y2=0
cc_254 N_A_117_297#_c_224_n N_X_c_630_n 0.002409f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_255 N_A_117_297#_c_222_n N_X_c_630_n 0.0246001f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_256 N_A_117_297#_c_223_n N_X_c_630_n 0.00753278f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_257 N_A_117_297#_c_224_n N_X_c_645_n 0.00855819f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_258 N_A_117_297#_M1001_g N_X_c_612_n 9.75885e-19 $X=2.4 $Y=0.445 $X2=0 $Y2=0
cc_259 N_A_117_297#_M1006_g N_X_c_612_n 9.75885e-19 $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_260 N_A_117_297#_c_221_n N_X_c_612_n 0.00463621f $X=1.67 $Y=0.445 $X2=0 $Y2=0
cc_261 N_A_117_297#_M1006_g N_X_c_613_n 0.0112224f $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_262 N_A_117_297#_M1010_g N_X_c_613_n 0.0112224f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_263 N_A_117_297#_c_222_n N_X_c_613_n 0.0482232f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_264 N_A_117_297#_c_223_n N_X_c_613_n 0.0050885f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_265 N_A_117_297#_M1001_g N_X_c_614_n 0.00346749f $X=2.4 $Y=0.445 $X2=0 $Y2=0
cc_266 N_A_117_297#_M1006_g N_X_c_614_n 0.00212617f $X=2.82 $Y=0.445 $X2=0 $Y2=0
cc_267 N_A_117_297#_c_222_n N_X_c_614_n 0.0220669f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_268 N_A_117_297#_c_271_n N_X_c_614_n 0.00506064f $X=1.67 $Y=0.81 $X2=0 $Y2=0
cc_269 N_A_117_297#_c_223_n N_X_c_614_n 0.00249422f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_270 N_A_117_297#_c_225_n N_X_c_631_n 0.0154866f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_271 N_A_117_297#_c_226_n N_X_c_631_n 0.0154866f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_272 N_A_117_297#_c_222_n N_X_c_631_n 0.0479857f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_117_297#_c_223_n N_X_c_631_n 0.00784151f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_274 N_A_117_297#_M1010_g N_X_c_615_n 9.75885e-19 $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_275 N_A_117_297#_M1011_g N_X_c_615_n 9.75885e-19 $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_276 N_A_117_297#_M1011_g N_X_c_616_n 0.0112224f $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_277 N_A_117_297#_M1012_g N_X_c_616_n 0.0112224f $X=4.28 $Y=0.445 $X2=0 $Y2=0
cc_278 N_A_117_297#_c_222_n N_X_c_616_n 0.0482232f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_279 N_A_117_297#_c_223_n N_X_c_616_n 0.0050885f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_280 N_A_117_297#_c_227_n N_X_c_632_n 0.0154866f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_281 N_A_117_297#_c_228_n N_X_c_632_n 0.0154866f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_282 N_A_117_297#_c_222_n N_X_c_632_n 0.0479857f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_283 N_A_117_297#_c_223_n N_X_c_632_n 0.00784151f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_284 N_A_117_297#_M1012_g N_X_c_617_n 9.75885e-19 $X=4.28 $Y=0.445 $X2=0 $Y2=0
cc_285 N_A_117_297#_M1014_g N_X_c_617_n 9.75885e-19 $X=4.7 $Y=0.445 $X2=0 $Y2=0
cc_286 N_A_117_297#_M1014_g N_X_c_618_n 0.0112224f $X=4.7 $Y=0.445 $X2=0 $Y2=0
cc_287 N_A_117_297#_M1017_g N_X_c_618_n 0.0112224f $X=5.22 $Y=0.445 $X2=0 $Y2=0
cc_288 N_A_117_297#_c_222_n N_X_c_618_n 0.0482232f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_289 N_A_117_297#_c_223_n N_X_c_618_n 0.0050885f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_290 N_A_117_297#_c_229_n N_X_c_633_n 0.0154866f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_291 N_A_117_297#_c_230_n N_X_c_633_n 0.0154866f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_292 N_A_117_297#_c_222_n N_X_c_633_n 0.0479857f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_293 N_A_117_297#_c_223_n N_X_c_633_n 0.00784151f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_294 N_A_117_297#_M1017_g N_X_c_619_n 9.75885e-19 $X=5.22 $Y=0.445 $X2=0 $Y2=0
cc_295 N_A_117_297#_M1018_g N_X_c_619_n 9.75885e-19 $X=5.64 $Y=0.445 $X2=0 $Y2=0
cc_296 N_A_117_297#_M1018_g N_X_c_620_n 0.0112224f $X=5.64 $Y=0.445 $X2=0 $Y2=0
cc_297 N_A_117_297#_M1020_g N_X_c_620_n 0.0112224f $X=6.16 $Y=0.445 $X2=0 $Y2=0
cc_298 N_A_117_297#_c_222_n N_X_c_620_n 0.0482232f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_299 N_A_117_297#_c_223_n N_X_c_620_n 0.0050885f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_300 N_A_117_297#_c_231_n N_X_c_634_n 0.0154866f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_301 N_A_117_297#_c_232_n N_X_c_634_n 0.0154866f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_302 N_A_117_297#_c_222_n N_X_c_634_n 0.0479857f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_303 N_A_117_297#_c_223_n N_X_c_634_n 0.00784151f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_304 N_A_117_297#_M1020_g N_X_c_621_n 9.75885e-19 $X=6.16 $Y=0.445 $X2=0 $Y2=0
cc_305 N_A_117_297#_M1024_g N_X_c_621_n 9.75885e-19 $X=6.58 $Y=0.445 $X2=0 $Y2=0
cc_306 N_A_117_297#_M1024_g N_X_c_622_n 0.0112224f $X=6.58 $Y=0.445 $X2=0 $Y2=0
cc_307 N_A_117_297#_c_222_n N_X_c_622_n 0.012676f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_308 N_A_117_297#_c_223_n N_X_c_622_n 0.00608873f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_309 N_A_117_297#_c_233_n N_X_c_635_n 0.0156082f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_310 N_A_117_297#_c_222_n N_X_c_635_n 0.0125956f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_311 N_A_117_297#_c_223_n N_X_c_635_n 0.00799345f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_312 N_A_117_297#_M1025_g N_X_c_623_n 9.75885e-19 $X=7.1 $Y=0.445 $X2=0 $Y2=0
cc_313 N_A_117_297#_M1030_g N_X_c_623_n 0.00169095f $X=7.52 $Y=0.445 $X2=0 $Y2=0
cc_314 N_A_117_297#_M1010_g N_X_c_624_n 0.00219873f $X=3.34 $Y=0.445 $X2=0 $Y2=0
cc_315 N_A_117_297#_M1011_g N_X_c_624_n 0.00219873f $X=3.76 $Y=0.445 $X2=0 $Y2=0
cc_316 N_A_117_297#_c_222_n N_X_c_624_n 0.0220669f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_317 N_A_117_297#_c_223_n N_X_c_624_n 0.00249422f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_318 N_A_117_297#_c_222_n N_X_c_636_n 0.0222213f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_319 N_A_117_297#_c_223_n N_X_c_636_n 0.00722373f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_320 N_A_117_297#_M1012_g N_X_c_625_n 0.00219873f $X=4.28 $Y=0.445 $X2=0 $Y2=0
cc_321 N_A_117_297#_M1014_g N_X_c_625_n 0.00219873f $X=4.7 $Y=0.445 $X2=0 $Y2=0
cc_322 N_A_117_297#_c_222_n N_X_c_625_n 0.0220669f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_323 N_A_117_297#_c_223_n N_X_c_625_n 0.00249422f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_324 N_A_117_297#_c_222_n N_X_c_637_n 0.0222213f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_325 N_A_117_297#_c_223_n N_X_c_637_n 0.00722373f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_326 N_A_117_297#_M1017_g N_X_c_626_n 0.00219873f $X=5.22 $Y=0.445 $X2=0 $Y2=0
cc_327 N_A_117_297#_M1018_g N_X_c_626_n 0.00219873f $X=5.64 $Y=0.445 $X2=0 $Y2=0
cc_328 N_A_117_297#_c_222_n N_X_c_626_n 0.0220669f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_329 N_A_117_297#_c_223_n N_X_c_626_n 0.00249422f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_330 N_A_117_297#_c_222_n N_X_c_638_n 0.0222213f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_331 N_A_117_297#_c_223_n N_X_c_638_n 0.00722373f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_332 N_A_117_297#_M1020_g N_X_c_627_n 0.00219873f $X=6.16 $Y=0.445 $X2=0 $Y2=0
cc_333 N_A_117_297#_M1024_g N_X_c_627_n 0.00219873f $X=6.58 $Y=0.445 $X2=0 $Y2=0
cc_334 N_A_117_297#_c_222_n N_X_c_627_n 0.0220669f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_335 N_A_117_297#_c_223_n N_X_c_627_n 0.00249422f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_336 N_A_117_297#_c_222_n N_X_c_639_n 0.0222213f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_337 N_A_117_297#_c_223_n N_X_c_639_n 0.00722373f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_338 N_A_117_297#_M1025_g N_X_c_628_n 0.0114186f $X=7.1 $Y=0.445 $X2=0 $Y2=0
cc_339 N_A_117_297#_M1030_g N_X_c_628_n 0.00640891f $X=7.52 $Y=0.445 $X2=0 $Y2=0
cc_340 N_A_117_297#_c_234_n N_X_c_728_n 0.0142154f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_341 N_A_117_297#_M1024_g X 9.86344e-19 $X=6.58 $Y=0.445 $X2=0 $Y2=0
cc_342 N_A_117_297#_c_233_n X 0.00146713f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_343 N_A_117_297#_c_234_n X 0.00196284f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_344 N_A_117_297#_M1025_g X 0.00132071f $X=7.1 $Y=0.445 $X2=0 $Y2=0
cc_345 N_A_117_297#_M1030_g X 0.00137081f $X=7.52 $Y=0.445 $X2=0 $Y2=0
cc_346 N_A_117_297#_c_235_n X 0.00179891f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_347 N_A_117_297#_c_222_n X 0.0127244f $X=6.52 $Y=1.16 $X2=0 $Y2=0
cc_348 N_A_117_297#_c_223_n X 0.0619784f $X=7.52 $Y=1.18 $X2=0 $Y2=0
cc_349 N_A_117_297#_c_220_n N_VGND_c_811_n 0.0230107f $X=1.535 $Y=0.81 $X2=0
+ $Y2=0
cc_350 N_A_117_297#_M1001_g N_VGND_c_812_n 0.00183908f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_351 N_A_117_297#_c_222_n N_VGND_c_812_n 0.0105308f $X=6.52 $Y=1.16 $X2=0
+ $Y2=0
cc_352 N_A_117_297#_M1001_g N_VGND_c_813_n 0.00585385f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_353 N_A_117_297#_M1006_g N_VGND_c_813_n 0.00436487f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_354 N_A_117_297#_M1006_g N_VGND_c_814_n 0.00183908f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_355 N_A_117_297#_M1010_g N_VGND_c_814_n 0.00183908f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_356 N_A_117_297#_M1010_g N_VGND_c_815_n 0.00436487f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_357 N_A_117_297#_M1011_g N_VGND_c_815_n 0.00436487f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_358 N_A_117_297#_M1011_g N_VGND_c_816_n 0.00183908f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_359 N_A_117_297#_M1012_g N_VGND_c_816_n 0.00183908f $X=4.28 $Y=0.445 $X2=0
+ $Y2=0
cc_360 N_A_117_297#_M1012_g N_VGND_c_817_n 0.00436487f $X=4.28 $Y=0.445 $X2=0
+ $Y2=0
cc_361 N_A_117_297#_M1014_g N_VGND_c_817_n 0.00436487f $X=4.7 $Y=0.445 $X2=0
+ $Y2=0
cc_362 N_A_117_297#_M1014_g N_VGND_c_818_n 0.00183908f $X=4.7 $Y=0.445 $X2=0
+ $Y2=0
cc_363 N_A_117_297#_M1017_g N_VGND_c_818_n 0.00183908f $X=5.22 $Y=0.445 $X2=0
+ $Y2=0
cc_364 N_A_117_297#_M1017_g N_VGND_c_819_n 0.00436487f $X=5.22 $Y=0.445 $X2=0
+ $Y2=0
cc_365 N_A_117_297#_M1018_g N_VGND_c_819_n 0.00436487f $X=5.64 $Y=0.445 $X2=0
+ $Y2=0
cc_366 N_A_117_297#_M1018_g N_VGND_c_820_n 0.00183908f $X=5.64 $Y=0.445 $X2=0
+ $Y2=0
cc_367 N_A_117_297#_M1020_g N_VGND_c_820_n 0.00183908f $X=6.16 $Y=0.445 $X2=0
+ $Y2=0
cc_368 N_A_117_297#_M1024_g N_VGND_c_821_n 0.00183908f $X=6.58 $Y=0.445 $X2=0
+ $Y2=0
cc_369 N_A_117_297#_M1025_g N_VGND_c_821_n 0.00183908f $X=7.1 $Y=0.445 $X2=0
+ $Y2=0
cc_370 N_A_117_297#_M1030_g N_VGND_c_822_n 0.00366311f $X=7.52 $Y=0.445 $X2=0
+ $Y2=0
cc_371 N_A_117_297#_M1020_g N_VGND_c_823_n 0.00436487f $X=6.16 $Y=0.445 $X2=0
+ $Y2=0
cc_372 N_A_117_297#_M1024_g N_VGND_c_823_n 0.00436487f $X=6.58 $Y=0.445 $X2=0
+ $Y2=0
cc_373 N_A_117_297#_M1025_g N_VGND_c_825_n 0.00436349f $X=7.1 $Y=0.445 $X2=0
+ $Y2=0
cc_374 N_A_117_297#_M1030_g N_VGND_c_825_n 0.00585385f $X=7.52 $Y=0.445 $X2=0
+ $Y2=0
cc_375 N_A_117_297#_c_219_n N_VGND_c_827_n 0.0128585f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_376 N_A_117_297#_c_220_n N_VGND_c_827_n 0.00236641f $X=1.535 $Y=0.81 $X2=0
+ $Y2=0
cc_377 N_A_117_297#_c_220_n N_VGND_c_828_n 0.00236641f $X=1.535 $Y=0.81 $X2=0
+ $Y2=0
cc_378 N_A_117_297#_c_221_n N_VGND_c_828_n 0.0129159f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_379 N_A_117_297#_M1009_s N_VGND_c_830_n 0.00216346f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_380 N_A_117_297#_M1028_s N_VGND_c_830_n 0.00216346f $X=1.535 $Y=0.235 $X2=0
+ $Y2=0
cc_381 N_A_117_297#_M1001_g N_VGND_c_830_n 0.0108765f $X=2.4 $Y=0.445 $X2=0
+ $Y2=0
cc_382 N_A_117_297#_M1006_g N_VGND_c_830_n 0.00612685f $X=2.82 $Y=0.445 $X2=0
+ $Y2=0
cc_383 N_A_117_297#_M1010_g N_VGND_c_830_n 0.00612685f $X=3.34 $Y=0.445 $X2=0
+ $Y2=0
cc_384 N_A_117_297#_M1011_g N_VGND_c_830_n 0.00612685f $X=3.76 $Y=0.445 $X2=0
+ $Y2=0
cc_385 N_A_117_297#_M1012_g N_VGND_c_830_n 0.00612685f $X=4.28 $Y=0.445 $X2=0
+ $Y2=0
cc_386 N_A_117_297#_M1014_g N_VGND_c_830_n 0.00612685f $X=4.7 $Y=0.445 $X2=0
+ $Y2=0
cc_387 N_A_117_297#_M1017_g N_VGND_c_830_n 0.00612685f $X=5.22 $Y=0.445 $X2=0
+ $Y2=0
cc_388 N_A_117_297#_M1018_g N_VGND_c_830_n 0.00612685f $X=5.64 $Y=0.445 $X2=0
+ $Y2=0
cc_389 N_A_117_297#_M1020_g N_VGND_c_830_n 0.00612685f $X=6.16 $Y=0.445 $X2=0
+ $Y2=0
cc_390 N_A_117_297#_M1024_g N_VGND_c_830_n 0.00612685f $X=6.58 $Y=0.445 $X2=0
+ $Y2=0
cc_391 N_A_117_297#_M1025_g N_VGND_c_830_n 0.00612437f $X=7.1 $Y=0.445 $X2=0
+ $Y2=0
cc_392 N_A_117_297#_M1030_g N_VGND_c_830_n 0.0117969f $X=7.52 $Y=0.445 $X2=0
+ $Y2=0
cc_393 N_A_117_297#_c_219_n N_VGND_c_830_n 0.0101718f $X=0.73 $Y=0.445 $X2=0
+ $Y2=0
cc_394 N_A_117_297#_c_220_n N_VGND_c_830_n 0.00886099f $X=1.535 $Y=0.81 $X2=0
+ $Y2=0
cc_395 N_A_117_297#_c_221_n N_VGND_c_830_n 0.0101963f $X=1.67 $Y=0.445 $X2=0
+ $Y2=0
cc_396 N_VPWR_c_478_n N_X_M1000_s 0.00265976f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_397 N_VPWR_c_478_n N_X_M1004_s 0.00300692f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_398 N_VPWR_c_478_n N_X_M1007_s 0.00300692f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_399 N_VPWR_c_478_n N_X_M1015_s 0.00300692f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_400 N_VPWR_c_478_n N_X_M1021_s 0.00300692f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_401 N_VPWR_c_478_n N_X_M1026_s 0.00300692f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_402 N_VPWR_c_482_n N_X_c_630_n 0.00837421f $X=2.14 $Y=1.64 $X2=0 $Y2=0
cc_403 N_VPWR_c_483_n N_X_c_645_n 0.0172937f $X=2.915 $Y=2.72 $X2=0 $Y2=0
cc_404 N_VPWR_c_478_n N_X_c_645_n 0.0113172f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_405 N_VPWR_M1003_d N_X_c_631_n 0.00187735f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_406 N_VPWR_c_484_n N_X_c_631_n 0.0172598f $X=3.08 $Y=1.96 $X2=0 $Y2=0
cc_407 N_VPWR_c_485_n N_X_c_748_n 0.0156407f $X=3.855 $Y=2.72 $X2=0 $Y2=0
cc_408 N_VPWR_c_478_n N_X_c_748_n 0.0103212f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_409 N_VPWR_M1005_d N_X_c_632_n 0.00187735f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_410 N_VPWR_c_486_n N_X_c_632_n 0.0172598f $X=4.02 $Y=1.96 $X2=0 $Y2=0
cc_411 N_VPWR_c_487_n N_X_c_752_n 0.0156407f $X=4.795 $Y=2.72 $X2=0 $Y2=0
cc_412 N_VPWR_c_478_n N_X_c_752_n 0.0103212f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_413 N_VPWR_M1008_d N_X_c_633_n 0.00187735f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_414 N_VPWR_c_488_n N_X_c_633_n 0.0172598f $X=4.96 $Y=1.96 $X2=0 $Y2=0
cc_415 N_VPWR_c_489_n N_X_c_756_n 0.0156407f $X=5.735 $Y=2.72 $X2=0 $Y2=0
cc_416 N_VPWR_c_478_n N_X_c_756_n 0.0103212f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_417 N_VPWR_M1016_d N_X_c_634_n 0.00187735f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_418 N_VPWR_c_490_n N_X_c_634_n 0.0172598f $X=5.9 $Y=1.96 $X2=0 $Y2=0
cc_419 N_VPWR_c_493_n N_X_c_760_n 0.0156407f $X=6.675 $Y=2.72 $X2=0 $Y2=0
cc_420 N_VPWR_c_478_n N_X_c_760_n 0.0103212f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_421 N_VPWR_M1023_d N_X_c_635_n 0.00187735f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_422 N_VPWR_c_491_n N_X_c_635_n 0.0158435f $X=6.84 $Y=1.96 $X2=0 $Y2=0
cc_423 N_VPWR_c_495_n N_X_c_764_n 0.0156407f $X=7.615 $Y=2.72 $X2=0 $Y2=0
cc_424 N_VPWR_c_478_n N_X_c_764_n 0.0103212f $X=8.05 $Y=2.72 $X2=0 $Y2=0
cc_425 N_VPWR_c_491_n N_X_c_728_n 0.00156604f $X=6.84 $Y=1.96 $X2=0 $Y2=0
cc_426 N_VPWR_c_492_n N_X_c_728_n 0.00758267f $X=7.78 $Y=1.63 $X2=0 $Y2=0
cc_427 N_VPWR_c_492_n X 7.72094e-19 $X=7.78 $Y=1.63 $X2=0 $Y2=0
cc_428 N_X_c_612_n N_VGND_c_813_n 0.0128585f $X=2.61 $Y=0.445 $X2=0 $Y2=0
cc_429 N_X_c_613_n N_VGND_c_813_n 0.00236641f $X=3.415 $Y=0.81 $X2=0 $Y2=0
cc_430 N_X_c_613_n N_VGND_c_814_n 0.0230108f $X=3.415 $Y=0.81 $X2=0 $Y2=0
cc_431 N_X_c_613_n N_VGND_c_815_n 0.00236641f $X=3.415 $Y=0.81 $X2=0 $Y2=0
cc_432 N_X_c_615_n N_VGND_c_815_n 0.0128585f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_433 N_X_c_616_n N_VGND_c_815_n 0.00236641f $X=4.355 $Y=0.81 $X2=0 $Y2=0
cc_434 N_X_c_616_n N_VGND_c_816_n 0.0230108f $X=4.355 $Y=0.81 $X2=0 $Y2=0
cc_435 N_X_c_616_n N_VGND_c_817_n 0.00236641f $X=4.355 $Y=0.81 $X2=0 $Y2=0
cc_436 N_X_c_617_n N_VGND_c_817_n 0.0128585f $X=4.49 $Y=0.445 $X2=0 $Y2=0
cc_437 N_X_c_618_n N_VGND_c_817_n 0.00236641f $X=5.295 $Y=0.81 $X2=0 $Y2=0
cc_438 N_X_c_618_n N_VGND_c_818_n 0.0230108f $X=5.295 $Y=0.81 $X2=0 $Y2=0
cc_439 N_X_c_618_n N_VGND_c_819_n 0.00236641f $X=5.295 $Y=0.81 $X2=0 $Y2=0
cc_440 N_X_c_619_n N_VGND_c_819_n 0.0128585f $X=5.43 $Y=0.445 $X2=0 $Y2=0
cc_441 N_X_c_620_n N_VGND_c_819_n 0.00236641f $X=6.235 $Y=0.81 $X2=0 $Y2=0
cc_442 N_X_c_620_n N_VGND_c_820_n 0.0230108f $X=6.235 $Y=0.81 $X2=0 $Y2=0
cc_443 N_X_c_622_n N_VGND_c_821_n 0.0210574f $X=6.96 $Y=0.81 $X2=0 $Y2=0
cc_444 N_X_c_628_n N_VGND_c_821_n 0.00226251f $X=7.202 $Y=0.81 $X2=0 $Y2=0
cc_445 N_X_c_620_n N_VGND_c_823_n 0.00236641f $X=6.235 $Y=0.81 $X2=0 $Y2=0
cc_446 N_X_c_621_n N_VGND_c_823_n 0.0128585f $X=6.37 $Y=0.445 $X2=0 $Y2=0
cc_447 N_X_c_622_n N_VGND_c_823_n 0.00236641f $X=6.96 $Y=0.81 $X2=0 $Y2=0
cc_448 N_X_c_623_n N_VGND_c_825_n 0.0129159f $X=7.31 $Y=0.445 $X2=0 $Y2=0
cc_449 N_X_c_628_n N_VGND_c_825_n 0.0025993f $X=7.202 $Y=0.81 $X2=0 $Y2=0
cc_450 N_X_M1001_d N_VGND_c_830_n 0.00216346f $X=2.475 $Y=0.235 $X2=0 $Y2=0
cc_451 N_X_M1010_d N_VGND_c_830_n 0.00216346f $X=3.415 $Y=0.235 $X2=0 $Y2=0
cc_452 N_X_M1012_d N_VGND_c_830_n 0.00216346f $X=4.355 $Y=0.235 $X2=0 $Y2=0
cc_453 N_X_M1017_d N_VGND_c_830_n 0.00216346f $X=5.295 $Y=0.235 $X2=0 $Y2=0
cc_454 N_X_M1020_d N_VGND_c_830_n 0.00216346f $X=6.235 $Y=0.235 $X2=0 $Y2=0
cc_455 N_X_M1025_d N_VGND_c_830_n 0.00216346f $X=7.175 $Y=0.235 $X2=0 $Y2=0
cc_456 N_X_c_612_n N_VGND_c_830_n 0.0101718f $X=2.61 $Y=0.445 $X2=0 $Y2=0
cc_457 N_X_c_613_n N_VGND_c_830_n 0.00886099f $X=3.415 $Y=0.81 $X2=0 $Y2=0
cc_458 N_X_c_615_n N_VGND_c_830_n 0.0101718f $X=3.55 $Y=0.445 $X2=0 $Y2=0
cc_459 N_X_c_616_n N_VGND_c_830_n 0.00886099f $X=4.355 $Y=0.81 $X2=0 $Y2=0
cc_460 N_X_c_617_n N_VGND_c_830_n 0.0101718f $X=4.49 $Y=0.445 $X2=0 $Y2=0
cc_461 N_X_c_618_n N_VGND_c_830_n 0.00886099f $X=5.295 $Y=0.81 $X2=0 $Y2=0
cc_462 N_X_c_619_n N_VGND_c_830_n 0.0101718f $X=5.43 $Y=0.445 $X2=0 $Y2=0
cc_463 N_X_c_620_n N_VGND_c_830_n 0.00886099f $X=6.235 $Y=0.81 $X2=0 $Y2=0
cc_464 N_X_c_621_n N_VGND_c_830_n 0.0101718f $X=6.37 $Y=0.445 $X2=0 $Y2=0
cc_465 N_X_c_622_n N_VGND_c_830_n 0.00489726f $X=6.96 $Y=0.81 $X2=0 $Y2=0
cc_466 N_X_c_623_n N_VGND_c_830_n 0.0101963f $X=7.31 $Y=0.445 $X2=0 $Y2=0
cc_467 N_X_c_628_n N_VGND_c_830_n 0.00424521f $X=7.202 $Y=0.81 $X2=0 $Y2=0
