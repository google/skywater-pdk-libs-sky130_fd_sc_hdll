* File: sky130_fd_sc_hdll__o221ai_1.spice
* Created: Wed Sep  2 08:44:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o221ai_1.pex.spice"
.subckt sky130_fd_sc_hdll__o221ai_1  VNB VPB C1 B1 B2 A2 A1 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* C1	C1
* VPB	VPB
* VNB	VNB
MM1004 N_A_123_47#_M1004_d N_C1_M1004_g N_Y_M1004_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.2145 PD=1.82 PS=1.96 NRD=0 NRS=11.988 M=1 R=4.33333 SA=75000.3
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1007 N_A_123_47#_M1007_d N_B1_M1007_g N_A_261_47#_M1007_s VNB NSHORT L=0.15
+ W=0.65 AD=0.104 AS=0.2015 PD=0.97 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1005 N_A_261_47#_M1005_d N_B2_M1005_g N_A_123_47#_M1007_d VNB NSHORT L=0.15
+ W=0.65 AD=0.13325 AS=0.104 PD=1.06 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_261_47#_M1005_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.13325 PD=0.92 PS=1.06 NRD=0 NRS=24.912 M=1 R=4.33333
+ SA=75001.3 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_A_261_47#_M1006_d N_A1_M1006_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_VPWR_M1001_d N_C1_M1001_g N_Y_M1001_s VPB PHIGHVT L=0.18 W=1 AD=0.485
+ AS=0.29 PD=1.97 PS=2.58 NRD=3.9203 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90002.8 A=0.18 P=2.36 MULT=1
MM1009 A_351_297# N_B1_M1009_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1 AD=0.13
+ AS=0.485 PD=1.26 PS=1.97 NRD=14.7553 NRS=3.9203 M=1 R=5.55556 SA=90001.3
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1000 N_Y_M1000_d N_B2_M1000_g A_351_297# VPB PHIGHVT L=0.18 W=1 AD=0.235
+ AS=0.13 PD=1.47 PS=1.26 NRD=0.9653 NRS=14.7553 M=1 R=5.55556 SA=90001.8
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1002 A_569_297# N_A2_M1002_g N_Y_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.235 PD=1.23 PS=1.47 NRD=11.8003 NRS=36.445 M=1 R=5.55556 SA=90002.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_569_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.115 PD=2.54 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90002.8
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
pX11_noxref noxref_15 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o221ai_1.pxi.spice"
*
.ends
*
*
