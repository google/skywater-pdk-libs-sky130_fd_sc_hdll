* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__inputiso0p_1 A SLEEP VGND VNB VPB VPWR X
X0 a_211_413# a_27_413# a_307_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 a_27_413# SLEEP VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X2 VGND a_211_413# X VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR a_211_413# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 VPWR a_27_413# a_211_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X5 VGND SLEEP a_27_413# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 a_211_413# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X7 a_307_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
