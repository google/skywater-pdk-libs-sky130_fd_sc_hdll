* File: sky130_fd_sc_hdll__nand3b_4.pex.spice
* Created: Thu Aug 27 19:14:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%A_N 3 5 7 8 17
c26 5 0 1.08454e-19 $X=0.495 $Y=1.41
r27 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.595
+ $Y=1.16 $X2=0.595 $Y2=1.16
r28 8 17 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.695 $Y2=1.175
r29 8 12 5.26818 $w=1.98e-07 $l=9.5e-08 $layer=LI1_cond $X=0.69 $Y=1.175
+ $X2=0.595 $Y2=1.175
r30 5 11 45.5843 $w=3.57e-07 $l=2.98747e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.602 $Y2=1.16
r31 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r32 1 11 36.1699 $w=3.57e-07 $l=2.00412e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.602 $Y2=1.16
r33 1 3 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=0.47 $Y=1.015
+ $X2=0.47 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%A_27_47# 1 2 7 9 12 14 16 19 21 23 26 28
+ 30 33 37 41 43 47 50 56 59 60 64 75
c109 56 0 1.39726e-19 $X=2.66 $Y=1.16
c110 33 0 1.99733e-19 $X=2.92 $Y=0.56
c111 12 0 1.08454e-19 $X=1.51 $Y=0.56
r112 75 76 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.895 $Y=1.217
+ $X2=2.92 $Y2=1.217
r113 72 73 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=2.425 $Y=1.217
+ $X2=2.45 $Y2=1.217
r114 71 72 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=1.98 $Y=1.217
+ $X2=2.425 $Y2=1.217
r115 70 71 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.955 $Y=1.217
+ $X2=1.98 $Y2=1.217
r116 67 68 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.217
+ $X2=1.51 $Y2=1.217
r117 64 67 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=1.385 $Y=1.16
+ $X2=1.485 $Y2=1.217
r118 63 64 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=1.22 $Y=1.16
+ $X2=1.385 $Y2=1.16
r119 62 63 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.22
+ $Y=1.16 $X2=1.22 $Y2=1.16
r120 57 75 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=2.66 $Y=1.217
+ $X2=2.895 $Y2=1.217
r121 57 73 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=2.66 $Y=1.217
+ $X2=2.45 $Y2=1.217
r122 56 57 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.66
+ $Y=1.16 $X2=2.66 $Y2=1.16
r123 54 70 34.6391 $w=3.27e-07 $l=2.35e-07 $layer=POLY_cond $X=1.72 $Y=1.217
+ $X2=1.955 $Y2=1.217
r124 54 68 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=1.72 $Y=1.217
+ $X2=1.51 $Y2=1.217
r125 53 56 52.1273 $w=1.98e-07 $l=9.4e-07 $layer=LI1_cond $X=1.72 $Y=1.175
+ $X2=2.66 $Y2=1.175
r126 53 54 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=1.72
+ $Y=1.16 $X2=1.72 $Y2=1.16
r127 51 62 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=1.335 $Y=1.175
+ $X2=1.195 $Y2=1.175
r128 51 53 21.35 $w=1.98e-07 $l=3.85e-07 $layer=LI1_cond $X=1.335 $Y=1.175
+ $X2=1.72 $Y2=1.175
r129 50 62 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=1.195 $Y=1.075
+ $X2=1.195 $Y2=1.175
r130 49 50 6.99698 $w=2.78e-07 $l=1.7e-07 $layer=LI1_cond $X=1.195 $Y=0.905
+ $X2=1.195 $Y2=1.075
r131 48 59 2.45687 $w=1.9e-07 $l=1.7e-07 $layer=LI1_cond $X=0.425 $Y=0.81
+ $X2=0.255 $Y2=0.81
r132 47 49 7.1467 $w=1.9e-07 $l=1.81384e-07 $layer=LI1_cond $X=1.055 $Y=0.81
+ $X2=1.195 $Y2=0.905
r133 47 48 36.7751 $w=1.88e-07 $l=6.3e-07 $layer=LI1_cond $X=1.055 $Y=0.81
+ $X2=0.425 $Y2=0.81
r134 43 45 23.0489 $w=3.38e-07 $l=6.8e-07 $layer=LI1_cond $X=0.255 $Y=1.66
+ $X2=0.255 $Y2=2.34
r135 41 60 8.46734 $w=3.38e-07 $l=1.7e-07 $layer=LI1_cond $X=0.255 $Y=1.615
+ $X2=0.255 $Y2=1.445
r136 41 43 1.52529 $w=3.38e-07 $l=4.5e-08 $layer=LI1_cond $X=0.255 $Y=1.615
+ $X2=0.255 $Y2=1.66
r137 39 59 3.98378 $w=2.57e-07 $l=1.30038e-07 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.255 $Y2=0.81
r138 39 60 34.2234 $w=1.73e-07 $l=5.4e-07 $layer=LI1_cond $X=0.172 $Y=0.905
+ $X2=0.172 $Y2=1.445
r139 35 59 3.98378 $w=2.57e-07 $l=9.5e-08 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.81
r140 35 37 11.355 $w=3.38e-07 $l=3.35e-07 $layer=LI1_cond $X=0.255 $Y=0.715
+ $X2=0.255 $Y2=0.38
r141 31 76 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=1.217
r142 31 33 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.92 $Y=1.025
+ $X2=2.92 $Y2=0.56
r143 28 75 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.217
r144 28 30 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.895 $Y=1.41
+ $X2=2.895 $Y2=1.985
r145 24 73 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=1.217
r146 24 26 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.45 $Y=1.025
+ $X2=2.45 $Y2=0.56
r147 21 72 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.217
r148 21 23 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.41
+ $X2=2.425 $Y2=1.985
r149 17 71 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=1.217
r150 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.98 $Y=1.025
+ $X2=1.98 $Y2=0.56
r151 14 70 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.217
r152 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
r153 10 68 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=1.217
r154 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.51 $Y=1.025
+ $X2=1.51 $Y2=0.56
r155 7 67 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.217
r156 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.485 $Y=1.41
+ $X2=1.485 $Y2=1.985
r157 2 45 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r158 2 43 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r159 1 37 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%B 3 5 7 10 12 14 17 19 21 22 24 27 29 30
+ 31 44 49 52 55
c73 44 0 1.39726e-19 $X=4.775 $Y=1.217
r74 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.775 $Y=1.217
+ $X2=4.8 $Y2=1.217
r75 43 55 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=4.515 $Y=1.175
+ $X2=4.8 $Y2=1.175
r76 43 52 6.65455 $w=1.98e-07 $l=1.2e-07 $layer=LI1_cond $X=4.515 $Y=1.175
+ $X2=4.395 $Y2=1.175
r77 42 44 38.3242 $w=3.27e-07 $l=2.6e-07 $layer=POLY_cond $X=4.515 $Y=1.217
+ $X2=4.775 $Y2=1.217
r78 42 43 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.515
+ $Y=1.16 $X2=4.515 $Y2=1.16
r79 40 42 30.9541 $w=3.27e-07 $l=2.1e-07 $layer=POLY_cond $X=4.305 $Y=1.217
+ $X2=4.515 $Y2=1.217
r80 39 40 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=4.28 $Y=1.217
+ $X2=4.305 $Y2=1.217
r81 38 39 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=3.835 $Y=1.217
+ $X2=4.28 $Y2=1.217
r82 37 38 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.81 $Y=1.217
+ $X2=3.835 $Y2=1.217
r83 36 37 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=3.365 $Y=1.217
+ $X2=3.81 $Y2=1.217
r84 35 36 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=3.34 $Y=1.217
+ $X2=3.365 $Y2=1.217
r85 31 55 1.66364 $w=1.98e-07 $l=3e-08 $layer=LI1_cond $X=4.83 $Y=1.175 $X2=4.8
+ $Y2=1.175
r86 30 52 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=4.37 $Y=1.175
+ $X2=4.395 $Y2=1.175
r87 30 49 24.1227 $w=1.98e-07 $l=4.35e-07 $layer=LI1_cond $X=4.37 $Y=1.175
+ $X2=3.935 $Y2=1.175
r88 29 49 1.38636 $w=1.98e-07 $l=2.5e-08 $layer=LI1_cond $X=3.91 $Y=1.175
+ $X2=3.935 $Y2=1.175
r89 25 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.8 $Y=1.025
+ $X2=4.8 $Y2=1.217
r90 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.8 $Y=1.025
+ $X2=4.8 $Y2=0.56
r91 22 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.217
r92 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.775 $Y=1.41
+ $X2=4.775 $Y2=1.985
r93 19 40 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.217
r94 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.305 $Y=1.41
+ $X2=4.305 $Y2=1.985
r95 15 39 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=1.217
r96 15 17 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.28 $Y=1.025
+ $X2=4.28 $Y2=0.56
r97 12 38 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.217
r98 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r99 8 37 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=1.217
r100 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.81 $Y=1.025
+ $X2=3.81 $Y2=0.56
r101 5 36 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.217
r102 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
r103 1 35 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=1.217
r104 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.34 $Y=1.025
+ $X2=3.34 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%C 1 3 6 8 10 13 15 17 20 22 24 27 29 30
+ 31 32 37 50 51 56 60 63 65
r77 63 65 22.4591 $w=1.98e-07 $l=4.05e-07 $layer=LI1_cond $X=6.255 $Y=1.175
+ $X2=6.66 $Y2=1.175
r78 51 52 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=7.175 $Y=1.217
+ $X2=7.2 $Y2=1.217
r79 49 51 35.3761 $w=3.27e-07 $l=2.4e-07 $layer=POLY_cond $X=6.935 $Y=1.217
+ $X2=7.175 $Y2=1.217
r80 49 50 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=6.935
+ $Y=1.16 $X2=6.935 $Y2=1.16
r81 47 49 30.2171 $w=3.27e-07 $l=2.05e-07 $layer=POLY_cond $X=6.73 $Y=1.217
+ $X2=6.935 $Y2=1.217
r82 46 47 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.705 $Y=1.217
+ $X2=6.73 $Y2=1.217
r83 45 46 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=6.26 $Y=1.217
+ $X2=6.705 $Y2=1.217
r84 44 45 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=6.235 $Y=1.217
+ $X2=6.26 $Y2=1.217
r85 43 44 65.5933 $w=3.27e-07 $l=4.45e-07 $layer=POLY_cond $X=5.79 $Y=1.217
+ $X2=6.235 $Y2=1.217
r86 42 43 3.68502 $w=3.27e-07 $l=2.5e-08 $layer=POLY_cond $X=5.765 $Y=1.217
+ $X2=5.79 $Y2=1.217
r87 40 56 9.15 $w=1.98e-07 $l=1.65e-07 $layer=LI1_cond $X=5.5 $Y=1.175 $X2=5.335
+ $Y2=1.175
r88 39 40 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.5 $Y=1.16
+ $X2=5.5 $Y2=1.16
r89 37 42 16.3472 $w=3.27e-07 $l=1.253e-07 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=5.765 $Y2=1.217
r90 37 39 36.6587 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=5.665 $Y=1.16
+ $X2=5.5 $Y2=1.16
r91 32 50 14.6955 $w=1.98e-07 $l=2.65e-07 $layer=LI1_cond $X=6.67 $Y=1.175
+ $X2=6.935 $Y2=1.175
r92 32 65 0.554545 $w=1.98e-07 $l=1e-08 $layer=LI1_cond $X=6.67 $Y=1.175
+ $X2=6.66 $Y2=1.175
r93 31 63 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=6.255 $Y2=1.175
r94 31 60 23.0136 $w=1.98e-07 $l=4.15e-07 $layer=LI1_cond $X=6.21 $Y=1.175
+ $X2=5.795 $Y2=1.175
r95 30 60 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.795 $Y2=1.175
r96 30 40 13.8636 $w=1.98e-07 $l=2.5e-07 $layer=LI1_cond $X=5.75 $Y=1.175
+ $X2=5.5 $Y2=1.175
r97 29 56 2.49545 $w=1.98e-07 $l=4.5e-08 $layer=LI1_cond $X=5.29 $Y=1.175
+ $X2=5.335 $Y2=1.175
r98 25 52 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=7.2 $Y=1.025
+ $X2=7.2 $Y2=1.217
r99 25 27 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=7.2 $Y=1.025
+ $X2=7.2 $Y2=0.56
r100 22 51 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.217
r101 22 24 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=7.175 $Y=1.41
+ $X2=7.175 $Y2=1.985
r102 18 47 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.73 $Y=1.025
+ $X2=6.73 $Y2=1.217
r103 18 20 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.73 $Y=1.025
+ $X2=6.73 $Y2=0.56
r104 15 46 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.217
r105 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.705 $Y=1.41
+ $X2=6.705 $Y2=1.985
r106 11 45 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=1.217
r107 11 13 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=6.26 $Y=1.025
+ $X2=6.26 $Y2=0.56
r108 8 44 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=6.235 $Y=1.41
+ $X2=6.235 $Y2=1.217
r109 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.235 $Y=1.41
+ $X2=6.235 $Y2=1.985
r110 4 43 21.0057 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.79 $Y=1.025
+ $X2=5.79 $Y2=1.217
r111 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.79 $Y=1.025
+ $X2=5.79 $Y2=0.56
r112 1 42 16.7191 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.765 $Y=1.41
+ $X2=5.765 $Y2=1.217
r113 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.765 $Y=1.41
+ $X2=5.765 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%VPWR 1 2 3 4 5 6 7 8 9 32 40 44 48 52 57
+ 59 61 66 67 69 70 72 73 75 76 77 89 97 102 107 111 113
r118 110 111 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=2.72
+ $X2=7.59 $Y2=2.72
r119 107 108 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r120 103 105 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r121 102 105 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r122 102 103 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r123 100 111 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=2.72
+ $X2=7.59 $Y2=2.72
r124 99 100 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=2.72
+ $X2=7.13 $Y2=2.72
r125 97 110 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.572 $Y2=2.72
r126 97 99 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.325 $Y=2.72
+ $X2=7.13 $Y2=2.72
r127 96 100 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=7.13 $Y2=2.72
r128 96 108 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.29 $Y2=2.72
r129 95 96 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r130 93 107 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=5.27 $Y2=2.72
r131 93 95 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=2.72
+ $X2=6.21 $Y2=2.72
r132 92 108 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.29 $Y2=2.72
r133 91 92 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r134 89 107 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=5.27 $Y2=2.72
r135 89 91 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=4.925 $Y=2.72
+ $X2=4.83 $Y2=2.72
r136 88 92 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.83 $Y2=2.72
r137 87 88 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r138 85 88 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r139 84 85 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r140 82 85 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r141 82 103 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r142 81 82 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r143 79 102 13.5574 $w=1.7e-07 $l=3.45e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=0.99 $Y2=2.72
r144 79 81 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r145 77 105 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.69 $Y2=2.72
r146 77 113 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=2.72
+ $X2=0.23 $Y2=2.72
r147 75 95 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.21 $Y2=2.72
r148 75 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=2.72
+ $X2=6.47 $Y2=2.72
r149 74 99 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=7.13 $Y2=2.72
r150 74 76 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=2.72
+ $X2=6.47 $Y2=2.72
r151 72 87 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=3.91 $Y2=2.72
r152 72 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.985 $Y=2.72
+ $X2=4.07 $Y2=2.72
r153 71 91 44.0374 $w=1.68e-07 $l=6.75e-07 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.83 $Y2=2.72
r154 71 73 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.155 $Y=2.72
+ $X2=4.07 $Y2=2.72
r155 69 84 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=2.99 $Y2=2.72
r156 69 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.045 $Y=2.72
+ $X2=3.13 $Y2=2.72
r157 68 87 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.91 $Y2=2.72
r158 68 70 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.215 $Y=2.72
+ $X2=3.13 $Y2=2.72
r159 66 81 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.07 $Y2=2.72
r160 66 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.105 $Y=2.72
+ $X2=2.19 $Y2=2.72
r161 65 84 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.99 $Y2=2.72
r162 65 67 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.275 $Y=2.72
+ $X2=2.19 $Y2=2.72
r163 61 64 23.7473 $w=3.28e-07 $l=6.8e-07 $layer=LI1_cond $X=7.49 $Y=1.66
+ $X2=7.49 $Y2=2.34
r164 59 110 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=7.49 $Y=2.635
+ $X2=7.572 $Y2=2.72
r165 59 64 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.49 $Y=2.635
+ $X2=7.49 $Y2=2.34
r166 55 76 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2.72
r167 55 57 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=6.47 $Y=2.635
+ $X2=6.47 $Y2=2
r168 50 107 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=2.72
r169 50 52 11.0074 $w=6.88e-07 $l=6.35e-07 $layer=LI1_cond $X=5.27 $Y=2.635
+ $X2=5.27 $Y2=2
r170 46 73 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2.72
r171 46 48 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=4.07 $Y=2.635
+ $X2=4.07 $Y2=2
r172 42 70 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.13 $Y=2.635
+ $X2=3.13 $Y2=2.72
r173 42 44 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=3.13 $Y=2.635
+ $X2=3.13 $Y2=2.34
r174 38 67 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r175 38 40 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r176 32 36 11.7874 $w=6.88e-07 $l=6.8e-07 $layer=LI1_cond $X=0.99 $Y=1.66
+ $X2=0.99 $Y2=2.34
r177 30 102 2.83173 $w=6.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.72
r178 30 36 5.11367 $w=6.88e-07 $l=2.95e-07 $layer=LI1_cond $X=0.99 $Y=2.635
+ $X2=0.99 $Y2=2.34
r179 9 64 400 $w=1.7e-07 $l=9.60937e-07 $layer=licon1_PDIFF $count=1 $X=7.265
+ $Y=1.485 $X2=7.49 $Y2=2.34
r180 9 61 400 $w=1.7e-07 $l=3e-07 $layer=licon1_PDIFF $count=1 $X=7.265 $Y=1.485
+ $X2=7.49 $Y2=1.66
r181 8 57 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=6.325
+ $Y=1.485 $X2=6.47 $Y2=2
r182 7 52 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=5.405
+ $Y=1.485 $X2=5.53 $Y2=2
r183 6 52 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=4.865
+ $Y=1.485 $X2=5.01 $Y2=2
r184 5 48 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.925
+ $Y=1.485 $X2=4.07 $Y2=2
r185 4 44 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.985
+ $Y=1.485 $X2=3.13 $Y2=2.34
r186 3 40 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.485 $X2=2.19 $Y2=2
r187 2 36 400 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=2.34
r188 2 32 400 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=1 $X=1.125
+ $Y=1.485 $X2=1.25 $Y2=1.66
r189 1 36 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
r190 1 32 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%Y 1 2 3 4 5 6 7 8 25 31 33 35 39 42 45 47
+ 48 51 53 57 59 61 63 68 70 73 84
c144 61 0 1.85528e-19 $X=6.915 $Y=1.665
r145 88 90 0.434473 $w=7.02e-07 $l=2.5e-08 $layer=LI1_cond $X=3.575 $Y=1.54
+ $X2=3.6 $Y2=1.54
r146 82 84 5.47436 $w=7.02e-07 $l=3.15e-07 $layer=LI1_cond $X=3.13 $Y=1.54
+ $X2=3.445 $Y2=1.54
r147 81 82 8.16809 $w=7.02e-07 $l=4.7e-07 $layer=LI1_cond $X=2.66 $Y=1.54
+ $X2=3.13 $Y2=1.54
r148 79 81 0.434473 $w=7.02e-07 $l=2.5e-08 $layer=LI1_cond $X=2.635 $Y=1.54
+ $X2=2.66 $Y2=1.54
r149 73 88 2.17236 $w=7.02e-07 $l=1.25e-07 $layer=LI1_cond $X=3.45 $Y=1.54
+ $X2=3.575 $Y2=1.54
r150 73 84 0.0868946 $w=7.02e-07 $l=5e-09 $layer=LI1_cond $X=3.45 $Y=1.54
+ $X2=3.445 $Y2=1.54
r151 61 72 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=6.915 $Y=1.665
+ $X2=6.915 $Y2=1.555
r152 61 63 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=6.915 $Y=1.665
+ $X2=6.915 $Y2=2.34
r153 60 70 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.165 $Y=1.555
+ $X2=5.975 $Y2=1.555
r154 59 72 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=6.725 $Y=1.555
+ $X2=6.915 $Y2=1.555
r155 59 60 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=6.725 $Y=1.555
+ $X2=6.165 $Y2=1.555
r156 55 70 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=1.555
r157 55 57 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=5.975 $Y=1.665
+ $X2=5.975 $Y2=2.34
r158 54 68 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.705 $Y=1.555
+ $X2=4.515 $Y2=1.555
r159 53 70 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=5.785 $Y=1.555
+ $X2=5.975 $Y2=1.555
r160 53 54 56.5745 $w=2.18e-07 $l=1.08e-06 $layer=LI1_cond $X=5.785 $Y=1.555
+ $X2=4.705 $Y2=1.555
r161 49 68 0.529033 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=4.515 $Y=1.665
+ $X2=4.515 $Y2=1.555
r162 49 51 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=4.515 $Y=1.665
+ $X2=4.515 $Y2=2.34
r163 48 90 9.13592 $w=7.02e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.765 $Y=1.555
+ $X2=3.6 $Y2=1.54
r164 47 68 7.92213 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=4.325 $Y=1.555
+ $X2=4.515 $Y2=1.555
r165 47 48 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=4.325 $Y=1.555
+ $X2=3.765 $Y2=1.555
r166 43 88 4.33065 $w=3.8e-07 $l=4.65e-07 $layer=LI1_cond $X=3.575 $Y=2.005
+ $X2=3.575 $Y2=1.54
r167 43 45 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=3.575 $Y=2.005
+ $X2=3.575 $Y2=2.34
r168 42 82 9.34032 $w=1.7e-07 $l=4.65e-07 $layer=LI1_cond $X=3.13 $Y=1.075
+ $X2=3.13 $Y2=1.54
r169 41 42 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.13 $Y=0.905
+ $X2=3.13 $Y2=1.075
r170 37 79 4.33065 $w=3.8e-07 $l=4.65e-07 $layer=LI1_cond $X=2.635 $Y=2.005
+ $X2=2.635 $Y2=1.54
r171 37 39 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=2.635 $Y=2.005
+ $X2=2.635 $Y2=2.34
r172 36 66 4.72888 $w=2.2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.885 $Y=1.555
+ $X2=1.695 $Y2=1.555
r173 35 79 9.57039 $w=7.02e-07 $l=1.97358e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=2.635 $Y2=1.54
r174 35 36 29.3349 $w=2.18e-07 $l=5.6e-07 $layer=LI1_cond $X=2.445 $Y=1.555
+ $X2=1.885 $Y2=1.555
r175 31 66 2.73777 $w=3.8e-07 $l=1.1e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=1.555
r176 31 33 20.471 $w=3.78e-07 $l=6.75e-07 $layer=LI1_cond $X=1.695 $Y=1.665
+ $X2=1.695 $Y2=2.34
r177 27 30 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=1.72 $Y=0.77
+ $X2=2.66 $Y2=0.77
r178 25 41 7.28469 $w=2.7e-07 $l=1.72337e-07 $layer=LI1_cond $X=3.045 $Y=0.77
+ $X2=3.13 $Y2=0.905
r179 25 30 16.433 $w=2.68e-07 $l=3.85e-07 $layer=LI1_cond $X=3.045 $Y=0.77
+ $X2=2.66 $Y2=0.77
r180 8 72 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.485 $X2=6.94 $Y2=1.66
r181 8 63 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=6.795
+ $Y=1.485 $X2=6.94 $Y2=2.34
r182 7 70 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.485 $X2=6 $Y2=1.66
r183 7 57 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.855
+ $Y=1.485 $X2=6 $Y2=2.34
r184 6 68 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=1.66
r185 6 51 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=4.395
+ $Y=1.485 $X2=4.54 $Y2=2.34
r186 5 90 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=1.66
r187 5 45 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=2.34
r188 4 81 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=1.66
r189 4 39 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.515
+ $Y=1.485 $X2=2.66 $Y2=2.34
r190 3 66 400 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=1.66
r191 3 33 400 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.575
+ $Y=1.485 $X2=1.72 $Y2=2.34
r192 2 30 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=2.525
+ $Y=0.235 $X2=2.66 $Y2=0.72
r193 1 27 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.235 $X2=1.72 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%VGND 1 2 3 4 17 21 25 27 29 32 33 35 36
+ 37 49 54 58 60
r87 57 58 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=7.59 $Y=0 $X2=7.59
+ $Y2=0
r88 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r89 52 58 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=7.13 $Y=0 $X2=7.59
+ $Y2=0
r90 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=7.13 $Y=0 $X2=7.13
+ $Y2=0
r91 49 57 4.63344 $w=1.7e-07 $l=2.47e-07 $layer=LI1_cond $X=7.325 $Y=0 $X2=7.572
+ $Y2=0
r92 49 51 12.7219 $w=1.68e-07 $l=1.95e-07 $layer=LI1_cond $X=7.325 $Y=0 $X2=7.13
+ $Y2=0
r93 48 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=7.13
+ $Y2=0
r94 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r95 45 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r96 44 45 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r97 42 45 1.178 $w=4.8e-07 $l=4.14e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=5.29
+ $Y2=0
r98 42 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r99 41 44 270.096 $w=1.68e-07 $l=4.14e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=5.29
+ $Y2=0
r100 41 42 1.86 $w=1.7e-07 $l=8.5e-07 $layer=mcon $count=5 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r101 39 54 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.77
+ $Y2=0
r102 39 41 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r103 37 55 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r104 37 60 0.00142271 $w=4.8e-07 $l=5e-09 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.23 $Y2=0
r105 35 47 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=6.385 $Y=0
+ $X2=6.21 $Y2=0
r106 35 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.385 $Y=0 $X2=6.47
+ $Y2=0
r107 34 51 37.5134 $w=1.68e-07 $l=5.75e-07 $layer=LI1_cond $X=6.555 $Y=0
+ $X2=7.13 $Y2=0
r108 34 36 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.555 $Y=0 $X2=6.47
+ $Y2=0
r109 32 44 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.29
+ $Y2=0
r110 32 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.365 $Y=0 $X2=5.49
+ $Y2=0
r111 31 47 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=5.615 $Y=0
+ $X2=6.21 $Y2=0
r112 31 33 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=5.615 $Y=0 $X2=5.49
+ $Y2=0
r113 27 57 3.13273 $w=3.3e-07 $l=1.19143e-07 $layer=LI1_cond $X=7.49 $Y=0.085
+ $X2=7.572 $Y2=0
r114 27 29 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=7.49 $Y=0.085
+ $X2=7.49 $Y2=0.38
r115 23 36 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0
r116 23 25 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.47 $Y=0.085
+ $X2=6.47 $Y2=0.38
r117 19 33 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=5.49 $Y=0.085
+ $X2=5.49 $Y2=0
r118 19 21 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=5.49 $Y=0.085
+ $X2=5.49 $Y2=0.38
r119 15 54 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0
r120 15 17 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=0.77 $Y=0.085
+ $X2=0.77 $Y2=0.38
r121 4 29 91 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_NDIFF $count=2 $X=7.275
+ $Y=0.235 $X2=7.49 $Y2=0.38
r122 3 25 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=6.335
+ $Y=0.235 $X2=6.47 $Y2=0.38
r123 2 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=5.405
+ $Y=0.235 $X2=5.53 $Y2=0.38
r124 1 17 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=0.545
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%A_225_47# 1 2 3 4 5 26
r34 24 26 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=4.07 $Y=0.36 $X2=5.01
+ $Y2=0.36
r35 22 24 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=3.13 $Y=0.36 $X2=4.07
+ $Y2=0.36
r36 20 22 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=2.19 $Y=0.36 $X2=3.13
+ $Y2=0.36
r37 17 20 49.645 $w=2.08e-07 $l=9.4e-07 $layer=LI1_cond $X=1.25 $Y=0.36 $X2=2.19
+ $Y2=0.36
r38 5 26 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.875
+ $Y=0.235 $X2=5.01 $Y2=0.38
r39 4 24 182 $w=1.7e-07 $l=2.47083e-07 $layer=licon1_NDIFF $count=1 $X=3.885
+ $Y=0.235 $X2=4.07 $Y2=0.38
r40 3 22 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.995
+ $Y=0.235 $X2=3.13 $Y2=0.38
r41 2 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.38
r42 1 17 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.125
+ $Y=0.235 $X2=1.25 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__NAND3B_4%A_683_47# 1 2 3 4 13 19 23 25 29 31 32
c56 25 0 1.85528e-19 $X=6.725 $Y=0.81
c57 13 0 1.99733e-19 $X=5.04 $Y=0.77
r58 27 29 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=6.915 $Y=0.715
+ $X2=6.915 $Y2=0.38
r59 26 32 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=6.165 $Y=0.81
+ $X2=5.975 $Y2=0.81
r60 25 27 7.85115 $w=1.9e-07 $l=2.32702e-07 $layer=LI1_cond $X=6.725 $Y=0.81
+ $X2=6.915 $Y2=0.715
r61 25 26 32.689 $w=1.88e-07 $l=5.6e-07 $layer=LI1_cond $X=6.725 $Y=0.81
+ $X2=6.165 $Y2=0.81
r62 21 32 0.987631 $w=3.8e-07 $l=9.5e-08 $layer=LI1_cond $X=5.975 $Y=0.715
+ $X2=5.975 $Y2=0.81
r63 21 23 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.975 $Y=0.715
+ $X2=5.975 $Y2=0.38
r64 19 32 8.79175 $w=1.9e-07 $l=1.9e-07 $layer=LI1_cond $X=5.785 $Y=0.81
+ $X2=5.975 $Y2=0.81
r65 19 31 35.6077 $w=1.88e-07 $l=6.1e-07 $layer=LI1_cond $X=5.785 $Y=0.81
+ $X2=5.175 $Y2=0.81
r66 15 18 40.1221 $w=2.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.6 $Y=0.77 $X2=4.54
+ $Y2=0.77
r67 13 31 6.78806 $w=2.68e-07 $l=1.35e-07 $layer=LI1_cond $X=5.04 $Y=0.77
+ $X2=5.175 $Y2=0.77
r68 13 18 21.3415 $w=2.68e-07 $l=5e-07 $layer=LI1_cond $X=5.04 $Y=0.77 $X2=4.54
+ $Y2=0.77
r69 4 29 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.805
+ $Y=0.235 $X2=6.94 $Y2=0.38
r70 3 23 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.865
+ $Y=0.235 $X2=6 $Y2=0.38
r71 2 18 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=4.355
+ $Y=0.235 $X2=4.54 $Y2=0.72
r72 1 15 182 $w=1.7e-07 $l=5.70044e-07 $layer=licon1_NDIFF $count=1 $X=3.415
+ $Y=0.235 $X2=3.6 $Y2=0.72
.ends

