* File: sky130_fd_sc_hdll__a31oi_1.pxi.spice
* Created: Thu Aug 27 18:55:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__A31OI_1%A3 N_A3_c_42_n N_A3_M1004_g N_A3_c_43_n
+ N_A3_M1005_g A3 N_A3_c_44_n PM_SKY130_FD_SC_HDLL__A31OI_1%A3
x_PM_SKY130_FD_SC_HDLL__A31OI_1%A2 N_A2_c_62_n N_A2_M1002_g N_A2_c_63_n
+ N_A2_M1000_g A2 A2 A2 PM_SKY130_FD_SC_HDLL__A31OI_1%A2
x_PM_SKY130_FD_SC_HDLL__A31OI_1%A1 N_A1_c_94_n N_A1_M1007_g N_A1_c_95_n
+ N_A1_M1001_g N_A1_c_96_n N_A1_c_99_n A1 A1 PM_SKY130_FD_SC_HDLL__A31OI_1%A1
x_PM_SKY130_FD_SC_HDLL__A31OI_1%B1 N_B1_c_132_n N_B1_M1003_g N_B1_c_136_n
+ N_B1_M1006_g N_B1_c_133_n B1 N_B1_c_135_n B1 PM_SKY130_FD_SC_HDLL__A31OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A31OI_1%VPWR N_VPWR_M1004_s N_VPWR_M1000_d
+ N_VPWR_c_167_n N_VPWR_c_168_n N_VPWR_c_169_n VPWR N_VPWR_c_170_n
+ N_VPWR_c_171_n N_VPWR_c_166_n N_VPWR_c_173_n
+ PM_SKY130_FD_SC_HDLL__A31OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A31OI_1%A_117_297# N_A_117_297#_M1004_d
+ N_A_117_297#_M1001_d N_A_117_297#_c_204_n N_A_117_297#_c_205_n
+ N_A_117_297#_c_207_n N_A_117_297#_c_211_n
+ PM_SKY130_FD_SC_HDLL__A31OI_1%A_117_297#
x_PM_SKY130_FD_SC_HDLL__A31OI_1%Y N_Y_M1007_d N_Y_M1006_d N_Y_c_232_n
+ N_Y_c_229_n N_Y_c_228_n Y Y PM_SKY130_FD_SC_HDLL__A31OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A31OI_1%VGND N_VGND_M1005_s N_VGND_M1003_d
+ N_VGND_c_265_n N_VGND_c_266_n N_VGND_c_267_n N_VGND_c_268_n VGND
+ N_VGND_c_269_n N_VGND_c_270_n PM_SKY130_FD_SC_HDLL__A31OI_1%VGND
cc_1 VNB N_A3_c_42_n 0.0333543f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A3_c_43_n 0.022189f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A3_c_44_n 0.0130035f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_4 VNB N_A2_c_62_n 0.0159401f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_A2_c_63_n 0.0201994f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB A2 0.0121097f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_7 VNB N_A1_c_94_n 0.0181102f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A1_c_95_n 0.0215418f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB N_A1_c_96_n 0.0039105f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_10 VNB N_B1_c_132_n 0.0210964f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_B1_c_133_n 0.0138256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB B1 0.0144946f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_13 VNB N_B1_c_135_n 0.040396f $X=-0.19 $Y=-0.24 $X2=0.23 $Y2=1.16
cc_14 VNB N_VPWR_c_166_n 0.117919f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_Y_c_228_n 0.00377889f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_265_n 0.0116117f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=1.105
cc_17 VNB N_VGND_c_266_n 0.0286227f $X=-0.19 $Y=-0.24 $X2=0.405 $Y2=1.16
cc_18 VNB N_VGND_c_267_n 0.0127572f $X=-0.19 $Y=-0.24 $X2=0.35 $Y2=1.16
cc_19 VNB N_VGND_c_268_n 0.018315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_269_n 0.0498888f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_VGND_c_270_n 0.164004f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VPB N_A3_c_42_n 0.0348612f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_23 VPB N_A3_c_44_n 0.00208732f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_24 VPB N_A2_c_63_n 0.0253031f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_25 VPB N_A1_c_95_n 0.0248614f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_26 VPB N_A1_c_96_n 0.00142353f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_27 VPB N_A1_c_99_n 0.00878239f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_28 VPB N_B1_c_136_n 0.0201868f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_29 VPB N_B1_c_133_n 0.00763397f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB B1 0.00462051f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_31 VPB N_B1_c_135_n 0.0162294f $X=-0.19 $Y=1.305 $X2=0.23 $Y2=1.16
cc_32 VPB N_VPWR_c_167_n 0.0102394f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=1.105
cc_33 VPB N_VPWR_c_168_n 0.0416087f $X=-0.19 $Y=1.305 $X2=0.405 $Y2=1.16
cc_34 VPB N_VPWR_c_169_n 0.00278317f $X=-0.19 $Y=1.305 $X2=0.35 $Y2=1.16
cc_35 VPB N_VPWR_c_170_n 0.0150949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_VPWR_c_171_n 0.0400865f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_VPWR_c_166_n 0.0539625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_173_n 0.00513543f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_Y_c_229_n 0.00874992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_Y_c_228_n 0.00549657f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB Y 0.0298621f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 N_A3_c_43_n N_A2_c_62_n 0.029553f $X=0.52 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_43 N_A3_c_42_n N_A2_c_63_n 0.064544f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_44 N_A3_c_44_n N_A2_c_63_n 4.25972e-19 $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_45 N_A3_c_43_n A2 0.00860769f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_46 N_A3_c_44_n A2 0.0232484f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_47 N_A3_c_42_n N_VPWR_c_168_n 0.0232094f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_48 N_A3_c_44_n N_VPWR_c_168_n 0.0250351f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_49 N_A3_c_42_n N_VPWR_c_169_n 6.36003e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_50 N_A3_c_42_n N_VPWR_c_170_n 0.00642146f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A3_c_42_n N_VPWR_c_166_n 0.0108123f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A3_c_42_n N_VGND_c_266_n 0.00493595f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A3_c_43_n N_VGND_c_266_n 0.00487766f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A3_c_44_n N_VGND_c_266_n 0.0255334f $X=0.35 $Y=1.16 $X2=0 $Y2=0
cc_55 N_A3_c_43_n N_VGND_c_269_n 0.00585385f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A3_c_43_n N_VGND_c_270_n 0.0115523f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_57 N_A2_c_62_n N_A1_c_94_n 0.0283137f $X=0.94 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_58 A2 N_A1_c_94_n 0.0103335f $X=0.66 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_59 N_A2_c_63_n N_A1_c_95_n 0.0544503f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A2_c_63_n N_A1_c_96_n 0.00190967f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_61 A2 N_A1_c_96_n 0.0200911f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_62 N_A2_c_63_n N_A1_c_99_n 0.00393488f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_63 A2 N_A1_c_99_n 0.00819259f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_64 N_A2_c_63_n N_VPWR_c_168_n 0.00209281f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A2_c_63_n N_VPWR_c_169_n 0.00812599f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_66 N_A2_c_63_n N_VPWR_c_170_n 0.00464801f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_67 N_A2_c_63_n N_VPWR_c_166_n 0.00541961f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_68 N_A2_c_63_n N_A_117_297#_c_204_n 0.00438908f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_69 N_A2_c_63_n N_A_117_297#_c_205_n 0.0156668f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_70 A2 N_A_117_297#_c_205_n 0.00646159f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_71 A2 N_A_117_297#_c_207_n 0.00668255f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_72 N_A2_c_62_n N_Y_c_232_n 6.28592e-19 $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_73 A2 N_Y_c_232_n 0.0260438f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_74 N_A2_c_62_n N_VGND_c_269_n 0.00373852f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_75 A2 N_VGND_c_269_n 0.0220321f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_76 N_A2_c_62_n N_VGND_c_270_n 0.0055679f $X=0.94 $Y=0.995 $X2=0 $Y2=0
cc_77 A2 N_VGND_c_270_n 0.0198829f $X=0.66 $Y=0.425 $X2=0 $Y2=0
cc_78 A2 A_119_47# 0.00280566f $X=0.66 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_79 A2 A_203_47# 0.00743603f $X=0.66 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_80 N_A1_c_94_n N_B1_c_132_n 0.00835782f $X=1.445 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_81 N_A1_c_95_n N_B1_c_136_n 0.0328402f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A1_c_96_n N_B1_c_136_n 2.61816e-19 $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_83 N_A1_c_99_n N_B1_c_136_n 0.00183333f $X=1.37 $Y=1.555 $X2=0 $Y2=0
cc_84 N_A1_c_95_n N_B1_c_133_n 0.0198762f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A1_c_96_n N_B1_c_133_n 0.00327917f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A1_c_99_n N_VPWR_M1000_d 0.00304699f $X=1.37 $Y=1.555 $X2=0 $Y2=0
cc_87 N_A1_c_95_n N_VPWR_c_169_n 0.00318096f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A1_c_95_n N_VPWR_c_171_n 0.00523784f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A1_c_95_n N_VPWR_c_166_n 0.00708275f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A1_c_99_n N_A_117_297#_M1001_d 0.00278382f $X=1.37 $Y=1.555 $X2=0 $Y2=0
cc_91 N_A1_c_95_n N_A_117_297#_c_205_n 0.0139738f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_92 N_A1_c_99_n N_A_117_297#_c_205_n 0.0361334f $X=1.37 $Y=1.555 $X2=0 $Y2=0
cc_93 N_A1_c_95_n N_A_117_297#_c_211_n 0.00465166f $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_94 N_A1_c_94_n N_Y_c_232_n 0.00898193f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A1_c_95_n N_Y_c_232_n 7.58557e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_96 N_A1_c_96_n N_Y_c_232_n 0.0158768f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_97 N_A1_c_95_n N_Y_c_229_n 8.88284e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A1_c_94_n N_Y_c_228_n 6.93201e-19 $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_99 N_A1_c_95_n N_Y_c_228_n 6.69813e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A1_c_96_n N_Y_c_228_n 0.022786f $X=1.505 $Y=1.16 $X2=0 $Y2=0
cc_101 N_A1_c_99_n N_Y_c_228_n 0.0120768f $X=1.37 $Y=1.555 $X2=0 $Y2=0
cc_102 N_A1_c_95_n Y 2.68909e-19 $X=1.47 $Y=1.41 $X2=0 $Y2=0
cc_103 N_A1_c_94_n N_VGND_c_269_n 0.00526912f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_104 N_A1_c_94_n N_VGND_c_270_n 0.00979147f $X=1.445 $Y=0.995 $X2=0 $Y2=0
cc_105 N_B1_c_136_n N_VPWR_c_171_n 0.00554913f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B1_c_136_n N_VPWR_c_166_n 0.0103036f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B1_c_136_n N_A_117_297#_c_205_n 0.0014443f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B1_c_136_n N_A_117_297#_c_211_n 0.00309878f $X=1.995 $Y=1.41 $X2=0
+ $Y2=0
cc_109 N_B1_c_132_n N_Y_c_232_n 0.0223611f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_110 N_B1_c_133_n N_Y_c_232_n 5.22569e-19 $X=1.995 $Y=1.202 $X2=0 $Y2=0
cc_111 N_B1_c_136_n N_Y_c_229_n 0.00428392f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_112 B1 N_Y_c_229_n 0.00701389f $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_113 N_B1_c_135_n N_Y_c_229_n 0.00951185f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_114 N_B1_c_132_n N_Y_c_228_n 0.0065307f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_115 N_B1_c_136_n N_Y_c_228_n 0.00270032f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B1_c_133_n N_Y_c_228_n 0.0107138f $X=1.995 $Y=1.202 $X2=0 $Y2=0
cc_117 B1 N_Y_c_228_n 0.0235173f $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_118 N_B1_c_135_n N_Y_c_228_n 0.00873736f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_119 N_B1_c_136_n Y 0.0142627f $X=1.995 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B1_c_132_n N_VGND_c_268_n 0.0063883f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_121 B1 N_VGND_c_268_n 0.0106263f $X=2.465 $Y=1.105 $X2=0 $Y2=0
cc_122 N_B1_c_135_n N_VGND_c_268_n 0.00430211f $X=2.41 $Y=1.16 $X2=0 $Y2=0
cc_123 N_B1_c_132_n N_VGND_c_269_n 0.00366111f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_124 N_B1_c_132_n N_VGND_c_270_n 0.00669912f $X=1.97 $Y=0.995 $X2=0 $Y2=0
cc_125 N_VPWR_c_166_n N_A_117_297#_M1004_d 0.00457543f $X=2.53 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_126 N_VPWR_c_166_n N_A_117_297#_M1001_d 0.00623459f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_127 N_VPWR_c_169_n N_A_117_297#_c_204_n 0.0145615f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_128 N_VPWR_c_170_n N_A_117_297#_c_204_n 0.00906681f $X=1.035 $Y=2.72 $X2=0
+ $Y2=0
cc_129 N_VPWR_c_166_n N_A_117_297#_c_204_n 0.00645867f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_130 N_VPWR_M1000_d N_A_117_297#_c_205_n 0.00440749f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_131 N_VPWR_c_169_n N_A_117_297#_c_205_n 0.01782f $X=1.2 $Y=2.34 $X2=0 $Y2=0
cc_132 N_VPWR_c_170_n N_A_117_297#_c_205_n 0.00265818f $X=1.035 $Y=2.72 $X2=0
+ $Y2=0
cc_133 N_VPWR_c_171_n N_A_117_297#_c_205_n 0.00305111f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_134 N_VPWR_c_166_n N_A_117_297#_c_205_n 0.0121722f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_135 N_VPWR_c_171_n N_A_117_297#_c_211_n 0.0101429f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_136 N_VPWR_c_166_n N_A_117_297#_c_211_n 0.00721179f $X=2.53 $Y=2.72 $X2=0
+ $Y2=0
cc_137 N_VPWR_c_166_n N_Y_M1006_d 0.00226583f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_138 N_VPWR_c_171_n Y 0.0244406f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_139 N_VPWR_c_166_n Y 0.0156038f $X=2.53 $Y=2.72 $X2=0 $Y2=0
cc_140 N_A_117_297#_c_205_n Y 0.0142914f $X=1.62 $Y=1.92 $X2=0 $Y2=0
cc_141 N_A_117_297#_c_211_n Y 0.0311525f $X=1.705 $Y=2.25 $X2=0 $Y2=0
cc_142 N_Y_c_232_n N_VGND_M1003_d 0.0153442f $X=2.07 $Y=0.56 $X2=0 $Y2=0
cc_143 N_Y_c_228_n N_VGND_M1003_d 0.00244197f $X=2.197 $Y=1.495 $X2=0 $Y2=0
cc_144 N_Y_c_232_n N_VGND_c_268_n 0.0225167f $X=2.07 $Y=0.56 $X2=0 $Y2=0
cc_145 N_Y_c_232_n N_VGND_c_269_n 0.0320104f $X=2.07 $Y=0.56 $X2=0 $Y2=0
cc_146 N_Y_M1007_d N_VGND_c_270_n 0.00302875f $X=1.52 $Y=0.235 $X2=0 $Y2=0
cc_147 N_Y_c_232_n N_VGND_c_270_n 0.0242483f $X=2.07 $Y=0.56 $X2=0 $Y2=0
cc_148 N_VGND_c_270_n A_119_47# 0.00261944f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
cc_149 N_VGND_c_270_n A_203_47# 0.010042f $X=2.53 $Y=0 $X2=-0.19 $Y2=-0.24
