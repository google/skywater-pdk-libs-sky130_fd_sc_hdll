* File: sky130_fd_sc_hdll__and2b_2.pex.spice
* Created: Wed Sep  2 08:21:57 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%A_N 2 3 5 8 10 13 18 23
c35 13 0 1.89169e-19 $X=0.365 $Y=1.16
r36 14 23 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=0.297 $Y=1.16
+ $X2=0.297 $Y2=1.19
r37 14 18 11.7134 $w=3.03e-07 $l=3.1e-07 $layer=LI1_cond $X=0.297 $Y=1.16
+ $X2=0.297 $Y2=0.85
r38 13 16 36.7604 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.397 $Y=1.16
+ $X2=0.397 $Y2=1.325
r39 13 15 45.5639 $w=3.95e-07 $l=1.65e-07 $layer=POLY_cond $X=0.397 $Y=1.16
+ $X2=0.397 $Y2=0.995
r40 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.365
+ $Y=1.16 $X2=0.365 $Y2=1.16
r41 10 23 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.297 $Y=1.53
+ $X2=0.297 $Y2=1.19
r42 8 15 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=0.52 $Y=0.445
+ $X2=0.52 $Y2=0.995
r43 3 5 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=0.495 $Y=1.99
+ $X2=0.495 $Y2=2.275
r44 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=0.495 $Y=1.89 $X2=0.495
+ $Y2=1.99
r45 2 16 187.341 $w=2e-07 $l=5.65e-07 $layer=POLY_cond $X=0.495 $Y=1.89
+ $X2=0.495 $Y2=1.325
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%A_27_413# 1 2 8 9 11 14 18 20 21 23 25 27
+ 34 35
c68 34 0 1.13894e-19 $X=1.14 $Y=0.97
c69 20 0 3.48245e-19 $X=0.67 $Y=1.9
c70 8 0 1.63008e-19 $X=1.06 $Y=1.89
r71 35 37 15.1216 $w=2.55e-07 $l=8e-08 $layer=POLY_cond $X=1.14 $Y=0.97 $X2=1.06
+ $Y2=0.97
r72 34 35 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.14
+ $Y=0.97 $X2=1.14 $Y2=0.97
r73 32 34 12.3276 $w=3.28e-07 $l=3.53e-07 $layer=LI1_cond $X=0.787 $Y=0.97
+ $X2=1.14 $Y2=0.97
r74 30 32 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=0.777 $Y=0.97
+ $X2=0.787 $Y2=0.97
r75 27 29 10.235 $w=2.38e-07 $l=2.1e-07 $layer=LI1_cond $X=0.765 $Y=0.445
+ $X2=0.765 $Y2=0.655
r76 24 32 2.74472 $w=2.35e-07 $l=1.65e-07 $layer=LI1_cond $X=0.787 $Y=1.135
+ $X2=0.787 $Y2=0.97
r77 24 25 31.8761 $w=2.33e-07 $l=6.5e-07 $layer=LI1_cond $X=0.787 $Y=1.135
+ $X2=0.787 $Y2=1.785
r78 23 30 3.26307 $w=2.15e-07 $l=1.65e-07 $layer=LI1_cond $X=0.777 $Y=0.805
+ $X2=0.777 $Y2=0.97
r79 23 29 8.0403 $w=2.13e-07 $l=1.5e-07 $layer=LI1_cond $X=0.777 $Y=0.805
+ $X2=0.777 $Y2=0.655
r80 20 25 6.81752 $w=2.3e-07 $l=1.64754e-07 $layer=LI1_cond $X=0.67 $Y=1.9
+ $X2=0.787 $Y2=1.785
r81 20 21 16.2845 $w=2.28e-07 $l=3.25e-07 $layer=LI1_cond $X=0.67 $Y=1.9
+ $X2=0.345 $Y2=1.9
r82 16 21 7.01789 $w=2.3e-07 $l=1.51658e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.345 $Y2=1.9
r83 16 18 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.26 $Y=2.015
+ $X2=0.26 $Y2=2.225
r84 12 35 79.3882 $w=2.55e-07 $l=4.95681e-07 $layer=POLY_cond $X=1.56 $Y=0.805
+ $X2=1.14 $Y2=0.97
r85 12 14 184.596 $w=1.5e-07 $l=3.6e-07 $layer=POLY_cond $X=1.56 $Y=0.805
+ $X2=1.56 $Y2=0.445
r86 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.06 $Y=1.99
+ $X2=1.06 $Y2=2.275
r87 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.06 $Y=1.89 $X2=1.06
+ $Y2=1.99
r88 7 37 8.54376 $w=2e-07 $l=1.65e-07 $layer=POLY_cond $X=1.06 $Y=1.135 $X2=1.06
+ $Y2=0.97
r89 7 8 250.341 $w=2e-07 $l=7.55e-07 $layer=POLY_cond $X=1.06 $Y=1.135 $X2=1.06
+ $Y2=1.89
r90 2 18 600 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=2.065 $X2=0.26 $Y2=2.225
r91 1 27 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%B 1 3 6 8
c31 8 0 1.63008e-19 $X=2.07 $Y=1.87
c32 6 0 2.45633e-19 $X=2.03 $Y=0.445
r33 11 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.82
+ $Y=1.73 $X2=1.82 $Y2=1.73
r34 8 12 9.29389 $w=3.08e-07 $l=2.5e-07 $layer=LI1_cond $X=2.07 $Y=1.8 $X2=1.82
+ $Y2=1.8
r35 4 11 81.466 $w=4.82e-07 $l=6.79831e-07 $layer=POLY_cond $X=2.03 $Y=1.165
+ $X2=1.777 $Y2=1.73
r36 4 6 369.191 $w=1.5e-07 $l=7.2e-07 $layer=POLY_cond $X=2.03 $Y=1.165 $X2=2.03
+ $Y2=0.445
r37 1 11 45.8181 $w=4.82e-07 $l=3.55837e-07 $layer=POLY_cond $X=1.55 $Y=1.99
+ $X2=1.777 $Y2=1.73
r38 1 3 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.55 $Y=1.99 $X2=1.55
+ $Y2=2.275
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%A_230_413# 1 2 7 9 10 12 13 14 15 17 18 20
+ 21 24 27 28 30 36
r82 39 40 3.08184 $w=3.91e-07 $l=2.5e-08 $layer=POLY_cond $X=2.545 $Y=1.197
+ $X2=2.57 $Y2=1.197
r83 36 37 12.494 $w=2.49e-07 $l=2.55e-07 $layer=LI1_cond $X=1.3 $Y=0.44
+ $X2=1.555 $Y2=0.44
r84 31 39 11.711 $w=3.91e-07 $l=9.5e-08 $layer=POLY_cond $X=2.45 $Y=1.197
+ $X2=2.545 $Y2=1.197
r85 30 31 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.45
+ $Y=1.16 $X2=2.45 $Y2=1.16
r86 28 34 16.6301 $w=4.05e-07 $l=5.86302e-07 $layer=LI1_cond $X=2.105 $Y=1.135
+ $X2=1.555 $Y2=1.21
r87 28 30 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=2.105 $Y=1.135
+ $X2=2.45 $Y2=1.135
r88 27 34 4.30998 $w=2.2e-07 $l=2.65e-07 $layer=LI1_cond $X=1.555 $Y=0.945
+ $X2=1.555 $Y2=1.21
r89 26 37 1.46089 $w=2.2e-07 $l=1.7e-07 $layer=LI1_cond $X=1.555 $Y=0.61
+ $X2=1.555 $Y2=0.44
r90 26 27 17.5486 $w=2.18e-07 $l=3.35e-07 $layer=LI1_cond $X=1.555 $Y=0.61
+ $X2=1.555 $Y2=0.945
r91 22 34 8.82617 $w=4.05e-07 $l=4.04344e-07 $layer=LI1_cond $X=1.262 $Y=1.475
+ $X2=1.555 $Y2=1.21
r92 22 24 25.801 $w=3.33e-07 $l=7.5e-07 $layer=LI1_cond $X=1.262 $Y=1.475
+ $X2=1.262 $Y2=2.225
r93 18 21 35.458 $w=1.65e-07 $l=2.24152e-07 $layer=POLY_cond $X=3.2 $Y=0.985
+ $X2=3.175 $Y2=1.197
r94 18 20 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=3.2 $Y=0.985
+ $X2=3.2 $Y2=0.56
r95 15 21 35.458 $w=1.65e-07 $l=2.13e-07 $layer=POLY_cond $X=3.175 $Y=1.41
+ $X2=3.175 $Y2=1.197
r96 15 17 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.175 $Y=1.41
+ $X2=3.175 $Y2=1.985
r97 14 40 10.1945 $w=3.91e-07 $l=9.3675e-08 $layer=POLY_cond $X=2.645 $Y=1.155
+ $X2=2.57 $Y2=1.197
r98 13 21 4.25972 $w=3.4e-07 $l=1.19164e-07 $layer=POLY_cond $X=3.075 $Y=1.155
+ $X2=3.175 $Y2=1.197
r99 13 14 72.9789 $w=3.4e-07 $l=4.3e-07 $layer=POLY_cond $X=3.075 $Y=1.155
+ $X2=2.645 $Y2=1.155
r100 10 40 25.3065 $w=1.5e-07 $l=2.12e-07 $layer=POLY_cond $X=2.57 $Y=0.985
+ $X2=2.57 $Y2=1.197
r101 10 12 136.567 $w=1.5e-07 $l=4.25e-07 $layer=POLY_cond $X=2.57 $Y=0.985
+ $X2=2.57 $Y2=0.56
r102 7 39 20.9208 $w=1.8e-07 $l=2.13e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.197
r103 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.545 $Y=1.41
+ $X2=2.545 $Y2=1.985
r104 2 24 600 $w=1.7e-07 $l=2.24499e-07 $layer=licon1_PDIFF $count=1 $X=1.15
+ $Y=2.065 $X2=1.305 $Y2=2.225
r105 1 36 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=1.175
+ $Y=0.235 $X2=1.3 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%VPWR 1 2 3 12 14 16 18 20 30 36 41 44 47
c44 41 0 1.59076e-19 $X=1.66 $Y=2.485
r45 46 47 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 43 44 10.5103 $w=6.38e-07 $l=1.7e-07 $layer=LI1_cond $X=2.225 $Y=2.485
+ $X2=2.395 $Y2=2.485
r47 39 43 2.89675 $w=6.38e-07 $l=1.55e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=2.225 $Y2=2.485
r48 39 41 14.9956 $w=6.38e-07 $l=4.1e-07 $layer=LI1_cond $X=2.07 $Y=2.485
+ $X2=1.66 $Y2=2.485
r49 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r50 36 37 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r51 34 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.45 $Y2=2.72
r52 34 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.07 $Y2=2.72
r53 33 44 38.8182 $w=1.68e-07 $l=5.95e-07 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=2.395 $Y2=2.72
r54 33 34 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r55 30 46 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.502 $Y2=2.72
r56 30 33 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=2.99 $Y2=2.72
r57 29 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.07 $Y2=2.72
r58 29 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=0.69 $Y2=2.72
r59 28 41 3.26203 $w=1.68e-07 $l=5e-08 $layer=LI1_cond $X=1.61 $Y=2.72 $X2=1.66
+ $Y2=2.72
r60 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r61 26 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r62 26 28 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.61 $Y2=2.72
r63 20 36 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r64 20 22 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r65 18 37 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r66 18 22 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r67 14 46 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.46 $Y=2.635
+ $X2=3.502 $Y2=2.72
r68 14 16 33.0794 $w=2.68e-07 $l=7.75e-07 $layer=LI1_cond $X=3.46 $Y=2.635
+ $X2=3.46 $Y2=1.86
r69 10 36 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.72
r70 10 12 11.0695 $w=3.78e-07 $l=3.65e-07 $layer=LI1_cond $X=0.705 $Y=2.635
+ $X2=0.705 $Y2=2.27
r71 3 16 300 $w=1.7e-07 $l=4.41588e-07 $layer=licon1_PDIFF $count=2 $X=3.265
+ $Y=1.485 $X2=3.41 $Y2=1.86
r72 2 43 300 $w=1.7e-07 $l=7.0516e-07 $layer=licon1_PDIFF $count=2 $X=1.64
+ $Y=2.065 $X2=2.225 $Y2=2.33
r73 1 12 600 $w=1.7e-07 $l=2.67862e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=2.065 $X2=0.73 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%X 1 2 10 13 14 20 26
c26 26 0 1.31739e-19 $X=2.832 $Y=1.58
r27 18 28 0.0464496 $w=5.13e-07 $l=2e-09 $layer=LI1_cond $X=2.832 $Y=1.837
+ $X2=2.832 $Y2=1.835
r28 18 20 0.766419 $w=5.13e-07 $l=3.3e-08 $layer=LI1_cond $X=2.832 $Y=1.837
+ $X2=2.832 $Y2=1.87
r29 13 28 0.557396 $w=5.13e-07 $l=2.4e-08 $layer=LI1_cond $X=2.832 $Y=1.811
+ $X2=2.832 $Y2=1.835
r30 13 26 6.82416 $w=5.13e-07 $l=2.31e-07 $layer=LI1_cond $X=2.832 $Y=1.811
+ $X2=2.832 $Y2=1.58
r31 13 14 7.29259 $w=5.13e-07 $l=3.14e-07 $layer=LI1_cond $X=2.832 $Y=1.896
+ $X2=2.832 $Y2=2.21
r32 13 20 0.603845 $w=5.13e-07 $l=2.6e-08 $layer=LI1_cond $X=2.832 $Y=1.896
+ $X2=2.832 $Y2=1.87
r33 12 26 27.693 $w=3.33e-07 $l=8.05e-07 $layer=LI1_cond $X=2.922 $Y=0.775
+ $X2=2.922 $Y2=1.58
r34 10 12 6.86365 $w=3.93e-07 $l=2.25e-07 $layer=LI1_cond $X=2.892 $Y=0.55
+ $X2=2.892 $Y2=0.775
r35 2 28 300 $w=1.7e-07 $l=4.16233e-07 $layer=licon1_PDIFF $count=2 $X=2.635
+ $Y=1.485 $X2=2.78 $Y2=1.835
r36 1 10 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=2.645
+ $Y=0.235 $X2=2.78 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__AND2B_2%VGND 1 2 3 10 12 16 18 20 23 24 25 34 43
r40 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r41 37 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=3.45
+ $Y2=0
r42 36 37 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r43 34 42 4.24142 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=3.325 $Y=0 $X2=3.502
+ $Y2=0
r44 34 36 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=3.325 $Y=0 $X2=2.99
+ $Y2=0
r45 33 37 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.99
+ $Y2=0
r46 32 33 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r47 30 33 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r48 29 32 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r49 29 30 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r50 27 39 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.212
+ $Y2=0
r51 27 29 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0 $X2=0.69
+ $Y2=0
r52 25 30 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r53 25 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r54 23 32 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.07
+ $Y2=0
r55 23 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.105 $Y=0 $X2=2.29
+ $Y2=0
r56 22 36 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.99
+ $Y2=0
r57 22 24 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=2.475 $Y=0 $X2=2.29
+ $Y2=0
r58 18 42 3.04328 $w=2.7e-07 $l=1.03899e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.502 $Y2=0
r59 18 20 19.8476 $w=2.68e-07 $l=4.65e-07 $layer=LI1_cond $X=3.46 $Y=0.085
+ $X2=3.46 $Y2=0.55
r60 14 24 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r61 14 16 11.9916 $w=3.68e-07 $l=3.85e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.47
r62 10 39 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r63 10 12 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.445
r64 3 20 182 $w=1.7e-07 $l=3.76497e-07 $layer=licon1_NDIFF $count=1 $X=3.275
+ $Y=0.235 $X2=3.41 $Y2=0.55
r65 2 16 182 $w=1.7e-07 $l=3.21559e-07 $layer=licon1_NDIFF $count=1 $X=2.105
+ $Y=0.235 $X2=2.31 $Y2=0.47
r66 1 12 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.445
.ends

