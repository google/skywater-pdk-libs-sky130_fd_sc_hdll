* File: sky130_fd_sc_hdll__dlrtn_2.pex.spice
* Created: Wed Sep  2 08:29:18 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%GATE_N 4 5 7 8 10 13 19 22 24
c39 19 0 2.42713e-19 $X=0.23 $Y=1.19
c40 13 0 3.98209e-20 $X=0.52 $Y=0.805
r41 22 25 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.4
r42 22 24 39.7811 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=0.3 $Y=1.235
+ $X2=0.3 $Y2=1.07
r43 19 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.3
+ $Y=1.235 $X2=0.3 $Y2=1.235
r44 8 13 2.83073 $w=1.5e-07 $l=7.5e-08 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.805
r45 8 10 91.58 $w=1.5e-07 $l=2.85e-07 $layer=POLY_cond $X=0.52 $Y=0.73 $X2=0.52
+ $Y2=0.445
r46 5 7 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.495 $Y=1.74
+ $X2=0.495 $Y2=2.135
r47 4 5 84.6064 $w=1.5e-07 $l=1.65e-07 $layer=POLY_cond $X=0.33 $Y=1.665
+ $X2=0.495 $Y2=1.665
r48 4 25 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=1.59 $X2=0.33
+ $Y2=1.4
r49 1 13 97.4255 $w=1.5e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.805
+ $X2=0.52 $Y2=0.805
r50 1 24 59.9997 $w=2.1e-07 $l=1.9e-07 $layer=POLY_cond $X=0.33 $Y=0.88 $X2=0.33
+ $Y2=1.07
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%A_27_363# 1 2 9 13 15 18 20 22 23 28 30 31
+ 32 36 37 39 42 44 45 48 50 52 53 59 60 64
c161 59 0 1.0603e-19 $X=3.365 $Y=1.87
c162 52 0 2.45073e-19 $X=3.22 $Y=1.87
c163 50 0 1.14507e-19 $X=3.21 $Y=0.915
c164 48 0 2.17725e-19 $X=2.945 $Y=0.9
c165 42 0 1.26282e-19 $X=3.21 $Y=1.575
c166 23 0 1.93796e-19 $X=0.965 $Y=1.59
c167 20 0 8.68433e-20 $X=3.42 $Y=1.99
c168 13 0 2.2873e-20 $X=0.965 $Y=1.74
c169 9 0 2.60437e-20 $X=0.94 $Y=0.445
r170 60 72 4.25306 $w=4.18e-07 $l=1.55e-07 $layer=LI1_cond $X=3.365 $Y=1.785
+ $X2=3.21 $Y2=1.785
r171 60 69 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.425
+ $Y=1.74 $X2=3.425 $Y2=1.74
r172 59 60 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.365 $Y=1.87
+ $X2=3.365 $Y2=1.87
r173 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.72 $Y=1.87
+ $X2=0.72 $Y2=1.87
r174 53 55 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=0.865 $Y=1.87
+ $X2=0.72 $Y2=1.87
r175 52 59 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=3.365 $Y2=1.87
r176 52 53 2.9146 $w=1.4e-07 $l=2.355e-06 $layer=MET1_cond $X=3.22 $Y=1.87
+ $X2=0.865 $Y2=1.87
r177 47 50 8.48326 $w=3.58e-07 $l=2.65e-07 $layer=LI1_cond $X=2.945 $Y=0.915
+ $X2=3.21 $Y2=0.915
r178 47 48 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.945
+ $Y=0.9 $X2=2.945 $Y2=0.9
r179 42 72 6.07598 $w=1.7e-07 $l=2.1e-07 $layer=LI1_cond $X=3.21 $Y=1.575
+ $X2=3.21 $Y2=1.785
r180 41 50 5.14255 $w=1.7e-07 $l=1.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=0.915
r181 41 42 31.3155 $w=1.68e-07 $l=4.8e-07 $layer=LI1_cond $X=3.21 $Y=1.095
+ $X2=3.21 $Y2=1.575
r182 40 64 28.8826 $w=2.7e-07 $l=1.3e-07 $layer=POLY_cond $X=0.81 $Y=1.235
+ $X2=0.94 $Y2=1.235
r183 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.81
+ $Y=1.235 $X2=0.81 $Y2=1.235
r184 37 56 2.74877 $w=2.9e-07 $l=8.5e-08 $layer=LI1_cond $X=0.75 $Y=1.795
+ $X2=0.75 $Y2=1.88
r185 37 39 22.2541 $w=2.88e-07 $l=5.6e-07 $layer=LI1_cond $X=0.75 $Y=1.795
+ $X2=0.75 $Y2=1.235
r186 36 45 7.71909 $w=2.88e-07 $l=1.45e-07 $layer=LI1_cond $X=0.75 $Y=1.215
+ $X2=0.75 $Y2=1.07
r187 36 39 0.794788 $w=2.88e-07 $l=2e-08 $layer=LI1_cond $X=0.75 $Y=1.215
+ $X2=0.75 $Y2=1.235
r188 34 45 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.69 $Y=0.805
+ $X2=0.69 $Y2=1.07
r189 33 44 4.90781 $w=1.7e-07 $l=1.55e-07 $layer=LI1_cond $X=0.395 $Y=1.88
+ $X2=0.24 $Y2=1.88
r190 32 56 4.68908 $w=1.7e-07 $l=1.45e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.75 $Y2=1.88
r191 32 33 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=1.88
+ $X2=0.395 $Y2=1.88
r192 30 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.69 $Y2=0.805
r193 30 31 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=0.605 $Y=0.72
+ $X2=0.395 $Y2=0.72
r194 26 31 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.395 $Y2=0.72
r195 26 28 12.3957 $w=1.68e-07 $l=1.9e-07 $layer=LI1_cond $X=0.31 $Y=0.635
+ $X2=0.31 $Y2=0.445
r196 20 69 48.3784 $w=2.91e-07 $l=2.52488e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.425 $Y2=1.74
r197 20 22 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.42 $Y=1.99
+ $X2=3.42 $Y2=2.275
r198 16 48 46.2115 $w=3.3e-07 $l=1.65e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.9
r199 16 18 164.085 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.945 $Y=0.735
+ $X2=2.945 $Y2=0.415
r200 13 23 60.4563 $w=1.8e-07 $l=1.5e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=1.59
r201 13 15 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=0.965 $Y=1.74
+ $X2=0.965 $Y2=2.135
r202 11 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.235
r203 11 23 112.809 $w=1.5e-07 $l=2.2e-07 $layer=POLY_cond $X=0.94 $Y=1.37
+ $X2=0.94 $Y2=1.59
r204 7 64 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=0.94 $Y=1.1
+ $X2=0.94 $Y2=1.235
r205 7 9 335.862 $w=1.5e-07 $l=6.55e-07 $layer=POLY_cond $X=0.94 $Y=1.1 $X2=0.94
+ $Y2=0.445
r206 2 44 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.815 $X2=0.26 $Y2=1.96
r207 1 28 182 $w=1.7e-07 $l=2.65236e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%D 2 3 5 8 10 11 12
c45 12 0 5.01492e-20 $X=1.61 $Y=1.19
c46 2 0 1.74491e-19 $X=1.955 $Y=1.67
r47 12 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.6
+ $Y=1.16 $X2=1.6 $Y2=1.16
r48 10 15 44.5896 $w=3.3e-07 $l=2.55e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.6 $Y2=1.16
r49 10 11 3.18546 $w=3.3e-07 $l=1e-07 $layer=POLY_cond $X=1.855 $Y=1.16
+ $X2=1.955 $Y2=1.16
r50 6 11 33.332 $w=1.75e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.955 $Y2=1.16
r51 6 8 282.021 $w=1.5e-07 $l=5.5e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.445
r52 3 5 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=1.955 $Y=1.77
+ $X2=1.955 $Y2=2.165
r53 2 3 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=1.955 $Y=1.67 $X2=1.955
+ $Y2=1.77
r54 1 11 33.332 $w=1.75e-07 $l=1.65e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.16
r55 1 2 114.394 $w=2e-07 $l=3.45e-07 $layer=POLY_cond $X=1.955 $Y=1.325
+ $X2=1.955 $Y2=1.67
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%A_319_369# 1 2 8 9 11 14 17 20 23 27 30 32
c78 32 0 1.14507e-19 $X=2.4 $Y=0.765
c79 30 0 1.2579e-19 $X=2.4 $Y=0.93
c80 17 0 1.74491e-19 $X=1.72 $Y=1.99
r81 30 33 40.8147 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=1.095
r82 30 32 48.4159 $w=2.7e-07 $l=1.65e-07 $layer=POLY_cond $X=2.4 $Y=0.93 $X2=2.4
+ $Y2=0.765
r83 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.4
+ $Y=0.93 $X2=2.4 $Y2=0.93
r84 27 29 12.2997 $w=3.67e-07 $l=4.63249e-07 $layer=LI1_cond $X=2.03 $Y=0.72
+ $X2=2.4 $Y2=0.93
r85 26 27 8.64305 $w=3.67e-07 $l=2.6e-07 $layer=LI1_cond $X=1.77 $Y=0.72
+ $X2=2.03 $Y2=0.72
r86 20 23 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.03 $Y=1.495
+ $X2=2.03 $Y2=1.58
r87 19 27 5.25812 $w=1.7e-07 $l=3.75e-07 $layer=LI1_cond $X=2.03 $Y=1.095
+ $X2=2.03 $Y2=0.72
r88 19 20 26.0963 $w=1.68e-07 $l=4e-07 $layer=LI1_cond $X=2.03 $Y=1.095 $X2=2.03
+ $Y2=1.495
r89 15 23 20.2246 $w=1.68e-07 $l=3.1e-07 $layer=LI1_cond $X=1.72 $Y=1.58
+ $X2=2.03 $Y2=1.58
r90 15 17 11.3498 $w=3.28e-07 $l=3.25e-07 $layer=LI1_cond $X=1.72 $Y=1.665
+ $X2=1.72 $Y2=1.99
r91 14 32 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.425 $Y=0.445
+ $X2=2.425 $Y2=0.765
r92 9 11 105.772 $w=1.8e-07 $l=3.95e-07 $layer=POLY_cond $X=2.425 $Y=1.77
+ $X2=2.425 $Y2=2.165
r93 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.425 $Y=1.67 $X2=2.425
+ $Y2=1.77
r94 8 33 190.657 $w=2e-07 $l=5.75e-07 $layer=POLY_cond $X=2.425 $Y=1.67
+ $X2=2.425 $Y2=1.095
r95 2 17 300 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_PDIFF $count=2 $X=1.595
+ $Y=1.845 $X2=1.72 $Y2=1.99
r96 1 26 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=1.645
+ $Y=0.235 $X2=1.77 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%A_203_47# 1 2 8 9 11 12 16 20 24 26 27 30
+ 33 36 40
c114 40 0 3.47682e-19 $X=2.87 $Y=1.44
c115 9 0 1.43299e-19 $X=2.95 $Y=1.99
c116 2 0 1.13552e-19 $X=1.055 $Y=1.815
r117 39 41 43.3814 $w=3.15e-07 $l=1.95e-07 $layer=POLY_cond $X=2.892 $Y=1.44
+ $X2=2.892 $Y2=1.635
r118 39 40 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.87
+ $Y=1.44 $X2=2.87 $Y2=1.44
r119 36 39 21.9826 $w=3.15e-07 $l=1.2e-07 $layer=POLY_cond $X=2.892 $Y=1.32
+ $X2=2.892 $Y2=1.44
r120 33 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.81 $Y=1.53
+ $X2=2.81 $Y2=1.53
r121 30 46 5.20126 $w=2.68e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=1.53 $X2=1.2
+ $Y2=1.445
r122 29 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.18 $Y=1.53
+ $X2=1.18 $Y2=1.53
r123 27 29 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.325 $Y=1.53
+ $X2=1.18 $Y2=1.53
r124 26 33 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=2.81 $Y2=1.53
r125 26 27 1.65841 $w=1.4e-07 $l=1.34e-06 $layer=MET1_cond $X=2.665 $Y=1.53
+ $X2=1.325 $Y2=1.53
r126 22 30 2.13415 $w=2.68e-07 $l=5e-08 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.2
+ $Y2=1.53
r127 22 24 16.2196 $w=2.68e-07 $l=3.8e-07 $layer=LI1_cond $X=1.2 $Y=1.58 $X2=1.2
+ $Y2=1.96
r128 20 46 65.2406 $w=1.68e-07 $l=1e-06 $layer=LI1_cond $X=1.15 $Y=0.445
+ $X2=1.15 $Y2=1.445
r129 14 16 410.213 $w=1.5e-07 $l=8e-07 $layer=POLY_cond $X=3.465 $Y=1.245
+ $X2=3.465 $Y2=0.445
r130 13 36 20.1192 $w=1.5e-07 $l=1.58e-07 $layer=POLY_cond $X=3.05 $Y=1.32
+ $X2=2.892 $Y2=1.32
r131 12 14 26.9307 $w=1.5e-07 $l=1.06066e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.465 $Y2=1.245
r132 12 13 174.34 $w=1.5e-07 $l=3.4e-07 $layer=POLY_cond $X=3.39 $Y=1.32
+ $X2=3.05 $Y2=1.32
r133 9 11 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.95 $Y=1.99
+ $X2=2.95 $Y2=2.275
r134 8 9 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.99
r135 8 41 84.5522 $w=2e-07 $l=2.55e-07 $layer=POLY_cond $X=2.95 $Y=1.89 $X2=2.95
+ $Y2=1.635
r136 2 24 300 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.815 $X2=1.2 $Y2=1.96
r137 1 20 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.15 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%A_750_21# 1 2 9 11 13 14 16 17 19 20 22 23
+ 25 26 33 36 39 41 44 45 50 54 61
c120 61 0 1.07771e-19 $X=6.19 $Y=1.202
c121 9 0 1.26282e-19 $X=3.825 $Y=0.445
r122 61 62 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=6.19 $Y=1.202
+ $X2=6.215 $Y2=1.202
r123 60 61 53.6976 $w=3.77e-07 $l=4.2e-07 $layer=POLY_cond $X=5.77 $Y=1.202
+ $X2=6.19 $Y2=1.202
r124 59 60 3.19629 $w=3.77e-07 $l=2.5e-08 $layer=POLY_cond $X=5.745 $Y=1.202
+ $X2=5.77 $Y2=1.202
r125 55 59 1.91777 $w=3.77e-07 $l=1.5e-08 $layer=POLY_cond $X=5.73 $Y=1.202
+ $X2=5.745 $Y2=1.202
r126 54 55 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.73
+ $Y=1.16 $X2=5.73 $Y2=1.16
r127 51 54 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=5.64 $Y=1.16 $X2=5.73
+ $Y2=1.16
r128 49 50 7.23989 $w=3.28e-07 $l=1.3e-07 $layer=LI1_cond $X=5.04 $Y=1.7
+ $X2=5.17 $Y2=1.7
r129 47 49 0.453993 $w=3.28e-07 $l=1.3e-08 $layer=LI1_cond $X=5.027 $Y=1.7
+ $X2=5.04 $Y2=1.7
r130 46 47 13.6896 $w=3.28e-07 $l=3.92e-07 $layer=LI1_cond $X=4.635 $Y=1.7
+ $X2=5.027 $Y2=1.7
r131 43 51 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.64 $Y2=1.16
r132 43 44 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=5.64 $Y=1.325
+ $X2=5.64 $Y2=1.535
r133 41 44 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.64 $Y2=1.535
r134 41 50 25.1176 $w=1.68e-07 $l=3.85e-07 $layer=LI1_cond $X=5.555 $Y=1.62
+ $X2=5.17 $Y2=1.62
r135 37 47 1.61437 $w=2.85e-07 $l=1.65e-07 $layer=LI1_cond $X=5.027 $Y=1.865
+ $X2=5.027 $Y2=1.7
r136 37 39 3.84148 $w=2.83e-07 $l=9.5e-08 $layer=LI1_cond $X=5.027 $Y=1.865
+ $X2=5.027 $Y2=1.96
r137 36 46 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=1.7
r138 36 45 46.3209 $w=1.68e-07 $l=7.1e-07 $layer=LI1_cond $X=4.635 $Y=1.535
+ $X2=4.635 $Y2=0.825
r139 31 45 7.25185 $w=3.28e-07 $l=1.65e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.825
r140 31 33 9.7783 $w=3.28e-07 $l=2.8e-07 $layer=LI1_cond $X=4.62 $Y=0.66
+ $X2=4.62 $Y2=0.38
r141 28 29 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.105
+ $Y=1.7 $X2=4.105 $Y2=1.7
r142 26 46 2.96841 $w=3.28e-07 $l=8.5e-08 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.635 $Y2=1.7
r143 26 28 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=4.55 $Y=1.7
+ $X2=4.105 $Y2=1.7
r144 23 62 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.202
r145 23 25 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=6.215 $Y=1.41
+ $X2=6.215 $Y2=1.985
r146 20 61 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=1.202
r147 20 22 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=6.19 $Y=0.995
+ $X2=6.19 $Y2=0.56
r148 17 60 24.4204 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=1.202
r149 17 19 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.77 $Y=0.995
+ $X2=5.77 $Y2=0.56
r150 14 59 20.0566 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.202
r151 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.745 $Y=1.41
+ $X2=5.745 $Y2=1.985
r152 11 29 53.3563 $w=3.12e-07 $l=3.38452e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=4.005 $Y2=1.7
r153 11 13 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=3.9 $Y=1.99
+ $X2=3.9 $Y2=2.275
r154 7 29 78.6992 $w=3.12e-07 $l=5.07075e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=4.005 $Y2=1.7
r155 7 9 425.596 $w=1.5e-07 $l=8.3e-07 $layer=POLY_cond $X=3.825 $Y=1.275
+ $X2=3.825 $Y2=0.445
r156 2 49 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=1.62
r157 2 39 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.895
+ $Y=1.485 $X2=5.04 $Y2=1.96
r158 1 33 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=4.495
+ $Y=0.235 $X2=4.62 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%A_604_47# 1 2 7 9 11 14 16 18 22 27 29 30
+ 32 33
c93 30 0 2.92347e-19 $X=3.85 $Y=1.16
c94 29 0 1.43299e-19 $X=3.765 $Y=2.165
r95 35 36 9.46122 $w=2.45e-07 $l=1.9e-07 $layer=LI1_cond $X=3.575 $Y=1.16
+ $X2=3.765 $Y2=1.16
r96 33 39 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=4.295 $Y=1.16
+ $X2=4.295 $Y2=1.25
r97 32 33 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.295
+ $Y=1.16 $X2=4.295 $Y2=1.16
r98 30 36 3.97745 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=3.765 $Y2=1.16
r99 30 32 15.5405 $w=3.28e-07 $l=4.45e-07 $layer=LI1_cond $X=3.85 $Y=1.16
+ $X2=4.295 $Y2=1.16
r100 28 36 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=1.16
r101 28 29 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=3.765 $Y=1.325
+ $X2=3.765 $Y2=2.165
r102 27 35 2.87745 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.575 $Y=0.995
+ $X2=3.575 $Y2=1.16
r103 26 27 28.0535 $w=1.68e-07 $l=4.3e-07 $layer=LI1_cond $X=3.575 $Y=0.565
+ $X2=3.575 $Y2=0.995
r104 22 26 7.39867 $w=2.85e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.575 $Y2=0.565
r105 22 24 11.5244 $w=2.83e-07 $l=2.85e-07 $layer=LI1_cond $X=3.49 $Y=0.422
+ $X2=3.205 $Y2=0.422
r106 18 29 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.765 $Y2=2.165
r107 18 20 25.93 $w=2.18e-07 $l=4.95e-07 $layer=LI1_cond $X=3.68 $Y=2.275
+ $X2=3.185 $Y2=2.275
r108 16 17 29.1618 $w=2e-07 $l=7.5e-08 $layer=POLY_cond $X=4.805 $Y=1.25
+ $X2=4.805 $Y2=1.175
r109 14 17 315.351 $w=1.5e-07 $l=6.15e-07 $layer=POLY_cond $X=4.83 $Y=0.56
+ $X2=4.83 $Y2=1.175
r110 9 16 53.8601 $w=2e-07 $l=1.6e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.25
r111 9 11 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.805 $Y=1.41
+ $X2=4.805 $Y2=1.985
r112 8 39 16.5046 $w=1.5e-07 $l=1.35e-07 $layer=POLY_cond $X=4.43 $Y=1.25
+ $X2=4.295 $Y2=1.25
r113 7 16 9.57678 $w=1.5e-07 $l=1e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.805 $Y2=1.25
r114 7 8 141.011 $w=1.5e-07 $l=2.75e-07 $layer=POLY_cond $X=4.705 $Y=1.25
+ $X2=4.43 $Y2=1.25
r115 2 20 600 $w=1.7e-07 $l=2.73038e-07 $layer=licon1_PDIFF $count=1 $X=3.04
+ $Y=2.065 $X2=3.185 $Y2=2.275
r116 1 24 182 $w=1.7e-07 $l=2.8801e-07 $layer=licon1_NDIFF $count=1 $X=3.02
+ $Y=0.235 $X2=3.205 $Y2=0.445
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%RESET_B 1 3 4 6 7
r33 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.25
+ $Y=1.16 $X2=5.25 $Y2=1.16
r34 4 10 51.486 $w=2.55e-07 $l=2.62202e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.25 $Y2=1.16
r35 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.275 $Y=1.41
+ $X2=5.275 $Y2=1.985
r36 1 10 39.2931 $w=2.55e-07 $l=1.72337e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.25 $Y2=1.16
r37 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%VPWR 1 2 3 4 5 18 22 27 30 35 39 40 42 43
+ 44 46 51 56 72 73 76 79 82
c103 35 0 1.07771e-19 $X=5.51 $Y=1.97
c104 18 0 1.31521e-19 $X=0.73 $Y=2.22
r105 79 80 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r106 76 77 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r107 72 73 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=2.72
+ $X2=6.67 $Y2=2.72
r108 70 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=6.67 $Y2=2.72
r109 69 70 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r110 67 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=6.21 $Y2=2.72
r111 67 86 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=4.37 $Y2=2.72
r112 66 67 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r113 64 66 42.7326 $w=1.68e-07 $l=6.55e-07 $layer=LI1_cond $X=4.635 $Y=2.72
+ $X2=5.29 $Y2=2.72
r114 63 86 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=4.37 $Y2=2.72
r115 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r116 60 63 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r117 60 80 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=2.07 $Y2=2.72
r118 59 62 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=2.72
+ $X2=3.91 $Y2=2.72
r119 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r120 57 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.19 $Y2=2.72
r121 57 59 13.3743 $w=1.68e-07 $l=2.05e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.53 $Y2=2.72
r122 56 64 8.15384 $w=1.7e-07 $l=2.93e-07 $layer=LI1_cond $X=4.342 $Y=2.72
+ $X2=4.635 $Y2=2.72
r123 56 86 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r124 56 82 8.58723 $w=5.83e-07 $l=4.2e-07 $layer=LI1_cond $X=4.342 $Y=2.72
+ $X2=4.342 $Y2=2.3
r125 56 62 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=4.05 $Y=2.72
+ $X2=3.91 $Y2=2.72
r126 55 80 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r127 55 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r128 54 55 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r129 52 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.73 $Y2=2.72
r130 52 54 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r131 51 79 7.44763 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=2.19 $Y2=2.72
r132 51 54 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=2.055 $Y=2.72
+ $X2=1.15 $Y2=2.72
r133 46 76 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.73 $Y2=2.72
r134 46 48 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=2.72
+ $X2=0.23 $Y2=2.72
r135 44 77 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r136 44 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r137 42 69 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=2.72
+ $X2=6.21 $Y2=2.72
r138 42 43 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=6.375 $Y=2.72
+ $X2=6.477 $Y2=2.72
r139 41 72 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=6.58 $Y=2.72 $X2=6.67
+ $Y2=2.72
r140 41 43 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=6.58 $Y=2.72
+ $X2=6.477 $Y2=2.72
r141 39 66 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.29 $Y2=2.72
r142 39 40 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.345 $Y=2.72
+ $X2=5.495 $Y2=2.72
r143 38 69 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=6.21 $Y2=2.72
r144 38 40 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=5.645 $Y=2.72
+ $X2=5.495 $Y2=2.72
r145 35 37 6.40424 $w=3.28e-07 $l=1.8e-07 $layer=LI1_cond $X=5.51 $Y=1.97
+ $X2=5.51 $Y2=2.15
r146 30 33 36.7894 $w=2.03e-07 $l=6.8e-07 $layer=LI1_cond $X=6.477 $Y=1.66
+ $X2=6.477 $Y2=2.34
r147 28 43 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=6.477 $Y=2.635
+ $X2=6.477 $Y2=2.72
r148 28 33 15.9601 $w=2.03e-07 $l=2.95e-07 $layer=LI1_cond $X=6.477 $Y=2.635
+ $X2=6.477 $Y2=2.34
r149 27 37 7.29881 $w=2.98e-07 $l=1.9e-07 $layer=LI1_cond $X=5.495 $Y=2.34
+ $X2=5.495 $Y2=2.15
r150 25 40 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.72
r151 25 27 11.3324 $w=2.98e-07 $l=2.95e-07 $layer=LI1_cond $X=5.495 $Y=2.635
+ $X2=5.495 $Y2=2.34
r152 20 79 0.256868 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2.72
r153 20 22 27.1038 $w=2.68e-07 $l=6.35e-07 $layer=LI1_cond $X=2.19 $Y=2.635
+ $X2=2.19 $Y2=2
r154 16 76 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.72
r155 16 18 14.4928 $w=3.28e-07 $l=4.15e-07 $layer=LI1_cond $X=0.73 $Y=2.635
+ $X2=0.73 $Y2=2.22
r156 5 33 400 $w=1.7e-07 $l=9.29274e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.485 $X2=6.46 $Y2=2.34
r157 5 30 400 $w=1.7e-07 $l=2.40312e-07 $layer=licon1_PDIFF $count=1 $X=6.305
+ $Y=1.485 $X2=6.46 $Y2=1.66
r158 4 35 600 $w=1.7e-07 $l=5.52766e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=1.97
r159 4 27 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.365
+ $Y=1.485 $X2=5.51 $Y2=2.34
r160 3 82 300 $w=1.7e-07 $l=6.62156e-07 $layer=licon1_PDIFF $count=2 $X=3.99
+ $Y=2.065 $X2=4.545 $Y2=2.3
r161 2 22 300 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=2 $X=2.045
+ $Y=1.845 $X2=2.19 $Y2=2
r162 1 18 600 $w=1.7e-07 $l=4.71964e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.815 $X2=0.73 $Y2=2.22
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%Q 1 2 7 10 16 20 23 24 27
r35 24 29 7.78328 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=1.19
+ $X2=6.235 $Y2=1.325
r36 24 27 7.78328 $w=3.98e-07 $l=1.35e-07 $layer=LI1_cond $X=6.235 $Y=1.19
+ $X2=6.235 $Y2=1.055
r37 23 29 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=6.12 $Y=1.495
+ $X2=6.12 $Y2=1.325
r38 20 21 3.0294 $w=3.88e-07 $l=8.5e-08 $layer=LI1_cond $X=6.01 $Y=2.34 $X2=6.01
+ $Y2=2.255
r39 18 27 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=6.12 $Y=0.825
+ $X2=6.12 $Y2=1.055
r40 16 18 16.8816 $w=3.88e-07 $l=4.45e-07 $layer=LI1_cond $X=6.01 $Y=0.38
+ $X2=6.01 $Y2=0.825
r41 10 21 22.1195 $w=3.08e-07 $l=5.95e-07 $layer=LI1_cond $X=6.05 $Y=1.66
+ $X2=6.05 $Y2=2.255
r42 7 23 8.09553 $w=3.08e-07 $l=1.55e-07 $layer=LI1_cond $X=6.05 $Y=1.65
+ $X2=6.05 $Y2=1.495
r43 7 10 0.371756 $w=3.08e-07 $l=1e-08 $layer=LI1_cond $X=6.05 $Y=1.65 $X2=6.05
+ $Y2=1.66
r44 2 20 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=2.34
r45 2 10 300 $w=1.7e-07 $l=2.36643e-07 $layer=licon1_PDIFF $count=2 $X=5.835
+ $Y=1.485 $X2=5.98 $Y2=1.66
r46 1 16 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=5.845
+ $Y=0.235 $X2=5.98 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__DLRTN_2%VGND 1 2 3 4 5 18 22 26 30 34 37 38 40 41
+ 42 44 49 54 70 71 74 77 80
c98 71 0 3.98209e-20 $X=6.67 $Y=0
r99 80 81 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r100 77 78 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r101 74 75 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r102 70 71 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.67 $Y=0 $X2=6.67
+ $Y2=0
r103 68 71 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=0 $X2=6.67
+ $Y2=0
r104 67 68 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r105 65 68 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=5.29 $Y=0 $X2=6.21
+ $Y2=0
r106 64 65 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r107 62 65 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r108 62 81 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=0 $X2=3.91
+ $Y2=0
r109 61 64 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=4.37 $Y=0 $X2=5.29
+ $Y2=0
r110 61 62 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=4.37 $Y=0 $X2=4.37
+ $Y2=0
r111 59 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.035
+ $Y2=0
r112 59 61 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=4.2 $Y=0 $X2=4.37
+ $Y2=0
r113 58 81 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0
+ $X2=3.91 $Y2=0
r114 58 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r115 57 58 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r116 55 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.355 $Y=0 $X2=2.19
+ $Y2=0
r117 55 57 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.355 $Y=0
+ $X2=2.53 $Y2=0
r118 54 80 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.87 $Y=0 $X2=4.035
+ $Y2=0
r119 54 57 87.4225 $w=1.68e-07 $l=1.34e-06 $layer=LI1_cond $X=3.87 $Y=0 $X2=2.53
+ $Y2=0
r120 53 78 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r121 53 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r122 52 53 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r123 50 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.895 $Y=0 $X2=0.73
+ $Y2=0
r124 50 52 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=0
+ $X2=1.15 $Y2=0
r125 49 77 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.025 $Y=0 $X2=2.19
+ $Y2=0
r126 49 52 57.0856 $w=1.68e-07 $l=8.75e-07 $layer=LI1_cond $X=2.025 $Y=0
+ $X2=1.15 $Y2=0
r127 44 74 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.565 $Y=0 $X2=0.73
+ $Y2=0
r128 44 46 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.565 $Y=0
+ $X2=0.23 $Y2=0
r129 42 75 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r130 42 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r131 40 67 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=6.375 $Y=0
+ $X2=6.21 $Y2=0
r132 40 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.375 $Y=0 $X2=6.48
+ $Y2=0
r133 39 70 5.54545 $w=1.68e-07 $l=8.5e-08 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.67
+ $Y2=0
r134 39 41 6.13603 $w=1.7e-07 $l=1.05e-07 $layer=LI1_cond $X=6.585 $Y=0 $X2=6.48
+ $Y2=0
r135 37 64 1.63102 $w=1.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.29
+ $Y2=0
r136 37 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.315 $Y=0 $X2=5.48
+ $Y2=0
r137 36 67 36.861 $w=1.68e-07 $l=5.65e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=6.21
+ $Y2=0
r138 36 38 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=5.645 $Y=0 $X2=5.48
+ $Y2=0
r139 32 41 0.593901 $w=2.1e-07 $l=8.5e-08 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.48 $Y2=0
r140 32 34 15.5801 $w=2.08e-07 $l=2.95e-07 $layer=LI1_cond $X=6.48 $Y=0.085
+ $X2=6.48 $Y2=0.38
r141 28 38 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0
r142 28 30 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=5.48 $Y=0.085
+ $X2=5.48 $Y2=0.38
r143 24 80 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0
r144 24 26 12.5721 $w=3.28e-07 $l=3.6e-07 $layer=LI1_cond $X=4.035 $Y=0.085
+ $X2=4.035 $Y2=0.445
r145 20 77 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0
r146 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.19 $Y=0.085
+ $X2=2.19 $Y2=0.36
r147 16 74 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r148 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r149 5 34 91 $w=1.7e-07 $l=2.57488e-07 $layer=licon1_NDIFF $count=2 $X=6.265
+ $Y=0.235 $X2=6.46 $Y2=0.38
r150 4 30 91 $w=1.7e-07 $l=2.31409e-07 $layer=licon1_NDIFF $count=2 $X=5.31
+ $Y=0.235 $X2=5.48 $Y2=0.38
r151 3 26 182 $w=1.7e-07 $l=2.69165e-07 $layer=licon1_NDIFF $count=1 $X=3.9
+ $Y=0.235 $X2=4.035 $Y2=0.445
r152 2 22 182 $w=1.7e-07 $l=1.8735e-07 $layer=licon1_NDIFF $count=1 $X=2.055
+ $Y=0.235 $X2=2.19 $Y2=0.36
r153 1 18 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

