* File: sky130_fd_sc_hdll__nand4bb_1.spice
* Created: Thu Aug 27 19:15:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand4bb_1.pex.spice"
.subckt sky130_fd_sc_hdll__nand4bb_1  VNB VPB B_N D C A_N VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1011 N_VGND_M1011_d N_B_N_M1011_g N_A_27_93#_M1011_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0894953 AS=0.1092 PD=0.820374 PS=1.36 NRD=45.156 NRS=0 M=1 R=2.8
+ SA=75000.2 SB=75002.3 A=0.063 P=1.14 MULT=1
MM1007 A_218_47# N_D_M1007_g N_VGND_M1011_d VNB NSHORT L=0.15 W=0.65 AD=0.13975
+ AS=0.138505 PD=1.08 PS=1.26963 NRD=29.532 NRS=0.912 M=1 R=4.33333 SA=75000.5
+ SB=75001.8 A=0.0975 P=1.6 MULT=1
MM1004 A_334_47# N_C_M1004_g A_218_47# VNB NSHORT L=0.15 W=0.65 AD=0.11375
+ AS=0.13975 PD=1 PS=1.08 NRD=22.152 NRS=29.532 M=1 R=4.33333 SA=75001.1
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1002 A_434_47# N_A_27_93#_M1002_g A_334_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.11375 PD=0.98 PS=1 NRD=20.304 NRS=22.152 M=1 R=4.33333
+ SA=75001.6 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1006 N_Y_M1006_d N_A_500_21#_M1006_g A_434_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.10725 PD=1.92 PS=0.98 NRD=8.304 NRS=20.304 M=1 R=4.33333
+ SA=75002.1 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_500_21#_M1010_d N_A_N_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1533 AS=0.1092 PD=1.57 PS=1.36 NRD=27.132 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.3 A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_B_N_M1000_g N_A_27_93#_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0933761 AS=0.1134 PD=0.807465 PS=1.38 NRD=34.0022 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90003.3 A=0.0756 P=1.2 MULT=1
MM1003 N_Y_M1003_d N_D_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.2
+ AS=0.222324 PD=1.4 PS=1.92254 NRD=9.8303 NRS=2.9353 M=1 R=5.55556 SA=90000.4
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1005_d N_C_M1005_g N_Y_M1003_d VPB PHIGHVT L=0.18 W=1 AD=0.16
+ AS=0.2 PD=1.32 PS=1.4 NRD=1.9503 NRS=13.7703 M=1 R=5.55556 SA=90001 SB=90001.6
+ A=0.18 P=2.36 MULT=1
MM1009 N_Y_M1009_d N_A_27_93#_M1009_g N_VPWR_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.16 PD=1.3 PS=1.32 NRD=0.9653 NRS=5.8903 M=1 R=5.55556 SA=90001.5
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_500_21#_M1001_g N_Y_M1009_d VPB PHIGHVT L=0.18 W=1
+ AD=0.349859 AS=0.15 PD=2.5493 PS=1.3 NRD=0.9653 NRS=2.9353 M=1 R=5.55556
+ SA=90002 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1008 N_A_500_21#_M1008_d N_A_N_M1008_g N_VPWR_M1001_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1365 AS=0.146941 PD=1.49 PS=1.0707 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90003.3 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
*
.include "sky130_fd_sc_hdll__nand4bb_1.pxi.spice"
*
.ends
*
*
