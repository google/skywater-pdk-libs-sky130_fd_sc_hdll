# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21o_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__a21o_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.865000 1.055000 1.535000 1.290000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.055000 0.695000 1.290000 ;
        RECT 0.525000 1.290000 0.695000 1.460000 ;
        RECT 0.525000 1.460000 1.875000 1.630000 ;
        RECT 1.705000 1.055000 2.045000 1.290000 ;
        RECT 1.705000 1.290000 1.875000 1.460000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.865000 1.055000 3.195000 1.615000 ;
    END
  END B1
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 8.010000 2.910000 ;
    END
  END VPB
  PIN X
    ANTENNADIFFAREA  1.862000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.905000 0.255000 4.235000 0.695000 ;
        RECT 3.905000 0.695000 7.055000 0.865000 ;
        RECT 3.935000 1.445000 7.025000 1.615000 ;
        RECT 3.935000 1.615000 4.205000 2.465000 ;
        RECT 4.845000 0.255000 5.175000 0.695000 ;
        RECT 4.875000 1.615000 5.145000 2.465000 ;
        RECT 5.785000 0.255000 6.115000 0.695000 ;
        RECT 5.815000 1.615000 6.085000 2.465000 ;
        RECT 6.545000 0.865000 6.795000 1.445000 ;
        RECT 6.725000 0.255000 7.055000 0.695000 ;
        RECT 6.755000 1.615000 7.025000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.820000 0.085000 ;
      RECT 0.000000  2.635000 7.820000 2.805000 ;
      RECT 0.095000  1.460000 0.355000 1.800000 ;
      RECT 0.095000  1.800000 2.275000 1.970000 ;
      RECT 0.095000  1.970000 0.425000 2.465000 ;
      RECT 0.205000  0.085000 0.535000 0.885000 ;
      RECT 0.595000  2.140000 0.865000 2.635000 ;
      RECT 1.035000  0.275000 1.365000 0.675000 ;
      RECT 1.035000  0.675000 3.735000 0.885000 ;
      RECT 1.035000  1.970000 1.365000 2.465000 ;
      RECT 1.535000  2.140000 1.805000 2.635000 ;
      RECT 1.945000  0.085000 2.275000 0.505000 ;
      RECT 1.975000  1.970000 2.275000 2.295000 ;
      RECT 1.975000  2.295000 3.245000 2.465000 ;
      RECT 2.045000  1.460000 2.275000 1.800000 ;
      RECT 2.445000  0.255000 2.745000 0.675000 ;
      RECT 2.445000  0.885000 2.695000 1.790000 ;
      RECT 2.445000  1.790000 2.745000 2.125000 ;
      RECT 2.915000  0.085000 3.735000 0.505000 ;
      RECT 2.915000  1.785000 3.245000 2.295000 ;
      RECT 3.485000  1.495000 3.735000 2.635000 ;
      RECT 3.565000  0.885000 3.735000 1.035000 ;
      RECT 3.565000  1.035000 6.135000 1.275000 ;
      RECT 4.375000  1.785000 4.705000 2.635000 ;
      RECT 4.405000  0.085000 4.675000 0.525000 ;
      RECT 5.315000  1.785000 5.645000 2.635000 ;
      RECT 5.345000  0.085000 5.615000 0.525000 ;
      RECT 6.255000  1.785000 6.585000 2.635000 ;
      RECT 6.285000  0.085000 6.555000 0.525000 ;
      RECT 7.215000  1.445000 7.525000 2.635000 ;
      RECT 7.225000  0.085000 7.475000 0.905000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21o_8
END LIBRARY
