# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o221ai_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.565000 1.075000  6.945000 1.445000 ;
        RECT 6.565000 1.445000  9.320000 1.615000 ;
        RECT 9.005000 1.075000 10.135000 1.275000 ;
        RECT 9.005000 1.275000  9.320000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.125000 1.075000 8.735000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.560000 1.075000 4.925000 1.275000 ;
        RECT 4.735000 1.275000 4.925000 1.445000 ;
        RECT 4.735000 1.445000 6.395000 1.615000 ;
        RECT 6.015000 1.075000 6.395000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.095000 0.995000 5.835000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 1.900000 1.275000 ;
    END
  END C1
  PIN VGND
    ANTENNADIFFAREA  0.767000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 10.770000 2.910000 ;
    END
  END VPB
  PIN VPWR
    ANTENNADIFFAREA  2.645000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  2.156000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.645000 2.325000 0.865000 ;
        RECT 0.625000 1.445000 4.565000 1.615000 ;
        RECT 0.625000 1.615000 0.875000 2.465000 ;
        RECT 1.565000 1.615000 2.325000 1.955000 ;
        RECT 1.565000 1.955000 1.815000 2.465000 ;
        RECT 2.120000 0.865000 2.325000 1.445000 ;
        RECT 4.345000 1.615000 4.565000 1.785000 ;
        RECT 4.345000 1.785000 8.565000 2.005000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 10.580000 0.085000 ;
      RECT  0.000000  2.635000 10.580000 2.805000 ;
      RECT  0.115000  0.255000  6.135000 0.475000 ;
      RECT  0.115000  0.475000  0.365000 0.895000 ;
      RECT  0.155000  1.485000  0.405000 2.635000 ;
      RECT  1.095000  1.825000  1.345000 2.635000 ;
      RECT  2.035000  2.125000  2.805000 2.635000 ;
      RECT  2.515000  0.645000  6.685000 0.735000 ;
      RECT  2.515000  0.735000 10.445000 0.820000 ;
      RECT  3.025000  1.785000  4.175000 1.955000 ;
      RECT  3.025000  1.955000  3.275000 2.465000 ;
      RECT  3.495000  2.125000  3.745000 2.635000 ;
      RECT  3.965000  1.955000  4.175000 2.265000 ;
      RECT  3.965000  2.265000  6.135000 2.465000 ;
      RECT  6.015000  0.820000 10.445000 0.905000 ;
      RECT  6.355000  0.255000  6.685000 0.645000 ;
      RECT  6.355000  2.175000  6.605000 2.635000 ;
      RECT  6.775000  2.265000  8.995000 2.465000 ;
      RECT  6.905000  0.085000  7.075000 0.555000 ;
      RECT  7.245000  0.255000  7.625000 0.725000 ;
      RECT  7.245000  0.725000  8.565000 0.735000 ;
      RECT  7.845000  0.085000  8.015000 0.555000 ;
      RECT  8.185000  0.255000  8.565000 0.725000 ;
      RECT  8.785000  0.085000  8.955000 0.555000 ;
      RECT  8.785000  1.785000  9.935000 1.955000 ;
      RECT  8.785000  1.955000  8.995000 2.265000 ;
      RECT  9.125000  0.255000  9.505000 0.725000 ;
      RECT  9.125000  0.725000 10.445000 0.735000 ;
      RECT  9.215000  2.125000  9.465000 2.635000 ;
      RECT  9.685000  1.445000  9.935000 1.785000 ;
      RECT  9.685000  1.955000  9.935000 2.465000 ;
      RECT  9.725000  0.085000  9.895000 0.555000 ;
      RECT 10.065000  0.255000 10.445000 0.725000 ;
      RECT 10.155000  1.445000 10.405000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221ai_4
END LIBRARY
