* File: sky130_fd_sc_hdll__o21a_4.pex.spice
* Created: Thu Aug 27 19:19:06 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O21A_4%A_80_21# 1 2 3 10 12 13 15 16 18 19 21 22
+ 24 25 27 28 30 31 33 34 41 43 46 48 49 52 54 56 61 62
c132 56 0 1.79518e-19 $X=2.44 $Y=0.762
c133 49 0 1.7149e-19 $X=2.565 $Y=1.957
c134 31 0 1.95549e-19 $X=2.31 $Y=1.41
r135 73 74 11.2865 $w=3.63e-07 $l=8.5e-08 $layer=POLY_cond $X=1.83 $Y=1.202
+ $X2=1.915 $Y2=1.202
r136 72 73 52.449 $w=3.63e-07 $l=3.95e-07 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.83 $Y2=1.202
r137 71 72 11.2865 $w=3.63e-07 $l=8.5e-08 $layer=POLY_cond $X=1.35 $Y=1.202
+ $X2=1.435 $Y2=1.202
r138 70 71 52.449 $w=3.63e-07 $l=3.95e-07 $layer=POLY_cond $X=0.955 $Y=1.202
+ $X2=1.35 $Y2=1.202
r139 69 70 11.2865 $w=3.63e-07 $l=8.5e-08 $layer=POLY_cond $X=0.87 $Y=1.202
+ $X2=0.955 $Y2=1.202
r140 62 65 0.909823 $w=3.78e-07 $l=3e-08 $layer=LI1_cond $X=4.685 $Y=1.99
+ $X2=4.685 $Y2=2.02
r141 55 61 5.12162 $w=2.42e-07 $l=1.30996e-07 $layer=LI1_cond $X=3.195 $Y=1.99
+ $X2=3.075 $Y2=1.967
r142 54 62 3.67462 $w=2.3e-07 $l=1.9e-07 $layer=LI1_cond $X=4.495 $Y=1.99
+ $X2=4.685 $Y2=1.99
r143 54 55 65.1381 $w=2.28e-07 $l=1.3e-06 $layer=LI1_cond $X=4.495 $Y=1.99
+ $X2=3.195 $Y2=1.99
r144 50 61 1.3799 $w=2.4e-07 $l=1.38e-07 $layer=LI1_cond $X=3.075 $Y=2.105
+ $X2=3.075 $Y2=1.967
r145 50 52 9.3636 $w=2.38e-07 $l=1.95e-07 $layer=LI1_cond $X=3.075 $Y=2.105
+ $X2=3.075 $Y2=2.3
r146 48 61 5.12162 $w=2.42e-07 $l=1.249e-07 $layer=LI1_cond $X=2.955 $Y=1.957
+ $X2=3.075 $Y2=1.967
r147 48 49 17.6256 $w=2.53e-07 $l=3.9e-07 $layer=LI1_cond $X=2.955 $Y=1.957
+ $X2=2.565 $Y2=1.957
r148 44 56 1.64524 $w=2.15e-07 $l=1.25e-07 $layer=LI1_cond $X=2.565 $Y=0.762
+ $X2=2.44 $Y2=0.762
r149 44 46 32.4292 $w=2.13e-07 $l=6.05e-07 $layer=LI1_cond $X=2.565 $Y=0.762
+ $X2=3.17 $Y2=0.762
r150 43 49 6.82464 $w=2.55e-07 $l=1.77113e-07 $layer=LI1_cond $X=2.445 $Y=1.83
+ $X2=2.565 $Y2=1.957
r151 43 59 23.7691 $w=2.38e-07 $l=4.95e-07 $layer=LI1_cond $X=2.445 $Y=1.83
+ $X2=2.445 $Y2=1.335
r152 41 76 15.27 $w=3.63e-07 $l=1.15e-07 $layer=POLY_cond $X=2.195 $Y=1.202
+ $X2=2.31 $Y2=1.202
r153 41 74 37.1791 $w=3.63e-07 $l=2.8e-07 $layer=POLY_cond $X=2.195 $Y=1.202
+ $X2=1.915 $Y2=1.202
r154 40 41 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=2.195
+ $Y=1.16 $X2=2.195 $Y2=1.16
r155 37 69 24.5647 $w=3.63e-07 $l=1.85e-07 $layer=POLY_cond $X=0.685 $Y=1.202
+ $X2=0.87 $Y2=1.202
r156 37 67 27.8843 $w=3.63e-07 $l=2.1e-07 $layer=POLY_cond $X=0.685 $Y=1.202
+ $X2=0.475 $Y2=1.202
r157 36 40 51.182 $w=3.38e-07 $l=1.51e-06 $layer=LI1_cond $X=0.685 $Y=1.165
+ $X2=2.195 $Y2=1.165
r158 36 37 58.112 $w=1.7e-07 $l=4.25e-07 $layer=licon1_POLY $count=2 $X=0.685
+ $Y=1.16 $X2=0.685 $Y2=1.16
r159 34 59 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.44 $Y=1.165
+ $X2=2.44 $Y2=1.335
r160 34 56 18.5774 $w=2.48e-07 $l=4.03e-07 $layer=LI1_cond $X=2.44 $Y=1.165
+ $X2=2.44 $Y2=0.762
r161 34 40 4.06745 $w=3.38e-07 $l=1.2e-07 $layer=LI1_cond $X=2.315 $Y=1.165
+ $X2=2.195 $Y2=1.165
r162 31 76 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.31 $Y=1.41
+ $X2=2.31 $Y2=1.202
r163 31 33 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.31 $Y=1.41
+ $X2=2.31 $Y2=1.985
r164 28 74 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=1.202
r165 28 30 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.915 $Y=0.995
+ $X2=1.915 $Y2=0.56
r166 25 73 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.83 $Y=1.41
+ $X2=1.83 $Y2=1.202
r167 25 27 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.83 $Y=1.41
+ $X2=1.83 $Y2=1.985
r168 22 72 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.435 $Y=0.995
+ $X2=1.435 $Y2=1.202
r169 22 24 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.435 $Y=0.995
+ $X2=1.435 $Y2=0.56
r170 19 71 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.35 $Y=1.41
+ $X2=1.35 $Y2=1.202
r171 19 21 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.35 $Y=1.41
+ $X2=1.35 $Y2=1.985
r172 16 70 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=1.202
r173 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.955 $Y=0.995
+ $X2=0.955 $Y2=0.56
r174 13 69 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.87 $Y=1.41
+ $X2=0.87 $Y2=1.202
r175 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.87 $Y=1.41
+ $X2=0.87 $Y2=1.985
r176 10 67 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=1.202
r177 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.475 $Y=0.995
+ $X2=0.475 $Y2=0.56
r178 3 65 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=4.56
+ $Y=1.485 $X2=4.71 $Y2=2.02
r179 2 61 600 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=1 $X=2.9
+ $Y=1.485 $X2=3.05 $Y2=1.96
r180 2 52 600 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=2.9
+ $Y=1.485 $X2=3.05 $Y2=2.3
r181 1 46 182 $w=1.7e-07 $l=5.88643e-07 $layer=licon1_NDIFF $count=1 $X=3.035
+ $Y=0.235 $X2=3.17 $Y2=0.76
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%B1 1 3 4 6 7 9 10 12 13 19 20
c51 19 0 1.95549e-19 $X=3.32 $Y=1.16
c52 10 0 1.04771e-19 $X=3.38 $Y=0.995
r53 20 21 5.14133 $w=3.75e-07 $l=4e-08 $layer=POLY_cond $X=3.34 $Y=1.202
+ $X2=3.38 $Y2=1.202
r54 18 20 2.57067 $w=3.75e-07 $l=2e-08 $layer=POLY_cond $X=3.32 $Y=1.202
+ $X2=3.34 $Y2=1.202
r55 18 19 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.32
+ $Y=1.16 $X2=3.32 $Y2=1.16
r56 16 18 46.272 $w=3.75e-07 $l=3.6e-07 $layer=POLY_cond $X=2.96 $Y=1.202
+ $X2=3.32 $Y2=1.202
r57 15 16 19.28 $w=3.75e-07 $l=1.5e-07 $layer=POLY_cond $X=2.81 $Y=1.202
+ $X2=2.96 $Y2=1.202
r58 13 19 5.90065 $w=7.48e-07 $l=3.7e-07 $layer=LI1_cond $X=3.11 $Y=1.53
+ $X2=3.11 $Y2=1.16
r59 10 21 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.38 $Y=0.995
+ $X2=3.38 $Y2=1.202
r60 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.38 $Y=0.995
+ $X2=3.38 $Y2=0.56
r61 7 20 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.34 $Y=1.41
+ $X2=3.34 $Y2=1.202
r62 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.34 $Y=1.41 $X2=3.34
+ $Y2=1.985
r63 4 16 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.96 $Y=0.995
+ $X2=2.96 $Y2=1.202
r64 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.96 $Y=0.995 $X2=2.96
+ $Y2=0.56
r65 1 15 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.81 $Y=1.41
+ $X2=2.81 $Y2=1.202
r66 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.81 $Y=1.41 $X2=2.81
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%A1 1 3 4 6 7 9 10 12 15 18 19 20 26 27
c69 15 0 3.10869e-19 $X=3.88 $Y=1.16
r70 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.495
+ $Y=1.16 $X2=5.495 $Y2=1.16
r71 20 27 2.53261 $w=4.7e-07 $l=1.05e-07 $layer=LI1_cond $X=5.645 $Y=1.6
+ $X2=5.645 $Y2=1.495
r72 20 27 0.636212 $w=4.68e-07 $l=2.5e-08 $layer=LI1_cond $X=5.645 $Y=1.47
+ $X2=5.645 $Y2=1.495
r73 20 26 7.88903 $w=4.68e-07 $l=3.1e-07 $layer=LI1_cond $X=5.645 $Y=1.47
+ $X2=5.645 $Y2=1.16
r74 18 20 5.66822 $w=2.1e-07 $l=2.35e-07 $layer=LI1_cond $X=5.41 $Y=1.6
+ $X2=5.645 $Y2=1.6
r75 18 19 68.3939 $w=2.08e-07 $l=1.295e-06 $layer=LI1_cond $X=5.41 $Y=1.6
+ $X2=4.115 $Y2=1.6
r76 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.88
+ $Y=1.16 $X2=3.88 $Y2=1.16
r77 13 19 7.41726 $w=2.1e-07 $l=2.24442e-07 $layer=LI1_cond $X=3.937 $Y=1.495
+ $X2=4.115 $Y2=1.6
r78 13 15 10.8752 $w=3.53e-07 $l=3.35e-07 $layer=LI1_cond $X=3.937 $Y=1.495
+ $X2=3.937 $Y2=1.16
r79 10 25 45.964 $w=3.43e-07 $l=2.91548e-07 $layer=POLY_cond $X=5.43 $Y=1.41
+ $X2=5.52 $Y2=1.16
r80 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.43 $Y=1.41
+ $X2=5.43 $Y2=1.985
r81 7 25 38.7084 $w=3.43e-07 $l=2.14942e-07 $layer=POLY_cond $X=5.405 $Y=0.995
+ $X2=5.52 $Y2=1.16
r82 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.405 $Y=0.995
+ $X2=5.405 $Y2=0.56
r83 4 16 45.167 $w=3.78e-07 $l=3.01247e-07 $layer=POLY_cond $X=4.04 $Y=1.41
+ $X2=3.927 $Y2=1.16
r84 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.04 $Y=1.41 $X2=4.04
+ $Y2=1.985
r85 1 16 39.1844 $w=3.78e-07 $l=1.9182e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.927 $Y2=1.16
r86 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.985 $Y=0.995
+ $X2=3.985 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%A2 1 3 4 6 7 9 10 12 13 19 20
c44 1 0 1.06187e-19 $X=4.445 $Y=0.995
r45 19 21 1.928 $w=3.75e-07 $l=1.5e-08 $layer=POLY_cond $X=4.935 $Y=1.202
+ $X2=4.95 $Y2=1.202
r46 19 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.935
+ $Y=1.16 $X2=4.935 $Y2=1.16
r47 17 19 1.28533 $w=3.75e-07 $l=1e-08 $layer=POLY_cond $X=4.925 $Y=1.202
+ $X2=4.935 $Y2=1.202
r48 16 17 58.4827 $w=3.75e-07 $l=4.55e-07 $layer=POLY_cond $X=4.47 $Y=1.202
+ $X2=4.925 $Y2=1.202
r49 15 16 3.21333 $w=3.75e-07 $l=2.5e-08 $layer=POLY_cond $X=4.445 $Y=1.202
+ $X2=4.47 $Y2=1.202
r50 13 20 3.84148 $w=3.28e-07 $l=1.1e-07 $layer=LI1_cond $X=4.825 $Y=1.16
+ $X2=4.935 $Y2=1.16
r51 10 21 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.95 $Y=1.41
+ $X2=4.95 $Y2=1.202
r52 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.95 $Y=1.41
+ $X2=4.95 $Y2=1.985
r53 7 17 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.925 $Y=0.995
+ $X2=4.925 $Y2=1.202
r54 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.925 $Y=0.995
+ $X2=4.925 $Y2=0.56
r55 4 16 19.9308 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.47 $Y=1.41
+ $X2=4.47 $Y2=1.202
r56 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.47 $Y=1.41 $X2=4.47
+ $Y2=1.985
r57 1 15 24.2915 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.445 $Y=0.995
+ $X2=4.445 $Y2=1.202
r58 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.445 $Y=0.995
+ $X2=4.445 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%VPWR 1 2 3 4 5 18 22 26 28 30 33 34 35 37
+ 42 47 56 64 67 70 78
c87 47 0 1.7149e-19 $X=2.335 $Y=2.72
c88 4 0 9.99115e-20 $X=3.43 $Y=1.485
r89 77 78 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r90 73 74 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r91 70 73 10.9482 $w=3.98e-07 $l=3.8e-07 $layer=LI1_cond $X=2.535 $Y=2.34
+ $X2=2.535 $Y2=2.72
r92 67 68 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r93 64 65 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 62 78 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 61 62 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r96 59 62 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r97 58 61 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r98 58 59 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r99 56 77 5.48516 $w=1.7e-07 $l=2.62e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.717 $Y2=2.72
r100 56 61 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=5.455 $Y=2.72
+ $X2=5.29 $Y2=2.72
r101 55 59 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r102 55 74 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r103 54 55 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 52 73 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=2.535 $Y2=2.72
r105 52 54 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.735 $Y=2.72
+ $X2=3.45 $Y2=2.72
r106 51 74 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r107 51 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.61 $Y2=2.72
r108 50 51 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r109 48 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=1.565 $Y2=2.72
r110 48 50 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=1.755 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 47 73 5.77842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.535 $Y2=2.72
r112 47 50 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=2.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r113 46 68 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r114 46 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r115 45 46 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r116 43 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.795 $Y=2.72
+ $X2=0.605 $Y2=2.72
r117 43 45 23.1604 $w=1.68e-07 $l=3.55e-07 $layer=LI1_cond $X=0.795 $Y=2.72
+ $X2=1.15 $Y2=2.72
r118 42 67 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.565 $Y2=2.72
r119 42 45 14.6791 $w=1.68e-07 $l=2.25e-07 $layer=LI1_cond $X=1.375 $Y=2.72
+ $X2=1.15 $Y2=2.72
r120 37 64 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.605 $Y2=2.72
r121 37 39 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=0.415 $Y=2.72
+ $X2=0.23 $Y2=2.72
r122 35 65 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r123 35 39 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r124 33 54 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.45 $Y2=2.72
r125 33 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.515 $Y=2.72
+ $X2=3.68 $Y2=2.72
r126 32 58 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=3.91 $Y2=2.72
r127 32 34 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.845 $Y=2.72
+ $X2=3.68 $Y2=2.72
r128 28 77 2.97287 $w=4.1e-07 $l=1.09864e-07 $layer=LI1_cond $X=5.66 $Y=2.635
+ $X2=5.717 $Y2=2.72
r129 28 30 17.2866 $w=4.08e-07 $l=6.15e-07 $layer=LI1_cond $X=5.66 $Y=2.635
+ $X2=5.66 $Y2=2.02
r130 24 34 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.68 $Y=2.635
+ $X2=3.68 $Y2=2.72
r131 24 26 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=3.68 $Y=2.635
+ $X2=3.68 $Y2=2.36
r132 20 67 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.565 $Y=2.635
+ $X2=1.565 $Y2=2.72
r133 20 22 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=1.565 $Y=2.635
+ $X2=1.565 $Y2=1.955
r134 16 64 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=0.605 $Y=2.635
+ $X2=0.605 $Y2=2.72
r135 16 18 20.6227 $w=3.78e-07 $l=6.8e-07 $layer=LI1_cond $X=0.605 $Y=2.635
+ $X2=0.605 $Y2=1.955
r136 5 30 300 $w=1.7e-07 $l=6.05372e-07 $layer=licon1_PDIFF $count=2 $X=5.52
+ $Y=1.485 $X2=5.67 $Y2=2.02
r137 4 26 600 $w=1.7e-07 $l=9.92157e-07 $layer=licon1_PDIFF $count=1 $X=3.43
+ $Y=1.485 $X2=3.68 $Y2=2.36
r138 3 70 600 $w=1.7e-07 $l=9.36149e-07 $layer=licon1_PDIFF $count=1 $X=2.4
+ $Y=1.485 $X2=2.57 $Y2=2.34
r139 2 22 300 $w=1.7e-07 $l=5.39815e-07 $layer=licon1_PDIFF $count=2 $X=1.44
+ $Y=1.485 $X2=1.59 $Y2=1.955
r140 1 18 300 $w=1.7e-07 $l=5.28819e-07 $layer=licon1_PDIFF $count=2 $X=0.455
+ $Y=1.485 $X2=0.58 $Y2=1.955
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%X 1 2 3 4 15 16 19 21 25 27 31 34 35 36 39
+ 41
c57 39 0 1.01803e-19 $X=0.22 $Y=0.805
r58 39 41 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=0.22 $Y=0.805
+ $X2=0.22 $Y2=0.85
r59 36 39 2.85134 $w=2.6e-07 $l=8.5e-08 $layer=LI1_cond $X=0.22 $Y=0.72 $X2=0.22
+ $Y2=0.805
r60 36 41 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=0.22 $Y=0.87 $X2=0.22
+ $Y2=0.85
r61 33 36 29.2543 $w=2.58e-07 $l=6.6e-07 $layer=LI1_cond $X=0.22 $Y=1.53
+ $X2=0.22 $Y2=0.87
r62 29 31 8.62626 $w=1.78e-07 $l=1.4e-07 $layer=LI1_cond $X=2.065 $Y=1.7
+ $X2=2.065 $Y2=1.84
r63 28 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.205 $Y=1.615
+ $X2=1.11 $Y2=1.615
r64 27 29 6.82373 $w=1.7e-07 $l=1.25499e-07 $layer=LI1_cond $X=1.975 $Y=1.615
+ $X2=2.065 $Y2=1.7
r65 27 28 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.975 $Y=1.615
+ $X2=1.205 $Y2=1.615
r66 23 35 0.945268 $w=1.9e-07 $l=8.5e-08 $layer=LI1_cond $X=1.11 $Y=1.7 $X2=1.11
+ $Y2=1.615
r67 23 25 8.17225 $w=1.88e-07 $l=1.4e-07 $layer=LI1_cond $X=1.11 $Y=1.7 $X2=1.11
+ $Y2=1.84
r68 19 34 5.69365 $w=1.88e-07 $l=9.5e-08 $layer=LI1_cond $X=0.74 $Y=0.71
+ $X2=0.645 $Y2=0.71
r69 19 21 56.0383 $w=1.88e-07 $l=9.6e-07 $layer=LI1_cond $X=0.74 $Y=0.71 $X2=1.7
+ $Y2=0.71
r70 16 33 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.35 $Y=1.615
+ $X2=0.22 $Y2=1.53
r71 15 35 5.66127 $w=1.7e-07 $l=9.5e-08 $layer=LI1_cond $X=1.015 $Y=1.615
+ $X2=1.11 $Y2=1.615
r72 15 16 43.385 $w=1.68e-07 $l=6.65e-07 $layer=LI1_cond $X=1.015 $Y=1.615
+ $X2=0.35 $Y2=1.615
r73 14 36 4.36088 $w=1.7e-07 $l=1.3e-07 $layer=LI1_cond $X=0.35 $Y=0.72 $X2=0.22
+ $Y2=0.72
r74 14 34 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.35 $Y=0.72
+ $X2=0.645 $Y2=0.72
r75 4 31 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=1.92
+ $Y=1.485 $X2=2.07 $Y2=1.84
r76 3 25 300 $w=1.7e-07 $l=4.23409e-07 $layer=licon1_PDIFF $count=2 $X=0.96
+ $Y=1.485 $X2=1.11 $Y2=1.84
r77 2 21 182 $w=1.7e-07 $l=5.62028e-07 $layer=licon1_NDIFF $count=1 $X=1.51
+ $Y=0.235 $X2=1.7 $Y2=0.71
r78 1 19 182 $w=1.7e-07 $l=5.72167e-07 $layer=licon1_NDIFF $count=1 $X=0.55
+ $Y=0.235 $X2=0.74 $Y2=0.72
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%VGND 1 2 3 4 5 16 18 22 24 28 32 35 36 37
+ 38 44 46 62 63 69 72
c89 16 0 1.01803e-19 $X=0.26 $Y=0.085
r90 72 73 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r91 70 73 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r92 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r93 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r94 60 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r95 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r96 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r97 56 57 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r98 54 57 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r99 54 73 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r100 53 56 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r101 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r102 51 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.345 $Y=0 $X2=2.18
+ $Y2=0
r103 51 53 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=2.345 $Y=0
+ $X2=2.53 $Y2=0
r104 50 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r105 49 50 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r106 47 66 4.78091 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.212 $Y2=0
r107 47 49 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.425 $Y=0
+ $X2=0.69 $Y2=0
r108 46 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.22
+ $Y2=0
r109 46 49 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0
+ $X2=0.69 $Y2=0
r110 44 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r111 44 66 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r112 40 62 25.7701 $w=1.68e-07 $l=3.95e-07 $layer=LI1_cond $X=5.355 $Y=0
+ $X2=5.75 $Y2=0
r113 38 59 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.975 $Y=0
+ $X2=4.83 $Y2=0
r114 37 42 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.165 $Y=0
+ $X2=5.165 $Y2=0.36
r115 37 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=5.355
+ $Y2=0
r116 37 38 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.165 $Y=0 $X2=4.975
+ $Y2=0
r117 35 56 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=4.055 $Y=0
+ $X2=3.91 $Y2=0
r118 35 36 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.055 $Y=0 $X2=4.225
+ $Y2=0
r119 34 59 28.3797 $w=1.68e-07 $l=4.35e-07 $layer=LI1_cond $X=4.395 $Y=0
+ $X2=4.83 $Y2=0
r120 34 36 8.79175 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=4.395 $Y=0 $X2=4.225
+ $Y2=0
r121 30 36 0.987631 $w=3.4e-07 $l=8.5e-08 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0
r122 30 32 9.32123 $w=3.38e-07 $l=2.75e-07 $layer=LI1_cond $X=4.225 $Y=0.085
+ $X2=4.225 $Y2=0.36
r123 26 72 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0
r124 26 28 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.18 $Y=0.085
+ $X2=2.18 $Y2=0.38
r125 25 69 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.385 $Y=0 $X2=1.22
+ $Y2=0
r126 24 72 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.18
+ $Y2=0
r127 24 25 41.1016 $w=1.68e-07 $l=6.3e-07 $layer=LI1_cond $X=2.015 $Y=0
+ $X2=1.385 $Y2=0
r128 20 69 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0
r129 20 22 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.22 $Y=0.085
+ $X2=1.22 $Y2=0.36
r130 16 66 2.98526 $w=3.3e-07 $l=1.06325e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.212 $Y2=0
r131 16 18 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.26 $Y=0.085
+ $X2=0.26 $Y2=0.38
r132 5 42 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=5
+ $Y=0.235 $X2=5.19 $Y2=0.36
r133 4 32 182 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=1 $X=4.06
+ $Y=0.235 $X2=4.22 $Y2=0.36
r134 3 28 182 $w=1.7e-07 $l=2.5229e-07 $layer=licon1_NDIFF $count=1 $X=1.99
+ $Y=0.235 $X2=2.18 $Y2=0.38
r135 2 22 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=1.03
+ $Y=0.235 $X2=1.22 $Y2=0.36
r136 1 18 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__O21A_4%A_525_47# 1 2 3 4 13 21 24
r39 26 27 11.5244 $w=3.28e-07 $l=3.3e-07 $layer=LI1_cond $X=3.72 $Y=0.37
+ $X2=3.72 $Y2=0.7
r40 24 26 0.349225 $w=3.28e-07 $l=1e-08 $layer=LI1_cond $X=3.72 $Y=0.36 $X2=3.72
+ $Y2=0.37
r41 19 21 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=4.71 $Y=0.7 $X2=5.67
+ $Y2=0.7
r42 17 27 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.885 $Y=0.7
+ $X2=3.72 $Y2=0.7
r43 17 19 53.8235 $w=1.68e-07 $l=8.25e-07 $layer=LI1_cond $X=3.885 $Y=0.7
+ $X2=4.71 $Y2=0.7
r44 13 26 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=3.555 $Y=0.37
+ $X2=3.72 $Y2=0.37
r45 13 15 40.3355 $w=2.28e-07 $l=8.05e-07 $layer=LI1_cond $X=3.555 $Y=0.37
+ $X2=2.75 $Y2=0.37
r46 4 21 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=5.48
+ $Y=0.235 $X2=5.67 $Y2=0.7
r47 3 19 182 $w=1.7e-07 $l=5.51883e-07 $layer=licon1_NDIFF $count=1 $X=4.52
+ $Y=0.235 $X2=4.71 $Y2=0.7
r48 2 24 91 $w=1.7e-07 $l=3.21481e-07 $layer=licon1_NDIFF $count=2 $X=3.455
+ $Y=0.235 $X2=3.72 $Y2=0.36
r49 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.75 $Y2=0.38
.ends

