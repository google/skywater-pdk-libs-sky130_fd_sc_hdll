* NGSPICE file created from sky130_fd_sc_hdll__o211ai_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
M1000 VGND A1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=2.145e+11p pd=1.96e+06u as=3.9325e+11p ps=3.81e+06u
M1001 a_27_47# A2 VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1002 Y A2 a_118_297# VPB phighvt w=1e+06u l=180000u
+  ad=9.2e+11p pd=5.84e+06u as=2.3e+11p ps=2.46e+06u
M1003 VPWR B1 Y VPB phighvt w=1e+06u l=180000u
+  ad=6.2e+11p pd=5.24e+06u as=0p ps=0u
M1004 Y C1 a_304_47# VNB nshort w=650000u l=150000u
+  ad=3.77e+11p pd=2.46e+06u as=2.4375e+11p ps=2.05e+06u
M1005 a_118_297# A1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 Y C1 VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_304_47# B1 a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

