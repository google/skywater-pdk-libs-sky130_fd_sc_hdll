* File: sky130_fd_sc_hdll__nor4b_1.pex.spice
* Created: Wed Sep  2 08:41:34 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%A_91_199# 1 2 7 9 10 12 15 18 19 23 25
r58 25 26 14.3668 $w=2.59e-07 $l=3.05e-07 $layer=LI1_cond $X=3.175 $Y=0.655
+ $X2=3.48 $Y2=0.655
r59 22 26 3.20129 $w=1.7e-07 $l=1.7e-07 $layer=LI1_cond $X=3.48 $Y=0.825
+ $X2=3.48 $Y2=0.655
r60 22 23 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=3.48 $Y=0.825
+ $X2=3.48 $Y2=1.795
r61 19 21 128.338 $w=2.08e-07 $l=2.43e-06 $layer=LI1_cond $X=0.745 $Y=1.9
+ $X2=3.175 $Y2=1.9
r62 18 23 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.395 $Y=1.9
+ $X2=3.48 $Y2=1.795
r63 18 21 11.619 $w=2.08e-07 $l=2.2e-07 $layer=LI1_cond $X=3.395 $Y=1.9
+ $X2=3.175 $Y2=1.9
r64 15 16 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.62
+ $Y=1.16 $X2=0.62 $Y2=1.16
r65 13 19 6.82129 $w=2.1e-07 $l=1.53786e-07 $layer=LI1_cond $X=0.635 $Y=1.795
+ $X2=0.745 $Y2=1.9
r66 13 15 33.2637 $w=2.18e-07 $l=6.35e-07 $layer=LI1_cond $X=0.635 $Y=1.795
+ $X2=0.635 $Y2=1.16
r67 10 16 38.8967 $w=3.59e-07 $l=2.18746e-07 $layer=POLY_cond $X=0.78 $Y=0.995
+ $X2=0.655 $Y2=1.16
r68 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.78 $Y=0.995
+ $X2=0.78 $Y2=0.56
r69 7 16 45.5371 $w=3.59e-07 $l=2.95804e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.655 $Y2=1.16
r70 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.755 $Y=1.41
+ $X2=0.755 $Y2=1.985
r71 2 21 600 $w=1.7e-07 $l=2.83373e-07 $layer=licon1_PDIFF $count=1 $X=3.03
+ $Y=1.68 $X2=3.175 $Y2=1.9
r72 1 25 182 $w=1.7e-07 $l=2.72213e-07 $layer=licon1_NDIFF $count=1 $X=2.99
+ $Y=0.465 $X2=3.175 $Y2=0.66
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%C 1 3 4 6 7 13
r28 7 13 0.578748 $w=6.18e-07 $l=3e-08 $layer=LI1_cond $X=1.18 $Y=1.305 $X2=1.15
+ $Y2=1.305
r29 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.2 $Y=1.16
+ $X2=1.2 $Y2=1.16
r30 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.25 $Y=0.995
+ $X2=1.225 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.25 $Y=0.995 $X2=1.25
+ $Y2=0.56
r32 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.225 $Y=1.41
+ $X2=1.225 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%B 1 3 4 6 7 13
r28 7 13 1.92916 $w=6.18e-07 $l=1e-07 $layer=LI1_cond $X=1.71 $Y=1.305 $X2=1.61
+ $Y2=1.305
r29 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.73
+ $Y=1.16 $X2=1.73 $Y2=1.16
r30 4 10 38.578 $w=2.95e-07 $l=1.77059e-07 $layer=POLY_cond $X=1.78 $Y=0.995
+ $X2=1.755 $Y2=1.16
r31 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.78 $Y=0.995 $X2=1.78
+ $Y2=0.56
r32 1 10 48.1208 $w=2.95e-07 $l=2.5e-07 $layer=POLY_cond $X=1.755 $Y=1.41
+ $X2=1.755 $Y2=1.16
r33 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.755 $Y=1.41
+ $X2=1.755 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%A 1 3 4 6 7 16
c28 16 0 3.59849e-20 $X=2.51 $Y=1.19
r29 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.26
+ $Y=1.16 $X2=2.26 $Y2=1.16
r30 7 16 0.0964579 $w=6.18e-07 $l=5e-09 $layer=LI1_cond $X=2.505 $Y=1.305
+ $X2=2.51 $Y2=1.305
r31 7 11 4.72644 $w=6.18e-07 $l=2.45e-07 $layer=LI1_cond $X=2.505 $Y=1.305
+ $X2=2.26 $Y2=1.305
r32 4 10 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=2.225 $Y=1.41
+ $X2=2.285 $Y2=1.16
r33 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.225 $Y=1.41
+ $X2=2.225 $Y2=1.985
r34 1 10 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=2.2 $Y=0.995
+ $X2=2.285 $Y2=1.16
r35 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.2 $Y=0.995 $X2=2.2
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%D_N 3 5 6 8 9 12 14
c31 6 0 3.59849e-20 $X=2.94 $Y=1.605
r32 12 15 37.8858 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.997 $Y=1.16
+ $X2=2.997 $Y2=1.325
r33 12 14 46.135 $w=3.15e-07 $l=1.65e-07 $layer=POLY_cond $X=2.997 $Y=1.16
+ $X2=2.997 $Y2=0.995
r34 9 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.975
+ $Y=1.16 $X2=2.975 $Y2=1.16
r35 6 8 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=2.94 $Y=1.605
+ $X2=2.94 $Y2=1.89
r36 5 6 33.5616 $w=2e-07 $l=1e-07 $layer=POLY_cond $X=2.94 $Y=1.505 $X2=2.94
+ $Y2=1.605
r37 5 15 59.6839 $w=2e-07 $l=1.8e-07 $layer=POLY_cond $X=2.94 $Y=1.505 $X2=2.94
+ $Y2=1.325
r38 3 14 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=2.915 $Y=0.675
+ $X2=2.915 $Y2=0.995
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%Y 1 2 3 10 11 14 16 20 23 24
c42 10 0 1.57721e-19 $X=0.905 $Y=0.74
r43 22 24 46.3193 $w=2.58e-07 $l=1.045e-06 $layer=LI1_cond $X=0.215 $Y=0.825
+ $X2=0.215 $Y2=1.87
r44 18 20 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=1.975 $Y=0.655
+ $X2=1.975 $Y2=0.495
r45 17 23 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=1.105 $Y=0.74 $X2=1.005
+ $Y2=0.74
r46 16 18 6.87494 $w=1.7e-07 $l=1.36015e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.975 $Y2=0.655
r47 16 17 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.875 $Y=0.74
+ $X2=1.105 $Y2=0.74
r48 12 23 0.764409 $w=2e-07 $l=8.5e-08 $layer=LI1_cond $X=1.005 $Y=0.655
+ $X2=1.005 $Y2=0.74
r49 12 14 8.87273 $w=1.98e-07 $l=1.6e-07 $layer=LI1_cond $X=1.005 $Y=0.655
+ $X2=1.005 $Y2=0.495
r50 11 22 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.345 $Y=0.74
+ $X2=0.215 $Y2=0.825
r51 10 23 5.90115 $w=1.7e-07 $l=1e-07 $layer=LI1_cond $X=0.905 $Y=0.74 $X2=1.005
+ $Y2=0.74
r52 10 11 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=0.905 $Y=0.74
+ $X2=0.345 $Y2=0.74
r53 3 24 300 $w=1.7e-07 $l=5.18748e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.945
r54 2 20 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=1.855
+ $Y=0.235 $X2=1.99 $Y2=0.495
r55 1 14 182 $w=1.7e-07 $l=3.20468e-07 $layer=licon1_NDIFF $count=1 $X=0.855
+ $Y=0.235 $X2=0.99 $Y2=0.495
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%VPWR 1 6 8 10 20 21 24
r32 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r33 21 25 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r34 20 21 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r35 18 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=2.515 $Y2=2.72
r36 18 20 48.6043 $w=1.68e-07 $l=7.45e-07 $layer=LI1_cond $X=2.705 $Y=2.72
+ $X2=3.45 $Y2=2.72
r37 17 25 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r38 16 17 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r39 12 16 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r40 10 24 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.515 $Y2=2.72
r41 10 16 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=2.325 $Y=2.72
+ $X2=2.07 $Y2=2.72
r42 8 17 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r43 8 12 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r44 4 24 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.515 $Y=2.635
+ $X2=2.515 $Y2=2.72
r45 4 6 11.0695 $w=3.78e-07 $l=3.65e-07 $layer=LI1_cond $X=2.515 $Y=2.635
+ $X2=2.515 $Y2=2.27
r46 1 6 600 $w=1.7e-07 $l=8.90421e-07 $layer=licon1_PDIFF $count=1 $X=2.315
+ $Y=1.485 $X2=2.54 $Y2=2.27
.ends

.subckt PM_SKY130_FD_SC_HDLL__NOR4B_1%VGND 1 2 3 12 16 20 23 24 26 27 28 37 43
+ 44 47
c50 23 0 1.57721e-19 $X=0.355 $Y=0
r51 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r52 44 48 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=2.53
+ $Y2=0
r53 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r54 41 47 11.1546 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=2.49
+ $Y2=0
r55 41 43 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=2.735 $Y=0 $X2=3.45
+ $Y2=0
r56 40 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r57 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r58 37 47 11.1546 $w=1.7e-07 $l=2.45e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.49
+ $Y2=0
r59 37 39 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=2.245 $Y=0 $X2=2.07
+ $Y2=0
r60 36 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r61 35 36 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r62 28 36 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r63 28 31 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r64 26 35 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.15
+ $Y2=0
r65 26 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.325 $Y=0 $X2=1.49
+ $Y2=0
r66 25 39 27.0749 $w=1.68e-07 $l=4.15e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=2.07
+ $Y2=0
r67 25 27 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.655 $Y=0 $X2=1.49
+ $Y2=0
r68 23 31 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.23
+ $Y2=0
r69 23 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.355 $Y=0 $X2=0.52
+ $Y2=0
r70 22 35 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.685 $Y=0 $X2=1.15
+ $Y2=0
r71 22 24 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=0.685 $Y=0 $X2=0.52
+ $Y2=0
r72 18 47 2.02226 $w=4.9e-07 $l=8.5e-08 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0
r73 18 20 7.44498 $w=4.88e-07 $l=3.05e-07 $layer=LI1_cond $X=2.49 $Y=0.085
+ $X2=2.49 $Y2=0.39
r74 14 27 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0
r75 14 16 10.6514 $w=3.28e-07 $l=3.05e-07 $layer=LI1_cond $X=1.49 $Y=0.085
+ $X2=1.49 $Y2=0.39
r76 10 24 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0
r77 10 12 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=0.52 $Y=0.085
+ $X2=0.52 $Y2=0.36
r78 3 20 91 $w=1.7e-07 $l=3.23342e-07 $layer=licon1_NDIFF $count=2 $X=2.275
+ $Y=0.235 $X2=2.53 $Y2=0.39
r79 2 16 182 $w=1.7e-07 $l=2.29783e-07 $layer=licon1_NDIFF $count=1 $X=1.325
+ $Y=0.235 $X2=1.49 $Y2=0.39
r80 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.375
+ $Y=0.235 $X2=0.52 $Y2=0.36
.ends

