* File: sky130_fd_sc_hdll__muxb4to1_2.spice
* Created: Thu Aug 27 19:11:52 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb4to1_2.pex.spice"
.subckt sky130_fd_sc_hdll__muxb4to1_2  VNB VPB D[0] S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[3]	D[3]
* S[3]	S[3]
* S[2]	S[2]
* D[2]	D[2]
* D[1]	D[1]
* S[1]	S[1]
* S[0]	S[0]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1013 N_A_27_47#_M1013_d N_D[0]_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1026 N_A_27_47#_M1026_d N_D[0]_M1026_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1011 N_A_27_47#_M1026_d N_S[0]_M1011_g N_Z_M1011_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1014 N_A_27_47#_M1014_d N_S[0]_M1014_g N_Z_M1011_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1021 N_VGND_M1021_d N_S[0]_M1021_g N_A_278_265#_M1021_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1018 N_A_701_47#_M1018_d N_S[1]_M1018_g N_VGND_M1021_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1010 N_A_845_69#_M1010_d N_S[1]_M1010_g N_Z_M1010_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1012 N_A_845_69#_M1012_d N_S[1]_M1012_g N_Z_M1010_s VNB NSHORT L=0.15 W=0.52
+ AD=0.102556 AS=0.0702 PD=0.906667 PS=0.79 NRD=16.728 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1019 N_VGND_M1019_d N_D[1]_M1019_g N_A_845_69#_M1012_d VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.128194 PD=0.92 PS=1.13333 NRD=0 NRS=3.684 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1024 N_VGND_M1019_d N_D[1]_M1024_g N_A_845_69#_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1028 N_A_1315_47#_M1028_d N_D[2]_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.4 A=0.0975 P=1.6 MULT=1
MM1033 N_A_1315_47#_M1033_d N_D[2]_M1033_g N_VGND_M1028_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1029 N_Z_M1029_d N_S[2]_M1029_g N_A_1315_47#_M1033_d VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75001.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1037 N_Z_M1029_d N_S[2]_M1037_g N_A_1315_47#_M1037_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.6
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1038 N_VGND_M1038_d N_S[2]_M1038_g N_A_1566_265#_M1038_s VNB NSHORT L=0.15
+ W=0.52 AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.2 SB=75000.6 A=0.078 P=1.34 MULT=1
MM1007 N_A_1989_47#_M1007_d N_S[3]_M1007_g N_VGND_M1038_d VNB NSHORT L=0.15
+ W=0.52 AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667
+ SA=75000.6 SB=75000.2 A=0.078 P=1.34 MULT=1
MM1025 N_Z_M1025_d N_S[3]_M1025_g N_A_2133_69#_M1025_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.6 A=0.078 P=1.34 MULT=1
MM1034 N_Z_M1025_d N_S[3]_M1034_g N_A_2133_69#_M1034_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.102556 PD=0.79 PS=0.906667 NRD=0 NRS=16.728 M=1 R=3.46667
+ SA=75000.6 SB=75001.2 A=0.078 P=1.34 MULT=1
MM1008 N_A_2133_69#_M1034_s N_D[3]_M1008_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.128194 AS=0.08775 PD=1.13333 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333
+ SA=75000.9 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1039 N_A_2133_69#_M1039_d N_D[3]_M1039_g N_VGND_M1008_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.4 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_27_297#_M1002_d N_D[0]_M1002_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1017 N_A_27_297#_M1017_d N_D[0]_M1017_g N_VPWR_M1002_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1005 N_A_27_297#_M1017_d N_A_278_265#_M1005_g N_Z_M1005_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1009 N_A_27_297#_M1009_d N_A_278_265#_M1009_g N_Z_M1005_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1006 N_VPWR_M1006_d N_S[0]_M1006_g N_A_278_265#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.7 A=0.18 P=2.36 MULT=1
MM1022 N_A_701_47#_M1022_d N_S[1]_M1022_g N_VPWR_M1006_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1020 N_A_824_333#_M1020_d N_A_701_47#_M1020_g N_Z_M1020_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1027 N_A_824_333#_M1027_d N_A_701_47#_M1027_g N_Z_M1020_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.148546 AS=0.1189 PD=1.21198 PS=1.11 NRD=14.4007 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1015 N_A_824_333#_M1027_d N_D[1]_M1015_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.181154 AS=0.145 PD=1.47802 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1023 N_A_824_333#_M1023_d N_D[1]_M1023_g N_VPWR_M1015_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1000 N_VPWR_M1000_d N_D[2]_M1000_g N_A_1315_297#_M1000_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.5 A=0.18 P=2.36 MULT=1
MM1030 N_VPWR_M1000_d N_D[2]_M1030_g N_A_1315_297#_M1030_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90000.6 SB=90001 A=0.18 P=2.36 MULT=1
MM1003 N_Z_M1003_d N_A_1566_265#_M1003_g N_A_1315_297#_M1030_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007
+ M=1 R=4.55556 SA=90001.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1031 N_Z_M1003_d N_A_1566_265#_M1031_g N_A_1315_297#_M1031_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1035 N_VPWR_M1035_d N_S[2]_M1035_g N_A_1566_265#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.18 AS=0.27 PD=1.36 PS=2.54 NRD=7.8603 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1016 N_A_1989_47#_M1016_d N_S[3]_M1016_g N_VPWR_M1035_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.18 PD=2.54 PS=1.36 NRD=0.9653 NRS=7.8603 M=1 R=5.55556 SA=90000.7
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1004 N_Z_M1004_d N_A_1989_47#_M1004_g N_A_2112_333#_M1004_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1032 N_Z_M1004_d N_A_1989_47#_M1032_g N_A_2112_333#_M1032_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.148546 PD=1.11 PS=1.21198 NRD=1.182 NRS=14.4007 M=1
+ R=4.55556 SA=90000.6 SB=90001.2 A=0.1476 P=2 MULT=1
MM1001 N_VPWR_M1001_d N_D[3]_M1001_g N_A_2112_333#_M1032_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.181154 PD=1.29 PS=1.47802 NRD=0.9653 NRS=0.9653 M=1
+ R=5.55556 SA=90001 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1036 N_VPWR_M1001_d N_D[3]_M1036_g N_A_2112_333#_M1036_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX40_noxref VNB VPB NWDIODE A=21.2823 P=29.73
c_129 VNB 0 7.27953e-19 $X=12.565 $Y=-0.085
*
.include "sky130_fd_sc_hdll__muxb4to1_2.pxi.spice"
*
.ends
*
*
