* File: sky130_fd_sc_hdll__o32ai_1.pxi.spice
* Created: Wed Sep  2 08:47:06 2020
* 
x_PM_SKY130_FD_SC_HDLL__O32AI_1%B1 N_B1_c_43_n N_B1_M1003_g N_B1_c_44_n
+ N_B1_M1006_g B1 B1 PM_SKY130_FD_SC_HDLL__O32AI_1%B1
x_PM_SKY130_FD_SC_HDLL__O32AI_1%B2 N_B2_c_66_n N_B2_M1002_g N_B2_c_67_n
+ N_B2_M1005_g B2 B2 PM_SKY130_FD_SC_HDLL__O32AI_1%B2
x_PM_SKY130_FD_SC_HDLL__O32AI_1%A3 N_A3_c_94_n N_A3_M1001_g N_A3_c_95_n
+ N_A3_M1009_g A3 A3 PM_SKY130_FD_SC_HDLL__O32AI_1%A3
x_PM_SKY130_FD_SC_HDLL__O32AI_1%A2 N_A2_c_120_n N_A2_M1004_g N_A2_c_121_n
+ N_A2_M1008_g A2 A2 A2 A2 PM_SKY130_FD_SC_HDLL__O32AI_1%A2
x_PM_SKY130_FD_SC_HDLL__O32AI_1%A1 N_A1_c_151_n N_A1_M1007_g N_A1_c_152_n
+ N_A1_M1000_g A1 N_A1_c_153_n A1 PM_SKY130_FD_SC_HDLL__O32AI_1%A1
x_PM_SKY130_FD_SC_HDLL__O32AI_1%VPWR N_VPWR_M1003_s N_VPWR_M1000_d
+ N_VPWR_c_172_n N_VPWR_c_173_n N_VPWR_c_174_n N_VPWR_c_175_n VPWR
+ N_VPWR_c_176_n N_VPWR_c_171_n PM_SKY130_FD_SC_HDLL__O32AI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__O32AI_1%Y N_Y_M1006_d N_Y_M1002_d N_Y_c_210_n Y Y Y Y
+ PM_SKY130_FD_SC_HDLL__O32AI_1%Y
x_PM_SKY130_FD_SC_HDLL__O32AI_1%A_27_47# N_A_27_47#_M1006_s N_A_27_47#_M1005_d
+ N_A_27_47#_M1008_d N_A_27_47#_c_240_n N_A_27_47#_c_249_n N_A_27_47#_c_264_p
+ PM_SKY130_FD_SC_HDLL__O32AI_1%A_27_47#
x_PM_SKY130_FD_SC_HDLL__O32AI_1%VGND N_VGND_M1001_d N_VGND_M1007_d
+ N_VGND_c_271_n N_VGND_c_272_n N_VGND_c_273_n N_VGND_c_274_n N_VGND_c_275_n
+ VGND N_VGND_c_276_n N_VGND_c_277_n PM_SKY130_FD_SC_HDLL__O32AI_1%VGND
cc_1 VNB N_B1_c_43_n 0.0378304f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_B1_c_44_n 0.0196949f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB B1 0.0238007f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_4 VNB N_B2_c_66_n 0.0259063f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B2_c_67_n 0.0175531f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB B2 0.00328264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A3_c_94_n 0.0192339f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_8 VNB N_A3_c_95_n 0.022688f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_9 VNB A3 0.00232616f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A2_c_120_n 0.0287236f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_A2_c_121_n 0.0190483f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB A2 0.0044374f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=0.765
cc_13 VNB N_A1_c_151_n 0.0213312f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_14 VNB N_A1_c_152_n 0.0309633f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_15 VNB N_A1_c_153_n 0.0179985f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_16 VNB N_VPWR_c_171_n 0.136896f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB Y 0.00292415f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_18 VNB N_A_27_47#_c_240_n 0.010655f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_VGND_c_271_n 0.00564356f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_VGND_c_272_n 0.0120624f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_21 VNB N_VGND_c_273_n 0.026729f $X=-0.19 $Y=-0.24 $X2=0.275 $Y2=1.16
cc_22 VNB N_VGND_c_274_n 0.0404603f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VGND_c_275_n 0.00631563f $X=-0.19 $Y=-0.24 $X2=0.225 $Y2=1.16
cc_24 VNB N_VGND_c_276_n 0.0197474f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_277_n 0.181457f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VPB N_B1_c_43_n 0.0386596f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_27 VPB B1 0.00323634f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_28 VPB N_B2_c_66_n 0.0279953f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_29 VPB B2 0.00110322f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_A3_c_95_n 0.0279271f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_31 VPB A3 0.00233114f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_A2_c_120_n 0.029669f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_33 VPB A2 0.00111582f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_34 VPB N_A1_c_152_n 0.0347378f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_35 VPB N_A1_c_153_n 0.00877135f $X=-0.19 $Y=1.305 $X2=0.352 $Y2=1.16
cc_36 VPB N_VPWR_c_172_n 0.0102356f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=0.765
cc_37 VPB N_VPWR_c_173_n 0.0430524f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_38 VPB N_VPWR_c_174_n 0.0104942f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_39 VPB N_VPWR_c_175_n 0.0436422f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_VPWR_c_176_n 0.0634444f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_41 VPB N_VPWR_c_171_n 0.0427625f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB Y 0.00104554f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_43 N_B1_c_43_n N_B2_c_66_n 0.0936988f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_44 N_B1_c_44_n N_B2_c_67_n 0.0222856f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_45 N_B1_c_43_n B2 4.86217e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_46 N_B1_c_43_n N_VPWR_c_173_n 0.00654458f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_47 B1 N_VPWR_c_173_n 0.022987f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_48 N_B1_c_43_n N_VPWR_c_176_n 0.00618965f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_49 N_B1_c_43_n N_VPWR_c_171_n 0.0112959f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_50 N_B1_c_44_n N_Y_c_210_n 0.00429437f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_51 B1 N_Y_c_210_n 0.0107598f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_52 N_B1_c_43_n Y 0.0395237f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_B1_c_44_n Y 0.00349401f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 B1 Y 0.0363777f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_55 B1 N_A_27_47#_M1006_s 0.0057692f $X=0.15 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_56 N_B1_c_43_n N_A_27_47#_c_240_n 0.00263424f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_B1_c_44_n N_A_27_47#_c_240_n 0.013234f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_58 B1 N_A_27_47#_c_240_n 0.0184592f $X=0.15 $Y=0.765 $X2=0 $Y2=0
cc_59 N_B1_c_44_n N_VGND_c_274_n 0.00357877f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_60 N_B1_c_44_n N_VGND_c_277_n 0.00648873f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_61 N_B2_c_67_n N_A3_c_94_n 0.0113112f $X=1.045 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_62 N_B2_c_66_n N_A3_c_95_n 0.0357264f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_63 B2 N_A3_c_95_n 0.00347605f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_64 N_B2_c_66_n A3 6.91453e-19 $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_65 B2 A3 0.0449473f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_66 N_B2_c_66_n N_VPWR_c_176_n 0.00429453f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_67 N_B2_c_66_n N_VPWR_c_171_n 0.00640061f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_68 B2 N_Y_M1002_d 0.00465833f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_69 N_B2_c_66_n N_Y_c_210_n 0.00370701f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B2_c_67_n N_Y_c_210_n 0.00140795f $X=1.045 $Y=0.995 $X2=0 $Y2=0
cc_71 N_B2_c_66_n Y 0.0082698f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_72 N_B2_c_67_n Y 0.00362768f $X=1.045 $Y=0.995 $X2=0 $Y2=0
cc_73 B2 Y 0.0479392f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_74 N_B2_c_66_n Y 0.0270246f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_75 B2 Y 0.0286885f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_76 N_B2_c_66_n N_A_27_47#_c_240_n 0.00161691f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_77 N_B2_c_67_n N_A_27_47#_c_240_n 0.0182139f $X=1.045 $Y=0.995 $X2=0 $Y2=0
cc_78 B2 N_A_27_47#_c_240_n 0.0222039f $X=1.155 $Y=1.19 $X2=0 $Y2=0
cc_79 N_B2_c_67_n N_VGND_c_274_n 0.00359319f $X=1.045 $Y=0.995 $X2=0 $Y2=0
cc_80 N_B2_c_67_n N_VGND_c_277_n 0.00556559f $X=1.045 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A3_c_95_n N_A2_c_120_n 0.045399f $X=1.6 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_82 A3 N_A2_c_120_n 0.00144443f $X=1.615 $Y=1.19 $X2=-0.19 $Y2=-0.24
cc_83 N_A3_c_94_n N_A2_c_121_n 0.0153097f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_84 N_A3_c_95_n A2 0.012378f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_85 A3 A2 0.0449492f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_86 N_A3_c_95_n N_VPWR_c_176_n 0.00672127f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A3_c_95_n N_VPWR_c_171_n 0.0128882f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A3_c_95_n Y 0.0253084f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_89 A3 Y 0.00166452f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_90 N_A3_c_94_n N_A_27_47#_c_240_n 0.0128794f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A3_c_94_n N_A_27_47#_c_249_n 0.0111456f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A3_c_95_n N_A_27_47#_c_249_n 0.00353687f $X=1.6 $Y=1.41 $X2=0 $Y2=0
cc_93 A3 N_A_27_47#_c_249_n 0.0188868f $X=1.615 $Y=1.19 $X2=0 $Y2=0
cc_94 N_A3_c_94_n N_VGND_c_271_n 0.00624423f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A3_c_94_n N_VGND_c_274_n 0.00415469f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A3_c_94_n N_VGND_c_277_n 0.00648583f $X=1.485 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A2_c_121_n N_A1_c_151_n 0.0217195f $X=2.26 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_98 N_A2_c_120_n N_A1_c_152_n 0.0718186f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_99 A2 N_A1_c_152_n 0.00414457f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_100 N_A2_c_120_n N_A1_c_153_n 0.00296713f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_101 A2 N_A1_c_153_n 0.0249348f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_102 N_A2_c_120_n N_VPWR_c_175_n 0.00378048f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_103 A2 N_VPWR_c_175_n 0.0263069f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_104 N_A2_c_120_n N_VPWR_c_176_n 0.00612893f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_105 A2 N_VPWR_c_176_n 0.0181402f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A2_c_120_n N_VPWR_c_171_n 0.0109872f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_107 A2 N_VPWR_c_171_n 0.0108216f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A2_c_120_n Y 5.25802e-19 $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_109 A2 Y 0.0293923f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_110 A2 A_338_297# 0.0158487f $X=1.97 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_111 N_A2_c_120_n N_A_27_47#_c_249_n 0.00149296f $X=2.235 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A2_c_121_n N_A_27_47#_c_249_n 0.0159805f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_113 A2 N_A_27_47#_c_249_n 0.0206881f $X=1.97 $Y=1.105 $X2=0 $Y2=0
cc_114 N_A2_c_121_n N_VGND_c_271_n 0.0071784f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_115 N_A2_c_121_n N_VGND_c_273_n 0.00184853f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_116 N_A2_c_121_n N_VGND_c_276_n 0.00428022f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_117 N_A2_c_121_n N_VGND_c_277_n 0.00665375f $X=2.26 $Y=0.995 $X2=0 $Y2=0
cc_118 N_A1_c_152_n N_VPWR_c_175_n 0.0275826f $X=2.705 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A1_c_153_n N_VPWR_c_175_n 0.0142419f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_120 N_A1_c_152_n N_VPWR_c_176_n 0.00661659f $X=2.705 $Y=1.41 $X2=0 $Y2=0
cc_121 N_A1_c_152_n N_VPWR_c_171_n 0.0111195f $X=2.705 $Y=1.41 $X2=0 $Y2=0
cc_122 N_A1_c_153_n N_A_27_47#_c_249_n 0.0131485f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_123 N_A1_c_151_n N_VGND_c_273_n 0.0137642f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_124 N_A1_c_152_n N_VGND_c_273_n 0.00535295f $X=2.705 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A1_c_153_n N_VGND_c_273_n 0.0191416f $X=2.8 $Y=1.16 $X2=0 $Y2=0
cc_126 N_A1_c_151_n N_VGND_c_276_n 0.0046653f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_127 N_A1_c_151_n N_VGND_c_277_n 0.00799591f $X=2.68 $Y=0.995 $X2=0 $Y2=0
cc_128 N_VPWR_c_171_n A_117_297# 0.00184694f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_129 N_VPWR_c_171_n N_Y_M1002_d 0.00415391f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_130 N_VPWR_c_176_n Y 0.0132994f $X=2.785 $Y=2.72 $X2=0 $Y2=0
cc_131 N_VPWR_c_171_n Y 0.0082112f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_132 N_VPWR_c_176_n Y 0.0480804f $X=2.785 $Y=2.72 $X2=0 $Y2=0
cc_133 N_VPWR_c_171_n Y 0.02903f $X=2.99 $Y=2.72 $X2=0 $Y2=0
cc_134 N_VPWR_c_171_n A_338_297# 0.0115153f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_135 N_VPWR_c_171_n A_465_297# 0.0123962f $X=2.99 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_136 N_VPWR_c_175_n N_VGND_c_273_n 0.0034085f $X=2.94 $Y=1.66 $X2=0 $Y2=0
cc_137 A_117_297# Y 0.00403556f $X=0.585 $Y=1.485 $X2=2.96 $Y2=2.635
cc_138 A_117_297# Y 3.84267e-19 $X=0.585 $Y=1.485 $X2=0 $Y2=0
cc_139 N_Y_M1006_d N_A_27_47#_c_240_n 0.0054624f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_140 N_Y_c_210_n N_A_27_47#_c_240_n 0.0348206f $X=0.73 $Y=0.74 $X2=0 $Y2=0
cc_141 N_Y_M1006_d N_VGND_c_277_n 0.00301157f $X=0.595 $Y=0.235 $X2=0 $Y2=0
cc_142 N_A_27_47#_c_249_n N_VGND_M1001_d 0.018488f $X=2.385 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_143 N_A_27_47#_c_240_n N_VGND_c_271_n 0.0156053f $X=1.065 $Y=0.37 $X2=0 $Y2=0
cc_144 N_A_27_47#_c_249_n N_VGND_c_271_n 0.0251797f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_145 N_A_27_47#_c_240_n N_VGND_c_274_n 0.0797104f $X=1.065 $Y=0.37 $X2=0 $Y2=0
cc_146 N_A_27_47#_c_249_n N_VGND_c_274_n 0.00286445f $X=2.385 $Y=0.74 $X2=0
+ $Y2=0
cc_147 N_A_27_47#_c_249_n N_VGND_c_276_n 0.00588563f $X=2.385 $Y=0.74 $X2=0
+ $Y2=0
cc_148 N_A_27_47#_c_264_p N_VGND_c_276_n 0.0062327f $X=2.47 $Y=0.54 $X2=0 $Y2=0
cc_149 N_A_27_47#_M1006_s N_VGND_c_277_n 0.00250339f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_150 N_A_27_47#_M1005_d N_VGND_c_277_n 0.00231261f $X=1.12 $Y=0.235 $X2=0
+ $Y2=0
cc_151 N_A_27_47#_M1008_d N_VGND_c_277_n 0.00421763f $X=2.335 $Y=0.235 $X2=0
+ $Y2=0
cc_152 N_A_27_47#_c_240_n N_VGND_c_277_n 0.0493289f $X=1.065 $Y=0.37 $X2=0 $Y2=0
cc_153 N_A_27_47#_c_249_n N_VGND_c_277_n 0.0172782f $X=2.385 $Y=0.74 $X2=0 $Y2=0
cc_154 N_A_27_47#_c_264_p N_VGND_c_277_n 0.00596842f $X=2.47 $Y=0.54 $X2=0 $Y2=0
