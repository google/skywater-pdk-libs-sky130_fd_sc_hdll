* File: sky130_fd_sc_hdll__a21boi_4.spice
* Created: Wed Sep  2 08:16:58 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21boi_4.pex.spice"
.subckt sky130_fd_sc_hdll__a21boi_4  VNB VPB B1_N A2 A1 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A1	A1
* A2	A2
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1015 N_VGND_M1015_d N_B1_N_M1015_g N_A_27_47#_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.30225 PD=1.03 PS=2.23 NRD=11.076 NRS=33.228 M=1 R=4.33333
+ SA=75000.4 SB=75006.4 A=0.0975 P=1.6 MULT=1
MM1002 N_VGND_M1015_d N_A_27_47#_M1002_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.10725 PD=1.03 PS=0.98 NRD=7.38 NRS=9.228 M=1 R=4.33333
+ SA=75000.9 SB=75005.9 A=0.0975 P=1.6 MULT=1
MM1018 N_VGND_M1018_d N_A_27_47#_M1018_g N_Y_M1002_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75001.4
+ SB=75005.4 A=0.0975 P=1.6 MULT=1
MM1019 N_VGND_M1018_d N_A_27_47#_M1019_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.10725 PD=0.98 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75001.9
+ SB=75004.9 A=0.0975 P=1.6 MULT=1
MM1025 N_VGND_M1025_d N_A_27_47#_M1025_g N_Y_M1019_s VNB NSHORT L=0.15 W=0.65
+ AD=0.24375 AS=0.10725 PD=1.4 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75002.4
+ SB=75004.4 A=0.0975 P=1.6 MULT=1
MM1000 N_A_724_47#_M1000_d N_A2_M1000_g N_VGND_M1025_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.24375 PD=0.92 PS=1.4 NRD=0 NRS=5.532 M=1 R=4.33333 SA=75003.3
+ SB=75003.5 A=0.0975 P=1.6 MULT=1
MM1007 N_Y_M1007_d N_A1_M1007_g N_A_724_47#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.08775 PD=1.01 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333 SA=75003.7
+ SB=75003.1 A=0.0975 P=1.6 MULT=1
MM1009 N_Y_M1007_d N_A1_M1009_g N_A_724_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.117 AS=0.10725 PD=1.01 PS=0.98 NRD=0 NRS=9.228 M=1 R=4.33333 SA=75004.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1013 N_Y_M1013_d N_A1_M1013_g N_A_724_47#_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.10725 PD=1 PS=0.98 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75004.7
+ SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1020 N_Y_M1013_d N_A1_M1020_g N_A_724_47#_M1020_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11375 AS=0.08775 PD=1 PS=0.92 NRD=3.684 NRS=0 M=1 R=4.33333 SA=75005.2
+ SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1001 N_A_724_47#_M1020_s N_A2_M1001_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=16.608 M=1 R=4.33333
+ SA=75005.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1004 N_A_724_47#_M1004_d N_A2_M1004_g N_VGND_M1001_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.12025 PD=0.98 PS=1.02 NRD=9.228 NRS=0 M=1 R=4.33333 SA=75006.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1012 N_A_724_47#_M1004_d N_A2_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.1755 PD=0.98 PS=1.84 NRD=0 NRS=0 M=1 R=4.33333 SA=75006.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_VPWR_M1010_d N_B1_N_M1010_g N_A_27_47#_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.275 PD=2.55 PS=2.55 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_227_297#_M1005_d N_A_27_47#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.325 AS=0.15 PD=2.65 PS=1.3 NRD=10.8153 NRS=1.9503 M=1 R=5.55556
+ SA=90000.2 SB=90005.5 A=0.18 P=2.36 MULT=1
MM1008 N_A_227_297#_M1008_d N_A_27_47#_M1008_g N_Y_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90000.7 SB=90005 A=0.18 P=2.36 MULT=1
MM1016 N_A_227_297#_M1008_d N_A_27_47#_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556
+ SA=90001.2 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1022 N_A_227_297#_M1022_d N_A_27_47#_M1022_g N_Y_M1016_s VPB PHIGHVT L=0.18
+ W=1 AD=0.165 AS=0.15 PD=1.33 PS=1.3 NRD=7.8603 NRS=1.9503 M=1 R=5.55556
+ SA=90001.7 SB=90004 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A2_M1003_g N_A_227_297#_M1022_d VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.165 PD=1.31 PS=1.33 NRD=3.9203 NRS=1.9503 M=1 R=5.55556
+ SA=90002.2 SB=90003.5 A=0.18 P=2.36 MULT=1
MM1014 N_VPWR_M1003_d N_A1_M1014_g N_A_227_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.155 AS=0.15 PD=1.31 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90002.7
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1017 N_VPWR_M1017_d N_A1_M1017_g N_A_227_297#_M1014_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.2
+ SB=90002.6 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1017_d N_A1_M1021_g N_A_227_297#_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.15 PD=1.3 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90003.6
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1024 N_VPWR_M1024_d N_A1_M1024_g N_A_227_297#_M1021_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.15 PD=1.29 PS=1.3 NRD=0.9653 NRS=1.9503 M=1 R=5.55556 SA=90004.1
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1024_d N_A2_M1006_g N_A_227_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A2_M1011_g N_A_227_297#_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1011_d N_A2_M1023_g N_A_227_297#_M1023_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.28 PD=1.29 PS=2.56 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90005.5 SB=90000.2 A=0.18 P=2.36 MULT=1
DX26_noxref VNB VPB NWDIODE A=12.4227 P=18.69
pX27_noxref noxref_12 A2 A2 PROBETYPE=1
c_47 VNB 0 1.09328e-19 $X=0.145 $Y=-0.085
c_90 VPB 0 3.14505e-20 $X=0.145 $Y=2.635
*
.include "sky130_fd_sc_hdll__a21boi_4.pxi.spice"
*
.ends
*
*
