* NGSPICE file created from sky130_fd_sc_hdll__sdfsbp_1.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__sdfsbp_1 CLK D SCD SCE SET_B VGND VNB VPB VPWR Q Q_N
M1000 VGND a_349_21# a_295_47# VNB nshort w=420000u l=150000u
+  ad=1.4601e+12p pd=1.494e+07u as=1.134e+11p ps=1.38e+06u
M1001 a_1930_295# a_1735_329# VGND VNB nshort w=420000u l=150000u
+  ad=1.092e+11p pd=1.36e+06u as=0p ps=0u
M1002 Q a_2632_47# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=1.9705e+12p ps=1.846e+07u
M1003 a_1930_295# a_1735_329# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.134e+11p pd=1.38e+06u as=0p ps=0u
M1004 a_1075_413# a_877_369# a_199_47# VPB phighvt w=420000u l=180000u
+  ad=1.218e+11p pd=1.42e+06u as=2.99e+11p ps=3.24e+06u
M1005 VGND SCE a_349_21# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.176e+11p ps=1.4e+06u
M1006 a_1735_329# a_877_369# a_1655_47# VNB nshort w=640000u l=150000u
+  ad=3.054e+11p pd=2.42e+06u as=4.736e+11p ps=2.76e+06u
M1007 VPWR SCD a_27_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=3.456e+11p ps=3.64e+06u
M1008 a_1219_21# a_1075_413# VPWR VPB phighvt w=420000u l=180000u
+  ad=1.701e+11p pd=1.65e+06u as=0p ps=0u
M1009 a_1870_413# a_877_369# a_1735_329# VPB phighvt w=420000u l=180000u
+  ad=1.302e+11p pd=1.46e+06u as=4.305e+11p ps=4.05e+06u
M1010 a_1655_47# a_1075_413# VGND VNB nshort w=640000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 Q a_2632_47# VGND VNB nshort w=650000u l=150000u
+  ad=1.69e+11p pd=1.82e+06u as=0p ps=0u
M1012 VPWR SCE a_349_21# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1013 a_1735_329# a_693_369# a_1652_329# VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=1.974e+11p ps=2.15e+06u
M1014 a_1735_329# SET_B VPWR VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1015 VGND CLK a_693_369# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1016 a_877_369# a_693_369# VGND VNB nshort w=420000u l=150000u
+  ad=1.218e+11p pd=1.42e+06u as=0p ps=0u
M1017 VPWR a_1930_295# a_1870_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_1467_47# a_1075_413# a_1219_21# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.512e+11p ps=1.56e+06u
M1019 a_27_369# a_349_21# a_199_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR SET_B a_1219_21# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_1177_47# a_877_369# a_1075_413# VNB nshort w=420000u l=150000u
+  ad=8.82e+10p pd=1.26e+06u as=1.344e+11p ps=1.48e+06u
M1022 VGND SET_B a_1467_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_877_369# a_693_369# VPWR VPB phighvt w=640000u l=180000u
+  ad=1.728e+11p pd=1.82e+06u as=0p ps=0u
M1024 a_199_47# SCE a_109_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.96e+06u as=1.26e+11p ps=1.44e+06u
M1025 VGND a_1219_21# a_1177_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1026 Q_N a_1735_329# VGND VNB nshort w=650000u l=150000u
+  ad=2.015e+11p pd=1.92e+06u as=0p ps=0u
M1027 a_1075_413# a_693_369# a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1028 a_295_47# D a_199_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_1652_329# a_1075_413# VPWR VPB phighvt w=840000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1030 VPWR a_1735_329# a_2632_47# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1031 a_211_369# SCE VPWR VPB phighvt w=640000u l=180000u
+  ad=1.472e+11p pd=1.74e+06u as=0p ps=0u
M1032 Q_N a_1735_329# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=2.7e+11p pd=2.54e+06u as=0p ps=0u
M1033 a_109_47# SCD VGND VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_2049_47# a_1930_295# a_1977_47# VNB nshort w=420000u l=150000u
+  ad=2.688e+11p pd=2.12e+06u as=8.82e+10p ps=1.26e+06u
M1035 VGND a_1735_329# a_2632_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=1.302e+11p ps=1.46e+06u
M1036 a_199_47# D a_211_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1037 a_1169_413# a_693_369# a_1075_413# VPB phighvt w=420000u l=180000u
+  ad=1.596e+11p pd=1.6e+06u as=0p ps=0u
M1038 VPWR a_1219_21# a_1169_413# VPB phighvt w=420000u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1039 VGND SET_B a_2049_47# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1040 VPWR CLK a_693_369# VPB phighvt w=640000u l=180000u
+  ad=0p pd=0u as=1.728e+11p ps=1.82e+06u
M1041 a_1977_47# a_693_369# a_1735_329# VNB nshort w=420000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends

