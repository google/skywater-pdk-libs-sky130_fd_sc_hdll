* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__muxb4to1_4 D[3] D[2] D[1] D[0] S[3] S[2] S[1] S[0] VGND
+ VNB VPB VPWR Z
X0 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X1 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X2 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X5 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 a_559_265# S[0] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_3135_265# S[2] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X9 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X10 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X11 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 VGND D[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_3135_265# S[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X16 VGND S[3] a_4006_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X17 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X18 a_1430_325# S[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X19 Z S[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X20 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X21 VPWR S[2] a_3135_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X22 VGND S[0] a_559_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X23 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X24 a_1693_66# D[1] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 a_4006_325# S[3] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X26 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X28 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_559_265# S[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X30 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X31 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X32 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X33 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X34 VPWR S[3] a_4006_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X35 VGND D[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X36 VPWR D[0] a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X37 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X38 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X39 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X40 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X41 VGND S[1] a_1430_325# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X42 a_1643_311# a_1430_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X43 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X44 Z S[2] a_2695_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X45 VGND S[2] a_3135_265# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X46 a_119_47# S[0] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X47 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X48 a_4269_66# S[3] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X49 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X50 VPWR D[2] a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X51 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X52 VPWR S[1] a_1430_325# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X53 VGND D[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X54 a_2695_47# S[2] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X55 Z S[0] a_119_47# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X56 VGND D[3] a_4269_66# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X57 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X58 a_119_47# D[0] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X59 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X60 VPWR S[0] a_559_265# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X61 Z a_1430_325# a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X62 a_4219_311# a_4006_325# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X63 Z S[1] a_1693_66# VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X64 a_117_297# D[0] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X65 a_2693_297# D[2] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X66 Z a_4006_325# a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X67 VPWR D[3] a_4219_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X68 a_4269_66# D[3] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X69 a_1430_325# S[1] VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X70 a_4219_311# D[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X71 Z a_3135_265# a_2693_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X72 a_1693_66# S[1] Z VNB sky130_fd_pr__nfet_01v8 w=520000u l=150000u
X73 Z a_559_265# a_117_297# VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X74 a_1643_311# D[1] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X75 a_4006_325# S[3] VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X76 a_2695_47# D[2] VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X77 a_2693_297# a_3135_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X78 a_117_297# a_559_265# Z VPB sky130_fd_pr__pfet_01v8_hvt w=820000u l=180000u
X79 VPWR D[1] a_1643_311# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
