* File: sky130_fd_sc_hdll__clkmux2_1.pxi.spice
* Created: Wed Sep  2 08:26:57 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_79_21# N_A_79_21#_M1002_d N_A_79_21#_M1009_d
+ N_A_79_21#_M1011_g N_A_79_21#_c_72_n N_A_79_21#_M1003_g N_A_79_21#_c_73_n
+ N_A_79_21#_c_74_n N_A_79_21#_c_120_p N_A_79_21#_c_75_n N_A_79_21#_c_83_p
+ N_A_79_21#_c_92_p N_A_79_21#_c_88_p PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_79_21#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%S N_S_c_146_n N_S_M1005_g N_S_M1000_g
+ N_S_c_148_n N_S_M1006_g N_S_M1007_g N_S_c_154_n N_S_c_170_n N_S_c_218_p
+ N_S_c_155_n N_S_c_193_p N_S_c_210_p N_S_c_150_n N_S_c_151_n S S
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_1%S
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A1 N_A1_M1002_g N_A1_c_240_n N_A1_M1004_g
+ N_A1_c_241_n N_A1_c_242_n N_A1_c_255_n N_A1_c_257_n A1 A1
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A1
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A0 N_A0_c_311_n N_A0_M1009_g N_A0_c_312_n
+ N_A0_c_313_n N_A0_M1001_g N_A0_c_308_n A0 N_A0_c_309_n N_A0_c_310_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A0
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_649_21# N_A_649_21#_M1007_d
+ N_A_649_21#_M1006_d N_A_649_21#_M1008_g N_A_649_21#_c_358_n
+ N_A_649_21#_c_367_n N_A_649_21#_M1010_g N_A_649_21#_c_359_n
+ N_A_649_21#_c_360_n N_A_649_21#_c_361_n N_A_649_21#_c_362_n
+ N_A_649_21#_c_363_n N_A_649_21#_c_368_n N_A_649_21#_c_364_n
+ N_A_649_21#_c_365_n PM_SKY130_FD_SC_HDLL__CLKMUX2_1%A_649_21#
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%X N_X_M1011_s N_X_M1003_s N_X_c_426_n X X X
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_1%X
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VPWR N_VPWR_M1003_d N_VPWR_M1010_d
+ N_VPWR_c_443_n N_VPWR_c_444_n N_VPWR_c_445_n N_VPWR_c_446_n VPWR
+ N_VPWR_c_447_n N_VPWR_c_442_n N_VPWR_c_449_n
+ PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VGND N_VGND_M1011_d N_VGND_M1008_d
+ N_VGND_c_496_n VGND N_VGND_c_497_n N_VGND_c_498_n N_VGND_c_499_n
+ N_VGND_c_500_n N_VGND_c_501_n PM_SKY130_FD_SC_HDLL__CLKMUX2_1%VGND
cc_1 VNB N_A_79_21#_M1011_g 0.0278942f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_2 VNB N_A_79_21#_c_72_n 0.0286882f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_A_79_21#_c_73_n 0.00195867f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_4 VNB N_A_79_21#_c_74_n 0.0193296f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.74
cc_5 VNB N_A_79_21#_c_75_n 0.0051489f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.955
cc_6 VNB N_S_c_146_n 0.0252834f $X=-0.19 $Y=-0.24 $X2=1.735 $Y2=0.235
cc_7 VNB N_S_M1000_g 0.0320387f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_S_c_148_n 0.0209544f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_9 VNB N_S_M1007_g 0.0335245f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_10 VNB N_S_c_150_n 5.74134e-19 $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=2.04
cc_11 VNB N_S_c_151_n 0.0037048f $X=-0.19 $Y=-0.24 $X2=2.67 $Y2=2.04
cc_12 VNB N_A1_M1002_g 0.0228368f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A1_c_240_n 0.0236121f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A1_c_241_n 0.00497376f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A1_c_242_n 0.0376981f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB A1 0.00997405f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_17 VNB N_A0_M1001_g 0.0254644f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_18 VNB N_A0_c_308_n 0.00955013f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_19 VNB N_A0_c_309_n 0.028761f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_20 VNB N_A0_c_310_n 0.00455985f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_21 VNB N_A_649_21#_M1008_g 0.02497f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_22 VNB N_A_649_21#_c_358_n 0.0070328f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_23 VNB N_A_649_21#_c_359_n 5.32232e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_649_21#_c_360_n 0.0308747f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.74
cc_25 VNB N_A_649_21#_c_361_n 0.00551271f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.825
cc_26 VNB N_A_649_21#_c_362_n 8.46441e-19 $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.955
cc_27 VNB N_A_649_21#_c_363_n 0.0158392f $X=-0.19 $Y=-0.24 $X2=2.67 $Y2=2.04
cc_28 VNB N_A_649_21#_c_364_n 0.0211382f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_649_21#_c_365_n 0.0166335f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.0472201f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_31 VNB N_VPWR_c_442_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_496_n 0.00309635f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.495
cc_33 VNB N_VGND_c_497_n 0.0151047f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_34 VNB N_VGND_c_498_n 0.0718072f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_499_n 0.0249556f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_VGND_c_500_n 0.24491f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.54
cc_37 VNB N_VGND_c_501_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0.565 $Y2=1.16
cc_38 VPB N_A_79_21#_c_72_n 0.0322083f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_39 VPB N_A_79_21#_c_73_n 0.0024294f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_40 VPB N_A_79_21#_c_75_n 0.00429564f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.955
cc_41 VPB N_S_c_146_n 0.0329644f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.235
cc_42 VPB N_S_c_148_n 0.0330042f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=0.495
cc_43 VPB N_S_c_154_n 0.0014488f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_44 VPB N_S_c_155_n 6.63611e-19 $X=-0.19 $Y=1.305 $X2=1.435 $Y2=0.74
cc_45 VPB N_S_c_150_n 6.16925e-19 $X=-0.19 $Y=1.305 $X2=1.61 $Y2=2.04
cc_46 VPB N_S_c_151_n 0.00125389f $X=-0.19 $Y=1.305 $X2=2.67 $Y2=2.04
cc_47 VPB S 0.00455426f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_48 VPB N_A1_c_240_n 0.0304527f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB N_A1_c_241_n 0.00280866f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB A1 0.00558813f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_51 VPB N_A0_c_311_n 0.020637f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.235
cc_52 VPB N_A0_c_312_n 0.0406981f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_53 VPB N_A0_c_313_n 0.00988758f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_54 VPB N_A0_c_308_n 8.40892e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB N_A0_c_310_n 0.0023903f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_56 VPB N_A_649_21#_c_358_n 0.00378234f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_57 VPB N_A_649_21#_c_367_n 0.0224682f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_58 VPB N_A_649_21#_c_368_n 0.0267191f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_59 VPB N_A_649_21#_c_364_n 0.0225129f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_60 VPB N_X_c_426_n 0.0065071f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB X 0.00942252f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_62 VPB X 0.0315701f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_63 VPB N_VPWR_c_443_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_64 VPB N_VPWR_c_444_n 0.00497347f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_65 VPB N_VPWR_c_445_n 0.0654208f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.74
cc_66 VPB N_VPWR_c_446_n 0.00439107f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.825
cc_67 VPB N_VPWR_c_447_n 0.0232568f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_68 VPB N_VPWR_c_442_n 0.0505956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_449_n 0.0226539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 N_A_79_21#_c_72_n N_S_c_146_n 0.0375189f $X=0.495 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_71 N_A_79_21#_c_73_n N_S_c_146_n 0.00107569f $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_72 N_A_79_21#_c_74_n N_S_c_146_n 0.00246858f $X=1.435 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_73 N_A_79_21#_c_75_n N_S_c_146_n 0.00361956f $X=1.525 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_79_21#_c_83_p N_S_c_146_n 6.54365e-19 $X=1.61 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_79_21#_M1011_g N_S_M1000_g 0.013677f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_73_n N_S_M1000_g 0.00297788f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_74_n N_S_M1000_g 0.0133748f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_75_n N_S_M1000_g 0.00343808f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_88_p N_S_M1000_g 0.00670281f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_72_n N_S_c_154_n 0.00114678f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_81 N_A_79_21#_M1009_d N_S_c_170_n 0.02385f $X=1.81 $Y=1.545 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_83_p N_S_c_170_n 0.0100943f $X=1.61 $Y=2.04 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_92_p N_S_c_170_n 0.0768599f $X=2.67 $Y=2.04 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_72_n N_S_c_151_n 0.00110986f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_73_n N_S_c_151_n 0.014361f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_74_n N_S_c_151_n 0.0211311f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_75_n N_S_c_151_n 0.0573317f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_75_n N_A1_M1002_g 2.53446e-19 $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_88_p N_A1_M1002_g 0.0200883f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_92_p N_A1_c_240_n 0.00495514f $X=2.67 $Y=2.04 $X2=0 $Y2=0
cc_91 N_A_79_21#_M1009_d N_A1_c_241_n 0.00263273f $X=1.81 $Y=1.545 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_75_n N_A1_c_241_n 0.053476f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_88_p N_A1_c_241_n 0.0138811f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_75_n N_A1_c_242_n 0.0072307f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_88_p N_A1_c_242_n 0.00134275f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_96 N_A_79_21#_M1009_d N_A1_c_255_n 0.0262928f $X=1.81 $Y=1.545 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_92_p N_A1_c_255_n 0.0639496f $X=2.67 $Y=2.04 $X2=0 $Y2=0
cc_98 N_A_79_21#_M1009_d N_A1_c_257_n 9.09665e-19 $X=1.81 $Y=1.545 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_92_p N_A1_c_257_n 0.00891696f $X=2.67 $Y=2.04 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_75_n N_A0_c_311_n 0.00341414f $X=1.525 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_101 N_A_79_21#_c_92_p N_A0_c_311_n 0.0138951f $X=2.67 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_102 N_A_79_21#_c_92_p N_A0_c_312_n 0.00104228f $X=2.67 $Y=2.04 $X2=0 $Y2=0
cc_103 N_A_79_21#_c_75_n N_A0_c_313_n 0.00178945f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_104 N_A_79_21#_c_88_p N_A0_c_313_n 3.50172e-19 $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_88_p N_A0_M1001_g 0.00400095f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_88_p N_A0_c_310_n 0.0174928f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_72_n N_X_c_426_n 0.00293198f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_79_21#_M1011_g X 0.0197284f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_72_n X 0.00327243f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_73_n X 0.0368837f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_120_p X 0.00993354f $X=0.685 $Y=0.74 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_72_n X 0.00974701f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_72_n N_VPWR_c_443_n 0.00846335f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_73_n N_VPWR_c_443_n 0.00331775f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_74_n N_VPWR_c_443_n 0.00388597f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_116 N_A_79_21#_M1009_d N_VPWR_c_442_n 0.00817943f $X=1.81 $Y=1.545 $X2=0
+ $Y2=0
cc_117 N_A_79_21#_c_72_n N_VPWR_c_442_n 0.0131124f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_72_n N_VPWR_c_449_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_75_n A_243_309# 0.00526835f $X=1.525 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_79_21#_c_83_p A_243_309# 0.00300196f $X=1.61 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_79_21#_c_74_n N_VGND_M1011_d 0.00244694f $X=1.435 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_79_21#_c_120_p N_VGND_M1011_d 8.75693e-19 $X=0.685 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_123 N_A_79_21#_M1011_g N_VGND_c_496_n 0.00910743f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_124 N_A_79_21#_c_72_n N_VGND_c_496_n 5.28725e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_74_n N_VGND_c_496_n 0.0160584f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_120_p N_VGND_c_496_n 0.00929542f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_127 N_A_79_21#_c_88_p N_VGND_c_496_n 0.00815458f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_128 N_A_79_21#_M1011_g N_VGND_c_497_n 0.0046653f $X=0.47 $Y=0.495 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_74_n N_VGND_c_498_n 0.00916117f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_88_p N_VGND_c_498_n 0.0313996f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_131 N_A_79_21#_M1002_d N_VGND_c_500_n 0.0122932f $X=1.735 $Y=0.235 $X2=0
+ $Y2=0
cc_132 N_A_79_21#_M1011_g N_VGND_c_500_n 0.00895857f $X=0.47 $Y=0.495 $X2=0
+ $Y2=0
cc_133 N_A_79_21#_c_74_n N_VGND_c_500_n 0.0152428f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_120_p N_VGND_c_500_n 8.0899e-19 $X=0.685 $Y=0.74 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_88_p N_VGND_c_500_n 0.0191349f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_88_p A_245_47# 0.00646653f $X=1.525 $Y=0.54 $X2=-0.19
+ $Y2=-0.24
cc_137 N_S_M1000_g N_A1_M1002_g 0.0156947f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_138 N_S_c_170_n N_A1_c_240_n 0.0140173f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_139 N_S_c_155_n N_A1_c_240_n 3.3557e-19 $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_140 N_S_c_146_n N_A1_c_242_n 0.0156947f $X=1.125 $Y=1.47 $X2=0 $Y2=0
cc_141 N_S_c_151_n N_A1_c_242_n 2.95407e-19 $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_142 N_S_c_170_n N_A1_c_255_n 0.00421347f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_143 N_S_c_155_n A1 0.0117446f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_144 N_S_c_146_n N_A0_c_311_n 0.0291584f $X=1.125 $Y=1.47 $X2=-0.19 $Y2=-0.24
cc_145 N_S_c_170_n N_A0_c_311_n 0.0135571f $X=3.245 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_146 N_S_c_146_n N_A0_c_313_n 0.00409565f $X=1.125 $Y=1.47 $X2=0 $Y2=0
cc_147 N_S_M1007_g N_A_649_21#_M1008_g 0.0166525f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_148 N_S_c_148_n N_A_649_21#_c_358_n 0.00791167f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_149 N_S_c_150_n N_A_649_21#_c_358_n 0.00114571f $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_150 N_S_c_148_n N_A_649_21#_c_367_n 0.0253237f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_151 N_S_c_170_n N_A_649_21#_c_367_n 0.00665392f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_152 N_S_c_155_n N_A_649_21#_c_367_n 0.00936369f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_153 N_S_c_193_p N_A_649_21#_c_367_n 0.0169742f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_154 N_S_c_150_n N_A_649_21#_c_367_n 9.61528e-19 $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_155 S N_A_649_21#_c_367_n 0.00468862f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_156 N_S_c_148_n N_A_649_21#_c_359_n 4.2108e-19 $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_157 N_S_M1007_g N_A_649_21#_c_359_n 0.00105012f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_158 N_S_c_155_n N_A_649_21#_c_359_n 0.00529971f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_159 N_S_c_150_n N_A_649_21#_c_359_n 0.00549551f $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_160 S N_A_649_21#_c_359_n 0.00442941f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_161 N_S_c_148_n N_A_649_21#_c_360_n 0.0078874f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_162 N_S_M1007_g N_A_649_21#_c_360_n 0.00773768f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_163 N_S_c_150_n N_A_649_21#_c_360_n 4.28614e-19 $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_164 S N_A_649_21#_c_360_n 0.00155646f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_165 N_S_c_148_n N_A_649_21#_c_361_n 0.00210123f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_166 N_S_M1007_g N_A_649_21#_c_361_n 0.0151946f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_167 N_S_c_150_n N_A_649_21#_c_361_n 0.0131349f $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_168 S N_A_649_21#_c_361_n 0.00986081f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_169 N_S_c_148_n N_A_649_21#_c_368_n 0.00747341f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_170 N_S_c_210_p N_A_649_21#_c_368_n 6.43652e-19 $X=3.9 $Y=1.44 $X2=0 $Y2=0
cc_171 N_S_c_148_n N_A_649_21#_c_364_n 0.0171101f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_172 N_S_M1007_g N_A_649_21#_c_364_n 0.00462428f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_173 N_S_c_210_p N_A_649_21#_c_364_n 0.0123401f $X=3.9 $Y=1.44 $X2=0 $Y2=0
cc_174 N_S_c_150_n N_A_649_21#_c_364_n 0.0228671f $X=3.89 $Y=1.22 $X2=0 $Y2=0
cc_175 S N_VPWR_M1010_d 0.00577639f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_176 N_S_c_146_n N_VPWR_c_443_n 0.00992112f $X=1.125 $Y=1.47 $X2=0 $Y2=0
cc_177 N_S_c_154_n N_VPWR_c_443_n 0.041629f $X=1.17 $Y=2.295 $X2=0 $Y2=0
cc_178 N_S_c_218_p N_VPWR_c_443_n 0.00976338f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_179 N_S_c_148_n N_VPWR_c_444_n 0.00324489f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_180 N_S_c_170_n N_VPWR_c_444_n 0.0136491f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_181 N_S_c_193_p N_VPWR_c_444_n 0.0330344f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_182 S N_VPWR_c_444_n 0.0129774f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_183 N_S_c_146_n N_VPWR_c_445_n 0.00482335f $X=1.125 $Y=1.47 $X2=0 $Y2=0
cc_184 N_S_c_170_n N_VPWR_c_445_n 0.127998f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_185 N_S_c_218_p N_VPWR_c_445_n 0.0118049f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_186 N_S_c_148_n N_VPWR_c_447_n 0.00673617f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_187 N_S_c_146_n N_VPWR_c_442_n 0.0080749f $X=1.125 $Y=1.47 $X2=0 $Y2=0
cc_188 N_S_c_148_n N_VPWR_c_442_n 0.0130085f $X=3.915 $Y=1.47 $X2=0 $Y2=0
cc_189 N_S_c_170_n N_VPWR_c_442_n 0.077726f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_190 N_S_c_218_p N_VPWR_c_442_n 0.00702939f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_191 N_S_c_170_n A_243_309# 0.0111518f $X=3.245 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_192 N_S_c_170_n A_599_309# 0.00646556f $X=3.245 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_193 N_S_M1000_g N_VGND_c_496_n 0.00593008f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_194 N_S_M1000_g N_VGND_c_498_n 0.00428022f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_195 N_S_M1007_g N_VGND_c_498_n 0.00646436f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_196 N_S_M1007_g N_VGND_c_499_n 0.00433717f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_197 N_S_M1000_g N_VGND_c_500_n 0.00672742f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_198 N_S_M1007_g N_VGND_c_500_n 0.00761805f $X=3.94 $Y=0.495 $X2=0 $Y2=0
cc_199 N_A1_c_241_n N_A0_c_311_n 0.00409325f $X=1.865 $Y=0.975 $X2=-0.19
+ $Y2=-0.24
cc_200 N_A1_c_257_n N_A0_c_311_n 0.00649866f $X=1.95 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_201 N_A1_c_240_n N_A0_c_312_n 0.00277644f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_202 N_A1_c_241_n N_A0_c_312_n 0.0101853f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_203 N_A1_c_255_n N_A0_c_312_n 0.016411f $X=2.785 $Y=1.7 $X2=0 $Y2=0
cc_204 A1 N_A0_c_312_n 0.00120799f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_205 N_A1_c_241_n N_A0_c_313_n 0.0020234f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_206 N_A1_c_242_n N_A0_c_313_n 0.0288992f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_207 N_A1_M1002_g N_A0_M1001_g 0.0106523f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A1_c_241_n N_A0_M1001_g 2.42785e-19 $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_209 A1 N_A0_M1001_g 0.00248702f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_210 N_A1_c_240_n N_A0_c_308_n 0.00936614f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_211 A1 N_A0_c_308_n 2.12428e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_212 N_A1_c_240_n N_A0_c_309_n 0.00503691f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_213 N_A1_c_241_n N_A0_c_309_n 0.00486025f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_214 N_A1_c_242_n N_A0_c_309_n 0.0169793f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_215 N_A1_c_255_n N_A0_c_309_n 2.70133e-19 $X=2.785 $Y=1.7 $X2=0 $Y2=0
cc_216 A1 N_A0_c_309_n 0.00144026f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_217 N_A1_M1002_g N_A0_c_310_n 9.93793e-19 $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_218 N_A1_c_240_n N_A0_c_310_n 0.00240846f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_219 N_A1_c_241_n N_A0_c_310_n 0.0256133f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_220 N_A1_c_242_n N_A0_c_310_n 9.69032e-19 $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_221 N_A1_c_255_n N_A0_c_310_n 0.0231818f $X=2.785 $Y=1.7 $X2=0 $Y2=0
cc_222 A1 N_A0_c_310_n 0.0929962f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_223 A1 N_A_649_21#_M1008_g 0.0260542f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_224 N_A1_c_240_n N_A_649_21#_c_367_n 0.0556404f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_225 N_A1_c_255_n N_A_649_21#_c_367_n 6.59428e-19 $X=2.785 $Y=1.7 $X2=0 $Y2=0
cc_226 A1 N_A_649_21#_c_367_n 5.7392e-19 $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_227 A1 N_A_649_21#_c_359_n 0.0179199f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_228 N_A1_c_240_n N_A_649_21#_c_360_n 0.0213383f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_229 A1 N_A_649_21#_c_362_n 0.0105375f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_230 N_A1_c_240_n N_VPWR_c_445_n 0.00429453f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_231 N_A1_c_240_n N_VPWR_c_442_n 0.0073872f $X=2.905 $Y=1.47 $X2=0 $Y2=0
cc_232 N_A1_c_255_n A_599_309# 0.0019065f $X=2.785 $Y=1.7 $X2=-0.19 $Y2=-0.24
cc_233 A1 A_599_309# 5.87758e-19 $X=2.905 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_234 N_A1_M1002_g N_VGND_c_498_n 0.00357668f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_235 A1 N_VGND_c_498_n 0.041242f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_236 N_A1_M1002_g N_VGND_c_500_n 0.00602486f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_237 N_A1_c_242_n N_VGND_c_500_n 0.00164284f $X=1.865 $Y=0.975 $X2=0 $Y2=0
cc_238 A1 N_VGND_c_500_n 0.0110914f $X=2.905 $Y=0.765 $X2=0 $Y2=0
cc_239 A1 A_478_47# 0.0167701f $X=2.905 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_240 N_A0_c_311_n N_VPWR_c_445_n 0.00429453f $X=1.72 $Y=1.47 $X2=0 $Y2=0
cc_241 N_A0_c_311_n N_VPWR_c_442_n 0.00774138f $X=1.72 $Y=1.47 $X2=0 $Y2=0
cc_242 N_A0_M1001_g N_VGND_c_498_n 0.00435091f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_243 N_A0_c_310_n N_VGND_c_498_n 0.0205158f $X=2.375 $Y=0.98 $X2=0 $Y2=0
cc_244 N_A0_M1001_g N_VGND_c_500_n 0.00904666f $X=2.315 $Y=0.445 $X2=0 $Y2=0
cc_245 N_A0_c_310_n N_VGND_c_500_n 0.0119866f $X=2.375 $Y=0.98 $X2=0 $Y2=0
cc_246 N_A0_c_310_n A_478_47# 0.00656391f $X=2.375 $Y=0.98 $X2=-0.19 $Y2=-0.24
cc_247 N_A_649_21#_c_367_n N_VPWR_c_444_n 0.00744201f $X=3.345 $Y=1.47 $X2=0
+ $Y2=0
cc_248 N_A_649_21#_c_367_n N_VPWR_c_445_n 0.00459563f $X=3.345 $Y=1.47 $X2=0
+ $Y2=0
cc_249 N_A_649_21#_c_368_n N_VPWR_c_447_n 0.0259839f $X=4.15 $Y=2 $X2=0 $Y2=0
cc_250 N_A_649_21#_M1006_d N_VPWR_c_442_n 0.00233913f $X=4.005 $Y=1.545 $X2=0
+ $Y2=0
cc_251 N_A_649_21#_c_367_n N_VPWR_c_442_n 0.00704825f $X=3.345 $Y=1.47 $X2=0
+ $Y2=0
cc_252 N_A_649_21#_c_368_n N_VPWR_c_442_n 0.0151509f $X=4.15 $Y=2 $X2=0 $Y2=0
cc_253 N_A_649_21#_c_361_n N_VGND_M1008_d 0.00234003f $X=4.035 $Y=0.78 $X2=0
+ $Y2=0
cc_254 N_A_649_21#_M1008_g N_VGND_c_498_n 0.023697f $X=3.32 $Y=0.445 $X2=0 $Y2=0
cc_255 N_A_649_21#_c_360_n N_VGND_c_498_n 6.87788e-19 $X=3.41 $Y=1.02 $X2=0
+ $Y2=0
cc_256 N_A_649_21#_c_361_n N_VGND_c_498_n 0.0210008f $X=4.035 $Y=0.78 $X2=0
+ $Y2=0
cc_257 N_A_649_21#_c_362_n N_VGND_c_498_n 0.0115145f $X=3.495 $Y=0.78 $X2=0
+ $Y2=0
cc_258 N_A_649_21#_c_361_n N_VGND_c_499_n 0.00345018f $X=4.035 $Y=0.78 $X2=0
+ $Y2=0
cc_259 N_A_649_21#_c_363_n N_VGND_c_499_n 0.0157596f $X=4.15 $Y=0.455 $X2=0
+ $Y2=0
cc_260 N_A_649_21#_c_365_n N_VGND_c_499_n 0.00189167f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_261 N_A_649_21#_M1007_d N_VGND_c_500_n 0.00218371f $X=4.015 $Y=0.235 $X2=0
+ $Y2=0
cc_262 N_A_649_21#_M1008_g N_VGND_c_500_n 0.00251647f $X=3.32 $Y=0.445 $X2=0
+ $Y2=0
cc_263 N_A_649_21#_c_361_n N_VGND_c_500_n 0.00766116f $X=4.035 $Y=0.78 $X2=0
+ $Y2=0
cc_264 N_A_649_21#_c_362_n N_VGND_c_500_n 7.21038e-19 $X=3.495 $Y=0.78 $X2=0
+ $Y2=0
cc_265 N_A_649_21#_c_363_n N_VGND_c_500_n 0.0093388f $X=4.15 $Y=0.455 $X2=0
+ $Y2=0
cc_266 N_A_649_21#_c_365_n N_VGND_c_500_n 0.00302259f $X=4.21 $Y=0.78 $X2=0
+ $Y2=0
cc_267 N_X_c_426_n N_VPWR_c_443_n 0.0587634f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_268 N_X_M1003_s N_VPWR_c_442_n 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_269 X N_VPWR_c_442_n 0.0126651f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_270 X N_VPWR_c_449_n 0.021418f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_271 X N_VGND_c_497_n 0.0176426f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_272 N_X_M1011_s N_VGND_c_500_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_273 X N_VGND_c_500_n 0.00974347f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_274 N_VPWR_c_442_n A_243_309# 0.003342f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_275 N_VPWR_c_442_n A_599_309# 0.00208801f $X=4.37 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_276 N_VGND_c_500_n A_245_47# 0.00371776f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_277 N_VGND_c_500_n A_478_47# 0.0188707f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
