* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__buf_12 A VGND VNB VPB VPWR X
M1000 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=2.61e+12p pd=2.322e+07u as=1.74e+12p ps=1.548e+07u
M1001 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=5.8e+11p ps=5.16e+06u
M1002 VGND A a_117_297# VNB nshort w=650000u l=150000u
+  ad=1.82e+12p pd=1.73e+07u as=4.16e+11p ps=3.88e+06u
M1003 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1004 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1005 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1006 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=1.2805e+12p ps=1.174e+07u
M1007 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1008 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1009 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1013 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1014 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1016 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 VPWR A a_117_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1020 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1021 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1022 VGND A a_117_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1023 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1024 VGND a_117_297# X VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1025 VPWR a_117_297# X VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1026 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1027 a_117_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1028 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1029 X a_117_297# VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1030 X a_117_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1031 a_117_297# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
.ends
