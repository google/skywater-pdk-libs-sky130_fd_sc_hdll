# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdlclkp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdlclkp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.455700 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.055000 1.075000 5.345000 1.120000 ;
        RECT 5.055000 1.120000 6.390000 1.260000 ;
        RECT 5.055000 1.260000 5.345000 1.305000 ;
        RECT 6.100000 1.075000 6.390000 1.120000 ;
        RECT 6.100000 1.260000 6.390000 1.305000 ;
    END
  END CLK
  PIN GATE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.905000 0.955000 1.295000 1.445000 ;
        RECT 0.905000 1.445000 1.340000 1.955000 ;
    END
  END GATE
  PIN GCLK
    ANTENNADIFFAREA  1.251250 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.000000 0.255000 7.380000 0.445000 ;
        RECT 7.130000 0.445000 7.380000 0.715000 ;
        RECT 7.130000 0.715000 7.820000 0.885000 ;
        RECT 7.130000 1.485000 7.820000 1.655000 ;
        RECT 7.130000 1.655000 7.380000 2.465000 ;
        RECT 7.650000 0.885000 7.820000 1.055000 ;
        RECT 7.650000 1.055000 9.055000 1.315000 ;
        RECT 7.650000 1.315000 7.820000 1.485000 ;
        RECT 8.205000 0.255000 8.595000 1.055000 ;
        RECT 8.205000 1.315000 8.595000 2.465000 ;
    END
  END GCLK
  PIN SCE
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.955000 0.345000 1.665000 ;
    END
  END SCE
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 9.390000 2.910000 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 9.200000 0.085000 ;
      RECT 0.000000  2.635000 9.200000 2.805000 ;
      RECT 0.085000  0.255000 0.345000 0.615000 ;
      RECT 0.085000  0.615000 1.295000 0.785000 ;
      RECT 0.085000  1.835000 0.345000 2.635000 ;
      RECT 0.515000  0.085000 0.895000 0.445000 ;
      RECT 0.515000  0.785000 0.735000 2.125000 ;
      RECT 0.515000  2.125000 1.360000 2.465000 ;
      RECT 1.115000  0.255000 1.295000 0.615000 ;
      RECT 1.465000  0.255000 2.700000 0.535000 ;
      RECT 1.465000  0.705000 1.855000 1.205000 ;
      RECT 1.465000  1.205000 2.015000 1.325000 ;
      RECT 1.510000  1.325000 2.015000 1.955000 ;
      RECT 1.530000  2.125000 2.405000 2.465000 ;
      RECT 2.025000  0.705000 2.360000 1.035000 ;
      RECT 2.235000  1.205000 3.265000 1.375000 ;
      RECT 2.235000  1.375000 2.405000 2.125000 ;
      RECT 2.530000  0.535000 2.700000 0.995000 ;
      RECT 2.530000  0.995000 3.265000 1.205000 ;
      RECT 2.575000  1.575000 2.795000 1.635000 ;
      RECT 2.575000  1.635000 3.705000 1.905000 ;
      RECT 2.575000  2.075000 3.265000 2.635000 ;
      RECT 2.920000  0.085000 3.265000 0.825000 ;
      RECT 3.485000  0.255000 3.705000 1.635000 ;
      RECT 3.485000  1.905000 3.705000 1.915000 ;
      RECT 3.485000  1.915000 5.915000 2.085000 ;
      RECT 3.485000  2.085000 3.705000 2.465000 ;
      RECT 3.895000  0.255000 4.225000 0.765000 ;
      RECT 3.895000  0.765000 4.320000 0.935000 ;
      RECT 3.895000  0.935000 4.065000 1.575000 ;
      RECT 3.895000  1.575000 4.305000 1.745000 ;
      RECT 3.895000  2.255000 5.915000 2.635000 ;
      RECT 4.235000  1.105000 4.830000 1.275000 ;
      RECT 4.395000  0.085000 4.775000 0.445000 ;
      RECT 4.525000  1.275000 4.830000 1.495000 ;
      RECT 4.525000  1.495000 5.375000 1.745000 ;
      RECT 4.540000  0.615000 5.245000 0.785000 ;
      RECT 4.540000  0.785000 4.830000 1.105000 ;
      RECT 4.995000  0.255000 5.245000 0.615000 ;
      RECT 5.055000  0.995000 5.345000 1.325000 ;
      RECT 5.415000  0.255000 5.835000 0.615000 ;
      RECT 5.415000  0.615000 6.910000 0.785000 ;
      RECT 5.565000  0.995000 5.915000 1.915000 ;
      RECT 6.005000  0.085000 6.830000 0.445000 ;
      RECT 6.135000  0.995000 6.565000 1.325000 ;
      RECT 6.135000  1.495000 6.910000 2.085000 ;
      RECT 6.135000  2.085000 6.305000 2.465000 ;
      RECT 6.555000  2.255000 6.885000 2.635000 ;
      RECT 6.740000  0.785000 6.910000 1.055000 ;
      RECT 6.740000  1.055000 7.430000 1.315000 ;
      RECT 6.740000  1.315000 6.910000 1.495000 ;
      RECT 7.600000  0.085000 7.850000 0.545000 ;
      RECT 7.600000  1.825000 7.850000 2.635000 ;
      RECT 8.765000  0.085000 9.035000 0.885000 ;
      RECT 8.765000  1.485000 9.035000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.680000  1.445000 1.850000 1.615000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.190000  0.765000 2.360000 0.935000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.150000  0.765000 4.320000 0.935000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.660000  1.445000 4.830000 1.615000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.115000  1.105000 5.285000 1.275000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.160000  1.105000 6.330000 1.275000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
      RECT 7.505000 -0.085000 7.675000 0.085000 ;
      RECT 7.505000  2.635000 7.675000 2.805000 ;
      RECT 7.965000 -0.085000 8.135000 0.085000 ;
      RECT 7.965000  2.635000 8.135000 2.805000 ;
      RECT 8.425000 -0.085000 8.595000 0.085000 ;
      RECT 8.425000  2.635000 8.595000 2.805000 ;
      RECT 8.885000 -0.085000 9.055000 0.085000 ;
      RECT 8.885000  2.635000 9.055000 2.805000 ;
    LAYER met1 ;
      RECT 1.620000 1.415000 1.910000 1.460000 ;
      RECT 1.620000 1.460000 4.890000 1.600000 ;
      RECT 1.620000 1.600000 1.910000 1.645000 ;
      RECT 2.130000 0.735000 2.420000 0.780000 ;
      RECT 2.130000 0.780000 4.380000 0.920000 ;
      RECT 2.130000 0.920000 2.420000 0.965000 ;
      RECT 4.090000 0.735000 4.380000 0.780000 ;
      RECT 4.090000 0.920000 4.380000 0.965000 ;
      RECT 4.600000 1.415000 4.890000 1.460000 ;
      RECT 4.600000 1.600000 4.890000 1.645000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdlclkp_4
END LIBRARY
