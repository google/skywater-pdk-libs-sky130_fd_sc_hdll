* File: sky130_fd_sc_hdll__a32oi_2.pex.spice
* Created: Wed Sep  2 08:21:02 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%B2 1 3 4 6 7 9 10 12 13 14 15 24 26
c49 15 0 1.31482e-19 $X=0.695 $Y=1.19
r50 24 25 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r51 22 24 33.4905 $w=3.67e-07 $l=2.55e-07 $layer=POLY_cond $X=0.71 $Y=1.202
+ $X2=0.965 $Y2=1.202
r52 20 22 24.9537 $w=3.67e-07 $l=1.9e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.71 $Y2=1.202
r53 19 20 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.52 $Y2=1.202
r54 15 30 19.5411 $w=2.08e-07 $l=3.7e-07 $layer=LI1_cond $X=0.695 $Y=1.18
+ $X2=0.325 $Y2=1.18
r55 15 22 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=0.71
+ $Y=1.16 $X2=0.71 $Y2=1.16
r56 14 26 15.096 $w=1.78e-07 $l=2.45e-07 $layer=LI1_cond $X=0.235 $Y=1.53
+ $X2=0.235 $Y2=1.285
r57 13 26 3.69874 $w=1.8e-07 $l=1.05e-07 $layer=LI1_cond $X=0.235 $Y=1.18
+ $X2=0.235 $Y2=1.285
r58 13 30 3.17035 $w=2.1e-07 $l=9e-08 $layer=LI1_cond $X=0.235 $Y=1.18 $X2=0.325
+ $Y2=1.18
r59 10 25 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r60 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r61 7 24 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r62 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r63 4 20 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=1.202
r64 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r65 1 19 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r66 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%B1 1 3 4 6 7 9 10 12 13 14 22 25
c53 22 0 1.31482e-19 $X=1.905 $Y=1.192
c54 7 0 1.74942e-19 $X=1.905 $Y=1.41
r55 22 23 3.10567 $w=3.88e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.192
+ $X2=1.93 $Y2=1.192
r56 20 22 42.2371 $w=3.88e-07 $l=3.4e-07 $layer=POLY_cond $X=1.565 $Y=1.192
+ $X2=1.905 $Y2=1.192
r57 18 20 16.1495 $w=3.88e-07 $l=1.3e-07 $layer=POLY_cond $X=1.435 $Y=1.192
+ $X2=1.565 $Y2=1.192
r58 17 18 3.10567 $w=3.88e-07 $l=2.5e-08 $layer=POLY_cond $X=1.41 $Y=1.192
+ $X2=1.435 $Y2=1.192
r59 14 20 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.565
+ $Y=1.16 $X2=1.565 $Y2=1.16
r60 13 14 20.0693 $w=2.08e-07 $l=3.8e-07 $layer=LI1_cond $X=1.185 $Y=1.18
+ $X2=1.565 $Y2=1.18
r61 13 25 1.58442 $w=2.08e-07 $l=3e-08 $layer=LI1_cond $X=1.185 $Y=1.18
+ $X2=1.155 $Y2=1.18
r62 10 23 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.93 $Y=0.975
+ $X2=1.93 $Y2=1.192
r63 10 12 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.93 $Y=0.975
+ $X2=1.93 $Y2=0.56
r64 7 22 20.7379 $w=1.8e-07 $l=2.18e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.192
r65 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r66 4 18 20.7379 $w=1.8e-07 $l=2.18e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.192
r67 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r68 1 17 25.1189 $w=1.5e-07 $l=2.17e-07 $layer=POLY_cond $X=1.41 $Y=0.975
+ $X2=1.41 $Y2=1.192
r69 1 3 133.353 $w=1.5e-07 $l=4.15e-07 $layer=POLY_cond $X=1.41 $Y=0.975
+ $X2=1.41 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A1 1 3 4 5 8 10 12 15 17 19 28 29 34 38
c51 28 0 2.96998e-19 $X=3 $Y=1.16
r52 29 30 3.8871 $w=3.1e-07 $l=2.5e-08 $layer=POLY_cond $X=3.265 $Y=1.217
+ $X2=3.29 $Y2=1.217
r53 28 38 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=3 $Y=1.35 $X2=2.995
+ $Y2=1.35
r54 27 29 41.2032 $w=3.1e-07 $l=2.65e-07 $layer=POLY_cond $X=3 $Y=1.217
+ $X2=3.265 $Y2=1.217
r55 27 28 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3 $Y=1.16
+ $X2=3 $Y2=1.16
r56 25 27 20.2129 $w=3.1e-07 $l=1.3e-07 $layer=POLY_cond $X=2.87 $Y=1.217 $X2=3
+ $Y2=1.217
r57 19 38 0.217469 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=2.985 $Y=1.35
+ $X2=2.995 $Y2=1.35
r58 19 34 9.7861 $w=5.48e-07 $l=4.5e-07 $layer=LI1_cond $X=2.985 $Y=1.35
+ $X2=2.535 $Y2=1.35
r59 17 34 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=2.53 $Y=1.35
+ $X2=2.535 $Y2=1.35
r60 13 30 19.7411 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=1.217
r61 13 15 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.29 $Y=1.025
+ $X2=3.29 $Y2=0.56
r62 10 29 15.4789 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.265 $Y=1.41
+ $X2=3.265 $Y2=1.217
r63 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.265 $Y=1.41
+ $X2=3.265 $Y2=1.985
r64 6 25 19.7411 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=1.217
r65 6 8 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.87 $Y=1.025
+ $X2=2.87 $Y2=0.56
r66 4 25 12.5919 $w=3.1e-07 $l=9.94987e-08 $layer=POLY_cond $X=2.795 $Y=1.16
+ $X2=2.87 $Y2=1.217
r67 4 5 71.0956 $w=2.7e-07 $l=3.2e-07 $layer=POLY_cond $X=2.795 $Y=1.16
+ $X2=2.475 $Y2=1.16
r68 1 5 28.3559 $w=2.7e-07 $l=2.95804e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.475 $Y2=1.16
r69 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A2 3 5 7 10 12 14 15 17 27 33 37
c44 37 0 9.24665e-20 $X=4.365 $Y=1.53
r45 27 29 41.3143 $w=3.15e-07 $l=2.7e-07 $layer=POLY_cond $X=4.275 $Y=1.217
+ $X2=4.545 $Y2=1.217
r46 25 27 14.5365 $w=3.15e-07 $l=9.5e-08 $layer=POLY_cond $X=4.18 $Y=1.217
+ $X2=4.275 $Y2=1.217
r47 24 25 68.0921 $w=3.15e-07 $l=4.45e-07 $layer=POLY_cond $X=3.735 $Y=1.217
+ $X2=4.18 $Y2=1.217
r48 23 24 3.8254 $w=3.15e-07 $l=2.5e-08 $layer=POLY_cond $X=3.71 $Y=1.217
+ $X2=3.735 $Y2=1.217
r49 17 37 1.95722 $w=5.48e-07 $l=9e-08 $layer=LI1_cond $X=4.275 $Y=1.35
+ $X2=4.365 $Y2=1.35
r50 17 33 7.82888 $w=5.48e-07 $l=3.6e-07 $layer=LI1_cond $X=4.275 $Y=1.35
+ $X2=3.915 $Y2=1.35
r51 17 27 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.275
+ $Y=1.16 $X2=4.275 $Y2=1.16
r52 15 33 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=3.91 $Y=1.35
+ $X2=3.915 $Y2=1.35
r53 12 29 15.85 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=4.545 $Y=1.41
+ $X2=4.545 $Y2=1.217
r54 12 14 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.545 $Y=1.41
+ $X2=4.545 $Y2=1.985
r55 8 25 20.1192 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=4.18 $Y=1.025
+ $X2=4.18 $Y2=1.217
r56 8 10 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=4.18 $Y=1.025
+ $X2=4.18 $Y2=0.56
r57 5 24 15.85 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=3.735 $Y=1.41
+ $X2=3.735 $Y2=1.217
r58 5 7 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.735 $Y=1.41
+ $X2=3.735 $Y2=1.985
r59 1 23 20.1192 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=3.71 $Y=1.025
+ $X2=3.71 $Y2=1.217
r60 1 3 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=3.71 $Y=1.025
+ $X2=3.71 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A3 1 3 6 8 10 13 15 18 20 21 22 23 30 35
+ 40
r48 37 38 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=6.155
+ $Y=1.16 $X2=6.155 $Y2=1.16
r49 35 37 26.7778 $w=3.33e-07 $l=1.85e-07 $layer=POLY_cond $X=5.97 $Y=1.212
+ $X2=6.155 $Y2=1.212
r50 34 35 3.61862 $w=3.33e-07 $l=2.5e-08 $layer=POLY_cond $X=5.945 $Y=1.212
+ $X2=5.97 $Y2=1.212
r51 33 38 8.48128 $w=5.48e-07 $l=3.9e-07 $layer=LI1_cond $X=5.765 $Y=1.35
+ $X2=6.155 $Y2=1.35
r52 32 33 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=5.765
+ $Y=1.16 $X2=5.765 $Y2=1.16
r53 30 34 16.3411 $w=3.33e-07 $l=1.23288e-07 $layer=POLY_cond $X=5.845 $Y=1.16
+ $X2=5.945 $Y2=1.212
r54 30 32 17.7739 $w=2.7e-07 $l=8e-08 $layer=POLY_cond $X=5.845 $Y=1.16
+ $X2=5.765 $Y2=1.16
r55 22 23 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=6.19 $Y=1.35
+ $X2=6.195 $Y2=1.35
r56 22 38 0.761141 $w=5.48e-07 $l=3.5e-08 $layer=LI1_cond $X=6.19 $Y=1.35
+ $X2=6.155 $Y2=1.35
r57 21 33 0.217469 $w=5.48e-07 $l=1e-08 $layer=LI1_cond $X=5.755 $Y=1.35
+ $X2=5.765 $Y2=1.35
r58 20 21 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=5.75 $Y=1.35
+ $X2=5.755 $Y2=1.35
r59 18 20 9.67736 $w=5.48e-07 $l=4.45e-07 $layer=LI1_cond $X=5.305 $Y=1.35
+ $X2=5.75 $Y2=1.35
r60 18 40 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=5.305 $Y=1.35 $X2=5.3
+ $Y2=1.35
r61 16 17 58.119 $w=3.11e-07 $l=3.75e-07 $layer=POLY_cond $X=5.025 $Y=1.217
+ $X2=5.4 $Y2=1.217
r62 15 32 64.4304 $w=2.7e-07 $l=2.9e-07 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.765 $Y2=1.16
r63 15 17 12.5913 $w=3.11e-07 $l=9.94987e-08 $layer=POLY_cond $X=5.475 $Y=1.16
+ $X2=5.4 $Y2=1.217
r64 11 35 21.4384 $w=1.5e-07 $l=1.97e-07 $layer=POLY_cond $X=5.97 $Y=1.015
+ $X2=5.97 $Y2=1.212
r65 11 13 233.309 $w=1.5e-07 $l=4.55e-07 $layer=POLY_cond $X=5.97 $Y=1.015
+ $X2=5.97 $Y2=0.56
r66 8 34 17.1428 $w=1.8e-07 $l=1.98e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.212
r67 8 10 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.945 $Y=1.41
+ $X2=5.945 $Y2=1.985
r68 4 17 19.8172 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=5.4 $Y=1.025 $X2=5.4
+ $Y2=1.217
r69 4 6 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=5.4 $Y=1.025 $X2=5.4
+ $Y2=0.56
r70 1 16 15.5536 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=5.025 $Y=1.41
+ $X2=5.025 $Y2=1.217
r71 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.025 $Y=1.41
+ $X2=5.025 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_297# 1 2 3 4 5 6 21 23 24 27 29 31 32
+ 33 37 41 45 49 51 53
r79 42 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.865 $Y=1.88
+ $X2=4.78 $Y2=1.88
r80 41 53 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=6.095 $Y=1.88
+ $X2=6.18 $Y2=1.88
r81 41 42 80.246 $w=1.68e-07 $l=1.23e-06 $layer=LI1_cond $X=6.095 $Y=1.88
+ $X2=4.865 $Y2=1.88
r82 38 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.585 $Y=1.88 $X2=3.5
+ $Y2=1.88
r83 37 51 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.695 $Y=1.88
+ $X2=4.78 $Y2=1.88
r84 37 38 72.4171 $w=1.68e-07 $l=1.11e-06 $layer=LI1_cond $X=4.695 $Y=1.88
+ $X2=3.585 $Y2=1.88
r85 34 47 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.225 $Y=1.88
+ $X2=2.14 $Y2=1.88
r86 33 49 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.415 $Y=1.88 $X2=3.5
+ $Y2=1.88
r87 33 34 77.6364 $w=1.68e-07 $l=1.19e-06 $layer=LI1_cond $X=3.415 $Y=1.88
+ $X2=2.225 $Y2=1.88
r88 31 47 3.40825 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.14 $Y=1.965
+ $X2=2.14 $Y2=1.88
r89 31 32 21.5294 $w=1.68e-07 $l=3.3e-07 $layer=LI1_cond $X=2.14 $Y=1.965
+ $X2=2.14 $Y2=2.295
r90 30 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.285 $Y=2.38 $X2=1.2
+ $Y2=2.38
r91 29 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.055 $Y=2.38
+ $X2=2.14 $Y2=2.295
r92 29 30 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=2.055 $Y=2.38
+ $X2=1.285 $Y2=2.38
r93 25 45 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.2 $Y=2.295 $X2=1.2
+ $Y2=2.38
r94 25 27 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.2 $Y=2.295
+ $X2=1.2 $Y2=1.96
r95 23 45 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.115 $Y=2.38 $X2=1.2
+ $Y2=2.38
r96 23 24 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.115 $Y=2.38
+ $X2=0.345 $Y2=2.38
r97 19 24 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.345 $Y2=2.38
r98 19 21 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=2.295
+ $X2=0.26 $Y2=1.96
r99 6 53 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=6.035
+ $Y=1.485 $X2=6.18 $Y2=1.96
r100 5 51 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.635
+ $Y=1.485 $X2=4.78 $Y2=1.96
r101 4 49 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=3.355
+ $Y=1.485 $X2=3.5 $Y2=1.96
r102 3 47 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=1.96
r103 2 27 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.96
r104 1 21 300 $w=1.7e-07 $l=5.33854e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%Y 1 2 3 4 15 17 18 19 25 27 31 33 34 35 36
+ 43 45
c87 43 0 1.92797e-19 $X=2.08 $Y=1.455
r88 42 45 1.25266 $w=2.28e-07 $l=2.5e-08 $layer=LI1_cond $X=2.08 $Y=0.825
+ $X2=2.08 $Y2=0.85
r89 36 43 2.9826 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=1.54 $X2=2.08
+ $Y2=1.455
r90 36 43 0.250531 $w=2.28e-07 $l=5e-09 $layer=LI1_cond $X=2.08 $Y=1.45 $X2=2.08
+ $Y2=1.455
r91 35 36 13.0276 $w=2.28e-07 $l=2.6e-07 $layer=LI1_cond $X=2.08 $Y=1.19
+ $X2=2.08 $Y2=1.45
r92 34 42 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.08 $Y=0.74
+ $X2=2.08 $Y2=0.825
r93 34 35 15.5329 $w=2.28e-07 $l=3.1e-07 $layer=LI1_cond $X=2.08 $Y=0.88
+ $X2=2.08 $Y2=1.19
r94 34 45 1.50319 $w=2.28e-07 $l=3e-08 $layer=LI1_cond $X=2.08 $Y=0.88 $X2=2.08
+ $Y2=0.85
r95 29 34 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.195 $Y=0.74
+ $X2=2.08 $Y2=0.74
r96 29 31 57.738 $w=1.68e-07 $l=8.85e-07 $layer=LI1_cond $X=2.195 $Y=0.74
+ $X2=3.08 $Y2=0.74
r97 28 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.755 $Y=1.54
+ $X2=1.67 $Y2=1.54
r98 27 36 4.03528 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.965 $Y=1.54
+ $X2=2.08 $Y2=1.54
r99 27 28 13.7005 $w=1.68e-07 $l=2.1e-07 $layer=LI1_cond $X=1.965 $Y=1.54
+ $X2=1.755 $Y2=1.54
r100 23 33 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.67 $Y=1.625
+ $X2=1.67 $Y2=1.54
r101 23 25 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=1.67 $Y=1.625
+ $X2=1.67 $Y2=1.96
r102 19 34 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=1.965 $Y=0.74
+ $X2=2.08 $Y2=0.74
r103 19 21 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=1.965 $Y=0.74
+ $X2=1.67 $Y2=0.74
r104 17 33 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.585 $Y=1.54
+ $X2=1.67 $Y2=1.54
r105 17 18 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.585 $Y=1.54
+ $X2=0.895 $Y2=1.54
r106 13 18 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.73 $Y=1.625
+ $X2=0.895 $Y2=1.54
r107 13 15 2.61919 $w=3.28e-07 $l=7.5e-08 $layer=LI1_cond $X=0.73 $Y=1.625
+ $X2=0.73 $Y2=1.7
r108 4 25 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=1.96
r109 3 15 300 $w=1.7e-07 $l=2.78209e-07 $layer=licon1_PDIFF $count=2 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=1.7
r110 2 31 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=2.945
+ $Y=0.235 $X2=3.08 $Y2=0.74
r111 1 21 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=1.485
+ $Y=0.235 $X2=1.67 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%VPWR 1 2 3 10 32 33 37 41 44 48 51 55
r82 53 55 8.3097 $w=5.48e-07 $l=9.5e-08 $layer=LI1_cond $X=5.75 $Y=2.53
+ $X2=5.845 $Y2=2.53
r83 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r84 50 53 1.52228 $w=5.48e-07 $l=7e-08 $layer=LI1_cond $X=5.68 $Y=2.53 $X2=5.75
+ $Y2=2.53
r85 50 51 18.3133 $w=5.48e-07 $l=5.55e-07 $layer=LI1_cond $X=5.68 $Y=2.53
+ $X2=5.125 $Y2=2.53
r86 46 48 9.61451 $w=5.48e-07 $l=1.55e-07 $layer=LI1_cond $X=4.37 $Y=2.53
+ $X2=4.525 $Y2=2.53
r87 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r88 43 46 1.30481 $w=5.48e-07 $l=6e-08 $layer=LI1_cond $X=4.31 $Y=2.53 $X2=4.37
+ $Y2=2.53
r89 43 44 17.9871 $w=5.48e-07 $l=5.4e-07 $layer=LI1_cond $X=4.31 $Y=2.53
+ $X2=3.77 $Y2=2.53
r90 39 41 10.0494 $w=5.48e-07 $l=1.75e-07 $layer=LI1_cond $X=2.99 $Y=2.53
+ $X2=3.165 $Y2=2.53
r91 39 40 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r92 36 39 0.108734 $w=5.48e-07 $l=5e-09 $layer=LI1_cond $X=2.985 $Y=2.53
+ $X2=2.99 $Y2=2.53
r93 36 37 17.9871 $w=5.48e-07 $l=5.4e-07 $layer=LI1_cond $X=2.985 $Y=2.53
+ $X2=2.445 $Y2=2.53
r94 33 54 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=6.21 $Y=2.72
+ $X2=5.75 $Y2=2.72
r95 32 55 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=6.21 $Y=2.72
+ $X2=5.845 $Y2=2.72
r96 32 33 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=2.72
+ $X2=6.21 $Y2=2.72
r97 29 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=5.75 $Y2=2.72
r98 29 47 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.83 $Y=2.72
+ $X2=4.37 $Y2=2.72
r99 28 51 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=5.125 $Y2=2.72
r100 28 48 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.83 $Y=2.72
+ $X2=4.525 $Y2=2.72
r101 28 29 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r102 24 47 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r103 24 40 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.99 $Y2=2.72
r104 23 44 20.877 $w=1.68e-07 $l=3.2e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.77 $Y2=2.72
r105 23 41 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=3.165 $Y2=2.72
r106 23 24 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r107 19 40 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.99 $Y2=2.72
r108 18 37 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.07 $Y=2.72
+ $X2=2.445 $Y2=2.72
r109 18 19 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r110 14 18 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r111 10 19 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=2.07 $Y2=2.72
r112 10 14 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r113 3 50 300 $w=1.7e-07 $l=1.10186e-06 $layer=licon1_PDIFF $count=2 $X=5.115
+ $Y=1.485 $X2=5.68 $Y2=2.34
r114 2 43 300 $w=1.7e-07 $l=1.07037e-06 $layer=licon1_PDIFF $count=2 $X=3.825
+ $Y=1.485 $X2=4.31 $Y2=2.34
r115 1 36 300 $w=1.7e-07 $l=1.08426e-06 $layer=licon1_PDIFF $count=2 $X=2.465
+ $Y=1.485 $X2=2.985 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A_27_47# 1 2 3 12 14 15 16 17 20
r44 18 23 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.285 $Y=0.38
+ $X2=1.16 $Y2=0.38
r45 18 20 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=1.285 $Y=0.38
+ $X2=2.14 $Y2=0.38
r46 17 25 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.715
+ $X2=1.16 $Y2=0.8
r47 16 23 2.89128 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.38
r48 16 17 11.5244 $w=2.48e-07 $l=2.5e-07 $layer=LI1_cond $X=1.16 $Y=0.465
+ $X2=1.16 $Y2=0.715
r49 14 25 4.25188 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=1.16 $Y2=0.8
r50 14 15 39.7968 $w=1.68e-07 $l=6.1e-07 $layer=LI1_cond $X=1.035 $Y=0.8
+ $X2=0.425 $Y2=0.8
r51 10 15 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.425 $Y2=0.8
r52 10 12 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.26 $Y=0.715
+ $X2=0.26 $Y2=0.38
r53 3 20 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.38
r54 2 25 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.72
r55 2 23 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.38
r56 1 12 91 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%VGND 1 2 3 14 16 18 21 27 36 41 45
r67 44 45 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=6.21 $Y=0 $X2=6.21
+ $Y2=0
r68 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r69 39 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.75 $Y=0 $X2=6.21
+ $Y2=0
r70 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r71 36 44 3.40825 $w=1.7e-07 $l=1.72e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=6.267
+ $Y2=0
r72 36 38 22.508 $w=1.68e-07 $l=3.45e-07 $layer=LI1_cond $X=6.095 $Y=0 $X2=5.75
+ $Y2=0
r73 35 39 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r74 34 35 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=4.83 $Y=0
+ $X2=4.83 $Y2=0
r75 32 35 1.04711 $w=4.8e-07 $l=3.68e-06 $layer=MET1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r76 32 42 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=0.69
+ $Y2=0
r77 31 34 240.086 $w=1.68e-07 $l=3.68e-06 $layer=LI1_cond $X=1.15 $Y=0 $X2=4.83
+ $Y2=0
r78 31 32 2.06667 $w=1.7e-07 $l=7.65e-07 $layer=mcon $count=4 $X=1.15 $Y=0
+ $X2=1.15 $Y2=0
r79 29 41 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.815 $Y=0 $X2=0.73
+ $Y2=0
r80 29 31 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=0.815 $Y=0 $X2=1.15
+ $Y2=0
r81 27 42 0.129466 $w=4.8e-07 $l=4.55e-07 $layer=MET1_cond $X=0.235 $Y=0
+ $X2=0.69 $Y2=0
r82 23 38 32.6203 $w=1.68e-07 $l=5e-07 $layer=LI1_cond $X=5.25 $Y=0 $X2=5.75
+ $Y2=0
r83 21 34 2.28342 $w=1.68e-07 $l=3.5e-08 $layer=LI1_cond $X=4.865 $Y=0 $X2=4.83
+ $Y2=0
r84 21 25 11.3748 $w=3.83e-07 $l=3.8e-07 $layer=LI1_cond $X=5.057 $Y=0 $X2=5.057
+ $Y2=0.38
r85 21 23 5.54671 $w=1.7e-07 $l=1.93e-07 $layer=LI1_cond $X=5.057 $Y=0 $X2=5.25
+ $Y2=0
r86 16 44 3.40825 $w=1.7e-07 $l=1.22327e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.267 $Y2=0
r87 16 18 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=6.18 $Y=0.085
+ $X2=6.18 $Y2=0.38
r88 12 41 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0
r89 12 14 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.73 $Y=0.085
+ $X2=0.73 $Y2=0.38
r90 3 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=6.045
+ $Y=0.235 $X2=6.18 $Y2=0.38
r91 2 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=4.91
+ $Y=0.235 $X2=5.035 $Y2=0.38
r92 1 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A_507_47# 1 2 3 16
r19 14 16 58.0642 $w=1.68e-07 $l=8.9e-07 $layer=LI1_cond $X=3.5 $Y=0.38 $X2=4.39
+ $Y2=0.38
r20 11 14 54.8021 $w=1.68e-07 $l=8.4e-07 $layer=LI1_cond $X=2.66 $Y=0.38 $X2=3.5
+ $Y2=0.38
r21 3 16 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=4.255
+ $Y=0.235 $X2=4.39 $Y2=0.38
r22 2 14 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.365
+ $Y=0.235 $X2=3.5 $Y2=0.38
r23 1 11 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.535
+ $Y=0.235 $X2=2.66 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A32OI_2%A_757_47# 1 2 7 12
r26 12 14 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=5.61 $Y=0.36
+ $X2=5.61 $Y2=0.72
r27 7 14 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=5.42 $Y=0.72 $X2=5.61
+ $Y2=0.72
r28 7 9 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=5.42 $Y=0.72 $X2=3.92
+ $Y2=0.72
r29 2 12 91 $w=1.7e-07 $l=2.13542e-07 $layer=licon1_NDIFF $count=2 $X=5.475
+ $Y=0.235 $X2=5.635 $Y2=0.36
r30 1 9 182 $w=1.7e-07 $l=5.48361e-07 $layer=licon1_NDIFF $count=1 $X=3.785
+ $Y=0.235 $X2=3.92 $Y2=0.72
.ends

