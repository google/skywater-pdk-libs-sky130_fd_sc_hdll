* File: sky130_fd_sc_hdll__a21bo_2.pxi.spice
* Created: Thu Aug 27 18:52:10 2020
* 
x_PM_SKY130_FD_SC_HDLL__A21BO_2%A_79_21# N_A_79_21#_M1011_d N_A_79_21#_M1005_s
+ N_A_79_21#_M1004_g N_A_79_21#_c_77_n N_A_79_21#_M1003_g N_A_79_21#_c_78_n
+ N_A_79_21#_M1007_g N_A_79_21#_M1010_g N_A_79_21#_c_73_n N_A_79_21#_c_74_n
+ N_A_79_21#_c_75_n N_A_79_21#_c_81_n N_A_79_21#_c_91_p N_A_79_21#_c_144_p
+ N_A_79_21#_c_92_p N_A_79_21#_c_82_n N_A_79_21#_c_83_n N_A_79_21#_c_84_n
+ N_A_79_21#_c_94_p N_A_79_21#_c_76_n N_A_79_21#_c_86_n N_A_79_21#_c_103_p
+ PM_SKY130_FD_SC_HDLL__A21BO_2%A_79_21#
x_PM_SKY130_FD_SC_HDLL__A21BO_2%B1_N N_B1_N_c_175_n N_B1_N_M1006_g
+ N_B1_N_c_176_n N_B1_N_M1008_g B1_N B1_N PM_SKY130_FD_SC_HDLL__A21BO_2%B1_N
x_PM_SKY130_FD_SC_HDLL__A21BO_2%A_317_93# N_A_317_93#_M1006_d
+ N_A_317_93#_M1008_d N_A_317_93#_c_213_n N_A_317_93#_M1005_g
+ N_A_317_93#_c_208_n N_A_317_93#_M1011_g N_A_317_93#_c_214_n
+ N_A_317_93#_c_209_n N_A_317_93#_c_215_n N_A_317_93#_c_210_n
+ N_A_317_93#_c_211_n N_A_317_93#_c_212_n
+ PM_SKY130_FD_SC_HDLL__A21BO_2%A_317_93#
x_PM_SKY130_FD_SC_HDLL__A21BO_2%A1 N_A1_c_263_n N_A1_M1001_g N_A1_c_264_n
+ N_A1_M1000_g A1 N_A1_c_265_n PM_SKY130_FD_SC_HDLL__A21BO_2%A1
x_PM_SKY130_FD_SC_HDLL__A21BO_2%A2 N_A2_c_294_n N_A2_M1002_g N_A2_c_295_n
+ N_A2_M1009_g A2 PM_SKY130_FD_SC_HDLL__A21BO_2%A2
x_PM_SKY130_FD_SC_HDLL__A21BO_2%VPWR N_VPWR_M1003_s N_VPWR_M1007_s
+ N_VPWR_M1001_d N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_325_n VPWR N_VPWR_c_326_n
+ N_VPWR_c_318_n N_VPWR_c_328_n PM_SKY130_FD_SC_HDLL__A21BO_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A21BO_2%X N_X_M1004_s N_X_M1003_d N_X_c_388_n
+ N_X_c_383_n N_X_c_392_n N_X_c_393_n N_X_c_398_n X N_X_c_386_n
+ PM_SKY130_FD_SC_HDLL__A21BO_2%X
x_PM_SKY130_FD_SC_HDLL__A21BO_2%A_523_297# N_A_523_297#_M1005_d
+ N_A_523_297#_M1009_d N_A_523_297#_c_430_n N_A_523_297#_c_425_n
+ N_A_523_297#_c_423_n PM_SKY130_FD_SC_HDLL__A21BO_2%A_523_297#
x_PM_SKY130_FD_SC_HDLL__A21BO_2%VGND N_VGND_M1004_d N_VGND_M1010_d
+ N_VGND_M1011_s N_VGND_M1002_d N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n N_VGND_c_460_n N_VGND_c_461_n
+ N_VGND_c_462_n VGND N_VGND_c_463_n N_VGND_c_464_n N_VGND_c_465_n
+ PM_SKY130_FD_SC_HDLL__A21BO_2%VGND
cc_1 VNB N_A_79_21#_M1004_g 0.0218602f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_2 VNB N_A_79_21#_M1010_g 0.0211558f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_3 VNB N_A_79_21#_c_73_n 0.0129982f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.217
cc_4 VNB N_A_79_21#_c_74_n 0.0207107f $X=-0.19 $Y=-0.24 $X2=0.875 $Y2=1.16
cc_5 VNB N_A_79_21#_c_75_n 0.0123912f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.217
cc_6 VNB N_A_79_21#_c_76_n 0.00298284f $X=-0.19 $Y=-0.24 $X2=2.605 $Y2=1.505
cc_7 VNB N_B1_N_c_175_n 0.0194307f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=0.235
cc_8 VNB N_B1_N_c_176_n 0.0246715f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB B1_N 0.00590379f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_10 VNB N_A_317_93#_c_208_n 0.0196384f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_317_93#_c_209_n 0.00397672f $X=-0.19 $Y=-0.24 $X2=1 $Y2=0.56
cc_12 VNB N_A_317_93#_c_210_n 0.00479358f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.217
cc_13 VNB N_A_317_93#_c_211_n 0.00553293f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_317_93#_c_212_n 0.0386752f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.895
cc_15 VNB N_A1_c_263_n 0.0230421f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=0.235
cc_16 VNB N_A1_c_264_n 0.0170058f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A1_c_265_n 0.00111037f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_18 VNB N_A2_c_294_n 0.0213299f $X=-0.19 $Y=-0.24 $X2=2.625 $Y2=0.235
cc_19 VNB N_A2_c_295_n 0.0270541f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB A2 0.0126724f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.025
cc_21 VNB N_VPWR_c_318_n 0.17485f $X=-0.19 $Y=-0.24 $X2=2.29 $Y2=2.11
cc_22 VNB N_X_c_383_n 0.0072777f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_23 VNB X 0.0217149f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.217
cc_24 VNB N_VGND_c_454_n 0.00994884f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_25 VNB N_VGND_c_455_n 0.017772f $X=-0.19 $Y=-0.24 $X2=0.975 $Y2=1.985
cc_26 VNB N_VGND_c_456_n 0.0181224f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.025
cc_27 VNB N_VGND_c_457_n 0.00815763f $X=-0.19 $Y=-0.24 $X2=0.595 $Y2=1.16
cc_28 VNB N_VGND_c_458_n 0.0118855f $X=-0.19 $Y=-0.24 $X2=0.785 $Y2=1.495
cc_29 VNB N_VGND_c_459_n 0.0167205f $X=-0.19 $Y=-0.24 $X2=0.785 $Y2=1.16
cc_30 VNB N_VGND_c_460_n 0.0277822f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_461_n 0.0211714f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.665
cc_32 VNB N_VGND_c_462_n 0.00631443f $X=-0.19 $Y=-0.24 $X2=1.3 $Y2=1.895
cc_33 VNB N_VGND_c_463_n 0.0300073f $X=-0.19 $Y=-0.24 $X2=2.29 $Y2=1.895
cc_34 VNB N_VGND_c_464_n 0.00525267f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_465_n 0.238309f $X=-0.19 $Y=-0.24 $X2=0.785 $Y2=1.16
cc_36 VPB N_A_79_21#_c_77_n 0.0183459f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_37 VPB N_A_79_21#_c_78_n 0.0189829f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_38 VPB N_A_79_21#_c_73_n 0.00694419f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.217
cc_39 VPB N_A_79_21#_c_75_n 0.00648954f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.217
cc_40 VPB N_A_79_21#_c_81_n 0.00119282f $X=-0.19 $Y=1.305 $X2=0.785 $Y2=1.16
cc_41 VPB N_A_79_21#_c_82_n 0.0139599f $X=-0.19 $Y=1.305 $X2=2.125 $Y2=2
cc_42 VPB N_A_79_21#_c_83_n 2.08527e-19 $X=-0.19 $Y=1.305 $X2=1.385 $Y2=2
cc_43 VPB N_A_79_21#_c_84_n 0.0100723f $X=-0.19 $Y=1.305 $X2=2.25 $Y2=2.105
cc_44 VPB N_A_79_21#_c_76_n 0.00109509f $X=-0.19 $Y=1.305 $X2=2.605 $Y2=1.505
cc_45 VPB N_A_79_21#_c_86_n 7.80569e-19 $X=-0.19 $Y=1.305 $X2=2.25 $Y2=2
cc_46 VPB N_B1_N_c_176_n 0.0276797f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB B1_N 0.00241926f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_48 VPB N_A_317_93#_c_213_n 0.0193149f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_49 VPB N_A_317_93#_c_214_n 0.00332605f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_50 VPB N_A_317_93#_c_215_n 0.00474693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_317_93#_c_211_n 0.00174522f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_52 VPB N_A_317_93#_c_212_n 0.015928f $X=-0.19 $Y=1.305 $X2=1.3 $Y2=1.895
cc_53 VPB N_A1_c_263_n 0.0247508f $X=-0.19 $Y=1.305 $X2=2.625 $Y2=0.235
cc_54 VPB N_A1_c_265_n 0.00100523f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_55 VPB N_A2_c_295_n 0.0292428f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_56 VPB A2 0.00717147f $X=-0.19 $Y=1.305 $X2=0.47 $Y2=1.025
cc_57 VPB N_VPWR_c_319_n 0.0102988f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_320_n 0.0127536f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_59 VPB N_VPWR_c_321_n 0.0185988f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.41
cc_60 VPB N_VPWR_c_322_n 0.00564356f $X=-0.19 $Y=1.305 $X2=1 $Y2=0.56
cc_61 VPB N_VPWR_c_323_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.217
cc_62 VPB N_VPWR_c_324_n 0.0434875f $X=-0.19 $Y=1.305 $X2=0.785 $Y2=1.495
cc_63 VPB N_VPWR_c_325_n 0.00323909f $X=-0.19 $Y=1.305 $X2=0.785 $Y2=1.16
cc_64 VPB N_VPWR_c_326_n 0.0237171f $X=-0.19 $Y=1.305 $X2=2.25 $Y2=2.11
cc_65 VPB N_VPWR_c_318_n 0.0579595f $X=-0.19 $Y=1.305 $X2=2.29 $Y2=2.11
cc_66 VPB N_VPWR_c_328_n 0.00631318f $X=-0.19 $Y=1.305 $X2=2.605 $Y2=1.505
cc_67 VPB X 0.0224901f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.217
cc_68 VPB N_X_c_386_n 0.00731822f $X=-0.19 $Y=1.305 $X2=0.785 $Y2=1.16
cc_69 VPB N_A_523_297#_c_423_n 0.0267021f $X=-0.19 $Y=1.305 $X2=0.975 $Y2=1.985
cc_70 N_A_79_21#_M1010_g N_B1_N_c_175_n 0.012429f $X=1 $Y=0.56 $X2=-0.19
+ $Y2=-0.24
cc_71 N_A_79_21#_c_78_n N_B1_N_c_176_n 0.0164349f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_72 N_A_79_21#_c_75_n N_B1_N_c_176_n 0.012429f $X=0.975 $Y=1.217 $X2=0 $Y2=0
cc_73 N_A_79_21#_c_81_n N_B1_N_c_176_n 0.00102591f $X=0.785 $Y=1.16 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_91_p N_B1_N_c_176_n 0.00196984f $X=1.215 $Y=1.58 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_92_p N_B1_N_c_176_n 0.00478166f $X=1.3 $Y=1.895 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_82_n N_B1_N_c_176_n 0.0139831f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_94_p N_B1_N_c_176_n 0.00260397f $X=2.29 $Y=1.77 $X2=0 $Y2=0
cc_78 N_A_79_21#_M1010_g B1_N 0.004792f $X=1 $Y=0.56 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_81_n B1_N 0.0142221f $X=0.785 $Y=1.16 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_91_p B1_N 0.0137558f $X=1.215 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_82_n B1_N 0.00398397f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_82_n N_A_317_93#_M1008_d 0.00229505f $X=2.125 $Y=2 $X2=0
+ $Y2=0
cc_83 N_A_79_21#_c_84_n N_A_317_93#_c_213_n 0.00425616f $X=2.25 $Y=2.105 $X2=0
+ $Y2=0
cc_84 N_A_79_21#_c_76_n N_A_317_93#_c_213_n 0.0173635f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_85 N_A_79_21#_c_76_n N_A_317_93#_c_208_n 0.0052026f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_86 N_A_79_21#_c_103_p N_A_317_93#_c_208_n 0.00860314f $X=2.775 $Y=0.73 $X2=0
+ $Y2=0
cc_87 N_A_79_21#_c_91_p N_A_317_93#_c_214_n 0.00928876f $X=1.215 $Y=1.58 $X2=0
+ $Y2=0
cc_88 N_A_79_21#_c_92_p N_A_317_93#_c_214_n 0.00447251f $X=1.3 $Y=1.895 $X2=0
+ $Y2=0
cc_89 N_A_79_21#_c_82_n N_A_317_93#_c_214_n 0.0320911f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_94_p N_A_317_93#_c_214_n 0.00403971f $X=2.29 $Y=1.77 $X2=0
+ $Y2=0
cc_91 N_A_79_21#_c_76_n N_A_317_93#_c_214_n 0.0104332f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_92 N_A_79_21#_c_76_n N_A_317_93#_c_209_n 0.00587043f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_93 N_A_79_21#_c_91_p N_A_317_93#_c_215_n 0.00223554f $X=1.215 $Y=1.58 $X2=0
+ $Y2=0
cc_94 N_A_79_21#_c_76_n N_A_317_93#_c_215_n 0.0101378f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_95 N_A_79_21#_c_103_p N_A_317_93#_c_210_n 0.00662477f $X=2.775 $Y=0.73 $X2=0
+ $Y2=0
cc_96 N_A_79_21#_c_82_n N_A_317_93#_c_211_n 0.00306578f $X=2.125 $Y=2 $X2=0
+ $Y2=0
cc_97 N_A_79_21#_c_76_n N_A_317_93#_c_211_n 0.0331168f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_98 N_A_79_21#_c_86_n N_A_317_93#_c_211_n 0.00260016f $X=2.25 $Y=2 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_82_n N_A_317_93#_c_212_n 3.30674e-19 $X=2.125 $Y=2 $X2=0
+ $Y2=0
cc_100 N_A_79_21#_c_76_n N_A_317_93#_c_212_n 0.0185631f $X=2.605 $Y=1.505 $X2=0
+ $Y2=0
cc_101 N_A_79_21#_c_86_n N_A_317_93#_c_212_n 0.00140592f $X=2.25 $Y=2 $X2=0
+ $Y2=0
cc_102 N_A_79_21#_c_76_n N_A1_c_263_n 0.00435796f $X=2.605 $Y=1.505 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_79_21#_c_103_p N_A1_c_263_n 0.00222594f $X=2.775 $Y=0.73 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_79_21#_c_76_n N_A1_c_264_n 0.0032701f $X=2.605 $Y=1.505 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_76_n N_A1_c_265_n 0.0375329f $X=2.605 $Y=1.505 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_103_p N_A1_c_265_n 0.00268802f $X=2.775 $Y=0.73 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_91_p N_VPWR_M1007_s 0.0107863f $X=1.215 $Y=1.58 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_92_p N_VPWR_M1007_s 0.00553291f $X=1.3 $Y=1.895 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_83_n N_VPWR_M1007_s 0.00444479f $X=1.385 $Y=2 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_77_n N_VPWR_c_320_n 0.009234f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_78_n N_VPWR_c_320_n 0.00114243f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_77_n N_VPWR_c_321_n 0.00464801f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_78_n N_VPWR_c_321_n 0.00681977f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_78_n N_VPWR_c_322_n 0.010433f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_91_p N_VPWR_c_322_n 0.00224709f $X=1.215 $Y=1.58 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_82_n N_VPWR_c_322_n 0.0065253f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_83_n N_VPWR_c_322_n 0.0141627f $X=1.385 $Y=2 $X2=0 $Y2=0
cc_118 N_A_79_21#_c_84_n N_VPWR_c_322_n 0.00572296f $X=2.25 $Y=2.105 $X2=0 $Y2=0
cc_119 N_A_79_21#_c_82_n N_VPWR_c_324_n 0.0126652f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_120 N_A_79_21#_c_84_n N_VPWR_c_324_n 0.0174202f $X=2.25 $Y=2.105 $X2=0 $Y2=0
cc_121 N_A_79_21#_M1005_s N_VPWR_c_318_n 0.00430086f $X=2.165 $Y=1.485 $X2=0
+ $Y2=0
cc_122 N_A_79_21#_c_77_n N_VPWR_c_318_n 0.00541979f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_78_n N_VPWR_c_318_n 0.0135443f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_82_n N_VPWR_c_318_n 0.0194284f $X=2.125 $Y=2 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_83_n N_VPWR_c_318_n 8.79686e-19 $X=1.385 $Y=2 $X2=0 $Y2=0
cc_126 N_A_79_21#_c_84_n N_VPWR_c_318_n 0.00953699f $X=2.25 $Y=2.105 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_144_p N_X_M1003_d 0.00252521f $X=0.95 $Y=1.58 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_77_n N_X_c_388_n 0.0184218f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_129 N_A_79_21#_M1004_g N_X_c_383_n 0.015561f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_130 N_A_79_21#_c_74_n N_X_c_383_n 0.0045056f $X=0.875 $Y=1.16 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_81_n N_X_c_383_n 0.0187691f $X=0.785 $Y=1.16 $X2=0 $Y2=0
cc_132 N_A_79_21#_M1004_g N_X_c_392_n 0.010295f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_78_n N_X_c_393_n 0.00250954f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_74_n N_X_c_393_n 7.5759e-19 $X=0.875 $Y=1.16 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_144_p N_X_c_393_n 0.0173589f $X=0.95 $Y=1.58 $X2=0 $Y2=0
cc_136 N_A_79_21#_c_92_p N_X_c_393_n 0.00290357f $X=1.3 $Y=1.895 $X2=0 $Y2=0
cc_137 N_A_79_21#_c_83_n N_X_c_393_n 0.00596625f $X=1.385 $Y=2 $X2=0 $Y2=0
cc_138 N_A_79_21#_c_78_n N_X_c_398_n 0.0105009f $X=0.975 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_79_21#_c_83_n N_X_c_398_n 0.00503008f $X=1.385 $Y=2 $X2=0 $Y2=0
cc_140 N_A_79_21#_M1004_g X 0.0187295f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_141 N_A_79_21#_c_77_n X 0.00908416f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_79_21#_c_81_n X 0.0254097f $X=0.785 $Y=1.16 $X2=0 $Y2=0
cc_143 N_A_79_21#_c_76_n N_A_523_297#_M1005_d 0.00261426f $X=2.605 $Y=1.505
+ $X2=-0.19 $Y2=-0.24
cc_144 N_A_79_21#_c_84_n N_A_523_297#_c_425_n 0.0276147f $X=2.25 $Y=2.105 $X2=0
+ $Y2=0
cc_145 N_A_79_21#_c_94_p N_A_523_297#_c_425_n 0.00389343f $X=2.29 $Y=1.77 $X2=0
+ $Y2=0
cc_146 N_A_79_21#_c_76_n N_A_523_297#_c_425_n 0.00868584f $X=2.605 $Y=1.505
+ $X2=0 $Y2=0
cc_147 N_A_79_21#_c_86_n N_A_523_297#_c_425_n 0.017956f $X=2.25 $Y=2 $X2=0 $Y2=0
cc_148 N_A_79_21#_M1004_g N_VGND_c_455_n 0.00450113f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_79_21#_M1004_g N_VGND_c_456_n 0.00425835f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A_79_21#_M1010_g N_VGND_c_456_n 0.00564095f $X=1 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_79_21#_M1004_g N_VGND_c_457_n 0.00103226f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_79_21#_M1010_g N_VGND_c_457_n 0.0108779f $X=1 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_79_21#_c_103_p N_VGND_c_463_n 0.00691282f $X=2.775 $Y=0.73 $X2=0
+ $Y2=0
cc_154 N_A_79_21#_M1011_d N_VGND_c_465_n 0.00431979f $X=2.625 $Y=0.235 $X2=0
+ $Y2=0
cc_155 N_A_79_21#_M1004_g N_VGND_c_465_n 0.0069606f $X=0.47 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_79_21#_M1010_g N_VGND_c_465_n 0.00969156f $X=1 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_79_21#_c_103_p N_VGND_c_465_n 0.0120006f $X=2.775 $Y=0.73 $X2=0 $Y2=0
cc_158 N_B1_N_c_176_n N_A_317_93#_c_214_n 0.00594348f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_159 B1_N N_A_317_93#_c_214_n 0.00633992f $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_160 N_B1_N_c_175_n N_A_317_93#_c_209_n 0.00421602f $X=1.51 $Y=0.995 $X2=0
+ $Y2=0
cc_161 N_B1_N_c_176_n N_A_317_93#_c_215_n 0.00567881f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_162 N_B1_N_c_176_n N_A_317_93#_c_210_n 0.00240199f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_163 B1_N N_A_317_93#_c_210_n 0.00530171f $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_164 N_B1_N_c_176_n N_A_317_93#_c_211_n 0.00266257f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_165 B1_N N_A_317_93#_c_211_n 0.0276068f $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_166 N_B1_N_c_176_n N_A_317_93#_c_212_n 0.00848927f $X=1.535 $Y=1.41 $X2=0
+ $Y2=0
cc_167 B1_N N_A_317_93#_c_212_n 2.86645e-19 $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_168 N_B1_N_c_176_n N_VPWR_c_324_n 5.44397e-19 $X=1.535 $Y=1.41 $X2=0 $Y2=0
cc_169 N_B1_N_c_175_n N_VGND_c_457_n 0.0054721f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_170 B1_N N_VGND_c_457_n 0.012136f $X=1.465 $Y=1.105 $X2=0 $Y2=0
cc_171 N_B1_N_c_175_n N_VGND_c_458_n 0.00327677f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B1_N_c_175_n N_VGND_c_461_n 0.00510437f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B1_N_c_175_n N_VGND_c_465_n 0.00512902f $X=1.51 $Y=0.995 $X2=0 $Y2=0
cc_174 N_A_317_93#_c_213_n N_A1_c_263_n 0.022612f $X=2.525 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_175 N_A_317_93#_c_212_n N_A1_c_263_n 0.0240867f $X=2.525 $Y=1.2 $X2=-0.19
+ $Y2=-0.24
cc_176 N_A_317_93#_c_208_n N_A1_c_264_n 0.0210761f $X=2.55 $Y=0.99 $X2=0 $Y2=0
cc_177 N_A_317_93#_c_213_n N_A1_c_265_n 2.06074e-19 $X=2.525 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_317_93#_c_212_n N_A1_c_265_n 5.39444e-19 $X=2.525 $Y=1.2 $X2=0 $Y2=0
cc_179 N_A_317_93#_c_213_n N_VPWR_c_324_n 0.00597712f $X=2.525 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_317_93#_c_213_n N_VPWR_c_318_n 0.0115507f $X=2.525 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_317_93#_c_213_n N_A_523_297#_c_425_n 0.0105415f $X=2.525 $Y=1.41
+ $X2=0 $Y2=0
cc_182 N_A_317_93#_c_208_n N_VGND_c_458_n 0.00482545f $X=2.55 $Y=0.99 $X2=0
+ $Y2=0
cc_183 N_A_317_93#_c_211_n N_VGND_c_458_n 0.00672869f $X=2.24 $Y=1.16 $X2=0
+ $Y2=0
cc_184 N_A_317_93#_c_212_n N_VGND_c_458_n 0.00694766f $X=2.525 $Y=1.2 $X2=0
+ $Y2=0
cc_185 N_A_317_93#_c_210_n N_VGND_c_461_n 0.00703609f $X=1.95 $Y=0.74 $X2=0
+ $Y2=0
cc_186 N_A_317_93#_c_208_n N_VGND_c_463_n 0.00446466f $X=2.55 $Y=0.99 $X2=0
+ $Y2=0
cc_187 N_A_317_93#_c_208_n N_VGND_c_465_n 0.00774817f $X=2.55 $Y=0.99 $X2=0
+ $Y2=0
cc_188 N_A_317_93#_c_210_n N_VGND_c_465_n 0.0119945f $X=1.95 $Y=0.74 $X2=0 $Y2=0
cc_189 N_A1_c_264_n N_A2_c_294_n 0.0300894f $X=3.03 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_190 N_A1_c_263_n N_A2_c_295_n 0.0694346f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A1_c_265_n N_A2_c_295_n 0.00173351f $X=2.97 $Y=1.16 $X2=0 $Y2=0
cc_192 N_A1_c_263_n A2 0.00237262f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A1_c_265_n A2 0.0260796f $X=2.97 $Y=1.16 $X2=0 $Y2=0
cc_194 N_A1_c_263_n N_VPWR_c_323_n 0.00403097f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A1_c_263_n N_VPWR_c_324_n 0.00518485f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A1_c_263_n N_VPWR_c_318_n 0.00687544f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A1_c_263_n N_A_523_297#_c_430_n 0.0119127f $X=3.005 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A1_c_265_n N_A_523_297#_c_430_n 0.00940041f $X=2.97 $Y=1.16 $X2=0 $Y2=0
cc_199 N_A1_c_263_n N_A_523_297#_c_425_n 0.00759714f $X=3.005 $Y=1.41 $X2=0
+ $Y2=0
cc_200 N_A1_c_265_n N_A_523_297#_c_425_n 6.21659e-19 $X=2.97 $Y=1.16 $X2=0 $Y2=0
cc_201 N_A1_c_263_n N_A_523_297#_c_423_n 5.73894e-19 $X=3.005 $Y=1.41 $X2=0
+ $Y2=0
cc_202 N_A1_c_264_n N_VGND_c_460_n 0.00359683f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_203 N_A1_c_264_n N_VGND_c_463_n 0.00585385f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_204 N_A1_c_264_n N_VGND_c_465_n 0.0110141f $X=3.03 $Y=0.995 $X2=0 $Y2=0
cc_205 N_A2_c_295_n N_VPWR_c_323_n 0.00378873f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A2_c_295_n N_VPWR_c_326_n 0.00487509f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A2_c_295_n N_VPWR_c_318_n 0.00754809f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_208 A2 N_A_523_297#_M1009_d 0.00582115f $X=3.42 $Y=1.105 $X2=0 $Y2=0
cc_209 N_A2_c_295_n N_A_523_297#_c_430_n 0.00820192f $X=3.475 $Y=1.41 $X2=0
+ $Y2=0
cc_210 A2 N_A_523_297#_c_430_n 0.00649519f $X=3.42 $Y=1.105 $X2=0 $Y2=0
cc_211 N_A2_c_295_n N_A_523_297#_c_425_n 5.29442e-19 $X=3.475 $Y=1.41 $X2=0
+ $Y2=0
cc_212 N_A2_c_295_n N_A_523_297#_c_423_n 0.0106652f $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_213 A2 N_A_523_297#_c_423_n 0.00752591f $X=3.42 $Y=1.105 $X2=0 $Y2=0
cc_214 N_A2_c_294_n N_VGND_c_460_n 0.0239315f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_215 N_A2_c_295_n N_VGND_c_460_n 7.72974e-19 $X=3.475 $Y=1.41 $X2=0 $Y2=0
cc_216 A2 N_VGND_c_460_n 0.0119779f $X=3.42 $Y=1.105 $X2=0 $Y2=0
cc_217 N_A2_c_294_n N_VGND_c_463_n 0.0046653f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_218 N_A2_c_294_n N_VGND_c_465_n 0.00799591f $X=3.45 $Y=0.995 $X2=0 $Y2=0
cc_219 N_VPWR_c_318_n N_X_M1003_d 0.00271101f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_220 N_VPWR_c_320_n N_X_c_388_n 9.31105e-19 $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_221 N_VPWR_c_321_n N_X_c_388_n 0.00265246f $X=1.14 $Y=2.72 $X2=0 $Y2=0
cc_222 N_VPWR_c_318_n N_X_c_388_n 0.00525658f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_223 N_VPWR_c_320_n N_X_c_398_n 0.0106235f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_224 N_VPWR_c_321_n N_X_c_398_n 0.0124337f $X=1.14 $Y=2.72 $X2=0 $Y2=0
cc_225 N_VPWR_c_322_n N_X_c_398_n 0.00877074f $X=1.305 $Y=2.36 $X2=0 $Y2=0
cc_226 N_VPWR_c_318_n N_X_c_398_n 0.00943451f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_227 N_VPWR_M1003_s X 0.00290274f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_228 N_VPWR_M1003_s N_X_c_386_n 0.00356271f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_229 N_VPWR_c_320_n N_X_c_386_n 0.0145189f $X=0.26 $Y=2.34 $X2=0 $Y2=0
cc_230 N_VPWR_c_318_n N_X_c_386_n 0.00144057f $X=3.91 $Y=2.72 $X2=0 $Y2=0
cc_231 N_VPWR_c_318_n N_A_523_297#_M1005_d 0.00239291f $X=3.91 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_232 N_VPWR_c_318_n N_A_523_297#_M1009_d 0.00217517f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_233 N_VPWR_M1001_d N_A_523_297#_c_430_n 0.00845322f $X=3.095 $Y=1.485 $X2=0
+ $Y2=0
cc_234 N_VPWR_c_323_n N_A_523_297#_c_430_n 0.0130812f $X=3.24 $Y=2.36 $X2=0
+ $Y2=0
cc_235 N_VPWR_c_324_n N_A_523_297#_c_430_n 0.0028731f $X=3.155 $Y=2.72 $X2=0
+ $Y2=0
cc_236 N_VPWR_c_326_n N_A_523_297#_c_430_n 0.00203428f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_237 N_VPWR_c_318_n N_A_523_297#_c_430_n 0.0099901f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_238 N_VPWR_c_323_n N_A_523_297#_c_425_n 0.0165641f $X=3.24 $Y=2.36 $X2=0
+ $Y2=0
cc_239 N_VPWR_c_324_n N_A_523_297#_c_425_n 0.0222543f $X=3.155 $Y=2.72 $X2=0
+ $Y2=0
cc_240 N_VPWR_c_318_n N_A_523_297#_c_425_n 0.0140211f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_241 N_VPWR_c_323_n N_A_523_297#_c_423_n 0.0209034f $X=3.24 $Y=2.36 $X2=0
+ $Y2=0
cc_242 N_VPWR_c_326_n N_A_523_297#_c_423_n 0.0243171f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_243 N_VPWR_c_318_n N_A_523_297#_c_423_n 0.0141345f $X=3.91 $Y=2.72 $X2=0
+ $Y2=0
cc_244 N_X_c_383_n N_VGND_M1004_d 0.00344693f $X=0.71 $Y=0.715 $X2=-0.19
+ $Y2=-0.24
cc_245 X N_VGND_M1004_d 6.00252e-19 $X=0.15 $Y=1.785 $X2=-0.19 $Y2=-0.24
cc_246 N_X_c_383_n N_VGND_c_455_n 0.0178745f $X=0.71 $Y=0.715 $X2=0 $Y2=0
cc_247 N_X_c_383_n N_VGND_c_456_n 0.00212146f $X=0.71 $Y=0.715 $X2=0 $Y2=0
cc_248 N_X_c_392_n N_VGND_c_456_n 0.0164101f $X=0.735 $Y=0.4 $X2=0 $Y2=0
cc_249 N_X_M1004_s N_VGND_c_465_n 0.00391907f $X=0.545 $Y=0.235 $X2=0 $Y2=0
cc_250 N_X_c_383_n N_VGND_c_465_n 0.00495188f $X=0.71 $Y=0.715 $X2=0 $Y2=0
cc_251 N_X_c_392_n N_VGND_c_465_n 0.0137078f $X=0.735 $Y=0.4 $X2=0 $Y2=0
cc_252 N_VGND_c_465_n A_621_47# 0.0115413f $X=3.91 $Y=0 $X2=-0.19 $Y2=-0.24
