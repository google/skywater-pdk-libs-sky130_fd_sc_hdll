# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o221a_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__o221a_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.305000 1.075000 3.955000 1.445000 ;
        RECT 3.305000 1.445000 5.225000 1.615000 ;
        RECT 4.975000 1.075000 5.535000 1.275000 ;
        RECT 4.975000 1.275000 5.225000 1.445000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.125000 1.075000 4.755000 1.275000 ;
    END
  END A2
  PIN B1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.065000 1.075000 1.730000 1.445000 ;
        RECT 1.065000 1.445000 3.045000 1.615000 ;
        RECT 2.665000 1.075000 3.045000 1.445000 ;
    END
  END B1
  PIN B2
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.075000 2.495000 1.275000 ;
    END
  END B2
  PIN C1
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.075000 0.440000 1.275000 ;
    END
  END C1
  PIN X
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.735000 0.255000 6.115000 0.725000 ;
        RECT 5.735000 0.725000 7.055000 0.735000 ;
        RECT 5.735000 0.735000 7.710000 0.905000 ;
        RECT 5.865000 1.785000 6.500000 1.955000 ;
        RECT 5.865000 1.955000 6.075000 2.465000 ;
        RECT 6.330000 1.445000 7.710000 1.615000 ;
        RECT 6.330000 1.615000 6.500000 1.785000 ;
        RECT 6.675000 0.255000 7.055000 0.725000 ;
        RECT 6.765000 1.615000 7.015000 2.465000 ;
        RECT 7.365000 0.905000 7.710000 1.445000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 3.435000  0.085000 3.765000 0.465000 ;
        RECT 4.455000  0.085000 4.625000 0.555000 ;
        RECT 5.395000  0.085000 5.565000 0.905000 ;
        RECT 6.335000  0.085000 6.505000 0.555000 ;
        RECT 7.275000  0.085000 7.530000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.145000 1.455000 0.395000 2.635000 ;
        RECT 1.085000 2.125000 1.335000 2.635000 ;
        RECT 2.965000 2.125000 3.725000 2.635000 ;
        RECT 5.355000 2.125000 5.605000 2.635000 ;
        RECT 6.295000 2.125000 6.545000 2.635000 ;
        RECT 7.235000 1.795000 7.485000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 3.255000 0.475000 ;
      RECT 0.085000 0.475000 0.345000 0.895000 ;
      RECT 0.515000 0.645000 0.895000 0.865000 ;
      RECT 0.615000 0.865000 0.895000 1.785000 ;
      RECT 0.615000 1.785000 5.645000 1.955000 ;
      RECT 0.615000 1.955000 0.865000 2.465000 ;
      RECT 1.115000 0.475000 1.285000 0.905000 ;
      RECT 1.455000 0.645000 4.235000 0.725000 ;
      RECT 1.455000 0.725000 5.175000 0.905000 ;
      RECT 1.555000 2.125000 1.805000 2.295000 ;
      RECT 1.555000 2.295000 2.745000 2.465000 ;
      RECT 2.495000 2.125000 2.745000 2.295000 ;
      RECT 3.945000 2.125000 4.195000 2.295000 ;
      RECT 3.945000 2.295000 5.135000 2.465000 ;
      RECT 3.985000 0.255000 4.235000 0.645000 ;
      RECT 4.795000 0.255000 5.175000 0.725000 ;
      RECT 4.885000 2.125000 5.135000 2.295000 ;
      RECT 5.475000 1.445000 5.925000 1.615000 ;
      RECT 5.475000 1.615000 5.645000 1.785000 ;
      RECT 5.705000 1.075000 7.055000 1.275000 ;
      RECT 5.705000 1.275000 5.925000 1.445000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o221a_4
