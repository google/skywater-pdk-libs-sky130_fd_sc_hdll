* File: sky130_fd_sc_hdll__a21bo_2.pex.spice
* Created: Thu Aug 27 18:52:10 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%A_79_21# 1 2 9 11 13 14 16 19 22 23 24 27
+ 30 31 33 34 35 36 42 44 45 53
c104 27 0 9.15276e-20 $X=0.785 $Y=1.16
c105 14 0 9.2021e-20 $X=0.975 $Y=1.41
r106 44 46 20.5508 $w=1.68e-07 $l=3.15e-07 $layer=LI1_cond $X=2.605 $Y=1.59
+ $X2=2.29 $Y2=1.59
r107 43 53 9.92344 $w=1.88e-07 $l=1.7e-07 $layer=LI1_cond $X=2.605 $Y=0.73
+ $X2=2.775 $Y2=0.73
r108 43 44 35.621 $w=2.18e-07 $l=6.8e-07 $layer=LI1_cond $X=2.605 $Y=0.825
+ $X2=2.605 $Y2=1.505
r109 40 45 5.16603 $w=2.1e-07 $l=1.2339e-07 $layer=LI1_cond $X=2.29 $Y=1.895
+ $X2=2.25 $Y2=2
r110 40 42 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=2.29 $Y=1.895
+ $X2=2.29 $Y2=1.77
r111 39 46 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=1.675
+ $X2=2.29 $Y2=1.59
r112 39 42 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=2.29 $Y=1.675
+ $X2=2.29 $Y2=1.77
r113 36 45 5.16603 $w=2.1e-07 $l=1.05e-07 $layer=LI1_cond $X=2.25 $Y=2.105
+ $X2=2.25 $Y2=2
r114 36 38 0.244 $w=2.5e-07 $l=5e-09 $layer=LI1_cond $X=2.25 $Y=2.105 $X2=2.25
+ $Y2=2.11
r115 34 45 1.34256 $w=2.1e-07 $l=1.25e-07 $layer=LI1_cond $X=2.125 $Y=2 $X2=2.25
+ $Y2=2
r116 34 35 39.0823 $w=2.08e-07 $l=7.4e-07 $layer=LI1_cond $X=2.125 $Y=2
+ $X2=1.385 $Y2=2
r117 33 35 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=1.3 $Y=1.895
+ $X2=1.385 $Y2=2
r118 32 33 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.3 $Y=1.665
+ $X2=1.3 $Y2=1.895
r119 30 32 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.215 $Y=1.58
+ $X2=1.3 $Y2=1.665
r120 30 31 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=1.215 $Y=1.58
+ $X2=0.95 $Y2=1.58
r121 27 28 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.785
+ $Y=1.16 $X2=0.785 $Y2=1.16
r122 25 31 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=0.785 $Y=1.495
+ $X2=0.95 $Y2=1.58
r123 25 27 11.699 $w=3.28e-07 $l=3.35e-07 $layer=LI1_cond $X=0.785 $Y=1.495
+ $X2=0.785 $Y2=1.16
r124 23 28 19.9956 $w=2.7e-07 $l=9e-08 $layer=POLY_cond $X=0.875 $Y=1.16
+ $X2=0.785 $Y2=1.16
r125 23 24 1.40033 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=0.875 $Y=1.16
+ $X2=0.975 $Y2=1.217
r126 21 28 42.213 $w=2.7e-07 $l=1.9e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.785 $Y2=1.16
r127 21 22 1.40033 $w=2.7e-07 $l=1.253e-07 $layer=POLY_cond $X=0.595 $Y=1.16
+ $X2=0.495 $Y2=1.217
r128 17 24 30.0832 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=1 $Y=1.025
+ $X2=0.975 $Y2=1.217
r129 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1 $Y=1.025 $X2=1
+ $Y2=0.56
r130 14 24 30.0832 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.217
r131 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.975 $Y=1.41
+ $X2=0.975 $Y2=1.985
r132 11 22 30.0832 $w=1.65e-07 $l=1.93e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.217
r133 11 13 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
r134 7 22 30.0832 $w=1.65e-07 $l=2.04118e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.495 $Y2=1.217
r135 7 9 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=0.47 $Y=1.025
+ $X2=0.47 $Y2=0.56
r136 2 42 600 $w=1.7e-07 $l=3.41833e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.485 $X2=2.29 $Y2=1.77
r137 2 38 600 $w=1.7e-07 $l=6.84653e-07 $layer=licon1_PDIFF $count=1 $X=2.165
+ $Y=1.485 $X2=2.29 $Y2=2.11
r138 1 53 182 $w=1.7e-07 $l=5.65044e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.775 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%B1_N 1 3 4 6 7 13
c33 4 0 2.82158e-19 $X=1.535 $Y=1.41
c34 1 0 7.10112e-20 $X=1.51 $Y=0.995
r35 7 13 3.49225 $w=3.28e-07 $l=1e-07 $layer=LI1_cond $X=1.55 $Y=1.16 $X2=1.45
+ $Y2=1.16
r36 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.57
+ $Y=1.16 $X2=1.57 $Y2=1.16
r37 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.57 $Y2=1.16
r38 4 6 76.3167 $w=1.8e-07 $l=2.85e-07 $layer=POLY_cond $X=1.535 $Y=1.41
+ $X2=1.535 $Y2=1.695
r39 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.51 $Y=0.995
+ $X2=1.57 $Y2=1.16
r40 1 3 102.827 $w=1.5e-07 $l=3.2e-07 $layer=POLY_cond $X=1.51 $Y=0.995 $X2=1.51
+ $Y2=0.675
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%A_317_93# 1 2 7 9 10 12 13 18 20 24 29 33
c55 33 0 7.10112e-20 $X=2.525 $Y=1.2
c56 13 0 9.2021e-20 $X=1.865 $Y=1.64
r57 33 34 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=2.525 $Y=1.2
+ $X2=2.55 $Y2=1.2
r58 30 33 37.4305 $w=3.67e-07 $l=2.85e-07 $layer=POLY_cond $X=2.24 $Y=1.2
+ $X2=2.525 $Y2=1.2
r59 29 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.24
+ $Y=1.16 $X2=2.24 $Y2=1.16
r60 26 29 10.1275 $w=3.28e-07 $l=2.9e-07 $layer=LI1_cond $X=1.95 $Y=1.16
+ $X2=2.24 $Y2=1.16
r61 22 24 11.7433 $w=1.68e-07 $l=1.8e-07 $layer=LI1_cond $X=1.77 $Y=0.74
+ $X2=1.95 $Y2=0.74
r62 19 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=1.325
+ $X2=1.95 $Y2=1.16
r63 19 20 15.0053 $w=1.68e-07 $l=2.3e-07 $layer=LI1_cond $X=1.95 $Y=1.325
+ $X2=1.95 $Y2=1.555
r64 18 26 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.95 $Y=0.995
+ $X2=1.95 $Y2=1.16
r65 17 24 0.716491 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=1.95 $Y=0.825
+ $X2=1.95 $Y2=0.74
r66 17 18 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.95 $Y=0.825
+ $X2=1.95 $Y2=0.995
r67 13 20 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.865 $Y=1.64
+ $X2=1.95 $Y2=1.555
r68 13 15 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=1.865 $Y=1.64
+ $X2=1.77 $Y2=1.64
r69 10 34 23.77 $w=1.5e-07 $l=2.1e-07 $layer=POLY_cond $X=2.55 $Y=0.99 $X2=2.55
+ $Y2=1.2
r70 10 12 138.173 $w=1.5e-07 $l=4.3e-07 $layer=POLY_cond $X=2.55 $Y=0.99
+ $X2=2.55 $Y2=0.56
r71 7 33 19.4219 $w=1.8e-07 $l=2.1e-07 $layer=POLY_cond $X=2.525 $Y=1.41
+ $X2=2.525 $Y2=1.2
r72 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.525 $Y=1.41
+ $X2=2.525 $Y2=1.985
r73 2 15 600 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_PDIFF $count=1 $X=1.625
+ $Y=1.485 $X2=1.77 $Y2=1.64
r74 1 22 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=1.585
+ $Y=0.465 $X2=1.77 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%A1 1 3 4 6 7 11
r31 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.97
+ $Y=1.16 $X2=2.97 $Y2=1.16
r32 7 11 20.5182 $w=1.98e-07 $l=3.7e-07 $layer=LI1_cond $X=2.985 $Y=1.53
+ $X2=2.985 $Y2=1.16
r33 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.03 $Y=0.995
+ $X2=2.97 $Y2=1.16
r34 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.03 $Y=0.995 $X2=3.03
+ $Y2=0.56
r35 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=2.97 $Y2=1.16
r36 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.005 $Y=1.41
+ $X2=3.005 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%A2 1 3 4 6 7
r24 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.51
+ $Y=1.16 $X2=3.51 $Y2=1.16
r25 4 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.475 $Y=1.41
+ $X2=3.51 $Y2=1.16
r26 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.475 $Y=1.41
+ $X2=3.475 $Y2=1.985
r27 1 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.45 $Y=0.995
+ $X2=3.51 $Y2=1.16
r28 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.45 $Y=0.995 $X2=3.45
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%VPWR 1 2 3 10 12 14 18 22 25 26 27 37 38
+ 44
c65 18 0 1.52452e-19 $X=1.305 $Y=2.36
r66 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r67 37 38 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r68 35 38 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=3.91 $Y2=2.72
r69 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r70 32 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r71 32 45 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=1.15 $Y2=2.72
r72 31 34 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=1.61 $Y=2.72
+ $X2=2.99 $Y2=2.72
r73 31 32 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 29 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.305 $Y2=2.72
r75 29 31 9.13369 $w=1.68e-07 $l=1.4e-07 $layer=LI1_cond $X=1.47 $Y=2.72
+ $X2=1.61 $Y2=2.72
r76 27 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r77 27 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r78 25 34 10.7647 $w=1.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=2.99 $Y2=2.72
r79 25 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.155 $Y=2.72
+ $X2=3.24 $Y2=2.72
r80 24 37 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.91 $Y2=2.72
r81 24 26 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.325 $Y=2.72
+ $X2=3.24 $Y2=2.72
r82 20 26 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=3.24 $Y=2.635
+ $X2=3.24 $Y2=2.72
r83 20 22 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=3.24 $Y=2.635
+ $X2=3.24 $Y2=2.36
r84 16 44 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.305 $Y=2.635
+ $X2=1.305 $Y2=2.72
r85 16 18 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.305 $Y=2.635
+ $X2=1.305 $Y2=2.36
r86 15 41 4.84905 $w=1.7e-07 $l=2.13e-07 $layer=LI1_cond $X=0.425 $Y=2.72
+ $X2=0.212 $Y2=2.72
r87 14 44 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.14 $Y=2.72
+ $X2=1.305 $Y2=2.72
r88 14 15 46.6471 $w=1.68e-07 $l=7.15e-07 $layer=LI1_cond $X=1.14 $Y=2.72
+ $X2=0.425 $Y2=2.72
r89 10 41 2.95951 $w=3.35e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.212 $Y2=2.72
r90 10 12 10.1484 $w=3.33e-07 $l=2.95e-07 $layer=LI1_cond $X=0.257 $Y=2.635
+ $X2=0.257 $Y2=2.34
r91 3 22 600 $w=1.7e-07 $l=9.44722e-07 $layer=licon1_PDIFF $count=1 $X=3.095
+ $Y=1.485 $X2=3.24 $Y2=2.36
r92 2 18 600 $w=1.7e-07 $l=9.87737e-07 $layer=licon1_PDIFF $count=1 $X=1.065
+ $Y=1.485 $X2=1.305 $Y2=2.36
r93 1 12 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%X 1 2 7 9 11 13 15 24 27
c40 15 0 2.28674e-20 $X=0.735 $Y=2.26
c41 13 0 1.06839e-19 $X=0.772 $Y=2.005
c42 2 0 2.64021e-20 $X=0.585 $Y=1.485
r43 24 27 2.81454 $w=2.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.245 $Y=1.92
+ $X2=0.245 $Y2=1.835
r44 24 27 1.06708 $w=2.68e-07 $l=2.5e-08 $layer=LI1_cond $X=0.245 $Y=1.81
+ $X2=0.245 $Y2=1.835
r45 18 24 39.4818 $w=2.68e-07 $l=9.25e-07 $layer=LI1_cond $X=0.245 $Y=0.885
+ $X2=0.245 $Y2=1.81
r46 13 23 2.87766 $w=2.55e-07 $l=8.5e-08 $layer=LI1_cond $X=0.772 $Y=2.005
+ $X2=0.772 $Y2=1.92
r47 13 15 11.5244 $w=2.53e-07 $l=2.55e-07 $layer=LI1_cond $X=0.772 $Y=2.005
+ $X2=0.772 $Y2=2.26
r48 9 18 30.3369 $w=1.68e-07 $l=4.65e-07 $layer=LI1_cond $X=0.71 $Y=0.8
+ $X2=0.245 $Y2=0.8
r49 9 11 9.55315 $w=3.78e-07 $l=3.15e-07 $layer=LI1_cond $X=0.71 $Y=0.715
+ $X2=0.71 $Y2=0.4
r50 8 24 4.47015 $w=1.7e-07 $l=1.35e-07 $layer=LI1_cond $X=0.38 $Y=1.92
+ $X2=0.245 $Y2=1.92
r51 7 23 4.29957 $w=1.7e-07 $l=1.27e-07 $layer=LI1_cond $X=0.645 $Y=1.92
+ $X2=0.772 $Y2=1.92
r52 7 8 17.2888 $w=1.68e-07 $l=2.65e-07 $layer=LI1_cond $X=0.645 $Y=1.92
+ $X2=0.38 $Y2=1.92
r53 2 23 600 $w=1.7e-07 $l=5.04455e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.735 $Y2=1.92
r54 2 15 600 $w=1.7e-07 $l=8.46685e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.735 $Y2=2.26
r55 1 11 91 $w=1.7e-07 $l=2.59711e-07 $layer=licon1_NDIFF $count=2 $X=0.545
+ $Y=0.235 $X2=0.735 $Y2=0.4
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%A_523_297# 1 2 9 14 16
r31 10 14 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.925 $Y=1.93
+ $X2=2.735 $Y2=1.93
r32 9 16 5.66317 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=3.495 $Y=1.93
+ $X2=3.685 $Y2=1.93
r33 9 10 37.1872 $w=1.68e-07 $l=5.7e-07 $layer=LI1_cond $X=3.495 $Y=1.93
+ $X2=2.925 $Y2=1.93
r34 2 16 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=3.565
+ $Y=1.485 $X2=3.71 $Y2=2
r35 1 14 300 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=2 $X=2.615
+ $Y=1.485 $X2=2.76 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21BO_2%VGND 1 2 3 4 13 15 17 21 25 27 29 32 33 34
+ 40 51 55
r51 54 55 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r52 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r53 46 55 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=0 $X2=3.91
+ $Y2=0
r54 45 46 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r55 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r56 42 45 60.0214 $w=1.68e-07 $l=9.2e-07 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r57 42 43 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r58 40 54 4.89672 $w=1.7e-07 $l=3.22e-07 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.817
+ $Y2=0
r59 40 45 2.93583 $w=1.68e-07 $l=4.5e-08 $layer=LI1_cond $X=3.495 $Y=0 $X2=3.45
+ $Y2=0
r60 39 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=2.53
+ $Y2=0
r61 39 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.15
+ $Y2=0
r62 38 39 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r63 36 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=1.235
+ $Y2=0
r64 36 38 43.7112 $w=1.68e-07 $l=6.7e-07 $layer=LI1_cond $X=1.4 $Y=0 $X2=2.07
+ $Y2=0
r65 34 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=1.15
+ $Y2=0
r66 34 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r67 32 38 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.07
+ $Y2=0
r68 32 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.125 $Y=0 $X2=2.29
+ $Y2=0
r69 31 42 4.89305 $w=1.68e-07 $l=7.5e-08 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.53
+ $Y2=0
r70 31 33 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.455 $Y=0 $X2=2.29
+ $Y2=0
r71 27 54 3.29997 $w=3.8e-07 $l=1.69245e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.817 $Y2=0
r72 27 29 19.8645 $w=3.78e-07 $l=6.55e-07 $layer=LI1_cond $X=3.685 $Y=0.085
+ $X2=3.685 $Y2=0.74
r73 23 33 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0
r74 23 25 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=2.29 $Y=0.085
+ $X2=2.29 $Y2=0.38
r75 19 51 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0
r76 19 21 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=1.235 $Y=0.085
+ $X2=1.235 $Y2=0.36
r77 18 48 4.09789 $w=1.7e-07 $l=1.73e-07 $layer=LI1_cond $X=0.345 $Y=0 $X2=0.172
+ $Y2=0
r78 17 51 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=1.235
+ $Y2=0
r79 17 18 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=1.07 $Y=0 $X2=0.345
+ $Y2=0
r80 13 48 3.07934 $w=2.55e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.172 $Y2=0
r81 13 15 13.3322 $w=2.53e-07 $l=2.95e-07 $layer=LI1_cond $X=0.217 $Y=0.085
+ $X2=0.217 $Y2=0.38
r82 4 29 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=3.525
+ $Y=0.235 $X2=3.71 $Y2=0.74
r83 3 25 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.165
+ $Y=0.235 $X2=2.29 $Y2=0.38
r84 2 21 91 $w=1.7e-07 $l=1.92614e-07 $layer=licon1_NDIFF $count=2 $X=1.075
+ $Y=0.235 $X2=1.215 $Y2=0.36
r85 1 15 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.38
.ends

