* File: sky130_fd_sc_hdll__a221oi_1.spice
* Created: Thu Aug 27 18:53:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a221oi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a221oi_1  VNB VPB C1 B2 B1 A1 A2 Y VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* Y	Y
* A2	A2
* A1	A1
* B1	B1
* B2	B2
* C1	C1
* VPB	VPB
* VNB	VNB
MM1008 N_VGND_M1008_d N_C1_M1008_g N_Y_M1008_s VNB NSHORT L=0.15 W=0.65
+ AD=0.1235 AS=0.2015 PD=1.03 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1002 A_225_47# N_B2_M1002_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65 AD=0.06825
+ AS=0.1235 PD=0.86 PS=1.03 NRD=9.228 NRS=19.38 M=1 R=4.33333 SA=75000.8
+ SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1003 N_Y_M1003_d N_B1_M1003_g A_225_47# VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.06825 PD=1.92 PS=0.86 NRD=8.304 NRS=9.228 M=1 R=4.33333 SA=75001.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1005 A_505_47# N_A1_M1005_g N_Y_M1005_s VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.2015 PD=1.03 PS=1.92 NRD=24.912 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_505_47# VNB NSHORT L=0.15 W=0.65 AD=0.18525
+ AS=0.1235 PD=1.87 PS=1.03 NRD=0 NRS=24.912 M=1 R=4.33333 SA=75000.8 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1006 N_A_117_297#_M1006_d N_C1_M1006_g N_Y_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1000 N_A_211_297#_M1000_d N_B2_M1000_g N_A_117_297#_M1006_d VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1009 N_A_117_297#_M1009_d N_B1_M1009_g N_A_211_297#_M1000_d VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1007 N_A_211_297#_M1007_d N_A1_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.175 AS=0.27 PD=1.35 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A2_M1001_g N_A_211_297#_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.29 AS=0.175 PD=2.58 PS=1.35 NRD=4.9053 NRS=12.7853 M=1 R=5.55556
+ SA=90000.7 SB=90000.2 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=6.5163 P=11.33
*
.include "sky130_fd_sc_hdll__a221oi_1.pxi.spice"
*
.ends
*
*
