# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__o21bai_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  7.360000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.145000 1.075000 7.250000 1.285000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.365000 1.075000 4.975000 1.275000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.510000 1.285000 ;
    END
  END B1_N
  PIN Y
    ANTENNADIFFAREA  1.576000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.035000 1.455000 4.765000 1.625000 ;
        RECT 1.035000 1.625000 1.375000 2.465000 ;
        RECT 1.520000 0.645000 2.925000 0.815000 ;
        RECT 2.065000 1.625000 2.315000 2.465000 ;
        RECT 2.695000 0.815000 2.925000 1.075000 ;
        RECT 2.695000 1.075000 3.195000 1.445000 ;
        RECT 2.695000 1.445000 4.765000 1.455000 ;
        RECT 3.575000 1.625000 3.825000 2.125000 ;
        RECT 4.515000 1.625000 4.765000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.360000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 7.360000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 7.360000 0.085000 ;
      RECT 0.000000  2.635000 7.360000 2.805000 ;
      RECT 0.145000  1.455000 0.850000 1.625000 ;
      RECT 0.145000  1.625000 0.475000 2.435000 ;
      RECT 0.225000  0.085000 0.395000 0.895000 ;
      RECT 0.565000  0.290000 0.945000 0.895000 ;
      RECT 0.680000  0.895000 0.945000 1.075000 ;
      RECT 0.680000  1.075000 2.525000 1.285000 ;
      RECT 0.680000  1.285000 0.850000 1.455000 ;
      RECT 0.695000  1.795000 0.865000 2.635000 ;
      RECT 1.180000  0.305000 3.395000 0.475000 ;
      RECT 1.595000  1.795000 1.845000 2.635000 ;
      RECT 2.535000  1.795000 2.785000 2.635000 ;
      RECT 3.025000  1.795000 3.355000 2.295000 ;
      RECT 3.025000  2.295000 5.235000 2.465000 ;
      RECT 3.145000  0.475000 3.395000 0.725000 ;
      RECT 3.145000  0.725000 7.155000 0.905000 ;
      RECT 3.615000  0.085000 3.785000 0.555000 ;
      RECT 3.955000  0.255000 4.335000 0.725000 ;
      RECT 4.045000  1.795000 4.295000 2.295000 ;
      RECT 4.555000  0.085000 4.725000 0.555000 ;
      RECT 4.895000  0.255000 5.275000 0.725000 ;
      RECT 4.985000  1.455000 7.115000 1.625000 ;
      RECT 4.985000  1.625000 5.235000 2.295000 ;
      RECT 5.455000  1.795000 5.705000 2.635000 ;
      RECT 5.495000  0.085000 5.665000 0.555000 ;
      RECT 5.835000  0.255000 6.215000 0.725000 ;
      RECT 5.925000  1.625000 6.175000 2.465000 ;
      RECT 6.395000  1.795000 6.645000 2.635000 ;
      RECT 6.435000  0.085000 6.605000 0.555000 ;
      RECT 6.775000  0.255000 7.155000 0.725000 ;
      RECT 6.865000  1.625000 7.115000 2.465000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
      RECT 6.125000 -0.085000 6.295000 0.085000 ;
      RECT 6.125000  2.635000 6.295000 2.805000 ;
      RECT 6.585000 -0.085000 6.755000 0.085000 ;
      RECT 6.585000  2.635000 6.755000 2.805000 ;
      RECT 7.045000 -0.085000 7.215000 0.085000 ;
      RECT 7.045000  2.635000 7.215000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__o21bai_4
