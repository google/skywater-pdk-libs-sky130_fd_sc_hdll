* File: sky130_fd_sc_hdll__a211oi_2.pex.spice
* Created: Wed Sep  2 08:16:09 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%C1 1 3 4 6 7 9 10 12 13 14 19 22
c41 1 0 8.90536e-20 $X=0.55 $Y=1.41
r42 22 23 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=1.03 $Y=1.202
+ $X2=1.055 $Y2=1.202
r43 21 22 60.0849 $w=3.65e-07 $l=4.55e-07 $layer=POLY_cond $X=0.575 $Y=1.202
+ $X2=1.03 $Y2=1.202
r44 20 21 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=0.55 $Y=1.202
+ $X2=0.575 $Y2=1.202
r45 18 20 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=0.315 $Y=1.202
+ $X2=0.55 $Y2=1.202
r46 18 19 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.315
+ $Y=1.16 $X2=0.315 $Y2=1.16
r47 13 14 12.8469 $w=3.03e-07 $l=3.4e-07 $layer=LI1_cond $X=0.252 $Y=1.19
+ $X2=0.252 $Y2=1.53
r48 13 19 1.13355 $w=3.03e-07 $l=3e-08 $layer=LI1_cond $X=0.252 $Y=1.19
+ $X2=0.252 $Y2=1.16
r49 10 23 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=1.202
r50 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.055 $Y=0.995
+ $X2=1.055 $Y2=0.56
r51 7 22 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.03 $Y=1.41
+ $X2=1.03 $Y2=1.202
r52 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.03 $Y=1.41 $X2=1.03
+ $Y2=1.985
r53 4 21 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.575 $Y=0.995
+ $X2=0.575 $Y2=1.202
r54 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.575 $Y=0.995
+ $X2=0.575 $Y2=0.56
r55 1 20 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.55 $Y=1.41
+ $X2=0.55 $Y2=1.202
r56 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.55 $Y=1.41 $X2=0.55
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%B1 1 3 4 6 7 9 10 12 13 14 15 24 26 32
c50 14 0 2.72215e-19 $X=1.165 $Y=1.53
r51 30 32 14.0598 $w=2.48e-07 $l=3.05e-07 $layer=LI1_cond $X=1.285 $Y=1.16
+ $X2=1.59 $Y2=1.16
r52 24 25 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.99 $Y=1.202
+ $X2=2.015 $Y2=1.202
r53 22 24 30.4421 $w=3.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.75 $Y=1.202
+ $X2=1.99 $Y2=1.202
r54 20 22 30.4421 $w=3.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.51 $Y=1.202
+ $X2=1.75 $Y2=1.202
r55 19 20 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.485 $Y=1.202
+ $X2=1.51 $Y2=1.202
r56 15 32 6.91466 $w=2.48e-07 $l=1.5e-07 $layer=LI1_cond $X=1.74 $Y=1.16
+ $X2=1.59 $Y2=1.16
r57 15 22 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.75
+ $Y=1.16 $X2=1.75 $Y2=1.16
r58 14 26 12.834 $w=2.18e-07 $l=2.45e-07 $layer=LI1_cond $X=1.175 $Y=1.53
+ $X2=1.175 $Y2=1.285
r59 13 26 3.64504 $w=2.2e-07 $l=1.25e-07 $layer=LI1_cond $X=1.175 $Y=1.16
+ $X2=1.175 $Y2=1.285
r60 13 30 3.20764 $w=2.5e-07 $l=1.1e-07 $layer=LI1_cond $X=1.175 $Y=1.16
+ $X2=1.285 $Y2=1.16
r61 10 25 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=1.202
r62 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.015 $Y=0.995
+ $X2=2.015 $Y2=0.56
r63 7 24 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.99 $Y=1.41
+ $X2=1.99 $Y2=1.202
r64 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.99 $Y=1.41 $X2=1.99
+ $Y2=1.985
r65 4 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.51 $Y=1.41
+ $X2=1.51 $Y2=1.202
r66 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.51 $Y=1.41 $X2=1.51
+ $Y2=1.985
r67 1 19 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=1.202
r68 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.485 $Y=0.995
+ $X2=1.485 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%A1 1 3 4 6 7 9 10 12 13 14 22 27 29
r39 27 29 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=3.005 $Y=1.16
+ $X2=3.23 $Y2=1.16
r40 22 23 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.47 $Y=1.202
+ $X2=3.495 $Y2=1.202
r41 20 22 8.24474 $w=3.8e-07 $l=6.5e-08 $layer=POLY_cond $X=3.405 $Y=1.202
+ $X2=3.47 $Y2=1.202
r42 18 20 52.6395 $w=3.8e-07 $l=4.15e-07 $layer=POLY_cond $X=2.99 $Y=1.202
+ $X2=3.405 $Y2=1.202
r43 17 18 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=2.965 $Y=1.202
+ $X2=2.99 $Y2=1.202
r44 14 29 8.0671 $w=2.48e-07 $l=1.75e-07 $layer=LI1_cond $X=3.405 $Y=1.16
+ $X2=3.23 $Y2=1.16
r45 14 20 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=3.405
+ $Y=1.16 $X2=3.405 $Y2=1.16
r46 13 27 1.61342 $w=2.48e-07 $l=3.5e-08 $layer=LI1_cond $X=2.97 $Y=1.16
+ $X2=3.005 $Y2=1.16
r47 10 23 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.495 $Y2=1.202
r48 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.495 $Y=0.995
+ $X2=3.495 $Y2=0.56
r49 7 22 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.47 $Y=1.41
+ $X2=3.47 $Y2=1.202
r50 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.47 $Y=1.41 $X2=3.47
+ $Y2=1.985
r51 4 18 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.99 $Y=1.41
+ $X2=2.99 $Y2=1.202
r52 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.99 $Y=1.41 $X2=2.99
+ $Y2=1.985
r53 1 17 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.965 $Y=0.995
+ $X2=2.965 $Y2=1.202
r54 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.965 $Y=0.995
+ $X2=2.965 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%A2 1 3 4 6 7 9 10 12 13 14 15 25 31 35
r43 25 26 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.43 $Y=1.202
+ $X2=4.455 $Y2=1.202
r44 24 31 10.372 $w=2.48e-07 $l=2.25e-07 $layer=LI1_cond $X=4.395 $Y=1.16
+ $X2=4.17 $Y2=1.16
r45 23 25 4.43947 $w=3.8e-07 $l=3.5e-08 $layer=POLY_cond $X=4.395 $Y=1.202
+ $X2=4.43 $Y2=1.202
r46 23 24 72.64 $w=1.7e-07 $l=3.4e-07 $layer=licon1_POLY $count=2 $X=4.395
+ $Y=1.16 $X2=4.395 $Y2=1.16
r47 21 23 56.4447 $w=3.8e-07 $l=4.45e-07 $layer=POLY_cond $X=3.95 $Y=1.202
+ $X2=4.395 $Y2=1.202
r48 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=3.925 $Y=1.202
+ $X2=3.95 $Y2=1.202
r49 15 35 12.276 $w=2.28e-07 $l=2.45e-07 $layer=LI1_cond $X=4.8 $Y=1.53 $X2=4.8
+ $Y2=1.285
r50 14 35 3.55828 $w=2.3e-07 $l=1.25e-07 $layer=LI1_cond $X=4.8 $Y=1.16 $X2=4.8
+ $Y2=1.285
r51 14 24 9.8303 $w=4.18e-07 $l=2.9e-07 $layer=LI1_cond $X=4.685 $Y=1.16
+ $X2=4.395 $Y2=1.16
r52 13 31 5.07075 $w=2.48e-07 $l=1.1e-07 $layer=LI1_cond $X=4.06 $Y=1.16
+ $X2=4.17 $Y2=1.16
r53 10 26 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.455 $Y=0.995
+ $X2=4.455 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.455 $Y=0.995
+ $X2=4.455 $Y2=0.56
r55 7 25 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.43 $Y=1.41
+ $X2=4.43 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.43 $Y=1.41 $X2=4.43
+ $Y2=1.985
r57 4 21 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.95 $Y=1.41
+ $X2=3.95 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.95 $Y=1.41 $X2=3.95
+ $Y2=1.985
r59 1 20 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.925 $Y=0.995
+ $X2=3.925 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.925 $Y=0.995
+ $X2=3.925 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%A_37_297# 1 2 3 12 14 15 18 20 22 24 26
r37 22 28 2.94404 $w=2.8e-07 $l=1e-07 $layer=LI1_cond $X=2.275 $Y=2.255
+ $X2=2.275 $Y2=2.355
r38 22 24 10.4955 $w=2.78e-07 $l=2.55e-07 $layer=LI1_cond $X=2.275 $Y=2.255
+ $X2=2.275 $Y2=2
r39 21 26 5.28167 $w=1.85e-07 $l=9.5e-08 $layer=LI1_cond $X=1.365 $Y=2.355
+ $X2=1.27 $Y2=2.355
r40 20 28 4.12165 $w=2e-07 $l=1.4e-07 $layer=LI1_cond $X=2.135 $Y=2.355
+ $X2=2.275 $Y2=2.355
r41 20 21 42.7 $w=1.98e-07 $l=7.7e-07 $layer=LI1_cond $X=2.135 $Y=2.355
+ $X2=1.365 $Y2=2.355
r42 16 26 1.24671 $w=1.9e-07 $l=1e-07 $layer=LI1_cond $X=1.27 $Y=2.255 $X2=1.27
+ $Y2=2.355
r43 16 18 17.8038 $w=1.88e-07 $l=3.05e-07 $layer=LI1_cond $X=1.27 $Y=2.255
+ $X2=1.27 $Y2=1.95
r44 14 26 5.28167 $w=1.85e-07 $l=1.02225e-07 $layer=LI1_cond $X=1.175 $Y=2.37
+ $X2=1.27 $Y2=2.355
r45 14 15 50.2353 $w=1.68e-07 $l=7.7e-07 $layer=LI1_cond $X=1.175 $Y=2.37
+ $X2=0.405 $Y2=2.37
r46 10 15 7.21222 $w=1.7e-07 $l=1.67183e-07 $layer=LI1_cond $X=0.275 $Y=2.285
+ $X2=0.405 $Y2=2.37
r47 10 12 14.8488 $w=2.58e-07 $l=3.35e-07 $layer=LI1_cond $X=0.275 $Y=2.285
+ $X2=0.275 $Y2=1.95
r48 3 28 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.23 $Y2=2.34
r49 3 24 600 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=2.08
+ $Y=1.485 $X2=2.23 $Y2=2
r50 2 18 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=1.12
+ $Y=1.485 $X2=1.27 $Y2=1.95
r51 1 12 300 $w=1.7e-07 $l=5.23784e-07 $layer=licon1_PDIFF $count=2 $X=0.185
+ $Y=1.485 $X2=0.31 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%Y 1 2 3 4 17 19 20 21 22 23 32 46
c46 20 0 1.85153e-19 $X=0.67 $Y=0.85
r47 23 46 0.720277 $w=3.18e-07 $l=2e-08 $layer=LI1_cond $X=0.735 $Y=1.85
+ $X2=0.735 $Y2=1.87
r48 23 43 8.64332 $w=3.18e-07 $l=2.4e-07 $layer=LI1_cond $X=0.735 $Y=1.85
+ $X2=0.735 $Y2=1.61
r49 22 43 2.88111 $w=3.18e-07 $l=8e-08 $layer=LI1_cond $X=0.735 $Y=1.53
+ $X2=0.735 $Y2=1.61
r50 21 22 12.2447 $w=3.18e-07 $l=3.4e-07 $layer=LI1_cond $X=0.735 $Y=1.19
+ $X2=0.735 $Y2=1.53
r51 20 30 3.48797 $w=3.15e-07 $l=1.0247e-07 $layer=LI1_cond $X=0.735 $Y=0.755
+ $X2=0.73 $Y2=0.655
r52 20 36 3.48797 $w=3.15e-07 $l=1e-07 $layer=LI1_cond $X=0.735 $Y=0.755
+ $X2=0.735 $Y2=0.855
r53 20 21 10.6241 $w=3.18e-07 $l=2.95e-07 $layer=LI1_cond $X=0.735 $Y=0.895
+ $X2=0.735 $Y2=1.19
r54 20 36 1.44055 $w=3.18e-07 $l=4e-08 $layer=LI1_cond $X=0.735 $Y=0.895
+ $X2=0.735 $Y2=0.855
r55 19 30 5.39046 $w=3.08e-07 $l=1.45e-07 $layer=LI1_cond $X=0.73 $Y=0.51
+ $X2=0.73 $Y2=0.655
r56 19 32 3.3458 $w=3.08e-07 $l=9e-08 $layer=LI1_cond $X=0.73 $Y=0.51 $X2=0.73
+ $Y2=0.42
r57 15 17 82.0727 $w=1.98e-07 $l=1.48e-06 $layer=LI1_cond $X=1.75 $Y=0.755
+ $X2=3.23 $Y2=0.755
r58 13 20 3.01902 $w=2e-07 $l=1.6e-07 $layer=LI1_cond $X=0.895 $Y=0.755
+ $X2=0.735 $Y2=0.755
r59 13 15 47.4136 $w=1.98e-07 $l=8.55e-07 $layer=LI1_cond $X=0.895 $Y=0.755
+ $X2=1.75 $Y2=0.755
r60 4 43 300 $w=1.7e-07 $l=2.03101e-07 $layer=licon1_PDIFF $count=2 $X=0.64
+ $Y=1.485 $X2=0.79 $Y2=1.61
r61 3 17 182 $w=1.7e-07 $l=6.07618e-07 $layer=licon1_NDIFF $count=1 $X=3.04
+ $Y=0.235 $X2=3.23 $Y2=0.755
r62 2 15 182 $w=1.7e-07 $l=6.07618e-07 $layer=licon1_NDIFF $count=1 $X=1.56
+ $Y=0.235 $X2=1.75 $Y2=0.755
r63 1 20 182 $w=1.7e-07 $l=5.90868e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.235 $X2=0.79 $Y2=0.76
r64 1 32 182 $w=1.7e-07 $l=2.45204e-07 $layer=licon1_NDIFF $count=1 $X=0.65
+ $Y=0.235 $X2=0.79 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%A_320_297# 1 2 3 12 16 18 20 22 25 27
r48 20 29 2.98511 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=4.19 $Y=1.655 $X2=4.19
+ $Y2=1.555
r49 20 22 27.5306 $w=2.68e-07 $l=6.45e-07 $layer=LI1_cond $X=4.19 $Y=1.655
+ $X2=4.19 $Y2=2.3
r50 19 27 6.58019 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=3.365 $Y=1.555
+ $X2=3.23 $Y2=1.555
r51 18 29 4.0299 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=4.055 $Y=1.555 $X2=4.19
+ $Y2=1.555
r52 18 19 38.2636 $w=1.98e-07 $l=6.9e-07 $layer=LI1_cond $X=4.055 $Y=1.555
+ $X2=3.365 $Y2=1.555
r53 14 27 0.287739 $w=2.7e-07 $l=1e-07 $layer=LI1_cond $X=3.23 $Y=1.655 $X2=3.23
+ $Y2=1.555
r54 14 16 27.5306 $w=2.68e-07 $l=6.45e-07 $layer=LI1_cond $X=3.23 $Y=1.655
+ $X2=3.23 $Y2=2.3
r55 13 25 5.04956 $w=2e-07 $l=1.9e-07 $layer=LI1_cond $X=1.915 $Y=1.555
+ $X2=1.725 $Y2=1.555
r56 12 27 6.58019 $w=2e-07 $l=1.35e-07 $layer=LI1_cond $X=3.095 $Y=1.555
+ $X2=3.23 $Y2=1.555
r57 12 13 65.4364 $w=1.98e-07 $l=1.18e-06 $layer=LI1_cond $X=3.095 $Y=1.555
+ $X2=1.915 $Y2=1.555
r58 3 29 400 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.485 $X2=4.19 $Y2=1.62
r59 3 22 400 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=4.04
+ $Y=1.485 $X2=4.19 $Y2=2.3
r60 2 27 400 $w=1.7e-07 $l=2.06761e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.23 $Y2=1.62
r61 2 16 400 $w=1.7e-07 $l=8.86834e-07 $layer=licon1_PDIFF $count=1 $X=3.08
+ $Y=1.485 $X2=3.23 $Y2=2.3
r62 1 25 300 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=2 $X=1.6
+ $Y=1.485 $X2=1.75 $Y2=1.65
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%VPWR 1 2 3 12 16 20 23 24 26 27 28 29 30
+ 31 48 52
r63 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.83 $Y=2.72
+ $X2=4.83 $Y2=2.72
r64 45 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=4.37 $Y=2.72
+ $X2=4.83 $Y2=2.72
r65 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.37 $Y=2.72
+ $X2=4.37 $Y2=2.72
r66 42 45 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=4.37 $Y2=2.72
r67 41 42 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r68 39 42 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r69 39 52 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=0.23 $Y2=2.72
r70 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r71 34 38 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=0.23 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 34 52 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r73 31 52 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=2.72
+ $X2=0.23 $Y2=2.72
r74 29 44 12.0695 $w=1.68e-07 $l=1.85e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.37 $Y2=2.72
r75 29 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.555 $Y=2.72
+ $X2=4.67 $Y2=2.72
r76 28 47 3.22941 $w=1.7e-07 $l=4.5e-08 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.83 $Y2=2.72
r77 28 30 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=4.785 $Y=2.72
+ $X2=4.67 $Y2=2.72
r78 26 41 9.45989 $w=1.68e-07 $l=1.45e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.45 $Y2=2.72
r79 26 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.595 $Y=2.72
+ $X2=3.71 $Y2=2.72
r80 25 44 35.5561 $w=1.68e-07 $l=5.45e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=4.37 $Y2=2.72
r81 25 27 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=3.825 $Y=2.72
+ $X2=3.71 $Y2=2.72
r82 23 38 6.85027 $w=1.68e-07 $l=1.05e-07 $layer=LI1_cond $X=2.635 $Y=2.72
+ $X2=2.53 $Y2=2.72
r83 23 24 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.635 $Y=2.72
+ $X2=2.75 $Y2=2.72
r84 22 41 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=3.45 $Y2=2.72
r85 22 24 6.59134 $w=1.7e-07 $l=1.15e-07 $layer=LI1_cond $X=2.865 $Y=2.72
+ $X2=2.75 $Y2=2.72
r86 18 30 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=4.67 $Y=2.635
+ $X2=4.67 $Y2=2.72
r87 18 20 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=4.67 $Y=2.635
+ $X2=4.67 $Y2=2
r88 14 27 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=3.71 $Y=2.635
+ $X2=3.71 $Y2=2.72
r89 14 16 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=3.71 $Y=2.635
+ $X2=3.71 $Y2=2
r90 10 24 0.280307 $w=2.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.72
r91 10 12 31.8174 $w=2.28e-07 $l=6.35e-07 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2
r92 3 20 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=4.52
+ $Y=1.485 $X2=4.67 $Y2=2
r93 2 16 300 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=2 $X=3.56
+ $Y=1.485 $X2=3.71 $Y2=2
r94 1 12 300 $w=1.7e-07 $l=5.74108e-07 $layer=licon1_PDIFF $count=2 $X=2.625
+ $Y=1.485 $X2=2.75 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%VGND 1 2 3 4 13 15 19 21 25 27 28 34 36
+ 49 50 56 59 64
c71 36 0 1.85153e-19 $X=1.055 $Y=0
r72 59 60 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r73 57 60 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=0 $X2=2.07
+ $Y2=0
r74 56 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=0 $X2=1.15
+ $Y2=0
r75 53 64 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r76 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r77 47 50 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r78 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r79 44 47 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r80 44 60 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r81 43 46 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r82 43 44 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r83 41 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.205
+ $Y2=0
r84 41 43 8.80749 $w=1.68e-07 $l=1.35e-07 $layer=LI1_cond $X=2.395 $Y=0 $X2=2.53
+ $Y2=0
r85 40 57 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.15
+ $Y2=0
r86 40 64 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=0.23
+ $Y2=0
r87 39 40 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r88 37 53 3.97288 $w=1.7e-07 $l=1.98e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.197
+ $Y2=0
r89 37 39 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.395 $Y=0 $X2=0.69
+ $Y2=0
r90 36 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=1.245
+ $Y2=0
r91 36 39 23.8128 $w=1.68e-07 $l=3.65e-07 $layer=LI1_cond $X=1.055 $Y=0 $X2=0.69
+ $Y2=0
r92 34 64 0.00569083 $w=4.8e-07 $l=2e-08 $layer=MET1_cond $X=0.21 $Y=0 $X2=0.23
+ $Y2=0
r93 30 49 30.9893 $w=1.68e-07 $l=4.75e-07 $layer=LI1_cond $X=4.355 $Y=0 $X2=4.83
+ $Y2=0
r94 28 46 4.24064 $w=1.68e-07 $l=6.5e-08 $layer=LI1_cond $X=3.975 $Y=0 $X2=3.91
+ $Y2=0
r95 27 32 10.9179 $w=3.78e-07 $l=3.6e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.165
+ $Y2=0.36
r96 27 30 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=4.355
+ $Y2=0
r97 27 28 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=4.165 $Y=0 $X2=3.975
+ $Y2=0
r98 23 59 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=0.085
+ $X2=2.205 $Y2=0
r99 23 25 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=2.205 $Y=0.085
+ $X2=2.205 $Y2=0.38
r100 22 56 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.435 $Y=0 $X2=1.245
+ $Y2=0
r101 21 59 9.48355 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=2.015 $Y=0 $X2=2.205
+ $Y2=0
r102 21 22 37.8396 $w=1.68e-07 $l=5.8e-07 $layer=LI1_cond $X=2.015 $Y=0
+ $X2=1.435 $Y2=0
r103 17 56 1.31983 $w=3.8e-07 $l=8.5e-08 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0
r104 17 19 8.9466 $w=3.78e-07 $l=2.95e-07 $layer=LI1_cond $X=1.245 $Y=0.085
+ $X2=1.245 $Y2=0.38
r105 13 53 3.17028 $w=2.5e-07 $l=1.15888e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.197 $Y2=0
r106 13 15 23.2793 $w=2.48e-07 $l=5.05e-07 $layer=LI1_cond $X=0.27 $Y=0.085
+ $X2=0.27 $Y2=0.59
r107 4 32 182 $w=1.7e-07 $l=2.44643e-07 $layer=licon1_NDIFF $count=1 $X=4
+ $Y=0.235 $X2=4.19 $Y2=0.36
r108 3 25 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=2.09
+ $Y=0.235 $X2=2.23 $Y2=0.38
r109 2 19 182 $w=1.7e-07 $l=2.03286e-07 $layer=licon1_NDIFF $count=1 $X=1.13
+ $Y=0.235 $X2=1.27 $Y2=0.38
r110 1 15 182 $w=1.7e-07 $l=4.12795e-07 $layer=licon1_NDIFF $count=1 $X=0.185
+ $Y=0.235 $X2=0.31 $Y2=0.59
.ends

.subckt PM_SKY130_FD_SC_HDLL__A211OI_2%A_525_47# 1 2 3 10 18 19 20
r29 20 22 4.148 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=4.71 $Y=0.635 $X2=4.71
+ $Y2=0.55
r30 18 20 6.85268 $w=2.2e-07 $l=1.71391e-07 $layer=LI1_cond $X=4.585 $Y=0.745
+ $X2=4.71 $Y2=0.635
r31 18 19 41.3832 $w=2.18e-07 $l=7.9e-07 $layer=LI1_cond $X=4.585 $Y=0.745
+ $X2=3.795 $Y2=0.745
r32 15 19 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=3.71 $Y=0.635
+ $X2=3.795 $Y2=0.745
r33 15 17 6.52406 $w=1.68e-07 $l=1e-07 $layer=LI1_cond $X=3.71 $Y=0.635 $X2=3.71
+ $Y2=0.535
r34 14 17 3.91444 $w=1.68e-07 $l=6e-08 $layer=LI1_cond $X=3.71 $Y=0.475 $X2=3.71
+ $Y2=0.535
r35 10 14 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=3.625 $Y=0.37
+ $X2=3.71 $Y2=0.475
r36 10 12 46.2121 $w=2.08e-07 $l=8.75e-07 $layer=LI1_cond $X=3.625 $Y=0.37
+ $X2=2.75 $Y2=0.37
r37 3 22 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=4.53
+ $Y=0.235 $X2=4.67 $Y2=0.55
r38 2 17 182 $w=1.7e-07 $l=3.63318e-07 $layer=licon1_NDIFF $count=1 $X=3.57
+ $Y=0.235 $X2=3.71 $Y2=0.535
r39 1 12 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=2.625
+ $Y=0.235 $X2=2.75 $Y2=0.38
.ends

