* File: sky130_fd_sc_hdll__o2bb2ai_2.spice
* Created: Wed Sep  2 08:46:28 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o2bb2ai_2.pex.spice"
.subckt sky130_fd_sc_hdll__o2bb2ai_2  VNB VPB A1_N A2_N B1 B2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B2	B2
* B1	B1
* A2_N	A2_N
* A1_N	A1_N
* VPB	VPB
* VNB	VNB
MM1004 N_VGND_M1004_d N_A1_N_M1004_g N_A_123_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2145 AS=0.08775 PD=1.96 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.3 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1001 N_A_121_297#_M1001_d N_A2_N_M1001_g N_A_123_47#_M1004_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1011 N_A_121_297#_M1001_d N_A2_N_M1011_g N_A_123_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.091 PD=1.02 PS=0.93 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A1_N_M1006_g N_A_123_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.091 PD=1.82 PS=0.93 NRD=0 NRS=0.912 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1010 N_A_503_47#_M1010_d N_A_121_297#_M1010_g N_Y_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.104 PD=1.92 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1012 N_A_503_47#_M1012_d N_A_121_297#_M1012_g N_Y_M1010_s VNB NSHORT L=0.15
+ W=0.65 AD=0.115375 AS=0.104 PD=1.005 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75002.1 A=0.0975 P=1.6 MULT=1
MM1013 N_A_503_47#_M1012_d N_B1_M1013_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.115375 AS=0.08775 PD=1.005 PS=0.92 NRD=14.76 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1002 N_A_503_47#_M1002_d N_B2_M1002_g N_VGND_M1013_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.6
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1017 N_A_503_47#_M1002_d N_B2_M1017_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1018 N_A_503_47#_M1018_d N_B1_M1018_g N_VGND_M1017_s VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75002.6
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_A_121_297#_M1000_d N_A1_N_M1000_g N_VPWR_M1000_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90004.9 A=0.18 P=2.36 MULT=1
MM1007 N_A_121_297#_M1000_d N_A2_N_M1007_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.7 SB=90004.5 A=0.18 P=2.36 MULT=1
MM1015 N_A_121_297#_M1015_d N_A2_N_M1015_g N_VPWR_M1007_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.145 PD=1.3 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90004 A=0.18 P=2.36 MULT=1
MM1003 N_A_121_297#_M1015_d N_A1_N_M1003_g N_VPWR_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.38 PD=1.3 PS=1.76 NRD=2.9353 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1009 N_VPWR_M1003_s N_A_121_297#_M1009_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.38 AS=0.145 PD=1.76 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1016_d N_A_121_297#_M1016_g N_Y_M1009_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1625 AS=0.145 PD=1.325 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90003 SB=90002.1 A=0.18 P=2.36 MULT=1
MM1014 N_A_788_297#_M1014_d N_B1_M1014_g N_VPWR_M1016_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1625 PD=1.29 PS=1.325 NRD=0.9653 NRS=7.8603 M=1 R=5.55556
+ SA=90003.5 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1005 N_A_788_297#_M1014_d N_B2_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1008 N_A_788_297#_M1008_d N_B2_M1008_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90004.5 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1019 N_A_788_297#_M1008_d N_B1_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.295 PD=1.29 PS=2.59 NRD=0.9653 NRS=1.9503 M=1 R=5.55556
+ SA=90004.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.2078 P=15.93
pX21_noxref noxref_14 A1_N A1_N PROBETYPE=1
pX22_noxref noxref_15 A2_N A2_N PROBETYPE=1
pX23_noxref noxref_16 B2 B2 PROBETYPE=1
*
.include "sky130_fd_sc_hdll__o2bb2ai_2.pxi.spice"
*
.ends
*
*
