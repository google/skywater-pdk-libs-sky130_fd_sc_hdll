* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__nand2_6 A B VGND VNB VPB VPWR Y
X0 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X15 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR A Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_27_47# A Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 a_27_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X20 Y A a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 VGND B a_27_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
.ends
