* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__a2bb2oi_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR Y
X0 a_27_297# a_455_21# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 a_695_297# A1_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 Y B2 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 Y a_455_21# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 VGND A2_N a_455_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X5 a_455_21# A2_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 a_455_21# A1_N VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 a_27_297# B1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X8 a_455_21# A2_N a_695_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 VGND a_455_21# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VPWR B1 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X11 a_27_297# B2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_119_47# B1 VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X13 a_119_47# B2 Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X14 a_695_297# A2_N a_455_21# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 VGND B1 a_119_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR B2 a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 Y a_455_21# a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 VPWR A1_N a_695_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 VGND A1_N a_455_21# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
