* File: sky130_fd_sc_hdll__bufbuf_16.pxi.spice
* Created: Wed Sep  2 08:24:44 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%A N_A_c_222_n N_A_M1022_g N_A_c_223_n
+ N_A_M1037_g A PM_SKY130_FD_SC_HDLL__BUFBUF_16%A
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_117_297# N_A_117_297#_M1037_d
+ N_A_117_297#_M1022_d N_A_117_297#_M1020_g N_A_117_297#_c_255_n
+ N_A_117_297#_M1027_g N_A_117_297#_M1038_g N_A_117_297#_c_256_n
+ N_A_117_297#_M1035_g N_A_117_297#_c_257_n N_A_117_297#_M1042_g
+ N_A_117_297#_M1050_g N_A_117_297#_c_248_n N_A_117_297#_c_258_n
+ N_A_117_297#_c_249_n N_A_117_297#_c_250_n N_A_117_297#_c_251_n
+ N_A_117_297#_c_259_n N_A_117_297#_c_252_n N_A_117_297#_c_253_n
+ N_A_117_297#_c_254_n PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_117_297#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_225_47# N_A_225_47#_M1020_s
+ N_A_225_47#_M1038_s N_A_225_47#_M1027_s N_A_225_47#_M1035_s
+ N_A_225_47#_M1012_g N_A_225_47#_c_358_n N_A_225_47#_M1005_g
+ N_A_225_47#_M1014_g N_A_225_47#_c_359_n N_A_225_47#_M1008_g
+ N_A_225_47#_M1023_g N_A_225_47#_c_360_n N_A_225_47#_M1010_g
+ N_A_225_47#_M1033_g N_A_225_47#_c_361_n N_A_225_47#_M1031_g
+ N_A_225_47#_M1045_g N_A_225_47#_c_362_n N_A_225_47#_M1039_g
+ N_A_225_47#_c_363_n N_A_225_47#_M1049_g N_A_225_47#_M1047_g
+ N_A_225_47#_c_348_n N_A_225_47#_c_364_n N_A_225_47#_c_349_n
+ N_A_225_47#_c_350_n N_A_225_47#_c_365_n N_A_225_47#_c_366_n
+ N_A_225_47#_c_396_n N_A_225_47#_c_398_n N_A_225_47#_c_351_n
+ N_A_225_47#_c_367_n N_A_225_47#_c_352_n N_A_225_47#_c_353_n
+ N_A_225_47#_c_354_n N_A_225_47#_c_355_n N_A_225_47#_c_369_n
+ N_A_225_47#_c_356_n N_A_225_47#_c_357_n
+ PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_225_47#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_589_47# N_A_589_47#_M1012_d
+ N_A_589_47#_M1023_d N_A_589_47#_M1045_d N_A_589_47#_M1005_s
+ N_A_589_47#_M1010_s N_A_589_47#_M1039_s N_A_589_47#_M1001_g
+ N_A_589_47#_c_583_n N_A_589_47#_M1000_g N_A_589_47#_M1002_g
+ N_A_589_47#_c_584_n N_A_589_47#_M1004_g N_A_589_47#_M1003_g
+ N_A_589_47#_c_585_n N_A_589_47#_M1009_g N_A_589_47#_M1006_g
+ N_A_589_47#_c_586_n N_A_589_47#_M1011_g N_A_589_47#_M1007_g
+ N_A_589_47#_c_587_n N_A_589_47#_M1013_g N_A_589_47#_M1015_g
+ N_A_589_47#_c_588_n N_A_589_47#_M1016_g N_A_589_47#_M1017_g
+ N_A_589_47#_c_589_n N_A_589_47#_M1019_g N_A_589_47#_M1018_g
+ N_A_589_47#_c_590_n N_A_589_47#_M1025_g N_A_589_47#_M1021_g
+ N_A_589_47#_c_591_n N_A_589_47#_M1029_g N_A_589_47#_M1024_g
+ N_A_589_47#_c_592_n N_A_589_47#_M1030_g N_A_589_47#_M1026_g
+ N_A_589_47#_c_593_n N_A_589_47#_M1032_g N_A_589_47#_M1028_g
+ N_A_589_47#_c_594_n N_A_589_47#_M1036_g N_A_589_47#_M1034_g
+ N_A_589_47#_c_595_n N_A_589_47#_M1040_g N_A_589_47#_M1043_g
+ N_A_589_47#_c_596_n N_A_589_47#_M1041_g N_A_589_47#_M1048_g
+ N_A_589_47#_c_597_n N_A_589_47#_M1044_g N_A_589_47#_c_598_n
+ N_A_589_47#_M1046_g N_A_589_47#_M1051_g N_A_589_47#_c_607_n
+ N_A_589_47#_c_608_n N_A_589_47#_c_572_n N_A_589_47#_c_573_n
+ N_A_589_47#_c_599_n N_A_589_47#_c_600_n N_A_589_47#_c_636_n
+ N_A_589_47#_c_640_n N_A_589_47#_c_574_n N_A_589_47#_c_601_n
+ N_A_589_47#_c_652_n N_A_589_47#_c_654_n N_A_589_47#_c_575_n
+ N_A_589_47#_c_602_n N_A_589_47#_c_576_n N_A_589_47#_c_577_n
+ N_A_589_47#_c_578_n N_A_589_47#_c_579_n N_A_589_47#_c_604_n
+ N_A_589_47#_c_580_n N_A_589_47#_c_605_n N_A_589_47#_c_581_n
+ N_A_589_47#_c_582_n PM_SKY130_FD_SC_HDLL__BUFBUF_16%A_589_47#
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%VPWR N_VPWR_M1022_s N_VPWR_M1027_d
+ N_VPWR_M1042_d N_VPWR_M1008_d N_VPWR_M1031_d N_VPWR_M1049_d N_VPWR_M1004_s
+ N_VPWR_M1011_s N_VPWR_M1016_s N_VPWR_M1025_s N_VPWR_M1030_s N_VPWR_M1036_s
+ N_VPWR_M1041_s N_VPWR_M1046_s N_VPWR_c_1019_n N_VPWR_c_1020_n N_VPWR_c_1021_n
+ N_VPWR_c_1022_n N_VPWR_c_1023_n N_VPWR_c_1024_n N_VPWR_c_1025_n
+ N_VPWR_c_1026_n N_VPWR_c_1027_n N_VPWR_c_1028_n N_VPWR_c_1029_n
+ N_VPWR_c_1030_n N_VPWR_c_1031_n N_VPWR_c_1032_n N_VPWR_c_1033_n
+ N_VPWR_c_1034_n N_VPWR_c_1035_n N_VPWR_c_1036_n N_VPWR_c_1037_n
+ N_VPWR_c_1038_n N_VPWR_c_1039_n N_VPWR_c_1040_n N_VPWR_c_1041_n
+ N_VPWR_c_1042_n N_VPWR_c_1043_n N_VPWR_c_1044_n N_VPWR_c_1045_n
+ N_VPWR_c_1046_n N_VPWR_c_1047_n N_VPWR_c_1048_n N_VPWR_c_1049_n
+ N_VPWR_c_1050_n N_VPWR_c_1051_n N_VPWR_c_1052_n N_VPWR_c_1053_n
+ N_VPWR_c_1054_n N_VPWR_c_1055_n N_VPWR_c_1056_n N_VPWR_c_1057_n
+ N_VPWR_c_1058_n VPWR N_VPWR_c_1059_n N_VPWR_c_1018_n VPWR
+ PM_SKY130_FD_SC_HDLL__BUFBUF_16%VPWR
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%X N_X_M1001_s N_X_M1003_s N_X_M1007_s
+ N_X_M1017_s N_X_M1021_s N_X_M1026_s N_X_M1034_s N_X_M1048_s N_X_M1000_d
+ N_X_M1009_d N_X_M1013_d N_X_M1019_d N_X_M1029_d N_X_M1032_d N_X_M1040_d
+ N_X_M1044_d N_X_c_1272_n N_X_c_1270_n N_X_c_1271_n N_X_c_1235_n N_X_c_1236_n
+ N_X_c_1252_n N_X_c_1253_n N_X_c_1299_n N_X_c_1301_n N_X_c_1305_n N_X_c_1237_n
+ N_X_c_1254_n N_X_c_1317_n N_X_c_1319_n N_X_c_1323_n N_X_c_1238_n N_X_c_1255_n
+ N_X_c_1335_n N_X_c_1339_n N_X_c_1239_n N_X_c_1256_n N_X_c_1351_n N_X_c_1355_n
+ N_X_c_1240_n N_X_c_1257_n N_X_c_1367_n N_X_c_1371_n N_X_c_1241_n N_X_c_1258_n
+ N_X_c_1383_n N_X_c_1387_n N_X_c_1242_n N_X_c_1259_n N_X_c_1399_n N_X_c_1401_n
+ N_X_c_1243_n N_X_c_1260_n N_X_c_1244_n N_X_c_1261_n N_X_c_1245_n N_X_c_1262_n
+ N_X_c_1246_n N_X_c_1263_n N_X_c_1247_n N_X_c_1264_n N_X_c_1248_n N_X_c_1265_n
+ N_X_c_1249_n N_X_c_1266_n N_X_c_1250_n N_X_c_1267_n X X
+ PM_SKY130_FD_SC_HDLL__BUFBUF_16%X
x_PM_SKY130_FD_SC_HDLL__BUFBUF_16%VGND N_VGND_M1037_s N_VGND_M1020_d
+ N_VGND_M1050_d N_VGND_M1014_s N_VGND_M1033_s N_VGND_M1047_s N_VGND_M1002_d
+ N_VGND_M1006_d N_VGND_M1015_d N_VGND_M1018_d N_VGND_M1024_d N_VGND_M1028_d
+ N_VGND_M1043_d N_VGND_M1051_d N_VGND_c_1598_n N_VGND_c_1599_n N_VGND_c_1600_n
+ N_VGND_c_1601_n N_VGND_c_1602_n N_VGND_c_1603_n N_VGND_c_1604_n
+ N_VGND_c_1605_n N_VGND_c_1606_n N_VGND_c_1607_n N_VGND_c_1608_n
+ N_VGND_c_1609_n N_VGND_c_1610_n N_VGND_c_1611_n N_VGND_c_1612_n
+ N_VGND_c_1613_n N_VGND_c_1614_n N_VGND_c_1615_n N_VGND_c_1616_n
+ N_VGND_c_1617_n N_VGND_c_1618_n N_VGND_c_1619_n N_VGND_c_1620_n
+ N_VGND_c_1621_n N_VGND_c_1622_n N_VGND_c_1623_n N_VGND_c_1624_n
+ N_VGND_c_1625_n N_VGND_c_1626_n N_VGND_c_1627_n N_VGND_c_1628_n
+ N_VGND_c_1629_n N_VGND_c_1630_n N_VGND_c_1631_n N_VGND_c_1632_n
+ N_VGND_c_1633_n N_VGND_c_1634_n N_VGND_c_1635_n N_VGND_c_1636_n
+ N_VGND_c_1637_n VGND N_VGND_c_1638_n N_VGND_c_1639_n VGND
+ PM_SKY130_FD_SC_HDLL__BUFBUF_16%VGND
cc_1 VNB N_A_c_222_n 0.0476248f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A_c_223_n 0.0247479f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB A 0.00738464f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_4 VNB N_A_117_297#_M1020_g 0.0221524f $X=-0.19 $Y=-0.24 $X2=0.352 $Y2=1.16
cc_5 VNB N_A_117_297#_M1038_g 0.0188756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_6 VNB N_A_117_297#_M1050_g 0.0185511f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_A_117_297#_c_248_n 0.00434074f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_8 VNB N_A_117_297#_c_249_n 0.00455418f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_117_297#_c_250_n 0.0210275f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A_117_297#_c_251_n 0.00261228f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_117_297#_c_252_n 7.96864e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_117_297#_c_253_n 0.00292873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_117_297#_c_254_n 0.0684039f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_225_47#_M1012_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_225_47#_M1014_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_225_47#_M1023_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_225_47#_M1033_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_225_47#_M1045_g 0.0188753f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_225_47#_M1047_g 0.0185509f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_225_47#_c_348_n 0.00451034f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_225_47#_c_349_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_225_47#_c_350_n 0.004399f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_A_225_47#_c_351_n 0.00102469f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_A_225_47#_c_352_n 0.00304777f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_A_225_47#_c_353_n 5.26104e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_A_225_47#_c_354_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_A_225_47#_c_355_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_A_225_47#_c_356_n 0.00153756f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_A_225_47#_c_357_n 0.13593f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_A_589_47#_M1001_g 0.0181991f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_A_589_47#_M1002_g 0.0183796f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_A_589_47#_M1003_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_A_589_47#_M1006_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_A_589_47#_M1007_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_A_589_47#_M1015_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VNB N_A_589_47#_M1017_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_A_589_47#_M1018_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_A_589_47#_M1021_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_589_47#_M1024_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_A_589_47#_M1026_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_A_589_47#_M1028_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_A_589_47#_M1034_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_A_589_47#_M1043_g 0.0183855f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_A_589_47#_M1048_g 0.0188758f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_A_589_47#_M1051_g 0.0218157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_A_589_47#_c_572_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_A_589_47#_c_573_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_A_589_47#_c_574_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_A_589_47#_c_575_n 9.58484e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_A_589_47#_c_576_n 0.00305698f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VNB N_A_589_47#_c_577_n 5.27693e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_52 VNB N_A_589_47#_c_578_n 0.00343466f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_53 VNB N_A_589_47#_c_579_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_54 VNB N_A_589_47#_c_580_n 0.00278347f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_55 VNB N_A_589_47#_c_581_n 0.00163661f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_56 VNB N_A_589_47#_c_582_n 0.376438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_57 VNB N_VPWR_c_1018_n 0.554392f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_58 VNB N_X_c_1235_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_59 VNB N_X_c_1236_n 0.00253087f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_60 VNB N_X_c_1237_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_61 VNB N_X_c_1238_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_62 VNB N_X_c_1239_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_63 VNB N_X_c_1240_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_64 VNB N_X_c_1241_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_65 VNB N_X_c_1242_n 0.00247798f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_66 VNB N_X_c_1243_n 0.00991015f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_67 VNB N_X_c_1244_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_68 VNB N_X_c_1245_n 0.00253075f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_69 VNB N_X_c_1246_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_70 VNB N_X_c_1247_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_71 VNB N_X_c_1248_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_72 VNB N_X_c_1249_n 0.0025306f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_73 VNB N_X_c_1250_n 0.00263423f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_74 VNB X 0.0213249f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_75 VNB N_VGND_c_1598_n 0.0110515f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_76 VNB N_VGND_c_1599_n 0.00656836f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_77 VNB N_VGND_c_1600_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_78 VNB N_VGND_c_1601_n 0.00467156f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_79 VNB N_VGND_c_1602_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_80 VNB N_VGND_c_1603_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_81 VNB N_VGND_c_1604_n 0.00466605f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_82 VNB N_VGND_c_1605_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_83 VNB N_VGND_c_1606_n 0.00467908f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_84 VNB N_VGND_c_1607_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_85 VNB N_VGND_c_1608_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_86 VNB N_VGND_c_1609_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_87 VNB N_VGND_c_1610_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_88 VNB N_VGND_c_1611_n 0.00468459f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_89 VNB N_VGND_c_1612_n 0.0130849f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_90 VNB N_VGND_c_1613_n 0.00472845f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_91 VNB N_VGND_c_1614_n 0.0334789f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_92 VNB N_VGND_c_1615_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_93 VNB N_VGND_c_1616_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_94 VNB N_VGND_c_1617_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_95 VNB N_VGND_c_1618_n 0.0200002f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_96 VNB N_VGND_c_1619_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_97 VNB N_VGND_c_1620_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_98 VNB N_VGND_c_1621_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_99 VNB N_VGND_c_1622_n 0.0193874f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_100 VNB N_VGND_c_1623_n 0.00323954f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_101 VNB N_VGND_c_1624_n 0.0198969f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_102 VNB N_VGND_c_1625_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_103 VNB N_VGND_c_1626_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_104 VNB N_VGND_c_1627_n 0.00324139f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_105 VNB N_VGND_c_1628_n 0.0193636f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_106 VNB N_VGND_c_1629_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_107 VNB N_VGND_c_1630_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_108 VNB N_VGND_c_1631_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_109 VNB N_VGND_c_1632_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_110 VNB N_VGND_c_1633_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_111 VNB N_VGND_c_1634_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_112 VNB N_VGND_c_1635_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_113 VNB N_VGND_c_1636_n 0.0193723f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_114 VNB N_VGND_c_1637_n 0.00324157f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_115 VNB N_VGND_c_1638_n 0.0194241f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_116 VNB N_VGND_c_1639_n 0.611674f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_117 VPB N_A_c_222_n 0.0442248f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_118 VPB N_A_117_297#_c_255_n 0.0194367f $X=-0.19 $Y=1.305 $X2=0.275 $Y2=1.16
cc_119 VPB N_A_117_297#_c_256_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_120 VPB N_A_117_297#_c_257_n 0.0159693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_121 VPB N_A_117_297#_c_258_n 0.00771792f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_122 VPB N_A_117_297#_c_259_n 0.00276992f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_123 VPB N_A_117_297#_c_252_n 0.00382457f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_124 VPB N_A_117_297#_c_254_n 0.0203235f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_125 VPB N_A_225_47#_c_358_n 0.0162292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_126 VPB N_A_225_47#_c_359_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_127 VPB N_A_225_47#_c_360_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_128 VPB N_A_225_47#_c_361_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_129 VPB N_A_225_47#_c_362_n 0.0158857f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_130 VPB N_A_225_47#_c_363_n 0.0159692f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_131 VPB N_A_225_47#_c_364_n 0.00788153f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_132 VPB N_A_225_47#_c_365_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_133 VPB N_A_225_47#_c_366_n 0.00454699f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_134 VPB N_A_225_47#_c_367_n 0.00100785f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_135 VPB N_A_225_47#_c_353_n 0.00252324f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_136 VPB N_A_225_47#_c_369_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_137 VPB N_A_225_47#_c_357_n 0.0384682f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_138 VPB N_A_589_47#_c_583_n 0.0162292f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_139 VPB N_A_589_47#_c_584_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_140 VPB N_A_589_47#_c_585_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_A_589_47#_c_586_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_A_589_47#_c_587_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_A_589_47#_c_588_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_A_589_47#_c_589_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_A_589_47#_c_590_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_A_589_47#_c_591_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_A_589_47#_c_592_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_A_589_47#_c_593_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_A_589_47#_c_594_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_A_589_47#_c_595_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_A_589_47#_c_596_n 0.0158869f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_A_589_47#_c_597_n 0.0158858f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_A_589_47#_c_598_n 0.0191645f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_A_589_47#_c_599_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_A_589_47#_c_600_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_A_589_47#_c_601_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_A_589_47#_c_602_n 9.4165e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_A_589_47#_c_577_n 0.0025308f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_A_589_47#_c_604_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_A_589_47#_c_605_n 0.00179747f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_A_589_47#_c_582_n 0.101888f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_1019_n 0.0110239f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_VPWR_c_1020_n 0.00749784f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB N_VPWR_c_1021_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 VPB N_VPWR_c_1022_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_166 VPB N_VPWR_c_1023_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_167 VPB N_VPWR_c_1024_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_168 VPB N_VPWR_c_1025_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_169 VPB N_VPWR_c_1026_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_170 VPB N_VPWR_c_1027_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_171 VPB N_VPWR_c_1028_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_172 VPB N_VPWR_c_1029_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_173 VPB N_VPWR_c_1030_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_174 VPB N_VPWR_c_1031_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_175 VPB N_VPWR_c_1032_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_176 VPB N_VPWR_c_1033_n 0.0135791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_177 VPB N_VPWR_c_1034_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_178 VPB N_VPWR_c_1035_n 0.03408f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_179 VPB N_VPWR_c_1036_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_180 VPB N_VPWR_c_1037_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_181 VPB N_VPWR_c_1038_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_182 VPB N_VPWR_c_1039_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_183 VPB N_VPWR_c_1040_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_184 VPB N_VPWR_c_1041_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_185 VPB N_VPWR_c_1042_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_186 VPB N_VPWR_c_1043_n 0.020564f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_187 VPB N_VPWR_c_1044_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_188 VPB N_VPWR_c_1045_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_189 VPB N_VPWR_c_1046_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_190 VPB N_VPWR_c_1047_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_191 VPB N_VPWR_c_1048_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_192 VPB N_VPWR_c_1049_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_193 VPB N_VPWR_c_1050_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_194 VPB N_VPWR_c_1051_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_195 VPB N_VPWR_c_1052_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_196 VPB N_VPWR_c_1053_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_197 VPB N_VPWR_c_1054_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_198 VPB N_VPWR_c_1055_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_199 VPB N_VPWR_c_1056_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_200 VPB N_VPWR_c_1057_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_201 VPB N_VPWR_c_1058_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_202 VPB N_VPWR_c_1059_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_203 VPB N_VPWR_c_1018_n 0.0599731f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_204 VPB N_X_c_1252_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_205 VPB N_X_c_1253_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_206 VPB N_X_c_1254_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_207 VPB N_X_c_1255_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_208 VPB N_X_c_1256_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_209 VPB N_X_c_1257_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_210 VPB N_X_c_1258_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_211 VPB N_X_c_1259_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_212 VPB N_X_c_1260_n 7.91715e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_213 VPB N_X_c_1261_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_214 VPB N_X_c_1262_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_215 VPB N_X_c_1263_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_216 VPB N_X_c_1264_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_217 VPB N_X_c_1265_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_218 VPB N_X_c_1266_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_219 VPB N_X_c_1267_n 0.00176159f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_220 VPB X 0.00742067f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_221 VPB X 0.0114825f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_222 N_A_c_223_n N_A_117_297#_c_248_n 0.00719164f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_223 N_A_c_222_n N_A_117_297#_c_258_n 0.0126029f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_223_n N_A_117_297#_c_249_n 0.00718626f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_225 N_A_c_223_n N_A_117_297#_c_251_n 0.00506895f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_226 N_A_c_222_n N_A_117_297#_c_259_n 0.00566585f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_227 N_A_c_222_n N_A_117_297#_c_252_n 0.00713327f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_228 N_A_c_222_n N_A_117_297#_c_253_n 0.00595469f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_229 A N_A_117_297#_c_253_n 0.0138154f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_230 N_A_c_223_n N_A_225_47#_c_350_n 3.65437e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_231 N_A_c_222_n N_A_225_47#_c_366_n 4.05342e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_232 N_A_c_222_n N_VPWR_c_1020_n 0.0124572f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_233 A N_VPWR_c_1020_n 0.0136987f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_234 N_A_c_222_n N_VPWR_c_1035_n 0.00597712f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_222_n N_VPWR_c_1018_n 0.0121883f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_c_222_n N_VGND_c_1599_n 0.00431355f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_237 N_A_c_223_n N_VGND_c_1599_n 0.00643264f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_238 A N_VGND_c_1599_n 0.0136981f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_239 N_A_c_223_n N_VGND_c_1614_n 0.00466005f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_240 N_A_c_223_n N_VGND_c_1639_n 0.0101005f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_241 N_A_117_297#_M1050_g N_A_225_47#_M1012_g 0.0207193f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_242 N_A_117_297#_c_257_n N_A_225_47#_c_358_n 0.0215651f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_243 N_A_117_297#_M1020_g N_A_225_47#_c_348_n 0.00693104f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_244 N_A_117_297#_M1038_g N_A_225_47#_c_348_n 5.47935e-19 $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_245 N_A_117_297#_c_248_n N_A_225_47#_c_348_n 0.0368926f $X=0.73 $Y=0.4 $X2=0
+ $Y2=0
cc_246 N_A_117_297#_c_255_n N_A_225_47#_c_364_n 0.0112091f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_247 N_A_117_297#_c_256_n N_A_225_47#_c_364_n 7.06303e-19 $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_248 N_A_117_297#_c_259_n N_A_225_47#_c_364_n 0.0660799f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_249 N_A_117_297#_M1020_g N_A_225_47#_c_349_n 0.00879805f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_250 N_A_117_297#_M1038_g N_A_225_47#_c_349_n 0.00879805f $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_251 N_A_117_297#_c_250_n N_A_225_47#_c_349_n 0.03957f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_252 N_A_117_297#_c_254_n N_A_225_47#_c_349_n 0.0031956f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_253 N_A_117_297#_M1020_g N_A_225_47#_c_350_n 0.00126794f $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_254 N_A_117_297#_c_250_n N_A_225_47#_c_350_n 0.0278128f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_255 N_A_117_297#_c_251_n N_A_225_47#_c_350_n 0.0140416f $X=0.705 $Y=0.905
+ $X2=0 $Y2=0
cc_256 N_A_117_297#_c_255_n N_A_225_47#_c_365_n 0.0137916f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_257 N_A_117_297#_c_256_n N_A_225_47#_c_365_n 0.0101048f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_258 N_A_117_297#_c_250_n N_A_225_47#_c_365_n 0.0394547f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_259 N_A_117_297#_c_254_n N_A_225_47#_c_365_n 0.00720931f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_260 N_A_117_297#_c_255_n N_A_225_47#_c_366_n 0.00138874f $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_261 N_A_117_297#_c_250_n N_A_225_47#_c_366_n 0.0279779f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_262 N_A_117_297#_c_259_n N_A_225_47#_c_366_n 0.0140417f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_263 N_A_117_297#_c_254_n N_A_225_47#_c_366_n 3.20658e-19 $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_264 N_A_117_297#_M1020_g N_A_225_47#_c_396_n 5.25882e-19 $X=1.46 $Y=0.56
+ $X2=0 $Y2=0
cc_265 N_A_117_297#_M1038_g N_A_225_47#_c_396_n 0.00657592f $X=1.93 $Y=0.56
+ $X2=0 $Y2=0
cc_266 N_A_117_297#_c_255_n N_A_225_47#_c_398_n 7.33057e-19 $X=1.485 $Y=1.41
+ $X2=0 $Y2=0
cc_267 N_A_117_297#_c_256_n N_A_225_47#_c_398_n 0.0137692f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_268 N_A_117_297#_c_257_n N_A_225_47#_c_398_n 0.0112091f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_269 N_A_117_297#_M1050_g N_A_225_47#_c_351_n 0.0116573f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_270 N_A_117_297#_c_257_n N_A_225_47#_c_367_n 0.0151183f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_271 N_A_117_297#_c_254_n N_A_225_47#_c_367_n 3.58038e-19 $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_272 N_A_117_297#_M1050_g N_A_225_47#_c_352_n 0.00410511f $X=2.45 $Y=0.56
+ $X2=0 $Y2=0
cc_273 N_A_117_297#_c_257_n N_A_225_47#_c_353_n 8.16926e-19 $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_274 N_A_117_297#_c_254_n N_A_225_47#_c_353_n 0.00327205f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_275 N_A_117_297#_M1038_g N_A_225_47#_c_355_n 0.0011682f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_276 N_A_117_297#_c_250_n N_A_225_47#_c_355_n 0.0307156f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_277 N_A_117_297#_c_254_n N_A_225_47#_c_355_n 0.00450461f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_278 N_A_117_297#_c_256_n N_A_225_47#_c_369_n 0.00259297f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_279 N_A_117_297#_c_257_n N_A_225_47#_c_369_n 0.00107777f $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_280 N_A_117_297#_c_250_n N_A_225_47#_c_369_n 0.0305808f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_281 N_A_117_297#_c_254_n N_A_225_47#_c_369_n 0.00723098f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_282 N_A_117_297#_c_250_n N_A_225_47#_c_356_n 0.014524f $X=2.06 $Y=1.16 $X2=0
+ $Y2=0
cc_283 N_A_117_297#_c_254_n N_A_225_47#_c_356_n 0.00220849f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_284 N_A_117_297#_c_254_n N_A_225_47#_c_357_n 0.0207193f $X=2.425 $Y=1.217
+ $X2=0 $Y2=0
cc_285 N_A_117_297#_M1050_g N_A_589_47#_c_607_n 5.33681e-19 $X=2.45 $Y=0.56
+ $X2=0 $Y2=0
cc_286 N_A_117_297#_c_257_n N_A_589_47#_c_608_n 7.33057e-19 $X=2.425 $Y=1.41
+ $X2=0 $Y2=0
cc_287 N_A_117_297#_c_259_n N_VPWR_c_1020_n 0.0761623f $X=0.73 $Y=1.63 $X2=0
+ $Y2=0
cc_288 N_A_117_297#_c_255_n N_VPWR_c_1021_n 0.00547044f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_289 N_A_117_297#_c_256_n N_VPWR_c_1021_n 0.00497803f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_290 N_A_117_297#_c_257_n N_VPWR_c_1022_n 0.00547044f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_291 N_A_117_297#_c_255_n N_VPWR_c_1035_n 0.00673617f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_292 N_A_117_297#_c_258_n N_VPWR_c_1035_n 0.0244686f $X=0.73 $Y=2.31 $X2=0
+ $Y2=0
cc_293 N_A_117_297#_c_256_n N_VPWR_c_1037_n 0.00597712f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_294 N_A_117_297#_c_257_n N_VPWR_c_1037_n 0.00673617f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_295 N_A_117_297#_M1022_d N_VPWR_c_1018_n 0.00217517f $X=0.585 $Y=1.485 $X2=0
+ $Y2=0
cc_296 N_A_117_297#_c_255_n N_VPWR_c_1018_n 0.0131262f $X=1.485 $Y=1.41 $X2=0
+ $Y2=0
cc_297 N_A_117_297#_c_256_n N_VPWR_c_1018_n 0.00999457f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_298 N_A_117_297#_c_257_n N_VPWR_c_1018_n 0.011869f $X=2.425 $Y=1.41 $X2=0
+ $Y2=0
cc_299 N_A_117_297#_c_258_n N_VPWR_c_1018_n 0.0141694f $X=0.73 $Y=2.31 $X2=0
+ $Y2=0
cc_300 N_A_117_297#_c_248_n N_VGND_c_1599_n 0.0481407f $X=0.73 $Y=0.4 $X2=0
+ $Y2=0
cc_301 N_A_117_297#_M1020_g N_VGND_c_1600_n 0.00390178f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_302 N_A_117_297#_M1038_g N_VGND_c_1600_n 0.00276126f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_303 N_A_117_297#_M1050_g N_VGND_c_1601_n 0.00268723f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_304 N_A_117_297#_M1020_g N_VGND_c_1614_n 0.00424619f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_305 N_A_117_297#_c_248_n N_VGND_c_1614_n 0.0236681f $X=0.73 $Y=0.4 $X2=0
+ $Y2=0
cc_306 N_A_117_297#_M1038_g N_VGND_c_1616_n 0.00424619f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_307 N_A_117_297#_M1050_g N_VGND_c_1616_n 0.00439206f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_308 N_A_117_297#_M1037_d N_VGND_c_1639_n 0.0020946f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_309 N_A_117_297#_M1020_g N_VGND_c_1639_n 0.00731205f $X=1.46 $Y=0.56 $X2=0
+ $Y2=0
cc_310 N_A_117_297#_M1038_g N_VGND_c_1639_n 0.00610552f $X=1.93 $Y=0.56 $X2=0
+ $Y2=0
cc_311 N_A_117_297#_M1050_g N_VGND_c_1639_n 0.00618081f $X=2.45 $Y=0.56 $X2=0
+ $Y2=0
cc_312 N_A_117_297#_c_248_n N_VGND_c_1639_n 0.0140809f $X=0.73 $Y=0.4 $X2=0
+ $Y2=0
cc_313 N_A_225_47#_M1047_g N_A_589_47#_M1001_g 0.0207158f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_314 N_A_225_47#_c_363_n N_A_589_47#_c_583_n 0.0216821f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_315 N_A_225_47#_M1012_g N_A_589_47#_c_607_n 0.0065059f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_316 N_A_225_47#_M1014_g N_A_589_47#_c_607_n 0.00693104f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_317 N_A_225_47#_M1023_g N_A_589_47#_c_607_n 5.47131e-19 $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_318 N_A_225_47#_c_358_n N_A_589_47#_c_608_n 0.0137692f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_319 N_A_225_47#_c_359_n N_A_589_47#_c_608_n 0.0115459f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_320 N_A_225_47#_c_360_n N_A_589_47#_c_608_n 7.68612e-19 $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_321 N_A_225_47#_c_398_n N_A_589_47#_c_608_n 0.00486061f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_322 N_A_225_47#_M1014_g N_A_589_47#_c_572_n 0.00879805f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_323 N_A_225_47#_M1023_g N_A_589_47#_c_572_n 0.00879805f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_324 N_A_225_47#_c_354_n N_A_589_47#_c_572_n 0.03957f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_325 N_A_225_47#_c_357_n N_A_589_47#_c_572_n 0.0031956f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_326 N_A_225_47#_M1012_g N_A_589_47#_c_573_n 0.00243606f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_327 N_A_225_47#_M1014_g N_A_589_47#_c_573_n 0.00113891f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_328 N_A_225_47#_c_351_n N_A_589_47#_c_573_n 0.00808484f $X=2.575 $Y=0.82
+ $X2=0 $Y2=0
cc_329 N_A_225_47#_c_354_n N_A_589_47#_c_573_n 0.030582f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_330 N_A_225_47#_c_357_n N_A_589_47#_c_573_n 0.00331919f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_331 N_A_225_47#_c_359_n N_A_589_47#_c_599_n 0.0137916f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_332 N_A_225_47#_c_360_n N_A_589_47#_c_599_n 0.0101048f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_333 N_A_225_47#_c_354_n N_A_589_47#_c_599_n 0.0394547f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_334 N_A_225_47#_c_357_n N_A_589_47#_c_599_n 0.00720931f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_335 N_A_225_47#_c_358_n N_A_589_47#_c_600_n 0.00386185f $X=2.895 $Y=1.41
+ $X2=0 $Y2=0
cc_336 N_A_225_47#_c_359_n N_A_589_47#_c_600_n 0.00107777f $X=3.365 $Y=1.41
+ $X2=0 $Y2=0
cc_337 N_A_225_47#_c_367_n N_A_589_47#_c_600_n 0.0149281f $X=2.575 $Y=1.53 $X2=0
+ $Y2=0
cc_338 N_A_225_47#_c_354_n N_A_589_47#_c_600_n 0.0305808f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_339 N_A_225_47#_c_357_n N_A_589_47#_c_600_n 0.0074788f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_340 N_A_225_47#_M1014_g N_A_589_47#_c_636_n 5.25882e-19 $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_341 N_A_225_47#_M1023_g N_A_589_47#_c_636_n 0.00657592f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_342 N_A_225_47#_M1033_g N_A_589_47#_c_636_n 0.00693104f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_343 N_A_225_47#_M1045_g N_A_589_47#_c_636_n 5.47131e-19 $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_344 N_A_225_47#_c_359_n N_A_589_47#_c_640_n 8.07084e-19 $X=3.365 $Y=1.41
+ $X2=0 $Y2=0
cc_345 N_A_225_47#_c_360_n N_A_589_47#_c_640_n 0.0141618f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_346 N_A_225_47#_c_361_n N_A_589_47#_c_640_n 0.0115459f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_347 N_A_225_47#_c_362_n N_A_589_47#_c_640_n 7.68612e-19 $X=4.775 $Y=1.41
+ $X2=0 $Y2=0
cc_348 N_A_225_47#_M1033_g N_A_589_47#_c_574_n 0.00879805f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_349 N_A_225_47#_M1045_g N_A_589_47#_c_574_n 0.00879805f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_350 N_A_225_47#_c_354_n N_A_589_47#_c_574_n 0.03957f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_351 N_A_225_47#_c_357_n N_A_589_47#_c_574_n 0.0031956f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_352 N_A_225_47#_c_361_n N_A_589_47#_c_601_n 0.0137916f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_353 N_A_225_47#_c_362_n N_A_589_47#_c_601_n 0.0101048f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_354 N_A_225_47#_c_354_n N_A_589_47#_c_601_n 0.0394547f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_355 N_A_225_47#_c_357_n N_A_589_47#_c_601_n 0.00720931f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_356 N_A_225_47#_M1033_g N_A_589_47#_c_652_n 5.25882e-19 $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_357 N_A_225_47#_M1045_g N_A_589_47#_c_652_n 0.00657592f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_358 N_A_225_47#_c_361_n N_A_589_47#_c_654_n 8.07084e-19 $X=4.305 $Y=1.41
+ $X2=0 $Y2=0
cc_359 N_A_225_47#_c_362_n N_A_589_47#_c_654_n 0.0141618f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_360 N_A_225_47#_c_363_n N_A_589_47#_c_654_n 0.0115459f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_361 N_A_225_47#_M1047_g N_A_589_47#_c_575_n 0.0116573f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_362 N_A_225_47#_c_363_n N_A_589_47#_c_602_n 0.0151183f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_363 N_A_225_47#_c_357_n N_A_589_47#_c_602_n 3.58038e-19 $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_364 N_A_225_47#_M1047_g N_A_589_47#_c_576_n 0.00415408f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_365 N_A_225_47#_c_363_n N_A_589_47#_c_577_n 8.26658e-19 $X=5.245 $Y=1.41
+ $X2=0 $Y2=0
cc_366 N_A_225_47#_c_357_n N_A_589_47#_c_577_n 0.00331109f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_367 N_A_225_47#_M1023_g N_A_589_47#_c_579_n 0.00113891f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_368 N_A_225_47#_M1033_g N_A_589_47#_c_579_n 0.00113891f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_369 N_A_225_47#_c_354_n N_A_589_47#_c_579_n 0.030582f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_370 N_A_225_47#_c_357_n N_A_589_47#_c_579_n 0.00331919f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_371 N_A_225_47#_c_360_n N_A_589_47#_c_604_n 0.00260297f $X=3.835 $Y=1.41
+ $X2=0 $Y2=0
cc_372 N_A_225_47#_c_361_n N_A_589_47#_c_604_n 0.00107777f $X=4.305 $Y=1.41
+ $X2=0 $Y2=0
cc_373 N_A_225_47#_c_354_n N_A_589_47#_c_604_n 0.0305808f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_374 N_A_225_47#_c_357_n N_A_589_47#_c_604_n 0.0074788f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_375 N_A_225_47#_M1045_g N_A_589_47#_c_580_n 0.0011682f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_376 N_A_225_47#_c_354_n N_A_589_47#_c_580_n 0.0274674f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_377 N_A_225_47#_c_357_n N_A_589_47#_c_580_n 0.00450461f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_378 N_A_225_47#_c_362_n N_A_589_47#_c_605_n 0.00259297f $X=4.775 $Y=1.41
+ $X2=0 $Y2=0
cc_379 N_A_225_47#_c_363_n N_A_589_47#_c_605_n 0.00128868f $X=5.245 $Y=1.41
+ $X2=0 $Y2=0
cc_380 N_A_225_47#_c_354_n N_A_589_47#_c_605_n 0.0274092f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_381 N_A_225_47#_c_357_n N_A_589_47#_c_605_n 0.00735453f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_382 N_A_225_47#_c_354_n N_A_589_47#_c_581_n 0.0130035f $X=4.9 $Y=1.16 $X2=0
+ $Y2=0
cc_383 N_A_225_47#_c_357_n N_A_589_47#_c_581_n 0.00237077f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_384 N_A_225_47#_c_357_n N_A_589_47#_c_582_n 0.0207158f $X=5.245 $Y=1.217
+ $X2=0 $Y2=0
cc_385 N_A_225_47#_c_365_n N_VPWR_M1027_d 0.00178587f $X=1.975 $Y=1.53 $X2=0
+ $Y2=0
cc_386 N_A_225_47#_c_367_n N_VPWR_M1042_d 0.00324655f $X=2.575 $Y=1.53 $X2=0
+ $Y2=0
cc_387 N_A_225_47#_c_364_n N_VPWR_c_1021_n 0.0411685f $X=1.25 $Y=1.63 $X2=0
+ $Y2=0
cc_388 N_A_225_47#_c_365_n N_VPWR_c_1021_n 0.0136682f $X=1.975 $Y=1.53 $X2=0
+ $Y2=0
cc_389 N_A_225_47#_c_398_n N_VPWR_c_1021_n 0.0507655f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_390 N_A_225_47#_c_358_n N_VPWR_c_1022_n 0.00497803f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_391 N_A_225_47#_c_398_n N_VPWR_c_1022_n 0.0416217f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_392 N_A_225_47#_c_367_n N_VPWR_c_1022_n 0.0151472f $X=2.575 $Y=1.53 $X2=0
+ $Y2=0
cc_393 N_A_225_47#_c_359_n N_VPWR_c_1023_n 0.0052072f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_394 N_A_225_47#_c_360_n N_VPWR_c_1023_n 0.004751f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_395 N_A_225_47#_c_361_n N_VPWR_c_1024_n 0.0052072f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_396 N_A_225_47#_c_362_n N_VPWR_c_1024_n 0.004751f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_397 N_A_225_47#_c_363_n N_VPWR_c_1025_n 0.0052072f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_398 N_A_225_47#_c_364_n N_VPWR_c_1035_n 0.0210596f $X=1.25 $Y=1.63 $X2=0
+ $Y2=0
cc_399 N_A_225_47#_c_398_n N_VPWR_c_1037_n 0.0223557f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_400 N_A_225_47#_c_358_n N_VPWR_c_1039_n 0.00597712f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_401 N_A_225_47#_c_359_n N_VPWR_c_1039_n 0.00673617f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_402 N_A_225_47#_c_360_n N_VPWR_c_1041_n 0.00597712f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_403 N_A_225_47#_c_361_n N_VPWR_c_1041_n 0.00673617f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_404 N_A_225_47#_c_362_n N_VPWR_c_1043_n 0.00597712f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_405 N_A_225_47#_c_363_n N_VPWR_c_1043_n 0.00673617f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_406 N_A_225_47#_M1027_s N_VPWR_c_1018_n 0.00217517f $X=1.125 $Y=1.485 $X2=0
+ $Y2=0
cc_407 N_A_225_47#_M1035_s N_VPWR_c_1018_n 0.00231261f $X=2.045 $Y=1.485 $X2=0
+ $Y2=0
cc_408 N_A_225_47#_c_358_n N_VPWR_c_1018_n 0.0100198f $X=2.895 $Y=1.41 $X2=0
+ $Y2=0
cc_409 N_A_225_47#_c_359_n N_VPWR_c_1018_n 0.0118438f $X=3.365 $Y=1.41 $X2=0
+ $Y2=0
cc_410 N_A_225_47#_c_360_n N_VPWR_c_1018_n 0.00999457f $X=3.835 $Y=1.41 $X2=0
+ $Y2=0
cc_411 N_A_225_47#_c_361_n N_VPWR_c_1018_n 0.0118438f $X=4.305 $Y=1.41 $X2=0
+ $Y2=0
cc_412 N_A_225_47#_c_362_n N_VPWR_c_1018_n 0.00999457f $X=4.775 $Y=1.41 $X2=0
+ $Y2=0
cc_413 N_A_225_47#_c_363_n N_VPWR_c_1018_n 0.011869f $X=5.245 $Y=1.41 $X2=0
+ $Y2=0
cc_414 N_A_225_47#_c_364_n N_VPWR_c_1018_n 0.0124725f $X=1.25 $Y=1.63 $X2=0
+ $Y2=0
cc_415 N_A_225_47#_c_398_n N_VPWR_c_1018_n 0.0140101f $X=2.19 $Y=1.63 $X2=0
+ $Y2=0
cc_416 N_A_225_47#_M1047_g N_X_c_1270_n 4.77587e-19 $X=5.27 $Y=0.56 $X2=0 $Y2=0
cc_417 N_A_225_47#_c_363_n N_X_c_1271_n 8.07084e-19 $X=5.245 $Y=1.41 $X2=0 $Y2=0
cc_418 N_A_225_47#_c_349_n N_VGND_M1020_d 0.00251598f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_419 N_A_225_47#_c_351_n N_VGND_M1050_d 0.00193551f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_420 N_A_225_47#_c_348_n N_VGND_c_1600_n 0.0184656f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_421 N_A_225_47#_c_349_n N_VGND_c_1600_n 0.0127122f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_422 N_A_225_47#_M1012_g N_VGND_c_1601_n 0.00268723f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_423 N_A_225_47#_c_351_n N_VGND_c_1601_n 0.0135251f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_424 N_A_225_47#_M1014_g N_VGND_c_1602_n 0.00390178f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_425 N_A_225_47#_M1023_g N_VGND_c_1602_n 0.00276126f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_426 N_A_225_47#_M1033_g N_VGND_c_1603_n 0.00390178f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_427 N_A_225_47#_M1045_g N_VGND_c_1603_n 0.00276126f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_428 N_A_225_47#_M1047_g N_VGND_c_1604_n 0.00268723f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_429 N_A_225_47#_c_348_n N_VGND_c_1614_n 0.020318f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_430 N_A_225_47#_c_349_n N_VGND_c_1614_n 0.00260082f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_431 N_A_225_47#_c_349_n N_VGND_c_1616_n 0.00193763f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_432 N_A_225_47#_c_396_n N_VGND_c_1616_n 0.022456f $X=2.19 $Y=0.4 $X2=0 $Y2=0
cc_433 N_A_225_47#_c_351_n N_VGND_c_1616_n 0.00248202f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_434 N_A_225_47#_M1012_g N_VGND_c_1618_n 0.00541562f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_435 N_A_225_47#_M1014_g N_VGND_c_1618_n 0.00424619f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_436 N_A_225_47#_M1023_g N_VGND_c_1620_n 0.00424619f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_437 N_A_225_47#_M1033_g N_VGND_c_1620_n 0.00424619f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_438 N_A_225_47#_M1045_g N_VGND_c_1622_n 0.00424619f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_439 N_A_225_47#_M1047_g N_VGND_c_1622_n 0.00439206f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_440 N_A_225_47#_M1020_s N_VGND_c_1639_n 0.0020946f $X=1.125 $Y=0.235 $X2=0
+ $Y2=0
cc_441 N_A_225_47#_M1038_s N_VGND_c_1639_n 0.00304616f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_442 N_A_225_47#_M1012_g N_VGND_c_1639_n 0.00965588f $X=2.87 $Y=0.56 $X2=0
+ $Y2=0
cc_443 N_A_225_47#_M1014_g N_VGND_c_1639_n 0.00611295f $X=3.34 $Y=0.56 $X2=0
+ $Y2=0
cc_444 N_A_225_47#_M1023_g N_VGND_c_1639_n 0.00599018f $X=3.81 $Y=0.56 $X2=0
+ $Y2=0
cc_445 N_A_225_47#_M1033_g N_VGND_c_1639_n 0.00611295f $X=4.28 $Y=0.56 $X2=0
+ $Y2=0
cc_446 N_A_225_47#_M1045_g N_VGND_c_1639_n 0.00610552f $X=4.75 $Y=0.56 $X2=0
+ $Y2=0
cc_447 N_A_225_47#_M1047_g N_VGND_c_1639_n 0.00618081f $X=5.27 $Y=0.56 $X2=0
+ $Y2=0
cc_448 N_A_225_47#_c_348_n N_VGND_c_1639_n 0.0123792f $X=1.25 $Y=0.4 $X2=0 $Y2=0
cc_449 N_A_225_47#_c_349_n N_VGND_c_1639_n 0.00961016f $X=1.975 $Y=0.82 $X2=0
+ $Y2=0
cc_450 N_A_225_47#_c_396_n N_VGND_c_1639_n 0.0142976f $X=2.19 $Y=0.4 $X2=0 $Y2=0
cc_451 N_A_225_47#_c_351_n N_VGND_c_1639_n 0.00561929f $X=2.575 $Y=0.82 $X2=0
+ $Y2=0
cc_452 N_A_589_47#_c_599_n N_VPWR_M1008_d 0.00199888f $X=3.855 $Y=1.53 $X2=0
+ $Y2=0
cc_453 N_A_589_47#_c_601_n N_VPWR_M1031_d 0.00199888f $X=4.795 $Y=1.53 $X2=0
+ $Y2=0
cc_454 N_A_589_47#_c_602_n N_VPWR_M1049_d 0.00347056f $X=5.39 $Y=1.53 $X2=0
+ $Y2=0
cc_455 N_A_589_47#_c_608_n N_VPWR_c_1022_n 0.0507655f $X=3.13 $Y=1.63 $X2=0
+ $Y2=0
cc_456 N_A_589_47#_c_608_n N_VPWR_c_1023_n 0.0385613f $X=3.13 $Y=1.63 $X2=0
+ $Y2=0
cc_457 N_A_589_47#_c_599_n N_VPWR_c_1023_n 0.0112848f $X=3.855 $Y=1.53 $X2=0
+ $Y2=0
cc_458 N_A_589_47#_c_640_n N_VPWR_c_1023_n 0.0470327f $X=4.07 $Y=1.63 $X2=0
+ $Y2=0
cc_459 N_A_589_47#_c_640_n N_VPWR_c_1024_n 0.0385613f $X=4.07 $Y=1.63 $X2=0
+ $Y2=0
cc_460 N_A_589_47#_c_601_n N_VPWR_c_1024_n 0.0112848f $X=4.795 $Y=1.53 $X2=0
+ $Y2=0
cc_461 N_A_589_47#_c_654_n N_VPWR_c_1024_n 0.0470327f $X=5.01 $Y=1.63 $X2=0
+ $Y2=0
cc_462 N_A_589_47#_c_583_n N_VPWR_c_1025_n 0.004751f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_463 N_A_589_47#_c_654_n N_VPWR_c_1025_n 0.0385613f $X=5.01 $Y=1.63 $X2=0
+ $Y2=0
cc_464 N_A_589_47#_c_602_n N_VPWR_c_1025_n 0.0124926f $X=5.39 $Y=1.53 $X2=0
+ $Y2=0
cc_465 N_A_589_47#_c_584_n N_VPWR_c_1026_n 0.0052072f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_466 N_A_589_47#_c_585_n N_VPWR_c_1026_n 0.004751f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_467 N_A_589_47#_c_586_n N_VPWR_c_1027_n 0.0052072f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_468 N_A_589_47#_c_587_n N_VPWR_c_1027_n 0.004751f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_469 N_A_589_47#_c_588_n N_VPWR_c_1028_n 0.0052072f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_470 N_A_589_47#_c_589_n N_VPWR_c_1028_n 0.004751f $X=8.535 $Y=1.41 $X2=0
+ $Y2=0
cc_471 N_A_589_47#_c_590_n N_VPWR_c_1029_n 0.0052072f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_472 N_A_589_47#_c_591_n N_VPWR_c_1029_n 0.004751f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_473 N_A_589_47#_c_592_n N_VPWR_c_1030_n 0.0052072f $X=9.945 $Y=1.41 $X2=0
+ $Y2=0
cc_474 N_A_589_47#_c_593_n N_VPWR_c_1030_n 0.004751f $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_475 N_A_589_47#_c_594_n N_VPWR_c_1031_n 0.0052072f $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_476 N_A_589_47#_c_595_n N_VPWR_c_1031_n 0.004751f $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_477 N_A_589_47#_c_596_n N_VPWR_c_1032_n 0.0052072f $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_478 N_A_589_47#_c_597_n N_VPWR_c_1032_n 0.004751f $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_479 N_A_589_47#_c_598_n N_VPWR_c_1034_n 0.00688901f $X=12.765 $Y=1.41 $X2=0
+ $Y2=0
cc_480 N_A_589_47#_c_608_n N_VPWR_c_1039_n 0.0223557f $X=3.13 $Y=1.63 $X2=0
+ $Y2=0
cc_481 N_A_589_47#_c_640_n N_VPWR_c_1041_n 0.0223557f $X=4.07 $Y=1.63 $X2=0
+ $Y2=0
cc_482 N_A_589_47#_c_654_n N_VPWR_c_1043_n 0.0223557f $X=5.01 $Y=1.63 $X2=0
+ $Y2=0
cc_483 N_A_589_47#_c_583_n N_VPWR_c_1045_n 0.00597712f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_484 N_A_589_47#_c_584_n N_VPWR_c_1045_n 0.00673617f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_485 N_A_589_47#_c_585_n N_VPWR_c_1047_n 0.00597712f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_486 N_A_589_47#_c_586_n N_VPWR_c_1047_n 0.00673617f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_487 N_A_589_47#_c_587_n N_VPWR_c_1049_n 0.00597712f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_488 N_A_589_47#_c_588_n N_VPWR_c_1049_n 0.00673617f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_489 N_A_589_47#_c_589_n N_VPWR_c_1051_n 0.00597712f $X=8.535 $Y=1.41 $X2=0
+ $Y2=0
cc_490 N_A_589_47#_c_590_n N_VPWR_c_1051_n 0.00673617f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_491 N_A_589_47#_c_591_n N_VPWR_c_1053_n 0.00597712f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_492 N_A_589_47#_c_592_n N_VPWR_c_1053_n 0.00673617f $X=9.945 $Y=1.41 $X2=0
+ $Y2=0
cc_493 N_A_589_47#_c_593_n N_VPWR_c_1055_n 0.00597712f $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_494 N_A_589_47#_c_594_n N_VPWR_c_1055_n 0.00673617f $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_495 N_A_589_47#_c_595_n N_VPWR_c_1057_n 0.00597712f $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_496 N_A_589_47#_c_596_n N_VPWR_c_1057_n 0.00673617f $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_497 N_A_589_47#_c_597_n N_VPWR_c_1059_n 0.00597712f $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_498 N_A_589_47#_c_598_n N_VPWR_c_1059_n 0.00673617f $X=12.765 $Y=1.41 $X2=0
+ $Y2=0
cc_499 N_A_589_47#_M1005_s N_VPWR_c_1018_n 0.00231261f $X=2.985 $Y=1.485 $X2=0
+ $Y2=0
cc_500 N_A_589_47#_M1010_s N_VPWR_c_1018_n 0.00231261f $X=3.925 $Y=1.485 $X2=0
+ $Y2=0
cc_501 N_A_589_47#_M1039_s N_VPWR_c_1018_n 0.00231261f $X=4.865 $Y=1.485 $X2=0
+ $Y2=0
cc_502 N_A_589_47#_c_583_n N_VPWR_c_1018_n 0.0100198f $X=5.715 $Y=1.41 $X2=0
+ $Y2=0
cc_503 N_A_589_47#_c_584_n N_VPWR_c_1018_n 0.0118438f $X=6.185 $Y=1.41 $X2=0
+ $Y2=0
cc_504 N_A_589_47#_c_585_n N_VPWR_c_1018_n 0.00999457f $X=6.655 $Y=1.41 $X2=0
+ $Y2=0
cc_505 N_A_589_47#_c_586_n N_VPWR_c_1018_n 0.0118438f $X=7.125 $Y=1.41 $X2=0
+ $Y2=0
cc_506 N_A_589_47#_c_587_n N_VPWR_c_1018_n 0.00999457f $X=7.595 $Y=1.41 $X2=0
+ $Y2=0
cc_507 N_A_589_47#_c_588_n N_VPWR_c_1018_n 0.0118438f $X=8.065 $Y=1.41 $X2=0
+ $Y2=0
cc_508 N_A_589_47#_c_589_n N_VPWR_c_1018_n 0.00999457f $X=8.535 $Y=1.41 $X2=0
+ $Y2=0
cc_509 N_A_589_47#_c_590_n N_VPWR_c_1018_n 0.0118438f $X=9.005 $Y=1.41 $X2=0
+ $Y2=0
cc_510 N_A_589_47#_c_591_n N_VPWR_c_1018_n 0.00999457f $X=9.475 $Y=1.41 $X2=0
+ $Y2=0
cc_511 N_A_589_47#_c_592_n N_VPWR_c_1018_n 0.0118438f $X=9.945 $Y=1.41 $X2=0
+ $Y2=0
cc_512 N_A_589_47#_c_593_n N_VPWR_c_1018_n 0.00999457f $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_513 N_A_589_47#_c_594_n N_VPWR_c_1018_n 0.0118438f $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_514 N_A_589_47#_c_595_n N_VPWR_c_1018_n 0.00999457f $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_515 N_A_589_47#_c_596_n N_VPWR_c_1018_n 0.0118438f $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_516 N_A_589_47#_c_597_n N_VPWR_c_1018_n 0.00999457f $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_517 N_A_589_47#_c_598_n N_VPWR_c_1018_n 0.0128216f $X=12.765 $Y=1.41 $X2=0
+ $Y2=0
cc_518 N_A_589_47#_c_608_n N_VPWR_c_1018_n 0.0140101f $X=3.13 $Y=1.63 $X2=0
+ $Y2=0
cc_519 N_A_589_47#_c_640_n N_VPWR_c_1018_n 0.0140101f $X=4.07 $Y=1.63 $X2=0
+ $Y2=0
cc_520 N_A_589_47#_c_654_n N_VPWR_c_1018_n 0.0140101f $X=5.01 $Y=1.63 $X2=0
+ $Y2=0
cc_521 N_A_589_47#_M1001_g N_X_c_1272_n 0.00229101f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_522 N_A_589_47#_M1002_g N_X_c_1272_n 0.00248233f $X=6.16 $Y=0.56 $X2=0 $Y2=0
cc_523 N_A_589_47#_M1001_g N_X_c_1270_n 0.00426764f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_524 N_A_589_47#_M1002_g N_X_c_1270_n 0.00445433f $X=6.16 $Y=0.56 $X2=0 $Y2=0
cc_525 N_A_589_47#_M1003_g N_X_c_1270_n 4.84753e-19 $X=6.63 $Y=0.56 $X2=0 $Y2=0
cc_526 N_A_589_47#_c_583_n N_X_c_1271_n 0.0141618f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_527 N_A_589_47#_c_584_n N_X_c_1271_n 0.0115459f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_528 N_A_589_47#_c_585_n N_X_c_1271_n 7.68612e-19 $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_529 N_A_589_47#_c_654_n N_X_c_1271_n 0.00629866f $X=5.01 $Y=1.63 $X2=0 $Y2=0
cc_530 N_A_589_47#_M1002_g N_X_c_1235_n 0.00879805f $X=6.16 $Y=0.56 $X2=0 $Y2=0
cc_531 N_A_589_47#_M1003_g N_X_c_1235_n 0.00879805f $X=6.63 $Y=0.56 $X2=0 $Y2=0
cc_532 N_A_589_47#_c_578_n N_X_c_1235_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_533 N_A_589_47#_c_582_n N_X_c_1235_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_534 N_A_589_47#_M1001_g N_X_c_1236_n 0.00245067f $X=5.69 $Y=0.56 $X2=0 $Y2=0
cc_535 N_A_589_47#_M1002_g N_X_c_1236_n 0.00115337f $X=6.16 $Y=0.56 $X2=0 $Y2=0
cc_536 N_A_589_47#_c_575_n N_X_c_1236_n 0.00808484f $X=5.39 $Y=0.82 $X2=0 $Y2=0
cc_537 N_A_589_47#_c_578_n N_X_c_1236_n 0.0305973f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_538 N_A_589_47#_c_582_n N_X_c_1236_n 0.00332f $X=12.765 $Y=1.217 $X2=0 $Y2=0
cc_539 N_A_589_47#_c_584_n N_X_c_1252_n 0.0137916f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_540 N_A_589_47#_c_585_n N_X_c_1252_n 0.0101048f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_541 N_A_589_47#_c_578_n N_X_c_1252_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_542 N_A_589_47#_c_582_n N_X_c_1252_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_543 N_A_589_47#_c_583_n N_X_c_1253_n 0.00386185f $X=5.715 $Y=1.41 $X2=0 $Y2=0
cc_544 N_A_589_47#_c_584_n N_X_c_1253_n 0.00107777f $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_545 N_A_589_47#_c_602_n N_X_c_1253_n 0.0149281f $X=5.39 $Y=1.53 $X2=0 $Y2=0
cc_546 N_A_589_47#_c_578_n N_X_c_1253_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_547 N_A_589_47#_c_582_n N_X_c_1253_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_548 N_A_589_47#_M1003_g N_X_c_1299_n 0.00226116f $X=6.63 $Y=0.56 $X2=0 $Y2=0
cc_549 N_A_589_47#_M1006_g N_X_c_1299_n 0.00248233f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_550 N_A_589_47#_M1002_g N_X_c_1301_n 4.7681e-19 $X=6.16 $Y=0.56 $X2=0 $Y2=0
cc_551 N_A_589_47#_M1003_g N_X_c_1301_n 0.0043216f $X=6.63 $Y=0.56 $X2=0 $Y2=0
cc_552 N_A_589_47#_M1006_g N_X_c_1301_n 0.00445433f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_553 N_A_589_47#_M1007_g N_X_c_1301_n 4.84753e-19 $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_554 N_A_589_47#_c_584_n N_X_c_1305_n 8.07084e-19 $X=6.185 $Y=1.41 $X2=0 $Y2=0
cc_555 N_A_589_47#_c_585_n N_X_c_1305_n 0.0141618f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_556 N_A_589_47#_c_586_n N_X_c_1305_n 0.0115459f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_557 N_A_589_47#_c_587_n N_X_c_1305_n 7.68612e-19 $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_558 N_A_589_47#_M1006_g N_X_c_1237_n 0.00879805f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_559 N_A_589_47#_M1007_g N_X_c_1237_n 0.00879805f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_560 N_A_589_47#_c_578_n N_X_c_1237_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_561 N_A_589_47#_c_582_n N_X_c_1237_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_562 N_A_589_47#_c_586_n N_X_c_1254_n 0.0137916f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_563 N_A_589_47#_c_587_n N_X_c_1254_n 0.0101048f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_564 N_A_589_47#_c_578_n N_X_c_1254_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_565 N_A_589_47#_c_582_n N_X_c_1254_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_566 N_A_589_47#_M1007_g N_X_c_1317_n 0.00226116f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_567 N_A_589_47#_M1015_g N_X_c_1317_n 0.00248233f $X=8.04 $Y=0.56 $X2=0 $Y2=0
cc_568 N_A_589_47#_M1006_g N_X_c_1319_n 4.7681e-19 $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_569 N_A_589_47#_M1007_g N_X_c_1319_n 0.0043216f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_570 N_A_589_47#_M1015_g N_X_c_1319_n 0.00445433f $X=8.04 $Y=0.56 $X2=0 $Y2=0
cc_571 N_A_589_47#_M1017_g N_X_c_1319_n 4.84753e-19 $X=8.51 $Y=0.56 $X2=0 $Y2=0
cc_572 N_A_589_47#_c_586_n N_X_c_1323_n 8.07084e-19 $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_573 N_A_589_47#_c_587_n N_X_c_1323_n 0.0141618f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_574 N_A_589_47#_c_588_n N_X_c_1323_n 0.0115459f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_575 N_A_589_47#_c_589_n N_X_c_1323_n 7.68612e-19 $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_576 N_A_589_47#_M1015_g N_X_c_1238_n 0.00879805f $X=8.04 $Y=0.56 $X2=0 $Y2=0
cc_577 N_A_589_47#_M1017_g N_X_c_1238_n 0.00879805f $X=8.51 $Y=0.56 $X2=0 $Y2=0
cc_578 N_A_589_47#_c_578_n N_X_c_1238_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_579 N_A_589_47#_c_582_n N_X_c_1238_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_580 N_A_589_47#_c_588_n N_X_c_1255_n 0.0137916f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_581 N_A_589_47#_c_589_n N_X_c_1255_n 0.0101048f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_582 N_A_589_47#_c_578_n N_X_c_1255_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_583 N_A_589_47#_c_582_n N_X_c_1255_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_584 N_A_589_47#_M1015_g N_X_c_1335_n 5.25882e-19 $X=8.04 $Y=0.56 $X2=0 $Y2=0
cc_585 N_A_589_47#_M1017_g N_X_c_1335_n 0.00657592f $X=8.51 $Y=0.56 $X2=0 $Y2=0
cc_586 N_A_589_47#_M1018_g N_X_c_1335_n 0.00693104f $X=8.98 $Y=0.56 $X2=0 $Y2=0
cc_587 N_A_589_47#_M1021_g N_X_c_1335_n 5.47131e-19 $X=9.45 $Y=0.56 $X2=0 $Y2=0
cc_588 N_A_589_47#_c_588_n N_X_c_1339_n 8.07084e-19 $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_589 N_A_589_47#_c_589_n N_X_c_1339_n 0.0141618f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_590 N_A_589_47#_c_590_n N_X_c_1339_n 0.0115459f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_591 N_A_589_47#_c_591_n N_X_c_1339_n 7.68612e-19 $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_592 N_A_589_47#_M1018_g N_X_c_1239_n 0.00879805f $X=8.98 $Y=0.56 $X2=0 $Y2=0
cc_593 N_A_589_47#_M1021_g N_X_c_1239_n 0.00879805f $X=9.45 $Y=0.56 $X2=0 $Y2=0
cc_594 N_A_589_47#_c_578_n N_X_c_1239_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_595 N_A_589_47#_c_582_n N_X_c_1239_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_596 N_A_589_47#_c_590_n N_X_c_1256_n 0.0137916f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_597 N_A_589_47#_c_591_n N_X_c_1256_n 0.0101048f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_598 N_A_589_47#_c_578_n N_X_c_1256_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_599 N_A_589_47#_c_582_n N_X_c_1256_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_600 N_A_589_47#_M1018_g N_X_c_1351_n 5.25882e-19 $X=8.98 $Y=0.56 $X2=0 $Y2=0
cc_601 N_A_589_47#_M1021_g N_X_c_1351_n 0.00657592f $X=9.45 $Y=0.56 $X2=0 $Y2=0
cc_602 N_A_589_47#_M1024_g N_X_c_1351_n 0.00693104f $X=9.92 $Y=0.56 $X2=0 $Y2=0
cc_603 N_A_589_47#_M1026_g N_X_c_1351_n 5.47131e-19 $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_604 N_A_589_47#_c_590_n N_X_c_1355_n 8.07084e-19 $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_605 N_A_589_47#_c_591_n N_X_c_1355_n 0.0141618f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_606 N_A_589_47#_c_592_n N_X_c_1355_n 0.0115459f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_607 N_A_589_47#_c_593_n N_X_c_1355_n 7.68612e-19 $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_608 N_A_589_47#_M1024_g N_X_c_1240_n 0.00879805f $X=9.92 $Y=0.56 $X2=0 $Y2=0
cc_609 N_A_589_47#_M1026_g N_X_c_1240_n 0.00879805f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_610 N_A_589_47#_c_578_n N_X_c_1240_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_611 N_A_589_47#_c_582_n N_X_c_1240_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_612 N_A_589_47#_c_592_n N_X_c_1257_n 0.0137916f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_613 N_A_589_47#_c_593_n N_X_c_1257_n 0.0101048f $X=10.415 $Y=1.41 $X2=0 $Y2=0
cc_614 N_A_589_47#_c_578_n N_X_c_1257_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_615 N_A_589_47#_c_582_n N_X_c_1257_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_616 N_A_589_47#_M1024_g N_X_c_1367_n 5.25882e-19 $X=9.92 $Y=0.56 $X2=0 $Y2=0
cc_617 N_A_589_47#_M1026_g N_X_c_1367_n 0.00657592f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_618 N_A_589_47#_M1028_g N_X_c_1367_n 0.00693104f $X=10.86 $Y=0.56 $X2=0 $Y2=0
cc_619 N_A_589_47#_M1034_g N_X_c_1367_n 5.47131e-19 $X=11.33 $Y=0.56 $X2=0 $Y2=0
cc_620 N_A_589_47#_c_592_n N_X_c_1371_n 8.07084e-19 $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_621 N_A_589_47#_c_593_n N_X_c_1371_n 0.0141618f $X=10.415 $Y=1.41 $X2=0 $Y2=0
cc_622 N_A_589_47#_c_594_n N_X_c_1371_n 0.0115459f $X=10.885 $Y=1.41 $X2=0 $Y2=0
cc_623 N_A_589_47#_c_595_n N_X_c_1371_n 7.68612e-19 $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_624 N_A_589_47#_M1028_g N_X_c_1241_n 0.00879805f $X=10.86 $Y=0.56 $X2=0 $Y2=0
cc_625 N_A_589_47#_M1034_g N_X_c_1241_n 0.00879805f $X=11.33 $Y=0.56 $X2=0 $Y2=0
cc_626 N_A_589_47#_c_578_n N_X_c_1241_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_627 N_A_589_47#_c_582_n N_X_c_1241_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_628 N_A_589_47#_c_594_n N_X_c_1258_n 0.0137916f $X=10.885 $Y=1.41 $X2=0 $Y2=0
cc_629 N_A_589_47#_c_595_n N_X_c_1258_n 0.0101048f $X=11.355 $Y=1.41 $X2=0 $Y2=0
cc_630 N_A_589_47#_c_578_n N_X_c_1258_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_631 N_A_589_47#_c_582_n N_X_c_1258_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_632 N_A_589_47#_M1028_g N_X_c_1383_n 5.25882e-19 $X=10.86 $Y=0.56 $X2=0 $Y2=0
cc_633 N_A_589_47#_M1034_g N_X_c_1383_n 0.00657592f $X=11.33 $Y=0.56 $X2=0 $Y2=0
cc_634 N_A_589_47#_M1043_g N_X_c_1383_n 0.00693104f $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_635 N_A_589_47#_M1048_g N_X_c_1383_n 5.47131e-19 $X=12.27 $Y=0.56 $X2=0 $Y2=0
cc_636 N_A_589_47#_c_594_n N_X_c_1387_n 8.07084e-19 $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_637 N_A_589_47#_c_595_n N_X_c_1387_n 0.0141618f $X=11.355 $Y=1.41 $X2=0 $Y2=0
cc_638 N_A_589_47#_c_596_n N_X_c_1387_n 0.0115459f $X=11.825 $Y=1.41 $X2=0 $Y2=0
cc_639 N_A_589_47#_c_597_n N_X_c_1387_n 7.68612e-19 $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_640 N_A_589_47#_M1043_g N_X_c_1242_n 0.00879805f $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_641 N_A_589_47#_M1048_g N_X_c_1242_n 0.00879805f $X=12.27 $Y=0.56 $X2=0 $Y2=0
cc_642 N_A_589_47#_c_578_n N_X_c_1242_n 0.03957f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_643 N_A_589_47#_c_582_n N_X_c_1242_n 0.0031956f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_644 N_A_589_47#_c_596_n N_X_c_1259_n 0.0137916f $X=11.825 $Y=1.41 $X2=0 $Y2=0
cc_645 N_A_589_47#_c_597_n N_X_c_1259_n 0.0101048f $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_646 N_A_589_47#_c_578_n N_X_c_1259_n 0.0394547f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_647 N_A_589_47#_c_582_n N_X_c_1259_n 0.00720931f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_648 N_A_589_47#_M1043_g N_X_c_1399_n 5.25882e-19 $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_649 N_A_589_47#_M1048_g N_X_c_1399_n 0.00657592f $X=12.27 $Y=0.56 $X2=0 $Y2=0
cc_650 N_A_589_47#_c_596_n N_X_c_1401_n 8.07084e-19 $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_651 N_A_589_47#_c_597_n N_X_c_1401_n 0.0141618f $X=12.295 $Y=1.41 $X2=0 $Y2=0
cc_652 N_A_589_47#_c_598_n N_X_c_1401_n 0.017566f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_653 N_A_589_47#_M1051_g N_X_c_1243_n 0.0137044f $X=12.79 $Y=0.56 $X2=0 $Y2=0
cc_654 N_A_589_47#_c_578_n N_X_c_1243_n 3.24343e-19 $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_655 N_A_589_47#_c_598_n N_X_c_1260_n 0.016975f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_656 N_A_589_47#_c_578_n N_X_c_1260_n 3.09302e-19 $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_657 N_A_589_47#_c_582_n N_X_c_1260_n 3.58038e-19 $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_658 N_A_589_47#_M1003_g N_X_c_1244_n 0.00115337f $X=6.63 $Y=0.56 $X2=0 $Y2=0
cc_659 N_A_589_47#_M1006_g N_X_c_1244_n 0.00115337f $X=7.1 $Y=0.56 $X2=0 $Y2=0
cc_660 N_A_589_47#_c_578_n N_X_c_1244_n 0.0305905f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_661 N_A_589_47#_c_582_n N_X_c_1244_n 0.00331994f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_662 N_A_589_47#_c_585_n N_X_c_1261_n 0.00260297f $X=6.655 $Y=1.41 $X2=0 $Y2=0
cc_663 N_A_589_47#_c_586_n N_X_c_1261_n 0.00107777f $X=7.125 $Y=1.41 $X2=0 $Y2=0
cc_664 N_A_589_47#_c_578_n N_X_c_1261_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_665 N_A_589_47#_c_582_n N_X_c_1261_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_666 N_A_589_47#_M1007_g N_X_c_1245_n 0.00115337f $X=7.57 $Y=0.56 $X2=0 $Y2=0
cc_667 N_A_589_47#_M1015_g N_X_c_1245_n 0.00115337f $X=8.04 $Y=0.56 $X2=0 $Y2=0
cc_668 N_A_589_47#_c_578_n N_X_c_1245_n 0.0305905f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_669 N_A_589_47#_c_582_n N_X_c_1245_n 0.00331994f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_670 N_A_589_47#_c_587_n N_X_c_1262_n 0.00260297f $X=7.595 $Y=1.41 $X2=0 $Y2=0
cc_671 N_A_589_47#_c_588_n N_X_c_1262_n 0.00107777f $X=8.065 $Y=1.41 $X2=0 $Y2=0
cc_672 N_A_589_47#_c_578_n N_X_c_1262_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_673 N_A_589_47#_c_582_n N_X_c_1262_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_674 N_A_589_47#_M1017_g N_X_c_1246_n 0.00113891f $X=8.51 $Y=0.56 $X2=0 $Y2=0
cc_675 N_A_589_47#_M1018_g N_X_c_1246_n 0.00113891f $X=8.98 $Y=0.56 $X2=0 $Y2=0
cc_676 N_A_589_47#_c_578_n N_X_c_1246_n 0.030582f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_677 N_A_589_47#_c_582_n N_X_c_1246_n 0.00331919f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_678 N_A_589_47#_c_589_n N_X_c_1263_n 0.00260297f $X=8.535 $Y=1.41 $X2=0 $Y2=0
cc_679 N_A_589_47#_c_590_n N_X_c_1263_n 0.00107777f $X=9.005 $Y=1.41 $X2=0 $Y2=0
cc_680 N_A_589_47#_c_578_n N_X_c_1263_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_681 N_A_589_47#_c_582_n N_X_c_1263_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_682 N_A_589_47#_M1021_g N_X_c_1247_n 0.00113891f $X=9.45 $Y=0.56 $X2=0 $Y2=0
cc_683 N_A_589_47#_M1024_g N_X_c_1247_n 0.00113891f $X=9.92 $Y=0.56 $X2=0 $Y2=0
cc_684 N_A_589_47#_c_578_n N_X_c_1247_n 0.030582f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_685 N_A_589_47#_c_582_n N_X_c_1247_n 0.00331919f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_686 N_A_589_47#_c_591_n N_X_c_1264_n 0.00260297f $X=9.475 $Y=1.41 $X2=0 $Y2=0
cc_687 N_A_589_47#_c_592_n N_X_c_1264_n 0.00107777f $X=9.945 $Y=1.41 $X2=0 $Y2=0
cc_688 N_A_589_47#_c_578_n N_X_c_1264_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_689 N_A_589_47#_c_582_n N_X_c_1264_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_690 N_A_589_47#_M1026_g N_X_c_1248_n 0.00113891f $X=10.39 $Y=0.56 $X2=0 $Y2=0
cc_691 N_A_589_47#_M1028_g N_X_c_1248_n 0.00113891f $X=10.86 $Y=0.56 $X2=0 $Y2=0
cc_692 N_A_589_47#_c_578_n N_X_c_1248_n 0.030582f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_693 N_A_589_47#_c_582_n N_X_c_1248_n 0.00331919f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_694 N_A_589_47#_c_593_n N_X_c_1265_n 0.00260297f $X=10.415 $Y=1.41 $X2=0
+ $Y2=0
cc_695 N_A_589_47#_c_594_n N_X_c_1265_n 0.00107777f $X=10.885 $Y=1.41 $X2=0
+ $Y2=0
cc_696 N_A_589_47#_c_578_n N_X_c_1265_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_697 N_A_589_47#_c_582_n N_X_c_1265_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_698 N_A_589_47#_M1034_g N_X_c_1249_n 0.00113891f $X=11.33 $Y=0.56 $X2=0 $Y2=0
cc_699 N_A_589_47#_M1043_g N_X_c_1249_n 0.00113891f $X=11.8 $Y=0.56 $X2=0 $Y2=0
cc_700 N_A_589_47#_c_578_n N_X_c_1249_n 0.030582f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_701 N_A_589_47#_c_582_n N_X_c_1249_n 0.00331919f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_702 N_A_589_47#_c_595_n N_X_c_1266_n 0.00260297f $X=11.355 $Y=1.41 $X2=0
+ $Y2=0
cc_703 N_A_589_47#_c_596_n N_X_c_1266_n 0.00107777f $X=11.825 $Y=1.41 $X2=0
+ $Y2=0
cc_704 N_A_589_47#_c_578_n N_X_c_1266_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_705 N_A_589_47#_c_582_n N_X_c_1266_n 0.0074788f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_706 N_A_589_47#_M1048_g N_X_c_1250_n 0.0011682f $X=12.27 $Y=0.56 $X2=0 $Y2=0
cc_707 N_A_589_47#_c_578_n N_X_c_1250_n 0.0307156f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_708 N_A_589_47#_c_582_n N_X_c_1250_n 0.00450461f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_709 N_A_589_47#_c_597_n N_X_c_1267_n 0.00260297f $X=12.295 $Y=1.41 $X2=0
+ $Y2=0
cc_710 N_A_589_47#_c_598_n N_X_c_1267_n 0.00107777f $X=12.765 $Y=1.41 $X2=0
+ $Y2=0
cc_711 N_A_589_47#_c_578_n N_X_c_1267_n 0.0305808f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_712 N_A_589_47#_c_582_n N_X_c_1267_n 0.00723098f $X=12.765 $Y=1.217 $X2=0
+ $Y2=0
cc_713 N_A_589_47#_c_598_n X 0.00142485f $X=12.765 $Y=1.41 $X2=0 $Y2=0
cc_714 N_A_589_47#_M1051_g X 0.0196725f $X=12.79 $Y=0.56 $X2=0 $Y2=0
cc_715 N_A_589_47#_c_578_n X 0.013577f $X=12.28 $Y=1.16 $X2=0 $Y2=0
cc_716 N_A_589_47#_c_572_n N_VGND_M1014_s 0.00251598f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_717 N_A_589_47#_c_574_n N_VGND_M1033_s 0.00251598f $X=4.795 $Y=0.82 $X2=0
+ $Y2=0
cc_718 N_A_589_47#_c_575_n N_VGND_M1047_s 0.00193551f $X=5.39 $Y=0.82 $X2=0
+ $Y2=0
cc_719 N_A_589_47#_c_607_n N_VGND_c_1602_n 0.0186688f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_720 N_A_589_47#_c_572_n N_VGND_c_1602_n 0.0127122f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_721 N_A_589_47#_c_636_n N_VGND_c_1603_n 0.0186688f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_722 N_A_589_47#_c_574_n N_VGND_c_1603_n 0.0127122f $X=4.795 $Y=0.82 $X2=0
+ $Y2=0
cc_723 N_A_589_47#_M1001_g N_VGND_c_1604_n 0.00268723f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_724 N_A_589_47#_c_575_n N_VGND_c_1604_n 0.0135251f $X=5.39 $Y=0.82 $X2=0
+ $Y2=0
cc_725 N_A_589_47#_M1002_g N_VGND_c_1605_n 0.00382673f $X=6.16 $Y=0.56 $X2=0
+ $Y2=0
cc_726 N_A_589_47#_M1003_g N_VGND_c_1605_n 0.00276126f $X=6.63 $Y=0.56 $X2=0
+ $Y2=0
cc_727 N_A_589_47#_M1006_g N_VGND_c_1606_n 0.00382673f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_728 N_A_589_47#_M1007_g N_VGND_c_1606_n 0.00276126f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_729 N_A_589_47#_M1015_g N_VGND_c_1607_n 0.00382673f $X=8.04 $Y=0.56 $X2=0
+ $Y2=0
cc_730 N_A_589_47#_M1017_g N_VGND_c_1607_n 0.00276126f $X=8.51 $Y=0.56 $X2=0
+ $Y2=0
cc_731 N_A_589_47#_M1018_g N_VGND_c_1608_n 0.00390178f $X=8.98 $Y=0.56 $X2=0
+ $Y2=0
cc_732 N_A_589_47#_M1021_g N_VGND_c_1608_n 0.00276126f $X=9.45 $Y=0.56 $X2=0
+ $Y2=0
cc_733 N_A_589_47#_M1024_g N_VGND_c_1609_n 0.00390178f $X=9.92 $Y=0.56 $X2=0
+ $Y2=0
cc_734 N_A_589_47#_M1026_g N_VGND_c_1609_n 0.00276126f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_735 N_A_589_47#_M1028_g N_VGND_c_1610_n 0.00390178f $X=10.86 $Y=0.56 $X2=0
+ $Y2=0
cc_736 N_A_589_47#_M1034_g N_VGND_c_1610_n 0.00276126f $X=11.33 $Y=0.56 $X2=0
+ $Y2=0
cc_737 N_A_589_47#_M1043_g N_VGND_c_1611_n 0.00390178f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_738 N_A_589_47#_M1048_g N_VGND_c_1611_n 0.00276126f $X=12.27 $Y=0.56 $X2=0
+ $Y2=0
cc_739 N_A_589_47#_M1051_g N_VGND_c_1613_n 0.00438629f $X=12.79 $Y=0.56 $X2=0
+ $Y2=0
cc_740 N_A_589_47#_c_607_n N_VGND_c_1618_n 0.0216617f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_741 N_A_589_47#_c_572_n N_VGND_c_1618_n 0.00260082f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_742 N_A_589_47#_c_572_n N_VGND_c_1620_n 0.00193763f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_743 N_A_589_47#_c_636_n N_VGND_c_1620_n 0.0216617f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_744 N_A_589_47#_c_574_n N_VGND_c_1620_n 0.00260082f $X=4.795 $Y=0.82 $X2=0
+ $Y2=0
cc_745 N_A_589_47#_c_574_n N_VGND_c_1622_n 0.00193763f $X=4.795 $Y=0.82 $X2=0
+ $Y2=0
cc_746 N_A_589_47#_c_652_n N_VGND_c_1622_n 0.022456f $X=5.01 $Y=0.4 $X2=0 $Y2=0
cc_747 N_A_589_47#_c_575_n N_VGND_c_1622_n 0.00245178f $X=5.39 $Y=0.82 $X2=0
+ $Y2=0
cc_748 N_A_589_47#_M1001_g N_VGND_c_1624_n 0.00539841f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_749 N_A_589_47#_M1002_g N_VGND_c_1624_n 0.00423108f $X=6.16 $Y=0.56 $X2=0
+ $Y2=0
cc_750 N_A_589_47#_M1003_g N_VGND_c_1626_n 0.00423108f $X=6.63 $Y=0.56 $X2=0
+ $Y2=0
cc_751 N_A_589_47#_M1006_g N_VGND_c_1626_n 0.00423108f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_752 N_A_589_47#_M1007_g N_VGND_c_1628_n 0.00423108f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_753 N_A_589_47#_M1015_g N_VGND_c_1628_n 0.00423108f $X=8.04 $Y=0.56 $X2=0
+ $Y2=0
cc_754 N_A_589_47#_M1017_g N_VGND_c_1630_n 0.00424619f $X=8.51 $Y=0.56 $X2=0
+ $Y2=0
cc_755 N_A_589_47#_M1018_g N_VGND_c_1630_n 0.00424619f $X=8.98 $Y=0.56 $X2=0
+ $Y2=0
cc_756 N_A_589_47#_M1021_g N_VGND_c_1632_n 0.00424619f $X=9.45 $Y=0.56 $X2=0
+ $Y2=0
cc_757 N_A_589_47#_M1024_g N_VGND_c_1632_n 0.00424619f $X=9.92 $Y=0.56 $X2=0
+ $Y2=0
cc_758 N_A_589_47#_M1026_g N_VGND_c_1634_n 0.00424619f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_759 N_A_589_47#_M1028_g N_VGND_c_1634_n 0.00424619f $X=10.86 $Y=0.56 $X2=0
+ $Y2=0
cc_760 N_A_589_47#_M1034_g N_VGND_c_1636_n 0.00424619f $X=11.33 $Y=0.56 $X2=0
+ $Y2=0
cc_761 N_A_589_47#_M1043_g N_VGND_c_1636_n 0.00424619f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_762 N_A_589_47#_M1048_g N_VGND_c_1638_n 0.00424619f $X=12.27 $Y=0.56 $X2=0
+ $Y2=0
cc_763 N_A_589_47#_M1051_g N_VGND_c_1638_n 0.00439206f $X=12.79 $Y=0.56 $X2=0
+ $Y2=0
cc_764 N_A_589_47#_M1012_d N_VGND_c_1639_n 0.00255524f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_765 N_A_589_47#_M1023_d N_VGND_c_1639_n 0.00255524f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_766 N_A_589_47#_M1045_d N_VGND_c_1639_n 0.00304616f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_767 N_A_589_47#_M1001_g N_VGND_c_1639_n 0.00961873f $X=5.69 $Y=0.56 $X2=0
+ $Y2=0
cc_768 N_A_589_47#_M1002_g N_VGND_c_1639_n 0.00612203f $X=6.16 $Y=0.56 $X2=0
+ $Y2=0
cc_769 N_A_589_47#_M1003_g N_VGND_c_1639_n 0.00599926f $X=6.63 $Y=0.56 $X2=0
+ $Y2=0
cc_770 N_A_589_47#_M1006_g N_VGND_c_1639_n 0.00612203f $X=7.1 $Y=0.56 $X2=0
+ $Y2=0
cc_771 N_A_589_47#_M1007_g N_VGND_c_1639_n 0.00599926f $X=7.57 $Y=0.56 $X2=0
+ $Y2=0
cc_772 N_A_589_47#_M1015_g N_VGND_c_1639_n 0.00612203f $X=8.04 $Y=0.56 $X2=0
+ $Y2=0
cc_773 N_A_589_47#_M1017_g N_VGND_c_1639_n 0.00599018f $X=8.51 $Y=0.56 $X2=0
+ $Y2=0
cc_774 N_A_589_47#_M1018_g N_VGND_c_1639_n 0.00611295f $X=8.98 $Y=0.56 $X2=0
+ $Y2=0
cc_775 N_A_589_47#_M1021_g N_VGND_c_1639_n 0.00599018f $X=9.45 $Y=0.56 $X2=0
+ $Y2=0
cc_776 N_A_589_47#_M1024_g N_VGND_c_1639_n 0.00611295f $X=9.92 $Y=0.56 $X2=0
+ $Y2=0
cc_777 N_A_589_47#_M1026_g N_VGND_c_1639_n 0.00599018f $X=10.39 $Y=0.56 $X2=0
+ $Y2=0
cc_778 N_A_589_47#_M1028_g N_VGND_c_1639_n 0.00611295f $X=10.86 $Y=0.56 $X2=0
+ $Y2=0
cc_779 N_A_589_47#_M1034_g N_VGND_c_1639_n 0.00599018f $X=11.33 $Y=0.56 $X2=0
+ $Y2=0
cc_780 N_A_589_47#_M1043_g N_VGND_c_1639_n 0.00611295f $X=11.8 $Y=0.56 $X2=0
+ $Y2=0
cc_781 N_A_589_47#_M1048_g N_VGND_c_1639_n 0.00610552f $X=12.27 $Y=0.56 $X2=0
+ $Y2=0
cc_782 N_A_589_47#_M1051_g N_VGND_c_1639_n 0.0071762f $X=12.79 $Y=0.56 $X2=0
+ $Y2=0
cc_783 N_A_589_47#_c_607_n N_VGND_c_1639_n 0.0140924f $X=3.13 $Y=0.4 $X2=0 $Y2=0
cc_784 N_A_589_47#_c_572_n N_VGND_c_1639_n 0.00961016f $X=3.855 $Y=0.82 $X2=0
+ $Y2=0
cc_785 N_A_589_47#_c_636_n N_VGND_c_1639_n 0.0140924f $X=4.07 $Y=0.4 $X2=0 $Y2=0
cc_786 N_A_589_47#_c_574_n N_VGND_c_1639_n 0.00961016f $X=4.795 $Y=0.82 $X2=0
+ $Y2=0
cc_787 N_A_589_47#_c_652_n N_VGND_c_1639_n 0.0142976f $X=5.01 $Y=0.4 $X2=0 $Y2=0
cc_788 N_A_589_47#_c_575_n N_VGND_c_1639_n 0.00565014f $X=5.39 $Y=0.82 $X2=0
+ $Y2=0
cc_789 N_VPWR_c_1018_n N_X_M1000_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_790 N_VPWR_c_1018_n N_X_M1009_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_791 N_VPWR_c_1018_n N_X_M1013_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_792 N_VPWR_c_1018_n N_X_M1019_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_793 N_VPWR_c_1018_n N_X_M1029_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_794 N_VPWR_c_1018_n N_X_M1032_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_795 N_VPWR_c_1018_n N_X_M1040_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_796 N_VPWR_c_1018_n N_X_M1044_d 0.00231261f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_797 N_VPWR_c_1025_n N_X_c_1271_n 0.0470327f $X=5.48 $Y=2 $X2=0 $Y2=0
cc_798 N_VPWR_c_1026_n N_X_c_1271_n 0.0385613f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_799 N_VPWR_c_1045_n N_X_c_1271_n 0.0223557f $X=6.335 $Y=2.72 $X2=0 $Y2=0
cc_800 N_VPWR_c_1018_n N_X_c_1271_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_801 N_VPWR_M1004_s N_X_c_1252_n 0.00199888f $X=6.275 $Y=1.485 $X2=0 $Y2=0
cc_802 N_VPWR_c_1026_n N_X_c_1252_n 0.0112848f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_803 N_VPWR_c_1026_n N_X_c_1305_n 0.0470327f $X=6.42 $Y=2 $X2=0 $Y2=0
cc_804 N_VPWR_c_1027_n N_X_c_1305_n 0.0385613f $X=7.36 $Y=2 $X2=0 $Y2=0
cc_805 N_VPWR_c_1047_n N_X_c_1305_n 0.0223557f $X=7.275 $Y=2.72 $X2=0 $Y2=0
cc_806 N_VPWR_c_1018_n N_X_c_1305_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_807 N_VPWR_M1011_s N_X_c_1254_n 0.00199888f $X=7.215 $Y=1.485 $X2=0 $Y2=0
cc_808 N_VPWR_c_1027_n N_X_c_1254_n 0.0112848f $X=7.36 $Y=2 $X2=0 $Y2=0
cc_809 N_VPWR_c_1027_n N_X_c_1323_n 0.0470327f $X=7.36 $Y=2 $X2=0 $Y2=0
cc_810 N_VPWR_c_1028_n N_X_c_1323_n 0.0385613f $X=8.3 $Y=2 $X2=0 $Y2=0
cc_811 N_VPWR_c_1049_n N_X_c_1323_n 0.0223557f $X=8.215 $Y=2.72 $X2=0 $Y2=0
cc_812 N_VPWR_c_1018_n N_X_c_1323_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_813 N_VPWR_M1016_s N_X_c_1255_n 0.00199888f $X=8.155 $Y=1.485 $X2=0 $Y2=0
cc_814 N_VPWR_c_1028_n N_X_c_1255_n 0.0112848f $X=8.3 $Y=2 $X2=0 $Y2=0
cc_815 N_VPWR_c_1028_n N_X_c_1339_n 0.0470327f $X=8.3 $Y=2 $X2=0 $Y2=0
cc_816 N_VPWR_c_1029_n N_X_c_1339_n 0.0385613f $X=9.24 $Y=2 $X2=0 $Y2=0
cc_817 N_VPWR_c_1051_n N_X_c_1339_n 0.0223557f $X=9.155 $Y=2.72 $X2=0 $Y2=0
cc_818 N_VPWR_c_1018_n N_X_c_1339_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_819 N_VPWR_M1025_s N_X_c_1256_n 0.00199888f $X=9.095 $Y=1.485 $X2=0 $Y2=0
cc_820 N_VPWR_c_1029_n N_X_c_1256_n 0.0112848f $X=9.24 $Y=2 $X2=0 $Y2=0
cc_821 N_VPWR_c_1029_n N_X_c_1355_n 0.0470327f $X=9.24 $Y=2 $X2=0 $Y2=0
cc_822 N_VPWR_c_1030_n N_X_c_1355_n 0.0385613f $X=10.18 $Y=2 $X2=0 $Y2=0
cc_823 N_VPWR_c_1053_n N_X_c_1355_n 0.0223557f $X=10.095 $Y=2.72 $X2=0 $Y2=0
cc_824 N_VPWR_c_1018_n N_X_c_1355_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_825 N_VPWR_M1030_s N_X_c_1257_n 0.00199888f $X=10.035 $Y=1.485 $X2=0 $Y2=0
cc_826 N_VPWR_c_1030_n N_X_c_1257_n 0.0112848f $X=10.18 $Y=2 $X2=0 $Y2=0
cc_827 N_VPWR_c_1030_n N_X_c_1371_n 0.0470327f $X=10.18 $Y=2 $X2=0 $Y2=0
cc_828 N_VPWR_c_1031_n N_X_c_1371_n 0.0385613f $X=11.12 $Y=2 $X2=0 $Y2=0
cc_829 N_VPWR_c_1055_n N_X_c_1371_n 0.0223557f $X=11.035 $Y=2.72 $X2=0 $Y2=0
cc_830 N_VPWR_c_1018_n N_X_c_1371_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_831 N_VPWR_M1036_s N_X_c_1258_n 0.00199888f $X=10.975 $Y=1.485 $X2=0 $Y2=0
cc_832 N_VPWR_c_1031_n N_X_c_1258_n 0.0112848f $X=11.12 $Y=2 $X2=0 $Y2=0
cc_833 N_VPWR_c_1031_n N_X_c_1387_n 0.0470327f $X=11.12 $Y=2 $X2=0 $Y2=0
cc_834 N_VPWR_c_1032_n N_X_c_1387_n 0.0385613f $X=12.06 $Y=2 $X2=0 $Y2=0
cc_835 N_VPWR_c_1057_n N_X_c_1387_n 0.0223557f $X=11.975 $Y=2.72 $X2=0 $Y2=0
cc_836 N_VPWR_c_1018_n N_X_c_1387_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_837 N_VPWR_M1041_s N_X_c_1259_n 0.00199888f $X=11.915 $Y=1.485 $X2=0 $Y2=0
cc_838 N_VPWR_c_1032_n N_X_c_1259_n 0.0112848f $X=12.06 $Y=2 $X2=0 $Y2=0
cc_839 N_VPWR_c_1032_n N_X_c_1401_n 0.0470327f $X=12.06 $Y=2 $X2=0 $Y2=0
cc_840 N_VPWR_c_1034_n N_X_c_1401_n 0.0385613f $X=13 $Y=2 $X2=0 $Y2=0
cc_841 N_VPWR_c_1059_n N_X_c_1401_n 0.0223557f $X=12.915 $Y=2.72 $X2=0 $Y2=0
cc_842 N_VPWR_c_1018_n N_X_c_1401_n 0.0140101f $X=13.11 $Y=2.72 $X2=0 $Y2=0
cc_843 N_VPWR_M1046_s N_X_c_1260_n 2.67089e-19 $X=12.855 $Y=1.485 $X2=0 $Y2=0
cc_844 N_VPWR_M1046_s X 0.00453067f $X=12.855 $Y=1.485 $X2=0 $Y2=0
cc_845 N_VPWR_c_1034_n X 0.0121952f $X=13 $Y=2 $X2=0 $Y2=0
cc_846 N_X_c_1235_n N_VGND_M1002_d 0.00251598f $X=6.675 $Y=0.82 $X2=0 $Y2=0
cc_847 N_X_c_1237_n N_VGND_M1006_d 0.00251598f $X=7.615 $Y=0.82 $X2=0 $Y2=0
cc_848 N_X_c_1238_n N_VGND_M1015_d 0.00251598f $X=8.555 $Y=0.82 $X2=0 $Y2=0
cc_849 N_X_c_1239_n N_VGND_M1018_d 0.00251598f $X=9.495 $Y=0.82 $X2=0 $Y2=0
cc_850 N_X_c_1240_n N_VGND_M1024_d 0.00251598f $X=10.435 $Y=0.82 $X2=0 $Y2=0
cc_851 N_X_c_1241_n N_VGND_M1028_d 0.00251598f $X=11.375 $Y=0.82 $X2=0 $Y2=0
cc_852 N_X_c_1242_n N_VGND_M1043_d 0.00251598f $X=12.315 $Y=0.82 $X2=0 $Y2=0
cc_853 N_X_c_1243_n N_VGND_M1051_d 0.00322906f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_854 N_X_c_1272_n N_VGND_c_1605_n 0.0116752f $X=5.925 $Y=0.45 $X2=0 $Y2=0
cc_855 N_X_c_1270_n N_VGND_c_1605_n 0.00700786f $X=5.925 $Y=0.735 $X2=0 $Y2=0
cc_856 N_X_c_1235_n N_VGND_c_1605_n 0.0127122f $X=6.675 $Y=0.82 $X2=0 $Y2=0
cc_857 N_X_c_1299_n N_VGND_c_1606_n 0.0116752f $X=6.865 $Y=0.45 $X2=0 $Y2=0
cc_858 N_X_c_1301_n N_VGND_c_1606_n 0.00700786f $X=6.865 $Y=0.735 $X2=0 $Y2=0
cc_859 N_X_c_1237_n N_VGND_c_1606_n 0.0127122f $X=7.615 $Y=0.82 $X2=0 $Y2=0
cc_860 N_X_c_1317_n N_VGND_c_1607_n 0.0116752f $X=7.805 $Y=0.45 $X2=0 $Y2=0
cc_861 N_X_c_1319_n N_VGND_c_1607_n 0.00700786f $X=7.805 $Y=0.735 $X2=0 $Y2=0
cc_862 N_X_c_1238_n N_VGND_c_1607_n 0.0127122f $X=8.555 $Y=0.82 $X2=0 $Y2=0
cc_863 N_X_c_1335_n N_VGND_c_1608_n 0.0186688f $X=8.77 $Y=0.4 $X2=0 $Y2=0
cc_864 N_X_c_1239_n N_VGND_c_1608_n 0.0127122f $X=9.495 $Y=0.82 $X2=0 $Y2=0
cc_865 N_X_c_1351_n N_VGND_c_1609_n 0.0186688f $X=9.71 $Y=0.4 $X2=0 $Y2=0
cc_866 N_X_c_1240_n N_VGND_c_1609_n 0.0127122f $X=10.435 $Y=0.82 $X2=0 $Y2=0
cc_867 N_X_c_1367_n N_VGND_c_1610_n 0.0186688f $X=10.65 $Y=0.4 $X2=0 $Y2=0
cc_868 N_X_c_1241_n N_VGND_c_1610_n 0.0127122f $X=11.375 $Y=0.82 $X2=0 $Y2=0
cc_869 N_X_c_1383_n N_VGND_c_1611_n 0.0186688f $X=11.59 $Y=0.4 $X2=0 $Y2=0
cc_870 N_X_c_1242_n N_VGND_c_1611_n 0.0127122f $X=12.315 $Y=0.82 $X2=0 $Y2=0
cc_871 N_X_c_1243_n N_VGND_c_1612_n 0.00222336f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_872 N_X_c_1243_n N_VGND_c_1613_n 0.0140453f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_873 N_X_c_1272_n N_VGND_c_1624_n 0.0223797f $X=5.925 $Y=0.45 $X2=0 $Y2=0
cc_874 N_X_c_1235_n N_VGND_c_1624_n 0.00260082f $X=6.675 $Y=0.82 $X2=0 $Y2=0
cc_875 N_X_c_1235_n N_VGND_c_1626_n 0.00193763f $X=6.675 $Y=0.82 $X2=0 $Y2=0
cc_876 N_X_c_1299_n N_VGND_c_1626_n 0.0221615f $X=6.865 $Y=0.45 $X2=0 $Y2=0
cc_877 N_X_c_1237_n N_VGND_c_1626_n 0.00260082f $X=7.615 $Y=0.82 $X2=0 $Y2=0
cc_878 N_X_c_1237_n N_VGND_c_1628_n 0.00193763f $X=7.615 $Y=0.82 $X2=0 $Y2=0
cc_879 N_X_c_1317_n N_VGND_c_1628_n 0.0221615f $X=7.805 $Y=0.45 $X2=0 $Y2=0
cc_880 N_X_c_1238_n N_VGND_c_1628_n 0.00260082f $X=8.555 $Y=0.82 $X2=0 $Y2=0
cc_881 N_X_c_1238_n N_VGND_c_1630_n 0.00193763f $X=8.555 $Y=0.82 $X2=0 $Y2=0
cc_882 N_X_c_1335_n N_VGND_c_1630_n 0.0216617f $X=8.77 $Y=0.4 $X2=0 $Y2=0
cc_883 N_X_c_1239_n N_VGND_c_1630_n 0.00260082f $X=9.495 $Y=0.82 $X2=0 $Y2=0
cc_884 N_X_c_1239_n N_VGND_c_1632_n 0.00193763f $X=9.495 $Y=0.82 $X2=0 $Y2=0
cc_885 N_X_c_1351_n N_VGND_c_1632_n 0.0216617f $X=9.71 $Y=0.4 $X2=0 $Y2=0
cc_886 N_X_c_1240_n N_VGND_c_1632_n 0.00260082f $X=10.435 $Y=0.82 $X2=0 $Y2=0
cc_887 N_X_c_1240_n N_VGND_c_1634_n 0.00193763f $X=10.435 $Y=0.82 $X2=0 $Y2=0
cc_888 N_X_c_1367_n N_VGND_c_1634_n 0.0216617f $X=10.65 $Y=0.4 $X2=0 $Y2=0
cc_889 N_X_c_1241_n N_VGND_c_1634_n 0.00260082f $X=11.375 $Y=0.82 $X2=0 $Y2=0
cc_890 N_X_c_1241_n N_VGND_c_1636_n 0.00193763f $X=11.375 $Y=0.82 $X2=0 $Y2=0
cc_891 N_X_c_1383_n N_VGND_c_1636_n 0.0216617f $X=11.59 $Y=0.4 $X2=0 $Y2=0
cc_892 N_X_c_1242_n N_VGND_c_1636_n 0.00260082f $X=12.315 $Y=0.82 $X2=0 $Y2=0
cc_893 N_X_c_1242_n N_VGND_c_1638_n 0.00193763f $X=12.315 $Y=0.82 $X2=0 $Y2=0
cc_894 N_X_c_1399_n N_VGND_c_1638_n 0.022456f $X=12.53 $Y=0.4 $X2=0 $Y2=0
cc_895 N_X_c_1243_n N_VGND_c_1638_n 0.00248202f $X=12.92 $Y=0.82 $X2=0 $Y2=0
cc_896 N_X_M1001_s N_VGND_c_1639_n 0.00255377f $X=5.765 $Y=0.235 $X2=0 $Y2=0
cc_897 N_X_M1003_s N_VGND_c_1639_n 0.00255431f $X=6.705 $Y=0.235 $X2=0 $Y2=0
cc_898 N_X_M1007_s N_VGND_c_1639_n 0.00255431f $X=7.645 $Y=0.235 $X2=0 $Y2=0
cc_899 N_X_M1017_s N_VGND_c_1639_n 0.00255524f $X=8.585 $Y=0.235 $X2=0 $Y2=0
cc_900 N_X_M1021_s N_VGND_c_1639_n 0.00255524f $X=9.525 $Y=0.235 $X2=0 $Y2=0
cc_901 N_X_M1026_s N_VGND_c_1639_n 0.00255524f $X=10.465 $Y=0.235 $X2=0 $Y2=0
cc_902 N_X_M1034_s N_VGND_c_1639_n 0.00255524f $X=11.405 $Y=0.235 $X2=0 $Y2=0
cc_903 N_X_M1048_s N_VGND_c_1639_n 0.00304616f $X=12.345 $Y=0.235 $X2=0 $Y2=0
cc_904 N_X_c_1272_n N_VGND_c_1639_n 0.0141899f $X=5.925 $Y=0.45 $X2=0 $Y2=0
cc_905 N_X_c_1235_n N_VGND_c_1639_n 0.00961016f $X=6.675 $Y=0.82 $X2=0 $Y2=0
cc_906 N_X_c_1299_n N_VGND_c_1639_n 0.0141768f $X=6.865 $Y=0.45 $X2=0 $Y2=0
cc_907 N_X_c_1237_n N_VGND_c_1639_n 0.00961016f $X=7.615 $Y=0.82 $X2=0 $Y2=0
cc_908 N_X_c_1317_n N_VGND_c_1639_n 0.0141768f $X=7.805 $Y=0.45 $X2=0 $Y2=0
cc_909 N_X_c_1238_n N_VGND_c_1639_n 0.00961016f $X=8.555 $Y=0.82 $X2=0 $Y2=0
cc_910 N_X_c_1335_n N_VGND_c_1639_n 0.0140924f $X=8.77 $Y=0.4 $X2=0 $Y2=0
cc_911 N_X_c_1239_n N_VGND_c_1639_n 0.00961016f $X=9.495 $Y=0.82 $X2=0 $Y2=0
cc_912 N_X_c_1351_n N_VGND_c_1639_n 0.0140924f $X=9.71 $Y=0.4 $X2=0 $Y2=0
cc_913 N_X_c_1240_n N_VGND_c_1639_n 0.00961016f $X=10.435 $Y=0.82 $X2=0 $Y2=0
cc_914 N_X_c_1367_n N_VGND_c_1639_n 0.0140924f $X=10.65 $Y=0.4 $X2=0 $Y2=0
cc_915 N_X_c_1241_n N_VGND_c_1639_n 0.00961016f $X=11.375 $Y=0.82 $X2=0 $Y2=0
cc_916 N_X_c_1383_n N_VGND_c_1639_n 0.0140924f $X=11.59 $Y=0.4 $X2=0 $Y2=0
cc_917 N_X_c_1242_n N_VGND_c_1639_n 0.00961016f $X=12.315 $Y=0.82 $X2=0 $Y2=0
cc_918 N_X_c_1399_n N_VGND_c_1639_n 0.0142976f $X=12.53 $Y=0.4 $X2=0 $Y2=0
cc_919 N_X_c_1243_n N_VGND_c_1639_n 0.00943502f $X=12.92 $Y=0.82 $X2=0 $Y2=0
