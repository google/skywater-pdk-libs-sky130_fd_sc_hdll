* File: sky130_fd_sc_hdll__clkinv_12.spice
* Created: Wed Sep  2 08:26:01 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__clkinv_12.pex.spice"
.subckt sky130_fd_sc_hdll__clkinv_12  VNB VPB A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1002 N_Y_M1002_d N_A_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.273 PD=0.69 PS=2.14 NRD=0 NRS=12.852 M=1 R=2.8 SA=75000.6 SB=75005.7
+ A=0.063 P=1.14 MULT=1
MM1006 N_Y_M1002_d N_A_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001 SB=75005.3
+ A=0.063 P=1.14 MULT=1
MM1009 N_Y_M1009_d N_A_M1009_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.5 SB=75004.8
+ A=0.063 P=1.14 MULT=1
MM1010 N_Y_M1009_d N_A_M1010_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75001.9 SB=75004.3
+ A=0.063 P=1.14 MULT=1
MM1013 N_Y_M1013_d N_A_M1013_g N_VGND_M1010_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75002.5 SB=75003.8
+ A=0.063 P=1.14 MULT=1
MM1014 N_Y_M1013_d N_A_M1014_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75002.9 SB=75003.4
+ A=0.063 P=1.14 MULT=1
MM1017 N_Y_M1017_d N_A_M1017_g N_VGND_M1014_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75003.4 SB=75002.9
+ A=0.063 P=1.14 MULT=1
MM1020 N_Y_M1017_d N_A_M1020_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75003.8 SB=75002.5
+ A=0.063 P=1.14 MULT=1
MM1024 N_Y_M1024_d N_A_M1024_g N_VGND_M1020_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75004.3 SB=75001.9
+ A=0.063 P=1.14 MULT=1
MM1026 N_Y_M1024_d N_A_M1026_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75004.8 SB=75001.5
+ A=0.063 P=1.14 MULT=1
MM1027 N_Y_M1027_d N_A_M1027_g N_VGND_M1026_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.0777 PD=0.69 PS=0.79 NRD=0 NRS=12.852 M=1 R=2.8 SA=75005.3 SB=75001
+ A=0.063 P=1.14 MULT=1
MM1028 N_Y_M1027_d N_A_M1028_g N_VGND_M1028_s VNB NSHORT L=0.15 W=0.42 AD=0.0567
+ AS=0.273 PD=0.69 PS=2.14 NRD=0 NRS=12.852 M=1 R=2.8 SA=75005.7 SB=75000.6
+ A=0.063 P=1.14 MULT=1
MM1000 N_VPWR_M1000_d N_A_M1000_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90008.2 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g N_Y_M1000_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.6
+ SB=90007.7 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1001_d N_A_M1003_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.1
+ SB=90007.2 A=0.18 P=2.36 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g N_Y_M1003_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90006.8 A=0.18 P=2.36 MULT=1
MM1005 N_VPWR_M1004_d N_A_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.1
+ SB=90006.3 A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90002.5
+ SB=90005.8 A=0.18 P=2.36 MULT=1
MM1008 N_VPWR_M1007_d N_A_M1008_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003
+ SB=90005.3 A=0.18 P=2.36 MULT=1
MM1011 N_VPWR_M1011_d N_A_M1011_g N_Y_M1008_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.5
+ SB=90004.9 A=0.18 P=2.36 MULT=1
MM1012 N_VPWR_M1011_d N_A_M1012_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90003.9
+ SB=90004.4 A=0.18 P=2.36 MULT=1
MM1015 N_VPWR_M1015_d N_A_M1015_g N_Y_M1012_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.4
+ SB=90003.9 A=0.18 P=2.36 MULT=1
MM1016 N_VPWR_M1015_d N_A_M1016_g N_Y_M1016_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90004.9
+ SB=90003.5 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_M1018_g N_Y_M1016_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.3
+ SB=90003 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1018_d N_A_M1019_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90005.8
+ SB=90002.5 A=0.18 P=2.36 MULT=1
MM1021 N_VPWR_M1021_d N_A_M1021_g N_Y_M1019_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.3
+ SB=90002.1 A=0.18 P=2.36 MULT=1
MM1022 N_VPWR_M1021_d N_A_M1022_g N_Y_M1022_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90006.8
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1023 N_VPWR_M1023_d N_A_M1023_g N_Y_M1022_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.2
+ SB=90001.1 A=0.18 P=2.36 MULT=1
MM1025 N_VPWR_M1023_d N_A_M1025_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90007.7
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1029 N_VPWR_M1029_d N_A_M1029_g N_Y_M1025_s VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90008.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX30_noxref VNB VPB NWDIODE A=15.3759 P=22.37
*
.include "sky130_fd_sc_hdll__clkinv_12.pxi.spice"
*
.ends
*
*
