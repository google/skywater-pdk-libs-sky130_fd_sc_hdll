* File: sky130_fd_sc_hdll__o22a_2.spice
* Created: Wed Sep  2 08:45:21 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__o22a_2.pex.spice"
.subckt sky130_fd_sc_hdll__o22a_2  VNB VPB B1 B2 A2 A1 VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A1	A1
* A2	A2
* B2	B2
* B1	B1
* VPB	VPB
* VNB	VNB
MM1006 N_X_M1006_d N_A_83_21#_M1006_g N_VGND_M1006_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.1755 PD=0.96 PS=1.84 NRD=6.456 NRS=0.912 M=1 R=4.33333
+ SA=75000.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1009 N_X_M1006_d N_A_83_21#_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10075 AS=0.2015 PD=0.96 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1011 N_A_83_21#_M1011_d N_B1_M1011_g N_A_321_47#_M1011_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.2 SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1000 N_A_321_47#_M1000_d N_B2_M1000_g N_A_83_21#_M1011_d VNB NSHORT L=0.15
+ W=0.65 AD=0.16575 AS=0.08775 PD=1.16 PS=0.92 NRD=23.988 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A2_M1008_g N_A_321_47#_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.09425 AS=0.16575 PD=0.94 PS=1.16 NRD=0 NRS=18.456 M=1 R=4.33333
+ SA=75001.3 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1004 N_A_321_47#_M1004_d N_A1_M1004_g N_VGND_M1008_d VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.09425 PD=1.82 PS=0.94 NRD=0 NRS=2.76 M=1 R=4.33333 SA=75001.8
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1001 N_X_M1001_d N_A_83_21#_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90003.1 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1001_d N_A_83_21#_M1010_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.4 PD=1.29 PS=1.8 NRD=0.9653 NRS=8.8453 M=1 R=5.55556 SA=90000.7
+ SB=90002.7 A=0.18 P=2.36 MULT=1
MM1005 A_411_297# N_B1_M1005_g N_VPWR_M1010_s VPB PHIGHVT L=0.18 W=1 AD=0.115
+ AS=0.4 PD=1.23 PS=1.8 NRD=11.8003 NRS=0.9653 M=1 R=5.55556 SA=90001.6
+ SB=90001.7 A=0.18 P=2.36 MULT=1
MM1007 N_A_83_21#_M1007_d N_B2_M1007_g A_411_297# VPB PHIGHVT L=0.18 W=1
+ AD=0.245 AS=0.115 PD=1.49 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556
+ SA=90002.1 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1002 A_627_297# N_A2_M1002_g N_A_83_21#_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.245 PD=1.23 PS=1.49 NRD=11.8003 NRS=40.3653 M=1 R=5.55556
+ SA=90002.7 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1003 N_VPWR_M1003_d N_A1_M1003_g A_627_297# VPB PHIGHVT L=0.18 W=1 AD=0.29
+ AS=0.115 PD=2.58 PS=1.23 NRD=0.9653 NRS=11.8003 M=1 R=5.55556 SA=90003.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_14 B2 B2 PROBETYPE=1
c_35 VNB 0 3.11972e-19 $X=0.13 $Y=-0.085
*
.include "sky130_fd_sc_hdll__o22a_2.pxi.spice"
*
.ends
*
*
