* NGSPICE file created from sky130_fd_sc_hdll__xnor2_2.ext - technology: sky130A

.subckt sky130_fd_sc_hdll__xnor2_2 A B VGND VNB VPB VPWR Y
M1000 a_514_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=8.5e+11p pd=7.7e+06u as=1.43e+12p ps=1.286e+07u
M1001 Y a_27_297# a_600_47# VNB nshort w=650000u l=150000u
+  ad=3.38e+11p pd=3.64e+06u as=7.4425e+11p ps=6.19e+06u
M1002 a_27_47# A VGND VNB nshort w=650000u l=150000u
+  ad=5.6875e+11p pd=5.65e+06u as=7.345e+11p ps=7.46e+06u
M1003 VGND A a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1004 VGND B a_600_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1005 VPWR B a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=8.65e+11p ps=7.73e+06u
M1006 VPWR A a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1007 a_27_47# B a_27_297# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=2.405e+11p ps=2.04e+06u
M1008 VPWR a_27_297# Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=6.15e+11p ps=5.23e+06u
M1009 a_27_297# A VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1010 Y a_27_297# VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1011 VGND A a_600_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1012 VPWR A a_27_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_600_47# a_27_297# Y VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1014 a_600_47# B VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1015 Y B a_514_297# VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1016 a_27_297# B VPWR VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
M1017 a_27_297# B a_27_47# VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1018 a_600_47# A VGND VNB nshort w=650000u l=150000u
+  ad=0p pd=0u as=0p ps=0u
M1019 a_514_297# B Y VPB phighvt w=1e+06u l=180000u
+  ad=0p pd=0u as=0p ps=0u
.ends

