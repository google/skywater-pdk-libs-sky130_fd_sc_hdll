* File: sky130_fd_sc_hdll__a21oi_1.pex.spice
* Created: Thu Aug 27 18:53:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%B1 1 3 4 6 7 8 14
r28 14 15 3.31956 $w=3.63e-07 $l=2.5e-08 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.54 $Y2=1.202
r29 12 14 36.5152 $w=3.63e-07 $l=2.75e-07 $layer=POLY_cond $X=0.24 $Y=1.202
+ $X2=0.515 $Y2=1.202
r30 8 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.24
+ $Y=1.16 $X2=0.24 $Y2=1.16
r31 7 8 14.8857 $w=2.38e-07 $l=3.1e-07 $layer=LI1_cond $X=0.215 $Y=0.85
+ $X2=0.215 $Y2=1.16
r32 4 15 23.5056 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.54 $Y2=1.202
r33 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r34 1 14 19.1638 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.202
r35 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%A1 1 3 4 6 7 8 9 25 27
r38 16 27 2.85155 $w=2.3e-07 $l=1.65e-07 $layer=LI1_cond $X=1.18 $Y=0.995
+ $X2=1.18 $Y2=1.16
r39 15 25 5.41299 $w=3.28e-07 $l=1.55e-07 $layer=LI1_cond $X=0.995 $Y=1.16
+ $X2=1.15 $Y2=1.16
r40 14 15 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.995
+ $Y=1.16 $X2=0.995 $Y2=1.16
r41 9 27 0.174613 $w=3.28e-07 $l=5e-09 $layer=LI1_cond $X=1.175 $Y=1.16 $X2=1.18
+ $Y2=1.16
r42 9 25 0.873063 $w=3.28e-07 $l=2.5e-08 $layer=LI1_cond $X=1.175 $Y=1.16
+ $X2=1.15 $Y2=1.16
r43 8 16 7.2654 $w=2.28e-07 $l=1.45e-07 $layer=LI1_cond $X=1.18 $Y=0.85 $X2=1.18
+ $Y2=0.995
r44 7 8 17.0361 $w=2.28e-07 $l=3.4e-07 $layer=LI1_cond $X=1.18 $Y=0.51 $X2=1.18
+ $Y2=0.85
r45 4 14 38.578 $w=2.95e-07 $l=1.65e-07 $layer=POLY_cond $X=1.02 $Y=0.995
+ $X2=1.02 $Y2=1.16
r46 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.02 $Y=0.995 $X2=1.02
+ $Y2=0.56
r47 1 14 48.1208 $w=2.95e-07 $l=2.62202e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=1.02 $Y2=1.16
r48 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.995 $Y=1.41
+ $X2=0.995 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%A2 1 3 4 6 7 10 15
r25 10 12 30.9481 $w=3.66e-07 $l=2.35e-07 $layer=POLY_cond $X=1.49 $Y=1.202
+ $X2=1.725 $Y2=1.202
r26 9 10 3.29235 $w=3.66e-07 $l=2.5e-08 $layer=POLY_cond $X=1.465 $Y=1.202
+ $X2=1.49 $Y2=1.202
r27 7 15 2.09535 $w=3.28e-07 $l=6e-08 $layer=LI1_cond $X=1.67 $Y=1.16 $X2=1.61
+ $Y2=1.16
r28 7 12 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.725
+ $Y=1.16 $X2=1.725 $Y2=1.16
r29 4 10 19.3576 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.49 $Y=1.41
+ $X2=1.49 $Y2=1.202
r30 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.49 $Y=1.41 $X2=1.49
+ $Y2=1.985
r31 1 9 23.7042 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=1.202
r32 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.465 $Y=0.995
+ $X2=1.465 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%Y 1 2 8 9 21 22
r24 21 22 16.7628 $w=2.73e-07 $l=4e-07 $layer=LI1_cond $X=0.232 $Y=1.81
+ $X2=0.232 $Y2=2.21
r25 13 21 5.23838 $w=2.73e-07 $l=1.25e-07 $layer=LI1_cond $X=0.232 $Y=1.685
+ $X2=0.232 $Y2=1.81
r26 9 11 5.15111 $w=2.25e-07 $l=9.5e-08 $layer=LI1_cond $X=0.772 $Y=0.645
+ $X2=0.772 $Y2=0.55
r27 8 13 22.4737 $w=1.88e-07 $l=3.85e-07 $layer=LI1_cond $X=0.617 $Y=1.59
+ $X2=0.232 $Y2=1.59
r28 7 9 9.5505 $w=1.78e-07 $l=1.55e-07 $layer=LI1_cond $X=0.617 $Y=0.735
+ $X2=0.772 $Y2=0.735
r29 7 8 34.3172 $w=2.23e-07 $l=6.7e-07 $layer=LI1_cond $X=0.617 $Y=0.825
+ $X2=0.617 $Y2=1.495
r30 2 21 300 $w=1.7e-07 $l=3.82426e-07 $layer=licon1_PDIFF $count=2 $X=0.15
+ $Y=1.485 $X2=0.275 $Y2=1.81
r31 1 11 182 $w=1.7e-07 $l=3.78583e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.755 $Y2=0.55
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%A_121_297# 1 2 7 8 9 11
r28 9 17 3.96742 $w=3.8e-07 $l=2.5e-07 $layer=LI1_cond $X=1.705 $Y=2.025
+ $X2=1.705 $Y2=1.775
r29 9 11 9.24987 $w=3.78e-07 $l=3.05e-07 $layer=LI1_cond $X=1.705 $Y=2.025
+ $X2=1.705 $Y2=2.33
r30 8 15 8.47222 $w=2.52e-07 $l=2.63344e-07 $layer=LI1_cond $X=0.92 $Y=1.775
+ $X2=0.73 $Y2=1.95
r31 7 17 3.01524 $w=5e-07 $l=1.9e-07 $layer=LI1_cond $X=1.515 $Y=1.775 $X2=1.705
+ $Y2=1.775
r32 7 8 14.2333 $w=4.98e-07 $l=5.95e-07 $layer=LI1_cond $X=1.515 $Y=1.775
+ $X2=0.92 $Y2=1.775
r33 2 17 400 $w=1.7e-07 $l=2.2798e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.485 $X2=1.73 $Y2=1.65
r34 2 11 400 $w=1.7e-07 $l=9.16938e-07 $layer=licon1_PDIFF $count=1 $X=1.58
+ $Y=1.485 $X2=1.73 $Y2=2.33
r35 1 15 300 $w=1.7e-07 $l=5.34766e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.755 $Y2=1.95
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%VPWR 1 6 8 10 17 18 21
r29 21 22 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r30 18 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=1.15 $Y2=2.72
r31 17 18 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r32 15 21 5.78184 $w=1.7e-07 $l=9.8e-08 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=1.237 $Y2=2.72
r33 15 17 47.9519 $w=1.68e-07 $l=7.35e-07 $layer=LI1_cond $X=1.335 $Y=2.72
+ $X2=2.07 $Y2=2.72
r34 10 21 5.78184 $w=1.7e-07 $l=9.7e-08 $layer=LI1_cond $X=1.14 $Y=2.72
+ $X2=1.237 $Y2=2.72
r35 10 12 59.369 $w=1.68e-07 $l=9.1e-07 $layer=LI1_cond $X=1.14 $Y=2.72 $X2=0.23
+ $Y2=2.72
r36 8 22 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r37 8 12 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r38 4 21 0.85348 $w=1.95e-07 $l=8.5e-08 $layer=LI1_cond $X=1.237 $Y=2.635
+ $X2=1.237 $Y2=2.72
r39 4 6 15.641 $w=1.93e-07 $l=2.75e-07 $layer=LI1_cond $X=1.237 $Y=2.635
+ $X2=1.237 $Y2=2.36
r40 1 6 600 $w=1.7e-07 $l=9.47035e-07 $layer=licon1_PDIFF $count=1 $X=1.085
+ $Y=1.485 $X2=1.235 $Y2=2.36
.ends

.subckt PM_SKY130_FD_SC_HDLL__A21OI_1%VGND 1 2 7 9 13 15 17 24 25 31
r28 31 32 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r29 25 32 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=0 $X2=1.61
+ $Y2=0
r30 24 25 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r31 22 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=1.745
+ $Y2=0
r32 22 24 11.4171 $w=1.68e-07 $l=1.75e-07 $layer=LI1_cond $X=1.895 $Y=0 $X2=2.07
+ $Y2=0
r33 21 32 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r34 20 21 6.2 $w=1.7e-07 $l=2.55e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r35 18 28 4.746 $w=1.7e-07 $l=2.2e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.22
+ $Y2=0
r36 18 20 16.3102 $w=1.68e-07 $l=2.5e-07 $layer=LI1_cond $X=0.44 $Y=0 $X2=0.69
+ $Y2=0
r37 17 31 8.04615 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=1.745
+ $Y2=0
r38 17 20 59.0428 $w=1.68e-07 $l=9.05e-07 $layer=LI1_cond $X=1.595 $Y=0 $X2=0.69
+ $Y2=0
r39 15 21 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r40 15 28 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r41 11 31 0.597483 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0
r42 11 13 17.0946 $w=2.98e-07 $l=4.45e-07 $layer=LI1_cond $X=1.745 $Y=0.085
+ $X2=1.745 $Y2=0.53
r43 7 28 3.02018 $w=3.3e-07 $l=1.09087e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.22 $Y2=0
r44 7 9 10.3021 $w=3.28e-07 $l=2.95e-07 $layer=LI1_cond $X=0.275 $Y=0.085
+ $X2=0.275 $Y2=0.38
r45 2 13 182 $w=1.7e-07 $l=3.78253e-07 $layer=licon1_NDIFF $count=1 $X=1.54
+ $Y=0.235 $X2=1.73 $Y2=0.53
r46 1 9 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=0.15
+ $Y=0.235 $X2=0.275 $Y2=0.38
.ends

