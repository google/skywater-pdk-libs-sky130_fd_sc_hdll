# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand4_1
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand4_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  2.760000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.175000 0.995000 2.640000 1.665000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.030000 0.300000 1.415000 0.825000 ;
        RECT 1.245000 0.825000 1.415000 0.995000 ;
        RECT 1.245000 0.995000 1.605000 1.325000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 0.300000 0.860000 0.995000 ;
        RECT 0.595000 0.995000 1.075000 1.325000 ;
    END
  END C
  PIN D
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 0.995000 0.395000 1.325000 ;
    END
  END D
  PIN VGND
    ANTENNADIFFAREA  0.201500 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 2.760000 0.240000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  0.870000 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 2.760000 2.960000 ;
    END
  END VPWR
  PIN Y
    ANTENNADIFFAREA  0.867500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 1.495000 1.945000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.535000 1.665000 1.865000 2.465000 ;
        RECT 1.670000 0.255000 2.415000 0.825000 ;
        RECT 1.775000 0.825000 1.945000 1.495000 ;
    END
  END Y
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 2.760000 0.085000 ;
      RECT 0.000000  2.635000 2.760000 2.805000 ;
      RECT 0.085000  1.495000 0.345000 2.635000 ;
      RECT 0.090000  0.085000 0.425000 0.825000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 2.115000  1.835000 2.395000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand4_1
END LIBRARY
