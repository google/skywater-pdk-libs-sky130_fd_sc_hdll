* File: sky130_fd_sc_hdll__clkinv_1.pxi.spice
* Created: Thu Aug 27 19:02:38 2020
* 
x_PM_SKY130_FD_SC_HDLL__CLKINV_1%A N_A_c_26_n N_A_M1001_g N_A_c_27_n N_A_M1002_g
+ N_A_M1000_g A A A N_A_c_25_n PM_SKY130_FD_SC_HDLL__CLKINV_1%A
x_PM_SKY130_FD_SC_HDLL__CLKINV_1%VPWR N_VPWR_M1001_s N_VPWR_M1002_s
+ N_VPWR_c_54_n N_VPWR_c_55_n N_VPWR_c_56_n N_VPWR_c_57_n VPWR N_VPWR_c_58_n
+ N_VPWR_c_53_n N_VPWR_c_60_n PM_SKY130_FD_SC_HDLL__CLKINV_1%VPWR
x_PM_SKY130_FD_SC_HDLL__CLKINV_1%Y N_Y_M1000_s N_Y_M1001_d N_Y_c_75_n Y Y Y Y Y
+ PM_SKY130_FD_SC_HDLL__CLKINV_1%Y
x_PM_SKY130_FD_SC_HDLL__CLKINV_1%VGND N_VGND_M1000_d N_VGND_c_99_n VGND
+ N_VGND_c_100_n N_VGND_c_101_n N_VGND_c_102_n N_VGND_c_103_n
+ PM_SKY130_FD_SC_HDLL__CLKINV_1%VGND
cc_1 VNB N_A_M1000_g 0.0419142f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.445
cc_2 VNB A 0.0441542f $X=-0.19 $Y=-0.24 $X2=0.145 $Y2=0.425
cc_3 VNB N_A_c_25_n 0.0776019f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.282
cc_4 VNB N_VPWR_c_53_n 0.079965f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.282
cc_5 VNB N_Y_c_75_n 0.01275f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.445
cc_6 VNB Y 0.0373569f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_7 VNB N_VGND_c_99_n 0.019189f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=2.065
cc_8 VNB N_VGND_c_100_n 0.0315538f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_VGND_c_101_n 0.0163041f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.282
cc_10 VNB N_VGND_c_102_n 0.147925f $X=-0.19 $Y=-0.24 $X2=0.24 $Y2=1.16
cc_11 VNB N_VGND_c_103_n 0.00535963f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.282
cc_12 VPB N_A_c_26_n 0.0207574f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.57
cc_13 VPB N_A_c_27_n 0.0207627f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.57
cc_14 VPB A 0.00366f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_15 VPB N_A_c_25_n 0.0581351f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.282
cc_16 VPB N_VPWR_c_54_n 0.00988417f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_17 VPB N_VPWR_c_55_n 0.036748f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.445
cc_18 VPB N_VPWR_c_56_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.145 $Y2=0.425
cc_19 VPB N_VPWR_c_57_n 0.0373169f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_20 VPB N_VPWR_c_58_n 0.0163041f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.282
cc_21 VPB N_VPWR_c_53_n 0.0569095f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=1.282
cc_22 VPB N_VPWR_c_60_n 0.00535984f $X=-0.19 $Y=1.305 $X2=0.205 $Y2=1.16
cc_23 N_A_c_26_n N_VPWR_c_55_n 0.00966062f $X=0.495 $Y=1.57 $X2=0 $Y2=0
cc_24 A N_VPWR_c_55_n 0.0123519f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_25 N_A_c_25_n N_VPWR_c_55_n 0.00232912f $X=0.965 $Y=1.282 $X2=0 $Y2=0
cc_26 N_A_c_26_n N_VPWR_c_56_n 0.00597712f $X=0.495 $Y=1.57 $X2=0 $Y2=0
cc_27 N_A_c_27_n N_VPWR_c_56_n 0.00673617f $X=0.965 $Y=1.57 $X2=0 $Y2=0
cc_28 N_A_c_27_n N_VPWR_c_57_n 0.0103794f $X=0.965 $Y=1.57 $X2=0 $Y2=0
cc_29 N_A_c_26_n N_VPWR_c_53_n 0.010906f $X=0.495 $Y=1.57 $X2=0 $Y2=0
cc_30 N_A_c_27_n N_VPWR_c_53_n 0.0131262f $X=0.965 $Y=1.57 $X2=0 $Y2=0
cc_31 N_A_M1000_g N_Y_c_75_n 0.00510869f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_32 A N_Y_c_75_n 0.029238f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_33 N_A_c_25_n N_Y_c_75_n 0.00147778f $X=0.965 $Y=1.282 $X2=0 $Y2=0
cc_34 N_A_c_26_n Y 0.0190937f $X=0.495 $Y=1.57 $X2=0 $Y2=0
cc_35 N_A_c_27_n Y 0.0165568f $X=0.965 $Y=1.57 $X2=0 $Y2=0
cc_36 A Y 0.00237165f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_37 N_A_c_25_n Y 0.0360099f $X=0.965 $Y=1.282 $X2=0 $Y2=0
cc_38 N_A_M1000_g Y 0.0170244f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_39 A Y 0.0396815f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_40 N_A_c_25_n Y 0.0431462f $X=0.965 $Y=1.282 $X2=0 $Y2=0
cc_41 N_A_M1000_g N_VGND_c_99_n 0.00452839f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_42 N_A_M1000_g N_VGND_c_100_n 0.00442535f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_43 A N_VGND_c_100_n 0.00966373f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_44 N_A_M1000_g N_VGND_c_102_n 0.00870582f $X=0.99 $Y=0.445 $X2=0 $Y2=0
cc_45 A N_VGND_c_102_n 0.00857725f $X=0.145 $Y=0.425 $X2=0 $Y2=0
cc_46 N_VPWR_c_53_n N_Y_M1001_d 0.00231261f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_47 N_VPWR_c_55_n Y 0.0616326f $X=0.26 $Y=1.83 $X2=0 $Y2=0
cc_48 N_VPWR_c_56_n Y 0.0223557f $X=1.115 $Y=2.72 $X2=0 $Y2=0
cc_49 N_VPWR_c_57_n Y 0.0508287f $X=1.2 $Y=1.83 $X2=0 $Y2=0
cc_50 N_VPWR_c_53_n Y 0.0140101f $X=1.61 $Y=2.72 $X2=0 $Y2=0
cc_51 N_VPWR_c_57_n Y 0.0142613f $X=1.2 $Y=1.83 $X2=0 $Y2=0
cc_52 Y N_VGND_c_99_n 0.023949f $X=1.165 $Y=0.765 $X2=0 $Y2=0
cc_53 N_Y_c_75_n N_VGND_c_100_n 0.0247439f $X=0.725 $Y=0.435 $X2=0 $Y2=0
cc_54 Y N_VGND_c_100_n 0.00321253f $X=1.165 $Y=0.765 $X2=0 $Y2=0
cc_55 N_Y_M1000_s N_VGND_c_102_n 0.00268143f $X=0.6 $Y=0.235 $X2=0 $Y2=0
cc_56 N_Y_c_75_n N_VGND_c_102_n 0.0142553f $X=0.725 $Y=0.435 $X2=0 $Y2=0
cc_57 Y N_VGND_c_102_n 0.00641982f $X=1.165 $Y=0.765 $X2=0 $Y2=0
