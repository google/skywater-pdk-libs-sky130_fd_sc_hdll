* File: sky130_fd_sc_hdll__nand2b_1.spice
* Created: Thu Aug 27 19:13:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nand2b_1.pex.spice"
.subckt sky130_fd_sc_hdll__nand2b_1  VNB VPB A_N B VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* B	B
* A_N	A_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_A_N_M1002_g N_A_27_93#_M1002_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0914579 AS=0.1302 PD=0.812523 PS=1.46 NRD=46.5 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.2 A=0.063 P=1.14 MULT=1
MM1005 A_226_47# N_B_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65 AD=0.08775
+ AS=0.141542 PD=0.92 PS=1.25748 NRD=14.76 NRS=8.304 M=1 R=4.33333 SA=75000.6
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_Y_M1004_d N_A_27_93#_M1004_g A_226_47# VNB NSHORT L=0.15 W=0.65
+ AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=14.76 M=1 R=4.33333
+ SA=75001 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_A_N_M1000_g N_A_27_93#_M1000_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0904183 AS=0.1134 PD=0.801549 PS=1.38 NRD=75.1752 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90001.2 A=0.0756 P=1.2 MULT=1
MM1003 N_Y_M1003_d N_B_M1003_g N_VPWR_M1000_d VPB PHIGHVT L=0.18 W=1 AD=0.145
+ AS=0.215282 PD=1.29 PS=1.90845 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.4
+ SB=90000.6 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_27_93#_M1001_g N_Y_M1003_d VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90000.2 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
pX7_noxref noxref_10 Y Y PROBETYPE=1
pX8_noxref noxref_11 Y Y PROBETYPE=1
pX9_noxref noxref_12 Y Y PROBETYPE=1
pX10_noxref noxref_13 Y Y PROBETYPE=1
pX11_noxref noxref_14 Y Y PROBETYPE=1
*
.include "sky130_fd_sc_hdll__nand2b_1.pxi.spice"
*
.ends
*
*
