* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__clkbuf_8 A VGND VNB VPB VPWR X
X0 VGND A a_118_297# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X1 X a_118_297# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X2 VPWR A a_118_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X3 X a_118_297# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X4 X a_118_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND a_118_297# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X6 VGND a_118_297# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X7 a_118_297# A VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_118_297# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X9 VPWR a_118_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND a_118_297# X VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 X a_118_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 VPWR a_118_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 X a_118_297# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X14 VPWR a_118_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 X a_118_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 a_118_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 VPWR a_118_297# X VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X18 X a_118_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X19 X a_118_297# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
.ends
