# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__sdfxtp_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__sdfxtp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.96000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN CLK
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN D
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.745000 1.355000 3.150000 1.685000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  1.028500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.030000 0.305000 10.410000 0.735000 ;
        RECT 10.030000 0.735000 11.850000 0.905000 ;
        RECT 10.030000 1.505000 11.850000 1.675000 ;
        RECT 10.030000 1.675000 10.410000 2.395000 ;
        RECT 10.980000 0.305000 11.360000 0.735000 ;
        RECT 10.980000 1.675000 11.360000 2.395000 ;
        RECT 11.550000 0.905000 11.850000 1.505000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.178200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.725000 1.035000 4.095000 1.655000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.356400 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.880000 0.615000 3.505000 0.785000 ;
        RECT 1.880000 0.785000 2.215000 1.685000 ;
        RECT 3.335000 0.785000 3.505000 1.115000 ;
    END
  END SCE
  PIN VNB
    PORT
      LAYER pwell ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
    END
  END VNB
  PIN VPB
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 12.150000 2.910000 ;
    END
  END VPB
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.960000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 11.960000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.000000 -0.085000 11.960000 0.085000 ;
      RECT  0.000000  2.635000 11.960000 2.805000 ;
      RECT  0.175000  0.345000  0.345000 0.635000 ;
      RECT  0.175000  0.635000  0.895000 0.805000 ;
      RECT  0.180000  1.795000  0.895000 1.965000 ;
      RECT  0.180000  1.965000  0.350000 2.465000 ;
      RECT  0.515000  0.085000  0.895000 0.465000 ;
      RECT  0.520000  2.135000  0.900000 2.635000 ;
      RECT  0.665000  0.805000  0.895000 1.795000 ;
      RECT  1.115000  0.345000  1.345000 2.465000 ;
      RECT  1.535000  0.275000  1.905000 0.445000 ;
      RECT  1.535000  0.445000  1.705000 1.860000 ;
      RECT  1.535000  1.860000  3.525000 2.075000 ;
      RECT  1.535000  2.075000  1.810000 2.445000 ;
      RECT  1.980000  2.245000  2.360000 2.635000 ;
      RECT  2.125000  0.085000  2.455000 0.445000 ;
      RECT  2.385000  0.955000  2.715000 1.125000 ;
      RECT  2.385000  1.125000  2.555000 1.860000 ;
      RECT  2.895000  2.245000  3.890000 2.415000 ;
      RECT  3.070000  0.275000  3.895000 0.445000 ;
      RECT  3.330000  1.355000  3.525000 1.860000 ;
      RECT  3.720000  1.825000  4.735000 1.995000 ;
      RECT  3.720000  1.995000  3.890000 2.245000 ;
      RECT  3.725000  0.445000  3.895000 0.695000 ;
      RECT  3.725000  0.695000  4.735000 0.865000 ;
      RECT  4.110000  2.165000  4.280000 2.635000 ;
      RECT  4.115000  0.085000  4.315000 0.525000 ;
      RECT  4.565000  0.365000  4.915000 0.535000 ;
      RECT  4.565000  0.535000  4.735000 0.695000 ;
      RECT  4.565000  0.865000  4.735000 1.825000 ;
      RECT  4.565000  1.995000  4.735000 2.065000 ;
      RECT  4.565000  2.065000  4.800000 2.440000 ;
      RECT  4.905000  0.705000  5.535000 1.035000 ;
      RECT  4.905000  1.035000  5.195000 1.905000 ;
      RECT  5.045000  2.190000  6.265000 2.360000 ;
      RECT  5.135000  0.365000  5.895000 0.535000 ;
      RECT  5.385000  1.655000  5.875000 2.010000 ;
      RECT  5.725000  0.535000  5.895000 1.245000 ;
      RECT  5.725000  1.245000  6.605000 1.485000 ;
      RECT  6.045000  1.485000  6.605000 1.575000 ;
      RECT  6.045000  1.575000  6.265000 2.190000 ;
      RECT  6.065000  0.765000  6.995000 1.065000 ;
      RECT  6.225000  0.085000  6.595000 0.585000 ;
      RECT  6.435000  1.835000  6.605000 2.635000 ;
      RECT  6.775000  0.365000  7.285000 0.535000 ;
      RECT  6.775000  0.535000  6.995000 0.765000 ;
      RECT  6.775000  1.065000  6.995000 2.135000 ;
      RECT  6.775000  2.135000  7.075000 2.465000 ;
      RECT  7.165000  0.705000  7.765000 1.035000 ;
      RECT  7.165000  1.245000  7.405000 1.965000 ;
      RECT  7.300000  2.165000  8.335000 2.335000 ;
      RECT  7.565000  0.365000  8.205000 0.535000 ;
      RECT  7.575000  1.035000  7.765000 1.575000 ;
      RECT  7.575000  1.575000  7.945000 1.905000 ;
      RECT  7.985000  0.535000  8.205000 0.995000 ;
      RECT  7.985000  0.995000  9.150000 1.325000 ;
      RECT  7.985000  1.325000  8.335000 1.405000 ;
      RECT  8.165000  1.405000  8.335000 2.165000 ;
      RECT  8.450000  0.085000  8.870000 0.615000 ;
      RECT  8.555000  1.575000  9.505000 1.905000 ;
      RECT  8.565000  2.135000  8.870000 2.635000 ;
      RECT  9.140000  0.300000  9.500000 0.825000 ;
      RECT  9.220000  1.905000  9.505000 2.455000 ;
      RECT  9.320000  0.825000  9.500000 1.075000 ;
      RECT  9.320000  1.075000 11.380000 1.325000 ;
      RECT  9.320000  1.325000  9.505000 1.575000 ;
      RECT  9.690000  0.085000  9.860000 0.695000 ;
      RECT  9.690000  1.625000  9.860000 2.635000 ;
      RECT 10.640000  0.085000 10.810000 0.565000 ;
      RECT 10.640000  1.845000 10.810000 2.635000 ;
      RECT 11.580000  0.085000 11.750000 0.565000 ;
      RECT 11.580000  1.845000 11.750000 2.635000 ;
    LAYER mcon ;
      RECT  0.145000 -0.085000  0.315000 0.085000 ;
      RECT  0.145000  2.635000  0.315000 2.805000 ;
      RECT  0.605000 -0.085000  0.775000 0.085000 ;
      RECT  0.605000  2.635000  0.775000 2.805000 ;
      RECT  0.665000  1.740000  0.835000 1.910000 ;
      RECT  1.065000 -0.085000  1.235000 0.085000 ;
      RECT  1.065000  2.635000  1.235000 2.805000 ;
      RECT  1.155000  0.720000  1.325000 0.890000 ;
      RECT  1.525000 -0.085000  1.695000 0.085000 ;
      RECT  1.525000  2.635000  1.695000 2.805000 ;
      RECT  1.985000 -0.085000  2.155000 0.085000 ;
      RECT  1.985000  2.635000  2.155000 2.805000 ;
      RECT  2.445000 -0.085000  2.615000 0.085000 ;
      RECT  2.445000  2.635000  2.615000 2.805000 ;
      RECT  2.905000 -0.085000  3.075000 0.085000 ;
      RECT  2.905000  2.635000  3.075000 2.805000 ;
      RECT  3.365000 -0.085000  3.535000 0.085000 ;
      RECT  3.365000  2.635000  3.535000 2.805000 ;
      RECT  3.825000 -0.085000  3.995000 0.085000 ;
      RECT  3.825000  2.635000  3.995000 2.805000 ;
      RECT  4.285000 -0.085000  4.455000 0.085000 ;
      RECT  4.285000  2.635000  4.455000 2.805000 ;
      RECT  4.745000 -0.085000  4.915000 0.085000 ;
      RECT  4.745000  2.635000  4.915000 2.805000 ;
      RECT  5.155000  0.720000  5.325000 0.890000 ;
      RECT  5.205000 -0.085000  5.375000 0.085000 ;
      RECT  5.205000  2.635000  5.375000 2.805000 ;
      RECT  5.665000 -0.085000  5.835000 0.085000 ;
      RECT  5.665000  1.740000  5.835000 1.910000 ;
      RECT  5.665000  2.635000  5.835000 2.805000 ;
      RECT  6.125000 -0.085000  6.295000 0.085000 ;
      RECT  6.125000  2.635000  6.295000 2.805000 ;
      RECT  6.585000 -0.085000  6.755000 0.085000 ;
      RECT  6.585000  2.635000  6.755000 2.805000 ;
      RECT  7.045000 -0.085000  7.215000 0.085000 ;
      RECT  7.045000  2.635000  7.215000 2.805000 ;
      RECT  7.225000  0.720000  7.395000 0.890000 ;
      RECT  7.225000  1.740000  7.395000 1.910000 ;
      RECT  7.505000 -0.085000  7.675000 0.085000 ;
      RECT  7.505000  2.635000  7.675000 2.805000 ;
      RECT  7.965000 -0.085000  8.135000 0.085000 ;
      RECT  7.965000  2.635000  8.135000 2.805000 ;
      RECT  8.425000 -0.085000  8.595000 0.085000 ;
      RECT  8.425000  2.635000  8.595000 2.805000 ;
      RECT  8.885000 -0.085000  9.055000 0.085000 ;
      RECT  8.885000  2.635000  9.055000 2.805000 ;
      RECT  9.345000 -0.085000  9.515000 0.085000 ;
      RECT  9.345000  2.635000  9.515000 2.805000 ;
      RECT  9.805000 -0.085000  9.975000 0.085000 ;
      RECT  9.805000  2.635000  9.975000 2.805000 ;
      RECT 10.265000 -0.085000 10.435000 0.085000 ;
      RECT 10.265000  2.635000 10.435000 2.805000 ;
      RECT 10.725000 -0.085000 10.895000 0.085000 ;
      RECT 10.725000  2.635000 10.895000 2.805000 ;
      RECT 11.185000 -0.085000 11.355000 0.085000 ;
      RECT 11.185000  2.635000 11.355000 2.805000 ;
      RECT 11.645000 -0.085000 11.815000 0.085000 ;
      RECT 11.645000  2.635000 11.815000 2.805000 ;
    LAYER met1 ;
      RECT 0.605000 1.710000 0.895000 1.800000 ;
      RECT 0.605000 1.800000 7.455000 1.940000 ;
      RECT 1.095000 0.690000 1.385000 0.780000 ;
      RECT 1.095000 0.780000 7.455000 0.920000 ;
      RECT 5.045000 0.690000 5.385000 0.780000 ;
      RECT 5.555000 1.710000 5.895000 1.800000 ;
      RECT 7.115000 0.690000 7.455000 0.780000 ;
      RECT 7.115000 1.710000 7.455000 1.800000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__sdfxtp_4
END LIBRARY
