# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__or3_4
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.600000 BY  2.720000 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.325000 1.075000 1.850000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.595000 1.075000 1.155000 1.325000 ;
        RECT 0.595000 1.325000 0.830000 2.050000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.425000 1.325000 ;
    END
  END C
  PIN VGND
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  PIN X
    ANTENNADIFFAREA  0.996000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.455000 0.265000 2.835000 0.735000 ;
        RECT 2.455000 0.735000 4.455000 0.905000 ;
        RECT 2.545000 1.445000 4.455000 1.615000 ;
        RECT 2.545000 1.615000 2.795000 2.465000 ;
        RECT 3.395000 0.265000 3.775000 0.735000 ;
        RECT 3.485000 1.615000 3.735000 2.465000 ;
        RECT 4.115000 0.905000 4.455000 1.445000 ;
    END
  END X
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.600000 0.085000 ;
      RECT 0.000000  2.635000 4.600000 2.805000 ;
      RECT 0.085000  0.255000 0.425000 0.725000 ;
      RECT 0.085000  0.725000 2.240000 0.905000 ;
      RECT 0.085000  1.495000 0.425000 2.295000 ;
      RECT 0.085000  2.295000 1.365000 2.465000 ;
      RECT 0.645000  0.085000 0.815000 0.555000 ;
      RECT 0.985000  0.255000 1.365000 0.725000 ;
      RECT 1.100000  1.495000 2.240000 1.665000 ;
      RECT 1.100000  1.665000 1.365000 2.295000 ;
      RECT 1.585000  0.085000 2.285000 0.555000 ;
      RECT 1.585000  1.835000 2.285000 2.635000 ;
      RECT 2.020000  0.905000 2.240000 1.075000 ;
      RECT 2.020000  1.075000 3.945000 1.245000 ;
      RECT 2.020000  1.245000 2.240000 1.495000 ;
      RECT 3.015000  1.795000 3.265000 2.635000 ;
      RECT 3.055000  0.085000 3.225000 0.555000 ;
      RECT 3.955000  1.795000 4.205000 2.635000 ;
      RECT 3.995000  0.085000 4.165000 0.555000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__or3_4
END LIBRARY
