# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__muxb8to1_4
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__muxb8to1_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  24.84000 BY  5.440000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D[0]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 1.055000 6.045000 1.325000 ;
    END
  END D[0]
  PIN D[1]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.655000 4.115000 6.045000 4.385000 ;
    END
  END D[1]
  PIN D[2]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.375000 1.055000 7.765000 1.325000 ;
    END
  END D[2]
  PIN D[3]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.375000 4.115000 7.765000 4.385000 ;
    END
  END D[3]
  PIN D[4]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.075000 1.055000 18.465000 1.325000 ;
    END
  END D[4]
  PIN D[5]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 17.075000 4.115000 18.465000 4.385000 ;
    END
  END D[5]
  PIN D[6]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.795000 1.055000 20.185000 1.325000 ;
    END
  END D[6]
  PIN D[7]
    ANTENNAGATEAREA  1.110000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 18.795000 4.115000 20.185000 4.385000 ;
    END
  END D[7]
  PIN S[0]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.995000 0.680000 1.325000 ;
    END
  END S[0]
  PIN S[1]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 4.115000 0.680000 4.445000 ;
    END
  END S[1]
  PIN S[2]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.740000 0.995000 12.335000 1.325000 ;
    END
  END S[2]
  PIN S[3]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 11.740000 4.115000 12.335000 4.445000 ;
    END
  END S[3]
  PIN S[4]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 0.995000 13.100000 1.325000 ;
    END
  END S[4]
  PIN S[5]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.505000 4.115000 13.100000 4.445000 ;
    END
  END S[5]
  PIN S[6]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.160000 0.995000 24.755000 1.325000 ;
    END
  END S[6]
  PIN S[7]
    ANTENNAGATEAREA  0.733200 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 24.160000 4.115000 24.755000 4.445000 ;
    END
  END S[7]
  PIN VGND
    ANTENNADIFFAREA  3.070600 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 24.840000 0.085000 ;
        RECT  0.270000  0.085000  0.560000 0.610000 ;
        RECT  1.190000  0.085000  1.480000 0.610000 ;
        RECT  4.185000  0.085000  4.435000 0.545000 ;
        RECT  5.105000  0.085000  5.375000 0.545000 ;
        RECT  6.045000  0.085000  6.375000 0.885000 ;
        RECT  7.045000  0.085000  7.315000 0.545000 ;
        RECT  7.985000  0.085000  8.235000 0.545000 ;
        RECT 10.940000  0.085000 11.230000 0.610000 ;
        RECT 11.860000  0.085000 12.150000 0.610000 ;
        RECT 12.690000  0.085000 12.980000 0.610000 ;
        RECT 13.610000  0.085000 13.900000 0.610000 ;
        RECT 16.605000  0.085000 16.855000 0.545000 ;
        RECT 17.525000  0.085000 17.795000 0.545000 ;
        RECT 18.465000  0.085000 18.795000 0.885000 ;
        RECT 19.465000  0.085000 19.735000 0.545000 ;
        RECT 20.405000  0.085000 20.655000 0.545000 ;
        RECT 23.360000  0.085000 23.650000 0.610000 ;
        RECT 24.280000  0.085000 24.570000 0.610000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
        RECT 14.405000 -0.085000 14.575000 0.085000 ;
        RECT 14.865000 -0.085000 15.035000 0.085000 ;
        RECT 15.325000 -0.085000 15.495000 0.085000 ;
        RECT 15.785000 -0.085000 15.955000 0.085000 ;
        RECT 16.245000 -0.085000 16.415000 0.085000 ;
        RECT 16.705000 -0.085000 16.875000 0.085000 ;
        RECT 17.165000 -0.085000 17.335000 0.085000 ;
        RECT 17.625000 -0.085000 17.795000 0.085000 ;
        RECT 18.085000 -0.085000 18.255000 0.085000 ;
        RECT 18.545000 -0.085000 18.715000 0.085000 ;
        RECT 19.005000 -0.085000 19.175000 0.085000 ;
        RECT 19.465000 -0.085000 19.635000 0.085000 ;
        RECT 19.925000 -0.085000 20.095000 0.085000 ;
        RECT 20.385000 -0.085000 20.555000 0.085000 ;
        RECT 20.845000 -0.085000 21.015000 0.085000 ;
        RECT 21.305000 -0.085000 21.475000 0.085000 ;
        RECT 21.765000 -0.085000 21.935000 0.085000 ;
        RECT 22.225000 -0.085000 22.395000 0.085000 ;
        RECT 22.685000 -0.085000 22.855000 0.085000 ;
        RECT 23.145000 -0.085000 23.315000 0.085000 ;
        RECT 23.605000 -0.085000 23.775000 0.085000 ;
        RECT 24.065000 -0.085000 24.235000 0.085000 ;
        RECT 24.525000 -0.085000 24.695000 0.085000 ;
    END
    PORT
      LAYER li1 ;
        RECT  0.000000 5.355000 24.840000 5.525000 ;
        RECT  0.270000 4.830000  0.560000 5.355000 ;
        RECT  1.190000 4.830000  1.480000 5.355000 ;
        RECT  4.185000 4.895000  4.435000 5.355000 ;
        RECT  5.105000 4.895000  5.375000 5.355000 ;
        RECT  6.045000 4.555000  6.375000 5.355000 ;
        RECT  7.045000 4.895000  7.315000 5.355000 ;
        RECT  7.985000 4.895000  8.235000 5.355000 ;
        RECT 10.940000 4.830000 11.230000 5.355000 ;
        RECT 11.860000 4.830000 12.150000 5.355000 ;
        RECT 12.690000 4.830000 12.980000 5.355000 ;
        RECT 13.610000 4.830000 13.900000 5.355000 ;
        RECT 16.605000 4.895000 16.855000 5.355000 ;
        RECT 17.525000 4.895000 17.795000 5.355000 ;
        RECT 18.465000 4.555000 18.795000 5.355000 ;
        RECT 19.465000 4.895000 19.735000 5.355000 ;
        RECT 20.405000 4.895000 20.655000 5.355000 ;
        RECT 23.360000 4.830000 23.650000 5.355000 ;
        RECT 24.280000 4.830000 24.570000 5.355000 ;
      LAYER mcon ;
        RECT  0.145000 5.355000  0.315000 5.525000 ;
        RECT  0.605000 5.355000  0.775000 5.525000 ;
        RECT  1.065000 5.355000  1.235000 5.525000 ;
        RECT  1.525000 5.355000  1.695000 5.525000 ;
        RECT  1.985000 5.355000  2.155000 5.525000 ;
        RECT  2.445000 5.355000  2.615000 5.525000 ;
        RECT  2.905000 5.355000  3.075000 5.525000 ;
        RECT  3.365000 5.355000  3.535000 5.525000 ;
        RECT  3.825000 5.355000  3.995000 5.525000 ;
        RECT  4.285000 5.355000  4.455000 5.525000 ;
        RECT  4.745000 5.355000  4.915000 5.525000 ;
        RECT  5.205000 5.355000  5.375000 5.525000 ;
        RECT  5.665000 5.355000  5.835000 5.525000 ;
        RECT  6.125000 5.355000  6.295000 5.525000 ;
        RECT  6.585000 5.355000  6.755000 5.525000 ;
        RECT  7.045000 5.355000  7.215000 5.525000 ;
        RECT  7.505000 5.355000  7.675000 5.525000 ;
        RECT  7.965000 5.355000  8.135000 5.525000 ;
        RECT  8.425000 5.355000  8.595000 5.525000 ;
        RECT  8.885000 5.355000  9.055000 5.525000 ;
        RECT  9.345000 5.355000  9.515000 5.525000 ;
        RECT  9.805000 5.355000  9.975000 5.525000 ;
        RECT 10.265000 5.355000 10.435000 5.525000 ;
        RECT 10.725000 5.355000 10.895000 5.525000 ;
        RECT 11.185000 5.355000 11.355000 5.525000 ;
        RECT 11.645000 5.355000 11.815000 5.525000 ;
        RECT 12.105000 5.355000 12.275000 5.525000 ;
        RECT 12.565000 5.355000 12.735000 5.525000 ;
        RECT 13.025000 5.355000 13.195000 5.525000 ;
        RECT 13.485000 5.355000 13.655000 5.525000 ;
        RECT 13.945000 5.355000 14.115000 5.525000 ;
        RECT 14.405000 5.355000 14.575000 5.525000 ;
        RECT 14.865000 5.355000 15.035000 5.525000 ;
        RECT 15.325000 5.355000 15.495000 5.525000 ;
        RECT 15.785000 5.355000 15.955000 5.525000 ;
        RECT 16.245000 5.355000 16.415000 5.525000 ;
        RECT 16.705000 5.355000 16.875000 5.525000 ;
        RECT 17.165000 5.355000 17.335000 5.525000 ;
        RECT 17.625000 5.355000 17.795000 5.525000 ;
        RECT 18.085000 5.355000 18.255000 5.525000 ;
        RECT 18.545000 5.355000 18.715000 5.525000 ;
        RECT 19.005000 5.355000 19.175000 5.525000 ;
        RECT 19.465000 5.355000 19.635000 5.525000 ;
        RECT 19.925000 5.355000 20.095000 5.525000 ;
        RECT 20.385000 5.355000 20.555000 5.525000 ;
        RECT 20.845000 5.355000 21.015000 5.525000 ;
        RECT 21.305000 5.355000 21.475000 5.525000 ;
        RECT 21.765000 5.355000 21.935000 5.525000 ;
        RECT 22.225000 5.355000 22.395000 5.525000 ;
        RECT 22.685000 5.355000 22.855000 5.525000 ;
        RECT 23.145000 5.355000 23.315000 5.525000 ;
        RECT 23.605000 5.355000 23.775000 5.525000 ;
        RECT 24.065000 5.355000 24.235000 5.525000 ;
        RECT 24.525000 5.355000 24.695000 5.525000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 24.840000 0.240000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 5.200000 24.840000 5.680000 ;
    END
  END VGND
  PIN VPWR
    ANTENNADIFFAREA  9.422400 ;
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 16.065000 2.635000 21.195000 2.805000 ;
        RECT 16.585000 1.835000 16.855000 2.635000 ;
        RECT 16.585000 2.805000 16.855000 3.605000 ;
        RECT 17.525000 1.835000 17.795000 2.635000 ;
        RECT 17.525000 2.805000 17.795000 3.605000 ;
        RECT 18.465000 1.495000 18.795000 2.635000 ;
        RECT 18.465000 2.805000 18.795000 3.945000 ;
        RECT 19.465000 1.835000 19.735000 2.635000 ;
        RECT 19.465000 2.805000 19.735000 3.605000 ;
        RECT 20.405000 1.835000 20.675000 2.635000 ;
        RECT 20.405000 2.805000 20.675000 3.605000 ;
      LAYER mcon ;
        RECT 16.245000 2.635000 16.415000 2.805000 ;
        RECT 16.705000 2.635000 16.875000 2.805000 ;
        RECT 17.165000 2.635000 17.335000 2.805000 ;
        RECT 17.625000 2.635000 17.795000 2.805000 ;
        RECT 18.085000 2.635000 18.255000 2.805000 ;
        RECT 18.545000 2.635000 18.715000 2.805000 ;
        RECT 19.005000 2.635000 19.175000 2.805000 ;
        RECT 19.465000 2.635000 19.635000 2.805000 ;
        RECT 19.925000 2.635000 20.095000 2.805000 ;
        RECT 20.385000 2.635000 20.555000 2.805000 ;
        RECT 20.845000 2.635000 21.015000 2.805000 ;
    END
    PORT
      LAYER li1 ;
        RECT 3.645000 2.635000 8.775000 2.805000 ;
        RECT 4.165000 1.835000 4.435000 2.635000 ;
        RECT 4.165000 2.805000 4.435000 3.605000 ;
        RECT 5.105000 1.835000 5.375000 2.635000 ;
        RECT 5.105000 2.805000 5.375000 3.605000 ;
        RECT 6.045000 1.495000 6.375000 2.635000 ;
        RECT 6.045000 2.805000 6.375000 3.945000 ;
        RECT 7.045000 1.835000 7.315000 2.635000 ;
        RECT 7.045000 2.805000 7.315000 3.605000 ;
        RECT 7.985000 1.835000 8.255000 2.635000 ;
        RECT 7.985000 2.805000 8.255000 3.605000 ;
      LAYER mcon ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 24.840000 2.960000 ;
    END
  END VPWR
  PIN Z
    ANTENNADIFFAREA  6.051200 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.205000 1.065000 3.475000 1.365000 ;
        RECT 2.205000 1.365000 2.535000 4.075000 ;
        RECT 2.205000 4.075000 3.475000 4.375000 ;
        RECT 2.405000 0.595000 2.735000 1.065000 ;
        RECT 2.405000 4.375000 2.735000 4.845000 ;
        RECT 3.145000 1.365000 3.475000 4.075000 ;
        RECT 3.245000 0.595000 3.575000 0.885000 ;
        RECT 3.245000 0.885000 3.475000 1.065000 ;
        RECT 3.245000 4.375000 3.475000 4.555000 ;
        RECT 3.245000 4.555000 3.575000 4.845000 ;
      LAYER mcon ;
        RECT 2.285000 1.785000 2.455000 1.955000 ;
        RECT 2.285000 3.485000 2.455000 3.655000 ;
        RECT 3.225000 1.785000 3.395000 1.955000 ;
        RECT 3.225000 3.485000 3.395000 3.655000 ;
    END
    PORT
      LAYER met1 ;
        RECT  2.225000 1.755000  2.515000 1.800000 ;
        RECT  2.225000 1.800000 22.615000 1.940000 ;
        RECT  2.225000 1.940000  2.515000 1.985000 ;
        RECT  2.225000 3.455000  2.515000 3.500000 ;
        RECT  2.225000 3.500000 22.615000 3.640000 ;
        RECT  2.225000 3.640000  2.515000 3.685000 ;
        RECT  3.165000 1.755000  3.455000 1.800000 ;
        RECT  3.165000 1.940000  3.455000 1.985000 ;
        RECT  3.165000 3.455000  3.455000 3.500000 ;
        RECT  3.165000 3.640000  3.455000 3.685000 ;
        RECT  8.965000 1.755000  9.255000 1.800000 ;
        RECT  8.965000 1.940000  9.255000 1.985000 ;
        RECT  8.965000 3.455000  9.255000 3.500000 ;
        RECT  8.965000 3.640000  9.255000 3.685000 ;
        RECT  9.905000 1.755000 10.195000 1.800000 ;
        RECT  9.905000 1.940000 10.195000 1.985000 ;
        RECT  9.905000 3.455000 10.195000 3.500000 ;
        RECT  9.905000 3.640000 10.195000 3.685000 ;
        RECT 14.645000 1.755000 14.935000 1.800000 ;
        RECT 14.645000 1.940000 14.935000 1.985000 ;
        RECT 14.645000 3.455000 14.935000 3.500000 ;
        RECT 14.645000 3.640000 14.935000 3.685000 ;
        RECT 15.585000 1.755000 15.875000 1.800000 ;
        RECT 15.585000 1.940000 15.875000 1.985000 ;
        RECT 15.585000 3.455000 15.875000 3.500000 ;
        RECT 15.585000 3.640000 15.875000 3.685000 ;
        RECT 21.385000 1.755000 21.675000 1.800000 ;
        RECT 21.385000 1.940000 21.675000 1.985000 ;
        RECT 21.385000 3.455000 21.675000 3.500000 ;
        RECT 21.385000 3.640000 21.675000 3.685000 ;
        RECT 22.325000 1.755000 22.615000 1.800000 ;
        RECT 22.325000 1.940000 22.615000 1.985000 ;
        RECT 22.325000 3.455000 22.615000 3.500000 ;
        RECT 22.325000 3.640000 22.615000 3.685000 ;
    END
  END Z
  OBS
    LAYER li1 ;
      RECT  0.000000 2.635000  2.035000 2.805000 ;
      RECT  0.220000 1.605000  0.520000 2.635000 ;
      RECT  0.220000 2.805000  0.520000 3.835000 ;
      RECT  0.690000 1.605000  1.020000 2.465000 ;
      RECT  0.690000 2.975000  1.020000 3.835000 ;
      RECT  0.770000 0.280000  1.020000 0.825000 ;
      RECT  0.770000 4.615000  1.020000 5.160000 ;
      RECT  0.850000 0.825000  1.020000 1.065000 ;
      RECT  0.850000 1.065000  2.035000 1.395000 ;
      RECT  0.850000 1.395000  1.020000 1.605000 ;
      RECT  0.850000 3.835000  1.020000 4.045000 ;
      RECT  0.850000 4.045000  2.035000 4.375000 ;
      RECT  0.850000 4.375000  1.020000 4.615000 ;
      RECT  1.215000 1.605000  1.490000 2.635000 ;
      RECT  1.215000 2.805000  1.490000 3.835000 ;
      RECT  1.735000 1.565000  2.035000 2.465000 ;
      RECT  1.735000 2.975000  2.035000 3.875000 ;
      RECT  1.985000 0.255000  4.015000 0.425000 ;
      RECT  1.985000 0.425000  2.235000 0.770000 ;
      RECT  1.985000 4.670000  2.235000 5.015000 ;
      RECT  1.985000 5.015000  4.015000 5.185000 ;
      RECT  2.705000 1.535000  2.975000 2.465000 ;
      RECT  2.705000 2.975000  2.975000 3.905000 ;
      RECT  2.905000 0.425000  3.075000 0.770000 ;
      RECT  2.905000 4.670000  3.075000 5.015000 ;
      RECT  3.645000 1.495000  5.875000 1.665000 ;
      RECT  3.645000 1.665000  3.945000 2.465000 ;
      RECT  3.645000 2.975000  3.945000 3.775000 ;
      RECT  3.645000 3.775000  5.875000 3.945000 ;
      RECT  3.745000 0.425000  4.015000 0.715000 ;
      RECT  3.745000 0.715000  5.875000 0.885000 ;
      RECT  3.745000 4.555000  5.875000 4.725000 ;
      RECT  3.745000 4.725000  4.015000 5.015000 ;
      RECT  4.605000 0.255000  4.935000 0.715000 ;
      RECT  4.605000 1.665000  4.935000 2.465000 ;
      RECT  4.605000 2.975000  4.935000 3.775000 ;
      RECT  4.605000 4.725000  4.935000 5.185000 ;
      RECT  5.545000 0.255000  5.875000 0.715000 ;
      RECT  5.545000 1.665000  5.875000 2.465000 ;
      RECT  5.545000 2.975000  5.875000 3.775000 ;
      RECT  5.545000 4.725000  5.875000 5.185000 ;
      RECT  6.545000 0.255000  6.875000 0.715000 ;
      RECT  6.545000 0.715000  8.675000 0.885000 ;
      RECT  6.545000 1.495000  8.775000 1.665000 ;
      RECT  6.545000 1.665000  6.875000 2.465000 ;
      RECT  6.545000 2.975000  6.875000 3.775000 ;
      RECT  6.545000 3.775000  8.775000 3.945000 ;
      RECT  6.545000 4.555000  8.675000 4.725000 ;
      RECT  6.545000 4.725000  6.875000 5.185000 ;
      RECT  7.485000 0.255000  7.815000 0.715000 ;
      RECT  7.485000 1.665000  7.815000 2.465000 ;
      RECT  7.485000 2.975000  7.815000 3.775000 ;
      RECT  7.485000 4.725000  7.815000 5.185000 ;
      RECT  8.405000 0.255000 10.435000 0.425000 ;
      RECT  8.405000 0.425000  8.675000 0.715000 ;
      RECT  8.405000 4.725000  8.675000 5.015000 ;
      RECT  8.405000 5.015000 10.435000 5.185000 ;
      RECT  8.475000 1.665000  8.775000 2.465000 ;
      RECT  8.475000 2.975000  8.775000 3.775000 ;
      RECT  8.845000 0.595000  9.175000 0.885000 ;
      RECT  8.845000 4.555000  9.175000 4.845000 ;
      RECT  8.945000 0.885000  9.175000 1.065000 ;
      RECT  8.945000 1.065000 10.215000 1.365000 ;
      RECT  8.945000 1.365000  9.275000 4.075000 ;
      RECT  8.945000 4.075000 10.215000 4.375000 ;
      RECT  8.945000 4.375000  9.175000 4.555000 ;
      RECT  9.345000 0.425000  9.515000 0.770000 ;
      RECT  9.345000 4.670000  9.515000 5.015000 ;
      RECT  9.445000 1.535000  9.715000 2.465000 ;
      RECT  9.445000 2.975000  9.715000 3.905000 ;
      RECT  9.685000 0.595000 10.015000 1.065000 ;
      RECT  9.685000 4.375000 10.015000 4.845000 ;
      RECT  9.885000 1.365000 10.215000 4.075000 ;
      RECT 10.185000 0.425000 10.435000 0.770000 ;
      RECT 10.185000 4.670000 10.435000 5.015000 ;
      RECT 10.385000 1.065000 11.570000 1.395000 ;
      RECT 10.385000 1.565000 10.685000 2.465000 ;
      RECT 10.385000 2.635000 14.455000 2.805000 ;
      RECT 10.385000 2.975000 10.685000 3.875000 ;
      RECT 10.385000 4.045000 11.570000 4.375000 ;
      RECT 10.930000 1.605000 11.205000 2.635000 ;
      RECT 10.930000 2.805000 11.205000 3.835000 ;
      RECT 11.400000 0.280000 11.650000 0.825000 ;
      RECT 11.400000 0.825000 11.570000 1.065000 ;
      RECT 11.400000 1.395000 11.570000 1.605000 ;
      RECT 11.400000 1.605000 11.730000 2.465000 ;
      RECT 11.400000 2.975000 11.730000 3.835000 ;
      RECT 11.400000 3.835000 11.570000 4.045000 ;
      RECT 11.400000 4.375000 11.570000 4.615000 ;
      RECT 11.400000 4.615000 11.650000 5.160000 ;
      RECT 11.900000 1.605000 12.200000 2.635000 ;
      RECT 11.900000 2.805000 12.200000 3.835000 ;
      RECT 12.640000 1.605000 12.940000 2.635000 ;
      RECT 12.640000 2.805000 12.940000 3.835000 ;
      RECT 13.110000 1.605000 13.440000 2.465000 ;
      RECT 13.110000 2.975000 13.440000 3.835000 ;
      RECT 13.190000 0.280000 13.440000 0.825000 ;
      RECT 13.190000 4.615000 13.440000 5.160000 ;
      RECT 13.270000 0.825000 13.440000 1.065000 ;
      RECT 13.270000 1.065000 14.455000 1.395000 ;
      RECT 13.270000 1.395000 13.440000 1.605000 ;
      RECT 13.270000 3.835000 13.440000 4.045000 ;
      RECT 13.270000 4.045000 14.455000 4.375000 ;
      RECT 13.270000 4.375000 13.440000 4.615000 ;
      RECT 13.635000 1.605000 13.910000 2.635000 ;
      RECT 13.635000 2.805000 13.910000 3.835000 ;
      RECT 14.155000 1.565000 14.455000 2.465000 ;
      RECT 14.155000 2.975000 14.455000 3.875000 ;
      RECT 14.405000 0.255000 16.435000 0.425000 ;
      RECT 14.405000 0.425000 14.655000 0.770000 ;
      RECT 14.405000 4.670000 14.655000 5.015000 ;
      RECT 14.405000 5.015000 16.435000 5.185000 ;
      RECT 14.625000 1.065000 15.895000 1.365000 ;
      RECT 14.625000 1.365000 14.955000 4.075000 ;
      RECT 14.625000 4.075000 15.895000 4.375000 ;
      RECT 14.825000 0.595000 15.155000 1.065000 ;
      RECT 14.825000 4.375000 15.155000 4.845000 ;
      RECT 15.125000 1.535000 15.395000 2.465000 ;
      RECT 15.125000 2.975000 15.395000 3.905000 ;
      RECT 15.325000 0.425000 15.495000 0.770000 ;
      RECT 15.325000 4.670000 15.495000 5.015000 ;
      RECT 15.565000 1.365000 15.895000 4.075000 ;
      RECT 15.665000 0.595000 15.995000 0.885000 ;
      RECT 15.665000 0.885000 15.895000 1.065000 ;
      RECT 15.665000 4.375000 15.895000 4.555000 ;
      RECT 15.665000 4.555000 15.995000 4.845000 ;
      RECT 16.065000 1.495000 18.295000 1.665000 ;
      RECT 16.065000 1.665000 16.365000 2.465000 ;
      RECT 16.065000 2.975000 16.365000 3.775000 ;
      RECT 16.065000 3.775000 18.295000 3.945000 ;
      RECT 16.165000 0.425000 16.435000 0.715000 ;
      RECT 16.165000 0.715000 18.295000 0.885000 ;
      RECT 16.165000 4.555000 18.295000 4.725000 ;
      RECT 16.165000 4.725000 16.435000 5.015000 ;
      RECT 17.025000 0.255000 17.355000 0.715000 ;
      RECT 17.025000 1.665000 17.355000 2.465000 ;
      RECT 17.025000 2.975000 17.355000 3.775000 ;
      RECT 17.025000 4.725000 17.355000 5.185000 ;
      RECT 17.965000 0.255000 18.295000 0.715000 ;
      RECT 17.965000 1.665000 18.295000 2.465000 ;
      RECT 17.965000 2.975000 18.295000 3.775000 ;
      RECT 17.965000 4.725000 18.295000 5.185000 ;
      RECT 18.965000 0.255000 19.295000 0.715000 ;
      RECT 18.965000 0.715000 21.095000 0.885000 ;
      RECT 18.965000 1.495000 21.195000 1.665000 ;
      RECT 18.965000 1.665000 19.295000 2.465000 ;
      RECT 18.965000 2.975000 19.295000 3.775000 ;
      RECT 18.965000 3.775000 21.195000 3.945000 ;
      RECT 18.965000 4.555000 21.095000 4.725000 ;
      RECT 18.965000 4.725000 19.295000 5.185000 ;
      RECT 19.905000 0.255000 20.235000 0.715000 ;
      RECT 19.905000 1.665000 20.235000 2.465000 ;
      RECT 19.905000 2.975000 20.235000 3.775000 ;
      RECT 19.905000 4.725000 20.235000 5.185000 ;
      RECT 20.825000 0.255000 22.855000 0.425000 ;
      RECT 20.825000 0.425000 21.095000 0.715000 ;
      RECT 20.825000 4.725000 21.095000 5.015000 ;
      RECT 20.825000 5.015000 22.855000 5.185000 ;
      RECT 20.895000 1.665000 21.195000 2.465000 ;
      RECT 20.895000 2.975000 21.195000 3.775000 ;
      RECT 21.265000 0.595000 21.595000 0.885000 ;
      RECT 21.265000 4.555000 21.595000 4.845000 ;
      RECT 21.365000 0.885000 21.595000 1.065000 ;
      RECT 21.365000 1.065000 22.635000 1.365000 ;
      RECT 21.365000 1.365000 21.695000 4.075000 ;
      RECT 21.365000 4.075000 22.635000 4.375000 ;
      RECT 21.365000 4.375000 21.595000 4.555000 ;
      RECT 21.765000 0.425000 21.935000 0.770000 ;
      RECT 21.765000 4.670000 21.935000 5.015000 ;
      RECT 21.865000 1.535000 22.135000 2.465000 ;
      RECT 21.865000 2.975000 22.135000 3.905000 ;
      RECT 22.105000 0.595000 22.435000 1.065000 ;
      RECT 22.105000 4.375000 22.435000 4.845000 ;
      RECT 22.305000 1.365000 22.635000 4.075000 ;
      RECT 22.605000 0.425000 22.855000 0.770000 ;
      RECT 22.605000 4.670000 22.855000 5.015000 ;
      RECT 22.805000 1.065000 23.990000 1.395000 ;
      RECT 22.805000 1.565000 23.105000 2.465000 ;
      RECT 22.805000 2.635000 24.840000 2.805000 ;
      RECT 22.805000 2.975000 23.105000 3.875000 ;
      RECT 22.805000 4.045000 23.990000 4.375000 ;
      RECT 23.350000 1.605000 23.625000 2.635000 ;
      RECT 23.350000 2.805000 23.625000 3.835000 ;
      RECT 23.820000 0.280000 24.070000 0.825000 ;
      RECT 23.820000 0.825000 23.990000 1.065000 ;
      RECT 23.820000 1.395000 23.990000 1.605000 ;
      RECT 23.820000 1.605000 24.150000 2.465000 ;
      RECT 23.820000 2.975000 24.150000 3.835000 ;
      RECT 23.820000 3.835000 23.990000 4.045000 ;
      RECT 23.820000 4.375000 23.990000 4.615000 ;
      RECT 23.820000 4.615000 24.070000 5.160000 ;
      RECT 24.320000 1.605000 24.620000 2.635000 ;
      RECT 24.320000 2.805000 24.620000 3.835000 ;
    LAYER mcon ;
      RECT  0.145000 2.635000  0.315000 2.805000 ;
      RECT  0.605000 2.635000  0.775000 2.805000 ;
      RECT  1.065000 2.635000  1.235000 2.805000 ;
      RECT  1.525000 2.635000  1.695000 2.805000 ;
      RECT  1.805000 2.140000  1.975000 2.310000 ;
      RECT  1.805000 3.130000  1.975000 3.300000 ;
      RECT  2.755000 2.140000  2.925000 2.310000 ;
      RECT  2.755000 3.130000  2.925000 3.300000 ;
      RECT  3.705000 2.140000  3.875000 2.310000 ;
      RECT  3.705000 3.130000  3.875000 3.300000 ;
      RECT  4.685000 2.140000  4.855000 2.310000 ;
      RECT  4.685000 3.130000  4.855000 3.300000 ;
      RECT  5.625000 2.140000  5.795000 2.310000 ;
      RECT  5.625000 3.130000  5.795000 3.300000 ;
      RECT  6.625000 2.140000  6.795000 2.310000 ;
      RECT  6.625000 3.130000  6.795000 3.300000 ;
      RECT  7.565000 2.140000  7.735000 2.310000 ;
      RECT  7.565000 3.130000  7.735000 3.300000 ;
      RECT  8.545000 2.140000  8.715000 2.310000 ;
      RECT  8.545000 3.130000  8.715000 3.300000 ;
      RECT  9.025000 1.785000  9.195000 1.955000 ;
      RECT  9.025000 3.485000  9.195000 3.655000 ;
      RECT  9.495000 2.140000  9.665000 2.310000 ;
      RECT  9.495000 3.130000  9.665000 3.300000 ;
      RECT  9.965000 1.785000 10.135000 1.955000 ;
      RECT  9.965000 3.485000 10.135000 3.655000 ;
      RECT 10.445000 2.140000 10.615000 2.310000 ;
      RECT 10.445000 3.130000 10.615000 3.300000 ;
      RECT 10.725000 2.635000 10.895000 2.805000 ;
      RECT 11.185000 2.635000 11.355000 2.805000 ;
      RECT 11.645000 2.635000 11.815000 2.805000 ;
      RECT 12.105000 2.635000 12.275000 2.805000 ;
      RECT 12.565000 2.635000 12.735000 2.805000 ;
      RECT 13.025000 2.635000 13.195000 2.805000 ;
      RECT 13.485000 2.635000 13.655000 2.805000 ;
      RECT 13.945000 2.635000 14.115000 2.805000 ;
      RECT 14.225000 2.140000 14.395000 2.310000 ;
      RECT 14.225000 3.130000 14.395000 3.300000 ;
      RECT 14.705000 1.785000 14.875000 1.955000 ;
      RECT 14.705000 3.485000 14.875000 3.655000 ;
      RECT 15.175000 2.140000 15.345000 2.310000 ;
      RECT 15.175000 3.130000 15.345000 3.300000 ;
      RECT 15.645000 1.785000 15.815000 1.955000 ;
      RECT 15.645000 3.485000 15.815000 3.655000 ;
      RECT 16.125000 2.140000 16.295000 2.310000 ;
      RECT 16.125000 3.130000 16.295000 3.300000 ;
      RECT 17.105000 2.140000 17.275000 2.310000 ;
      RECT 17.105000 3.130000 17.275000 3.300000 ;
      RECT 18.045000 2.140000 18.215000 2.310000 ;
      RECT 18.045000 3.130000 18.215000 3.300000 ;
      RECT 19.045000 2.140000 19.215000 2.310000 ;
      RECT 19.045000 3.130000 19.215000 3.300000 ;
      RECT 19.985000 2.140000 20.155000 2.310000 ;
      RECT 19.985000 3.130000 20.155000 3.300000 ;
      RECT 20.965000 2.140000 21.135000 2.310000 ;
      RECT 20.965000 3.130000 21.135000 3.300000 ;
      RECT 21.445000 1.785000 21.615000 1.955000 ;
      RECT 21.445000 3.485000 21.615000 3.655000 ;
      RECT 21.915000 2.140000 22.085000 2.310000 ;
      RECT 21.915000 3.130000 22.085000 3.300000 ;
      RECT 22.385000 1.785000 22.555000 1.955000 ;
      RECT 22.385000 3.485000 22.555000 3.655000 ;
      RECT 22.865000 2.140000 23.035000 2.310000 ;
      RECT 22.865000 3.130000 23.035000 3.300000 ;
      RECT 23.145000 2.635000 23.315000 2.805000 ;
      RECT 23.605000 2.635000 23.775000 2.805000 ;
      RECT 24.065000 2.635000 24.235000 2.805000 ;
      RECT 24.525000 2.635000 24.695000 2.805000 ;
    LAYER met1 ;
      RECT  1.745000 2.110000  2.035000 2.155000 ;
      RECT  1.745000 2.155000  5.855000 2.295000 ;
      RECT  1.745000 2.295000  2.035000 2.340000 ;
      RECT  1.745000 3.100000  2.035000 3.145000 ;
      RECT  1.745000 3.145000  5.855000 3.285000 ;
      RECT  1.745000 3.285000  2.035000 3.330000 ;
      RECT  2.695000 2.110000  2.985000 2.155000 ;
      RECT  2.695000 2.295000  2.985000 2.340000 ;
      RECT  2.695000 3.100000  2.985000 3.145000 ;
      RECT  2.695000 3.285000  2.985000 3.330000 ;
      RECT  3.645000 2.110000  3.935000 2.155000 ;
      RECT  3.645000 2.295000  3.935000 2.340000 ;
      RECT  3.645000 3.100000  3.935000 3.145000 ;
      RECT  3.645000 3.285000  3.935000 3.330000 ;
      RECT  4.625000 2.110000  4.915000 2.155000 ;
      RECT  4.625000 2.295000  4.915000 2.340000 ;
      RECT  4.625000 3.100000  4.915000 3.145000 ;
      RECT  4.625000 3.285000  4.915000 3.330000 ;
      RECT  5.565000 2.110000  5.855000 2.155000 ;
      RECT  5.565000 2.295000  5.855000 2.340000 ;
      RECT  5.565000 3.100000  5.855000 3.145000 ;
      RECT  5.565000 3.285000  5.855000 3.330000 ;
      RECT  6.565000 2.110000  6.855000 2.155000 ;
      RECT  6.565000 2.155000 10.675000 2.295000 ;
      RECT  6.565000 2.295000  6.855000 2.340000 ;
      RECT  6.565000 3.100000  6.855000 3.145000 ;
      RECT  6.565000 3.145000 10.675000 3.285000 ;
      RECT  6.565000 3.285000  6.855000 3.330000 ;
      RECT  7.505000 2.110000  7.795000 2.155000 ;
      RECT  7.505000 2.295000  7.795000 2.340000 ;
      RECT  7.505000 3.100000  7.795000 3.145000 ;
      RECT  7.505000 3.285000  7.795000 3.330000 ;
      RECT  8.485000 2.110000  8.775000 2.155000 ;
      RECT  8.485000 2.295000  8.775000 2.340000 ;
      RECT  8.485000 3.100000  8.775000 3.145000 ;
      RECT  8.485000 3.285000  8.775000 3.330000 ;
      RECT  9.435000 2.110000  9.725000 2.155000 ;
      RECT  9.435000 2.295000  9.725000 2.340000 ;
      RECT  9.435000 3.100000  9.725000 3.145000 ;
      RECT  9.435000 3.285000  9.725000 3.330000 ;
      RECT 10.385000 2.110000 10.675000 2.155000 ;
      RECT 10.385000 2.295000 10.675000 2.340000 ;
      RECT 10.385000 3.100000 10.675000 3.145000 ;
      RECT 10.385000 3.285000 10.675000 3.330000 ;
      RECT 14.165000 2.110000 14.455000 2.155000 ;
      RECT 14.165000 2.155000 18.275000 2.295000 ;
      RECT 14.165000 2.295000 14.455000 2.340000 ;
      RECT 14.165000 3.100000 14.455000 3.145000 ;
      RECT 14.165000 3.145000 18.275000 3.285000 ;
      RECT 14.165000 3.285000 14.455000 3.330000 ;
      RECT 15.115000 2.110000 15.405000 2.155000 ;
      RECT 15.115000 2.295000 15.405000 2.340000 ;
      RECT 15.115000 3.100000 15.405000 3.145000 ;
      RECT 15.115000 3.285000 15.405000 3.330000 ;
      RECT 16.065000 2.110000 16.355000 2.155000 ;
      RECT 16.065000 2.295000 16.355000 2.340000 ;
      RECT 16.065000 3.100000 16.355000 3.145000 ;
      RECT 16.065000 3.285000 16.355000 3.330000 ;
      RECT 17.045000 2.110000 17.335000 2.155000 ;
      RECT 17.045000 2.295000 17.335000 2.340000 ;
      RECT 17.045000 3.100000 17.335000 3.145000 ;
      RECT 17.045000 3.285000 17.335000 3.330000 ;
      RECT 17.985000 2.110000 18.275000 2.155000 ;
      RECT 17.985000 2.295000 18.275000 2.340000 ;
      RECT 17.985000 3.100000 18.275000 3.145000 ;
      RECT 17.985000 3.285000 18.275000 3.330000 ;
      RECT 18.985000 2.110000 19.275000 2.155000 ;
      RECT 18.985000 2.155000 23.095000 2.295000 ;
      RECT 18.985000 2.295000 19.275000 2.340000 ;
      RECT 18.985000 3.100000 19.275000 3.145000 ;
      RECT 18.985000 3.145000 23.095000 3.285000 ;
      RECT 18.985000 3.285000 19.275000 3.330000 ;
      RECT 19.925000 2.110000 20.215000 2.155000 ;
      RECT 19.925000 2.295000 20.215000 2.340000 ;
      RECT 19.925000 3.100000 20.215000 3.145000 ;
      RECT 19.925000 3.285000 20.215000 3.330000 ;
      RECT 20.905000 2.110000 21.195000 2.155000 ;
      RECT 20.905000 2.295000 21.195000 2.340000 ;
      RECT 20.905000 3.100000 21.195000 3.145000 ;
      RECT 20.905000 3.285000 21.195000 3.330000 ;
      RECT 21.855000 2.110000 22.145000 2.155000 ;
      RECT 21.855000 2.295000 22.145000 2.340000 ;
      RECT 21.855000 3.100000 22.145000 3.145000 ;
      RECT 21.855000 3.285000 22.145000 3.330000 ;
      RECT 22.805000 2.110000 23.095000 2.155000 ;
      RECT 22.805000 2.295000 23.095000 2.340000 ;
      RECT 22.805000 3.100000 23.095000 3.145000 ;
      RECT 22.805000 3.285000 23.095000 3.330000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__muxb8to1_4
END LIBRARY
