* File: sky130_fd_sc_hdll__mux2_1.pxi.spice
* Created: Wed Sep  2 08:34:23 2020
* 
x_PM_SKY130_FD_SC_HDLL__MUX2_1%A_79_21# N_A_79_21#_M1004_d N_A_79_21#_M1002_d
+ N_A_79_21#_c_75_n N_A_79_21#_M1010_g N_A_79_21#_c_76_n N_A_79_21#_M1005_g
+ N_A_79_21#_c_77_n N_A_79_21#_c_78_n N_A_79_21#_c_130_p N_A_79_21#_c_79_n
+ N_A_79_21#_c_85_p N_A_79_21#_c_93_p N_A_79_21#_c_90_p
+ PM_SKY130_FD_SC_HDLL__MUX2_1%A_79_21#
x_PM_SKY130_FD_SC_HDLL__MUX2_1%S N_S_c_149_n N_S_c_150_n N_S_M1009_g N_S_M1000_g
+ N_S_c_151_n N_S_M1011_g N_S_M1008_g N_S_c_153_n N_S_c_154_n N_S_c_155_n
+ N_S_c_156_n N_S_c_157_n N_S_c_147_n N_S_c_148_n S S S
+ PM_SKY130_FD_SC_HDLL__MUX2_1%S
x_PM_SKY130_FD_SC_HDLL__MUX2_1%A1 N_A1_M1004_g N_A1_c_240_n N_A1_M1003_g
+ N_A1_c_237_n N_A1_c_238_n N_A1_c_242_n N_A1_c_243_n A1 A1
+ PM_SKY130_FD_SC_HDLL__MUX2_1%A1
x_PM_SKY130_FD_SC_HDLL__MUX2_1%A0 N_A0_c_302_n N_A0_M1002_g N_A0_c_303_n
+ N_A0_c_304_n N_A0_M1007_g N_A0_c_299_n A0 N_A0_c_300_n N_A0_c_301_n
+ PM_SKY130_FD_SC_HDLL__MUX2_1%A0
x_PM_SKY130_FD_SC_HDLL__MUX2_1%A_657_21# N_A_657_21#_M1008_d N_A_657_21#_M1011_d
+ N_A_657_21#_M1001_g N_A_657_21#_c_346_n N_A_657_21#_c_353_n
+ N_A_657_21#_M1006_g N_A_657_21#_c_347_n N_A_657_21#_c_348_n
+ N_A_657_21#_c_349_n N_A_657_21#_c_350_n N_A_657_21#_c_351_n
+ N_A_657_21#_c_355_n PM_SKY130_FD_SC_HDLL__MUX2_1%A_657_21#
x_PM_SKY130_FD_SC_HDLL__MUX2_1%X N_X_M1010_s N_X_M1005_s N_X_c_395_n X X X
+ PM_SKY130_FD_SC_HDLL__MUX2_1%X
x_PM_SKY130_FD_SC_HDLL__MUX2_1%VPWR N_VPWR_M1005_d N_VPWR_M1006_d N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n VPWR N_VPWR_c_415_n
+ N_VPWR_c_410_n N_VPWR_c_417_n PM_SKY130_FD_SC_HDLL__MUX2_1%VPWR
x_PM_SKY130_FD_SC_HDLL__MUX2_1%VGND N_VGND_M1010_d N_VGND_M1001_d N_VGND_c_452_n
+ N_VGND_c_453_n VGND N_VGND_c_454_n N_VGND_c_455_n N_VGND_c_456_n
+ N_VGND_c_457_n N_VGND_c_458_n N_VGND_c_459_n PM_SKY130_FD_SC_HDLL__MUX2_1%VGND
cc_1 VNB N_A_79_21#_c_75_n 0.0203674f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_A_79_21#_c_76_n 0.0286882f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_3 VNB N_A_79_21#_c_77_n 0.00127487f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_4 VNB N_A_79_21#_c_78_n 0.0158219f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=0.74
cc_5 VNB N_A_79_21#_c_79_n 0.00504946f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=1.955
cc_6 VNB N_S_M1000_g 0.0320387f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_7 VNB N_S_M1008_g 0.0525446f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_8 VNB N_S_c_147_n 0.00360945f $X=-0.19 $Y=-0.24 $X2=2.535 $Y2=2.04
cc_9 VNB N_S_c_148_n 0.0248526f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_A1_M1004_g 0.0221567f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A1_c_237_n 0.00411936f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_12 VNB N_A1_c_238_n 0.0454385f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_13 VNB A1 0.0150165f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A0_M1007_g 0.0252073f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_15 VNB N_A0_c_299_n 0.0124763f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_16 VNB N_A0_c_300_n 0.0348785f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_17 VNB N_A0_c_301_n 0.00979231f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_18 VNB N_A_657_21#_M1001_g 0.0244915f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_19 VNB N_A_657_21#_c_346_n 0.0129448f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_20 VNB N_A_657_21#_c_347_n 0.00985669f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=1.16
cc_21 VNB N_A_657_21#_c_348_n 0.0280367f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=0.74
cc_22 VNB N_A_657_21#_c_349_n 0.0251039f $X=-0.19 $Y=-0.24 $X2=2.535 $Y2=2.04
cc_23 VNB N_A_657_21#_c_350_n 0.0137474f $X=-0.19 $Y=-0.24 $X2=1.525 $Y2=0.54
cc_24 VNB N_A_657_21#_c_351_n 0.0248547f $X=-0.19 $Y=-0.24 $X2=1.87 $Y2=0.54
cc_25 VNB X 0.045502f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.985
cc_26 VNB N_VPWR_c_410_n 0.193827f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_452_n 0.00309635f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.56
cc_28 VNB N_VGND_c_453_n 0.00465782f $X=-0.19 $Y=-0.24 $X2=0.6 $Y2=0.825
cc_29 VNB N_VGND_c_454_n 0.0151047f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB N_VGND_c_455_n 0.0614079f $X=-0.19 $Y=-0.24 $X2=1.61 $Y2=2.04
cc_31 VNB N_VGND_c_456_n 0.0265797f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_457_n 0.247995f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_458_n 0.00603371f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_459_n 0.00772189f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VPB N_A_79_21#_c_76_n 0.0340517f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_36 VPB N_A_79_21#_c_77_n 0.0024294f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_37 VPB N_A_79_21#_c_79_n 0.0108875f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.955
cc_38 VPB N_S_c_149_n 0.0268063f $X=-0.19 $Y=1.305 $X2=1.81 $Y2=1.87
cc_39 VPB N_S_c_150_n 0.0246517f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_40 VPB N_S_c_151_n 0.0612273f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_41 VPB N_S_M1008_g 0.0045419f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_42 VPB N_S_c_153_n 0.00442737f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=0.74
cc_43 VPB N_S_c_154_n 0.0427435f $X=-0.19 $Y=1.305 $X2=0.685 $Y2=0.74
cc_44 VPB N_S_c_155_n 0.00182422f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.825
cc_45 VPB N_S_c_156_n 0.00278937f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.955
cc_46 VPB N_S_c_157_n 0.00173472f $X=-0.19 $Y=1.305 $X2=1.61 $Y2=2.04
cc_47 VPB N_S_c_147_n 0.00126685f $X=-0.19 $Y=1.305 $X2=2.535 $Y2=2.04
cc_48 VPB N_S_c_148_n 0.00492931f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_49 VPB S 0.00986479f $X=-0.19 $Y=1.305 $X2=0.565 $Y2=1.16
cc_50 VPB N_A1_c_240_n 0.0545586f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A1_c_237_n 0.00640998f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_52 VPB N_A1_c_242_n 0.0218398f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.825
cc_53 VPB N_A1_c_243_n 2.25457e-19 $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_54 VPB A1 0.00130976f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB N_A0_c_302_n 0.0204961f $X=-0.19 $Y=1.305 $X2=1.735 $Y2=0.235
cc_56 VPB N_A0_c_303_n 0.0445243f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_A0_c_304_n 0.0118266f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_A0_c_299_n 0.0231504f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_59 VPB N_A0_c_301_n 0.00328657f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.16
cc_60 VPB N_A_657_21#_c_346_n 0.0192975f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_61 VPB N_A_657_21#_c_353_n 0.0215405f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.825
cc_62 VPB N_A_657_21#_c_350_n 0.0324779f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.54
cc_63 VPB N_A_657_21#_c_355_n 0.0215259f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_X_c_395_n 0.0065071f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_65 VPB X 0.00942252f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_66 VPB X 0.0315701f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=0.825
cc_67 VPB N_VPWR_c_411_n 0.00474148f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.985
cc_68 VPB N_VPWR_c_412_n 0.0109087f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_413_n 0.0660484f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=0.825
cc_70 VPB N_VPWR_c_414_n 0.00324402f $X=-0.19 $Y=1.305 $X2=1.525 $Y2=1.955
cc_71 VPB N_VPWR_c_415_n 0.0259916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_410_n 0.0887972f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_417_n 0.0226539f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 N_A_79_21#_c_76_n N_S_c_149_n 0.00709235f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_75 N_A_79_21#_c_79_n N_S_c_150_n 4.89657e-19 $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_76 N_A_79_21#_c_85_p N_S_c_150_n 6.54365e-19 $X=1.61 $Y=2.04 $X2=0 $Y2=0
cc_77 N_A_79_21#_c_75_n N_S_M1000_g 0.013677f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_78 N_A_79_21#_c_77_n N_S_M1000_g 0.00297788f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_79 N_A_79_21#_c_78_n N_S_M1000_g 0.0133748f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_80 N_A_79_21#_c_79_n N_S_M1000_g 0.00343808f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_81 N_A_79_21#_c_90_p N_S_M1000_g 0.00670281f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_82 N_A_79_21#_c_76_n N_S_c_153_n 0.0011476f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_79_21#_c_85_p N_S_c_154_n 0.0116702f $X=1.61 $Y=2.04 $X2=0 $Y2=0
cc_84 N_A_79_21#_c_93_p N_S_c_154_n 0.0759798f $X=2.535 $Y=2.04 $X2=0 $Y2=0
cc_85 N_A_79_21#_c_76_n N_S_c_147_n 0.00110986f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_86 N_A_79_21#_c_77_n N_S_c_147_n 0.014361f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_87 N_A_79_21#_c_78_n N_S_c_147_n 0.0211311f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_88 N_A_79_21#_c_79_n N_S_c_147_n 0.0703039f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_89 N_A_79_21#_c_76_n N_S_c_148_n 0.0202694f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_79_21#_c_77_n N_S_c_148_n 0.00107569f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_91 N_A_79_21#_c_78_n N_S_c_148_n 0.00246808f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_92 N_A_79_21#_c_79_n N_S_c_148_n 0.00405008f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_93 N_A_79_21#_c_90_p N_A1_M1004_g 0.0269722f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_94 N_A_79_21#_c_93_p N_A1_c_240_n 0.00448094f $X=2.535 $Y=2.04 $X2=0 $Y2=0
cc_95 N_A_79_21#_c_79_n N_A1_c_237_n 0.0570095f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_96 N_A_79_21#_c_90_p N_A1_c_237_n 0.0124631f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_97 N_A_79_21#_c_79_n N_A1_c_238_n 0.00856035f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_98 N_A_79_21#_c_90_p N_A1_c_238_n 0.00174897f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_99 N_A_79_21#_c_93_p N_A1_c_242_n 0.0568676f $X=2.535 $Y=2.04 $X2=0 $Y2=0
cc_100 N_A_79_21#_c_79_n N_A1_c_243_n 0.0137204f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_101 N_A_79_21#_c_93_p N_A1_c_243_n 0.0111679f $X=2.535 $Y=2.04 $X2=0 $Y2=0
cc_102 N_A_79_21#_c_79_n N_A0_c_302_n 0.00256066f $X=1.525 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_103 N_A_79_21#_c_93_p N_A0_c_302_n 0.0176382f $X=2.535 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_104 N_A_79_21#_c_93_p N_A0_c_303_n 0.0155064f $X=2.535 $Y=2.04 $X2=0 $Y2=0
cc_105 N_A_79_21#_c_79_n N_A0_c_304_n 0.00196313f $X=1.525 $Y=1.955 $X2=0 $Y2=0
cc_106 N_A_79_21#_c_90_p N_A0_M1007_g 0.00161075f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_107 N_A_79_21#_c_76_n N_X_c_395_n 0.00292963f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_108 N_A_79_21#_c_75_n X 0.0193288f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_109 N_A_79_21#_c_76_n X 0.00327243f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_79_21#_c_77_n X 0.0344429f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_111 N_A_79_21#_c_76_n X 0.00976225f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_112 N_A_79_21#_c_76_n N_VPWR_c_411_n 0.009924f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_79_21#_c_77_n N_VPWR_c_411_n 0.00331775f $X=0.6 $Y=1.16 $X2=0 $Y2=0
cc_114 N_A_79_21#_c_78_n N_VPWR_c_411_n 0.00369736f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_115 N_A_79_21#_c_76_n N_VPWR_c_410_n 0.0140376f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_116 N_A_79_21#_c_76_n N_VPWR_c_417_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_79_21#_c_79_n A_243_374# 7.59015e-19 $X=1.525 $Y=1.955 $X2=-0.19
+ $Y2=-0.24
cc_118 N_A_79_21#_c_85_p A_243_374# 0.00300196f $X=1.61 $Y=2.04 $X2=-0.19
+ $Y2=-0.24
cc_119 N_A_79_21#_c_77_n N_VGND_M1010_d 8.23133e-19 $X=0.6 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_120 N_A_79_21#_c_78_n N_VGND_M1010_d 0.00683237f $X=1.435 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_121 N_A_79_21#_c_130_p N_VGND_M1010_d 8.75693e-19 $X=0.685 $Y=0.74 $X2=-0.19
+ $Y2=-0.24
cc_122 N_A_79_21#_c_75_n N_VGND_c_452_n 0.00910743f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_123 N_A_79_21#_c_76_n N_VGND_c_452_n 5.28725e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_79_21#_c_78_n N_VGND_c_452_n 0.0160584f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_125 N_A_79_21#_c_130_p N_VGND_c_452_n 0.00929542f $X=0.685 $Y=0.74 $X2=0
+ $Y2=0
cc_126 N_A_79_21#_c_90_p N_VGND_c_452_n 0.00815458f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_127 N_A_79_21#_c_75_n N_VGND_c_454_n 0.0046653f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_128 N_A_79_21#_c_78_n N_VGND_c_455_n 0.00916117f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_129 N_A_79_21#_c_90_p N_VGND_c_455_n 0.0313996f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_130 N_A_79_21#_M1004_d N_VGND_c_457_n 0.015588f $X=1.735 $Y=0.235 $X2=0 $Y2=0
cc_131 N_A_79_21#_c_75_n N_VGND_c_457_n 0.00895857f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_132 N_A_79_21#_c_78_n N_VGND_c_457_n 0.0152428f $X=1.435 $Y=0.74 $X2=0 $Y2=0
cc_133 N_A_79_21#_c_130_p N_VGND_c_457_n 8.0899e-19 $X=0.685 $Y=0.74 $X2=0 $Y2=0
cc_134 N_A_79_21#_c_90_p N_VGND_c_457_n 0.0191349f $X=1.525 $Y=0.54 $X2=0 $Y2=0
cc_135 N_A_79_21#_c_90_p A_245_47# 0.00646653f $X=1.525 $Y=0.54 $X2=-0.19
+ $Y2=-0.24
cc_136 N_S_M1000_g N_A1_M1004_g 0.0162658f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_137 N_S_c_154_n N_A1_c_240_n 0.0142103f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_138 N_S_c_156_n N_A1_c_240_n 0.00110572f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_139 N_S_c_157_n N_A1_c_240_n 0.00339969f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_140 N_S_c_147_n N_A1_c_238_n 3.855e-19 $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_141 N_S_c_148_n N_A1_c_238_n 0.0162658f $X=1.08 $Y=1.16 $X2=0 $Y2=0
cc_142 N_S_c_154_n N_A1_c_242_n 0.0106963f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_143 N_S_c_156_n N_A1_c_242_n 0.00133732f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_144 N_S_c_157_n N_A1_c_242_n 0.0123492f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_145 N_S_c_156_n A1 0.0143252f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_146 N_S_c_150_n N_A0_c_302_n 0.0156044f $X=1.125 $Y=1.795 $X2=-0.19 $Y2=-0.24
cc_147 N_S_c_153_n N_A0_c_302_n 7.57284e-19 $X=1.17 $Y=2.295 $X2=-0.19 $Y2=-0.24
cc_148 N_S_c_154_n N_A0_c_302_n 0.0121952f $X=3.245 $Y=2.38 $X2=-0.19 $Y2=-0.24
cc_149 N_S_c_149_n N_A0_c_304_n 0.00408375f $X=1.125 $Y=1.695 $X2=0 $Y2=0
cc_150 N_S_M1008_g N_A_657_21#_M1001_g 0.0147771f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_151 N_S_c_151_n N_A_657_21#_c_346_n 0.02165f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_152 N_S_M1008_g N_A_657_21#_c_346_n 0.0104002f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_153 N_S_c_156_n N_A_657_21#_c_346_n 0.00571499f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_154 N_S_c_157_n N_A_657_21#_c_346_n 0.00174484f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_155 S N_A_657_21#_c_346_n 0.00741113f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_156 N_S_c_151_n N_A_657_21#_c_353_n 0.0109261f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_157 N_S_c_154_n N_A_657_21#_c_353_n 0.0052034f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_158 N_S_c_157_n N_A_657_21#_c_353_n 0.0141277f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_159 N_S_c_151_n N_A_657_21#_c_347_n 0.00366753f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_160 N_S_M1008_g N_A_657_21#_c_347_n 0.0177096f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_161 N_S_c_156_n N_A_657_21#_c_347_n 0.00522993f $X=3.33 $Y=1.63 $X2=0 $Y2=0
cc_162 S N_A_657_21#_c_347_n 0.0243329f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_163 N_S_M1008_g N_A_657_21#_c_348_n 0.0144241f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_164 S N_A_657_21#_c_348_n 0.00257432f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_165 N_S_M1008_g N_A_657_21#_c_349_n 0.0101674f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_166 N_S_c_151_n N_A_657_21#_c_350_n 0.0102106f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_167 N_S_M1008_g N_A_657_21#_c_350_n 0.0134138f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_168 S N_A_657_21#_c_350_n 0.0164556f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_169 S N_A_657_21#_c_351_n 4.91502e-19 $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_170 N_S_c_149_n N_VPWR_c_411_n 0.00234447f $X=1.125 $Y=1.695 $X2=0 $Y2=0
cc_171 N_S_c_150_n N_VPWR_c_411_n 0.00478183f $X=1.125 $Y=1.795 $X2=0 $Y2=0
cc_172 N_S_c_153_n N_VPWR_c_411_n 0.0415786f $X=1.17 $Y=2.295 $X2=0 $Y2=0
cc_173 N_S_c_155_n N_VPWR_c_411_n 0.00997526f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_174 N_S_c_151_n N_VPWR_c_412_n 0.00679996f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_175 N_S_c_154_n N_VPWR_c_412_n 0.0137895f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_176 N_S_c_157_n N_VPWR_c_412_n 0.0294586f $X=3.33 $Y=2.295 $X2=0 $Y2=0
cc_177 S N_VPWR_c_412_n 0.010519f $X=3.805 $Y=1.445 $X2=0 $Y2=0
cc_178 N_S_c_150_n N_VPWR_c_413_n 0.00206875f $X=1.125 $Y=1.795 $X2=0 $Y2=0
cc_179 N_S_c_154_n N_VPWR_c_413_n 0.139371f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_180 N_S_c_155_n N_VPWR_c_413_n 0.0143028f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_181 N_S_c_151_n N_VPWR_c_415_n 0.00641313f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_182 N_S_c_150_n N_VPWR_c_410_n 0.00122187f $X=1.125 $Y=1.795 $X2=0 $Y2=0
cc_183 N_S_c_151_n N_VPWR_c_410_n 0.0062839f $X=3.915 $Y=1.795 $X2=0 $Y2=0
cc_184 N_S_c_154_n N_VPWR_c_410_n 0.0800988f $X=3.245 $Y=2.38 $X2=0 $Y2=0
cc_185 N_S_c_155_n N_VPWR_c_410_n 0.00769712f $X=1.27 $Y=2.38 $X2=0 $Y2=0
cc_186 N_S_M1000_g N_VGND_c_452_n 0.00593008f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_187 N_S_M1008_g N_VGND_c_453_n 0.0059679f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_188 N_S_M1000_g N_VGND_c_455_n 0.00428022f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_189 N_S_M1008_g N_VGND_c_456_n 0.00585385f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_190 N_S_M1000_g N_VGND_c_457_n 0.00672742f $X=1.15 $Y=0.445 $X2=0 $Y2=0
cc_191 N_S_M1008_g N_VGND_c_457_n 0.0123317f $X=3.94 $Y=0.445 $X2=0 $Y2=0
cc_192 N_A1_c_240_n N_A0_c_303_n 0.00326777f $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_193 N_A1_c_242_n N_A0_c_303_n 0.0179077f $X=2.855 $Y=1.7 $X2=0 $Y2=0
cc_194 N_A1_c_243_n N_A0_c_303_n 0.00497621f $X=1.95 $Y=1.7 $X2=0 $Y2=0
cc_195 N_A1_c_238_n N_A0_c_304_n 0.0102357f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_196 N_A1_c_243_n N_A0_c_304_n 0.00262213f $X=1.95 $Y=1.7 $X2=0 $Y2=0
cc_197 N_A1_M1004_g N_A0_M1007_g 0.00777686f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_198 A1 N_A0_M1007_g 0.00294405f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_199 N_A1_c_240_n N_A0_c_299_n 0.016746f $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_200 N_A1_c_237_n N_A0_c_299_n 0.00704662f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_201 N_A1_c_242_n N_A0_c_299_n 0.00445205f $X=2.855 $Y=1.7 $X2=0 $Y2=0
cc_202 A1 N_A0_c_299_n 0.00257547f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_203 N_A1_c_237_n N_A0_c_300_n 3.66295e-19 $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_204 N_A1_c_238_n N_A0_c_300_n 0.0111748f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_205 N_A1_c_242_n N_A0_c_300_n 0.00166378f $X=2.855 $Y=1.7 $X2=0 $Y2=0
cc_206 A1 N_A0_c_300_n 0.00347787f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_207 N_A1_M1004_g N_A0_c_301_n 0.00268799f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_208 N_A1_c_240_n N_A0_c_301_n 2.37679e-19 $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_209 N_A1_c_237_n N_A0_c_301_n 0.0281261f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_210 N_A1_c_238_n N_A0_c_301_n 0.00258381f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_211 N_A1_c_242_n N_A0_c_301_n 0.0226282f $X=2.855 $Y=1.7 $X2=0 $Y2=0
cc_212 A1 N_A0_c_301_n 0.0707809f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_213 A1 N_A_657_21#_M1001_g 0.0109694f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_214 N_A1_c_240_n N_A_657_21#_c_346_n 0.026158f $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_215 A1 N_A_657_21#_c_346_n 6.15513e-19 $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_216 N_A1_c_240_n N_A_657_21#_c_353_n 0.0337616f $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_217 A1 N_A_657_21#_c_347_n 0.0116592f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_218 A1 N_A_657_21#_c_348_n 0.0108957f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_219 N_A1_c_240_n N_VPWR_c_413_n 0.00102161f $X=2.975 $Y=1.795 $X2=0 $Y2=0
cc_220 N_A1_M1004_g N_VGND_c_455_n 0.00357668f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_221 A1 N_VGND_c_455_n 0.0153299f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_222 N_A1_M1004_g N_VGND_c_457_n 0.00618492f $X=1.66 $Y=0.445 $X2=0 $Y2=0
cc_223 N_A1_c_238_n N_VGND_c_457_n 0.00102921f $X=1.865 $Y=0.98 $X2=0 $Y2=0
cc_224 A1 N_VGND_c_457_n 0.00839556f $X=2.895 $Y=0.765 $X2=0 $Y2=0
cc_225 A1 A_499_47# 0.0147234f $X=2.895 $Y=0.765 $X2=-0.19 $Y2=-0.24
cc_226 N_A0_c_300_n N_A_657_21#_M1001_g 0.00397499f $X=2.48 $Y=0.98 $X2=0 $Y2=0
cc_227 N_A0_c_302_n N_VPWR_c_413_n 0.00102161f $X=1.72 $Y=1.795 $X2=0 $Y2=0
cc_228 N_A0_M1007_g N_VGND_c_455_n 0.00357668f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_229 N_A0_c_301_n N_VGND_c_455_n 0.0185253f $X=2.48 $Y=0.98 $X2=0 $Y2=0
cc_230 N_A0_M1007_g N_VGND_c_457_n 0.00732049f $X=2.42 $Y=0.445 $X2=0 $Y2=0
cc_231 N_A0_c_300_n N_VGND_c_457_n 0.00116644f $X=2.48 $Y=0.98 $X2=0 $Y2=0
cc_232 N_A0_c_301_n N_VGND_c_457_n 0.0117533f $X=2.48 $Y=0.98 $X2=0 $Y2=0
cc_233 N_A0_c_301_n A_499_47# 0.00527918f $X=2.48 $Y=0.98 $X2=-0.19 $Y2=-0.24
cc_234 N_A_657_21#_c_353_n N_VPWR_c_412_n 0.00223023f $X=3.385 $Y=1.795 $X2=0
+ $Y2=0
cc_235 N_A_657_21#_c_353_n N_VPWR_c_413_n 0.00281778f $X=3.385 $Y=1.795 $X2=0
+ $Y2=0
cc_236 N_A_657_21#_c_355_n N_VPWR_c_415_n 0.0141376f $X=4.357 $Y=2.08 $X2=0
+ $Y2=0
cc_237 N_A_657_21#_c_353_n N_VPWR_c_410_n 0.00209463f $X=3.385 $Y=1.795 $X2=0
+ $Y2=0
cc_238 N_A_657_21#_c_355_n N_VPWR_c_410_n 0.0156259f $X=4.357 $Y=2.08 $X2=0
+ $Y2=0
cc_239 N_A_657_21#_M1001_g N_VGND_c_453_n 0.0275028f $X=3.36 $Y=0.445 $X2=0
+ $Y2=0
cc_240 N_A_657_21#_c_347_n N_VGND_c_453_n 0.0245813f $X=4.035 $Y=0.98 $X2=0
+ $Y2=0
cc_241 N_A_657_21#_c_348_n N_VGND_c_453_n 0.00403031f $X=3.45 $Y=0.98 $X2=0
+ $Y2=0
cc_242 N_A_657_21#_c_349_n N_VGND_c_456_n 0.0129431f $X=4.15 $Y=0.455 $X2=0
+ $Y2=0
cc_243 N_A_657_21#_M1008_d N_VGND_c_457_n 0.0028471f $X=4.015 $Y=0.235 $X2=0
+ $Y2=0
cc_244 N_A_657_21#_c_349_n N_VGND_c_457_n 0.00919761f $X=4.15 $Y=0.455 $X2=0
+ $Y2=0
cc_245 N_X_c_395_n N_VPWR_c_411_n 0.0587634f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_246 N_X_M1005_s N_VPWR_c_410_n 0.00217517f $X=0.135 $Y=1.485 $X2=0 $Y2=0
cc_247 X N_VPWR_c_410_n 0.0126651f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_248 X N_VPWR_c_417_n 0.021418f $X=0.15 $Y=1.785 $X2=0 $Y2=0
cc_249 X N_VGND_c_454_n 0.0176426f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_250 N_X_M1010_s N_VGND_c_457_n 0.00387172f $X=0.135 $Y=0.235 $X2=0 $Y2=0
cc_251 X N_VGND_c_457_n 0.00974347f $X=0.15 $Y=0.425 $X2=0 $Y2=0
cc_252 N_VGND_c_457_n A_245_47# 0.00371776f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
cc_253 N_VGND_c_457_n A_499_47# 0.0194586f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
