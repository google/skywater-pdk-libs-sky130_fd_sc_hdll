* File: sky130_fd_sc_hdll__buf_2.spice
* Created: Wed Sep  2 08:24:16 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__buf_2.pex.spice"
.subckt sky130_fd_sc_hdll__buf_2  VNB VPB A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_M1000_g N_A_27_47#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1302 PD=0.765421 PS=1.46 NRD=11.424 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75001.4 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_47#_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.154375 AS=0.11785 PD=1.125 PS=1.18458 NRD=26.76 NRS=0.912 M=1 R=4.33333
+ SA=75000.5 SB=75000.9 A=0.0975 P=1.6 MULT=1
MM1005 N_X_M1001_d N_A_27_47#_M1005_g N_VGND_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.154375 AS=0.25025 PD=1.125 PS=2.07 NRD=9.228 NRS=21.228 M=1 R=4.33333
+ SA=75001.1 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1002 N_VPWR_M1002_d N_A_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.64
+ AD=0.122693 AS=0.1728 PD=1.04976 PS=1.82 NRD=12.2928 NRS=1.5366 M=1 R=3.55556
+ SA=90000.2 SB=90001.4 A=0.1152 P=1.64 MULT=1
MM1003 N_X_M1003_d N_A_27_47#_M1003_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1975 AS=0.191707 PD=1.395 PS=1.64024 NRD=20.685 NRS=4.9053 M=1 R=5.55556
+ SA=90000.5 SB=90000.9 A=0.18 P=2.36 MULT=1
MM1004 N_X_M1003_d N_A_27_47#_M1004_g N_VPWR_M1004_s VPB PHIGHVT L=0.18 W=1
+ AD=0.1975 AS=0.395 PD=1.395 PS=2.79 NRD=1.9503 NRS=24.6053 M=1 R=5.55556
+ SA=90001.1 SB=90000.3 A=0.18 P=2.36 MULT=1
DX6_noxref VNB VPB NWDIODE A=4.3014 P=8.57
*
.include "sky130_fd_sc_hdll__buf_2.pxi.spice"
*
.ends
*
*
