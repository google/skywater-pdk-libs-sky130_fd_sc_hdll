# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__nand3_2
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__nand3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.140000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.995000 0.330000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.170000 1.075000 2.615000 1.275000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.555000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.785000 1.075000 4.000000 1.275000 ;
    END
  END C
  PIN Y
    ANTENNADIFFAREA  1.078000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.515000 0.635000 0.895000 1.445000 ;
        RECT 0.515000 1.445000 3.295000 1.665000 ;
        RECT 0.515000 1.665000 0.895000 2.465000 ;
        RECT 1.455000 1.665000 1.835000 2.465000 ;
        RECT 2.915000 1.665000 3.295000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 4.330000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.090000  0.295000 2.305000 0.465000 ;
      RECT 0.090000  0.465000 0.345000 0.785000 ;
      RECT 0.090000  1.495000 0.345000 2.635000 ;
      RECT 1.115000  1.835000 1.285000 2.635000 ;
      RECT 1.455000  0.635000 3.295000 0.905000 ;
      RECT 2.055000  1.835000 2.745000 2.635000 ;
      RECT 2.495000  0.085000 2.825000 0.465000 ;
      RECT 3.515000  0.085000 3.895000 0.885000 ;
      RECT 3.515000  1.445000 3.895000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__nand3_2
END LIBRARY
