* File: sky130_fd_sc_hdll__a21boi_1.spice
* Created: Wed Sep  2 08:16:45 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21boi_1.pex.spice"
.subckt sky130_fd_sc_hdll__a21boi_1  VNB VPB B1_N A1 A2 VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A2	A2
* A1	A1
* B1_N	B1_N
* VPB	VPB
* VNB	VNB
MM1002 N_VGND_M1002_d N_B1_N_M1002_g N_A_27_413#_M1002_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0927336 AS=0.1533 PD=0.816449 PS=1.57 NRD=17.856 NRS=28.56 M=1
+ R=2.8 SA=75000.3 SB=75002 A=0.063 P=1.14 MULT=1
MM1005 N_Y_M1005_d N_A_27_413#_M1005_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.1755 AS=0.143516 PD=1.19 PS=1.26355 NRD=9.228 NRS=9.228 M=1 R=4.33333
+ SA=75000.6 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1003 A_434_47# N_A1_M1003_g N_Y_M1005_d VNB NSHORT L=0.15 W=0.65 AD=0.13325
+ AS=0.1755 PD=1.06 PS=1.19 NRD=27.684 NRS=38.76 M=1 R=4.33333 SA=75001.3
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_434_47# VNB NSHORT L=0.15 W=0.65 AD=0.19825
+ AS=0.13325 PD=1.91 PS=1.06 NRD=7.38 NRS=27.684 M=1 R=4.33333 SA=75001.9
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VPWR_M1000_d N_B1_N_M1000_g N_A_27_413#_M1000_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1155 AS=0.1155 PD=1.39 PS=1.39 NRD=4.6886 NRS=4.6886 M=1 R=2.33333
+ SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1007 N_A_338_297#_M1007_d N_A_27_413#_M1007_g N_Y_M1007_s VPB PHIGHVT L=0.18
+ W=1 AD=0.15 AS=0.325 PD=1.3 PS=2.65 NRD=1.9503 NRS=11.8003 M=1 R=5.55556
+ SA=90000.2 SB=90001.3 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A1_M1001_g N_A_338_297#_M1007_d VPB PHIGHVT L=0.18 W=1
+ AD=0.21 AS=0.15 PD=1.42 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90000.7
+ SB=90000.8 A=0.18 P=2.36 MULT=1
MM1006 N_A_338_297#_M1006_d N_A2_M1006_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.21 PD=2.55 PS=1.42 NRD=1.9503 NRS=25.5903 M=1 R=5.55556
+ SA=90001.3 SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hdll__a21boi_1.pxi.spice"
*
.ends
*
*
