* File: sky130_fd_sc_hdll__diode_8.pxi.spice
* Created: Thu Aug 27 19:05:25 2020
* 
x_PM_SKY130_FD_SC_HDLL__DIODE_8%DIODE N_DIODE_D0_noxref_neg DIODE DIODE
+ N_DIODE_c_8_n PM_SKY130_FD_SC_HDLL__DIODE_8%DIODE
x_PM_SKY130_FD_SC_HDLL__DIODE_8%VGND VGND N_VGND_c_15_n N_VGND_c_16_n
+ PM_SKY130_FD_SC_HDLL__DIODE_8%VGND
x_PM_SKY130_FD_SC_HDLL__DIODE_8%VPWR VPWR N_VPWR_c_21_n N_VPWR_c_20_n
+ PM_SKY130_FD_SC_HDLL__DIODE_8%VPWR
cc_1 VNB N_DIODE_c_8_n 0.166226f $X=-0.19 $Y=-0.24 $X2=3.37 $Y2=0.37
cc_2 VNB N_VGND_c_15_n 0.0884987f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_3 VNB N_VGND_c_16_n 0.20018f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_4 VNB N_VPWR_c_20_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_5 VPB N_DIODE_c_8_n 0.203133f $X=-0.19 $Y=1.305 $X2=3.37 $Y2=0.37
cc_6 VPB N_VPWR_c_21_n 0.0884987f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_7 VPB N_VPWR_c_20_n 0.0720925f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_8 N_DIODE_c_8_n N_VGND_c_15_n 0.245391f $X=3.37 $Y=0.37 $X2=0 $Y2=0
cc_9 N_DIODE_D0_noxref_neg N_VGND_c_16_n 0.0325442f $X=0.135 $Y=0.195 $X2=0
+ $Y2=0
cc_10 N_DIODE_c_8_n N_VGND_c_16_n 0.135113f $X=3.37 $Y=0.37 $X2=0 $Y2=0
cc_11 N_DIODE_c_8_n N_VPWR_c_21_n 0.250074f $X=3.37 $Y=0.37 $X2=0 $Y2=0
cc_12 N_DIODE_c_8_n N_VPWR_c_20_n 0.135113f $X=3.37 $Y=0.37 $X2=0 $Y2=0
