* File: sky130_fd_sc_hdll__buf_8.pxi.spice
* Created: Thu Aug 27 19:00:43 2020
* 
x_PM_SKY130_FD_SC_HDLL__BUF_8%A N_A_c_103_n N_A_M1001_g N_A_M1002_g N_A_c_104_n
+ N_A_M1008_g N_A_M1015_g N_A_c_105_n N_A_M1019_g N_A_M1021_g A A A N_A_c_102_n
+ A A PM_SKY130_FD_SC_HDLL__BUF_8%A
x_PM_SKY130_FD_SC_HDLL__BUF_8%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1015_d
+ N_A_27_47#_M1001_d N_A_27_47#_M1008_d N_A_27_47#_M1004_g N_A_27_47#_c_183_n
+ N_A_27_47#_M1000_g N_A_27_47#_M1005_g N_A_27_47#_c_184_n N_A_27_47#_M1003_g
+ N_A_27_47#_M1009_g N_A_27_47#_c_185_n N_A_27_47#_M1006_g N_A_27_47#_M1011_g
+ N_A_27_47#_c_186_n N_A_27_47#_M1007_g N_A_27_47#_M1014_g N_A_27_47#_c_187_n
+ N_A_27_47#_M1010_g N_A_27_47#_M1017_g N_A_27_47#_c_188_n N_A_27_47#_M1012_g
+ N_A_27_47#_M1018_g N_A_27_47#_c_189_n N_A_27_47#_M1013_g N_A_27_47#_c_190_n
+ N_A_27_47#_M1016_g N_A_27_47#_M1020_g N_A_27_47#_c_191_n N_A_27_47#_c_202_n
+ N_A_27_47#_c_174_n N_A_27_47#_c_175_n N_A_27_47#_c_192_n N_A_27_47#_c_193_n
+ N_A_27_47#_c_216_n N_A_27_47#_c_219_n N_A_27_47#_c_176_n N_A_27_47#_c_194_n
+ N_A_27_47#_c_177_n N_A_27_47#_c_178_n N_A_27_47#_c_179_n N_A_27_47#_c_196_n
+ N_A_27_47#_c_180_n N_A_27_47#_c_181_n N_A_27_47#_c_182_n
+ PM_SKY130_FD_SC_HDLL__BUF_8%A_27_47#
x_PM_SKY130_FD_SC_HDLL__BUF_8%VPWR N_VPWR_M1001_s N_VPWR_M1019_s N_VPWR_M1003_s
+ N_VPWR_M1007_s N_VPWR_M1012_s N_VPWR_M1016_s N_VPWR_c_396_n N_VPWR_c_397_n
+ N_VPWR_c_398_n N_VPWR_c_399_n N_VPWR_c_400_n N_VPWR_c_401_n N_VPWR_c_402_n
+ N_VPWR_c_403_n VPWR VPWR N_VPWR_c_404_n N_VPWR_c_405_n N_VPWR_c_406_n
+ N_VPWR_c_407_n N_VPWR_c_395_n N_VPWR_c_409_n N_VPWR_c_410_n N_VPWR_c_411_n
+ N_VPWR_c_412_n N_VPWR_c_413_n N_VPWR_c_414_n N_VPWR_c_415_n
+ PM_SKY130_FD_SC_HDLL__BUF_8%VPWR
x_PM_SKY130_FD_SC_HDLL__BUF_8%X N_X_M1004_d N_X_M1009_d N_X_M1014_d N_X_M1018_d
+ N_X_M1000_d N_X_M1006_d N_X_M1010_d N_X_M1013_d N_X_c_513_n N_X_c_514_n
+ N_X_c_498_n N_X_c_499_n N_X_c_505_n N_X_c_506_n N_X_c_532_n N_X_c_533_n
+ N_X_c_500_n N_X_c_507_n N_X_c_543_n N_X_c_544_n N_X_c_501_n N_X_c_508_n
+ N_X_c_554_n N_X_c_502_n N_X_c_509_n N_X_c_503_n N_X_c_510_n X X X N_X_c_573_n
+ PM_SKY130_FD_SC_HDLL__BUF_8%X
x_PM_SKY130_FD_SC_HDLL__BUF_8%VGND N_VGND_M1002_s N_VGND_M1021_s N_VGND_M1005_s
+ N_VGND_M1011_s N_VGND_M1017_s N_VGND_M1020_s N_VGND_c_637_n N_VGND_c_638_n
+ N_VGND_c_639_n N_VGND_c_640_n N_VGND_c_641_n N_VGND_c_642_n N_VGND_c_643_n
+ VGND VGND N_VGND_c_644_n VGND N_VGND_c_645_n N_VGND_c_646_n N_VGND_c_647_n
+ N_VGND_c_648_n N_VGND_c_649_n N_VGND_c_650_n N_VGND_c_651_n N_VGND_c_652_n
+ N_VGND_c_653_n N_VGND_c_654_n N_VGND_c_655_n N_VGND_c_656_n
+ PM_SKY130_FD_SC_HDLL__BUF_8%VGND
cc_1 VNB N_A_M1002_g 0.0231077f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.56
cc_2 VNB N_A_M1015_g 0.0183641f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_3 VNB N_A_M1021_g 0.0175026f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=0.56
cc_4 VNB A 0.00806404f $X=-0.19 $Y=-0.24 $X2=1.065 $Y2=1.105
cc_5 VNB N_A_c_102_n 0.0861762f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.212
cc_6 VNB N_A_27_47#_M1004_g 0.0180221f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.41
cc_7 VNB N_A_27_47#_M1005_g 0.0181352f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_47#_M1009_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_9 VNB N_A_27_47#_M1011_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_10 VNB N_A_27_47#_M1014_g 0.0181597f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.175
cc_11 VNB N_A_27_47#_M1017_g 0.0181268f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_A_27_47#_M1018_g 0.0181187f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB N_A_27_47#_M1020_g 0.0241264f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_A_27_47#_c_174_n 0.00350914f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_A_27_47#_c_175_n 0.00185814f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_A_27_47#_c_176_n 0.00166201f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_A_27_47#_c_177_n 0.00305801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_A_27_47#_c_178_n 0.00103736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_A_27_47#_c_179_n 0.00274061f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_180_n 0.00114159f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_21 VNB N_A_27_47#_c_181_n 0.00142427f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_A_27_47#_c_182_n 0.199381f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_23 VNB N_VPWR_c_395_n 0.250759f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_X_c_498_n 0.00380791f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.212
cc_25 VNB N_X_c_499_n 0.00129721f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.212
cc_26 VNB N_X_c_500_n 0.00380791f $X=-0.19 $Y=-0.24 $X2=0.695 $Y2=1.19
cc_27 VNB N_X_c_501_n 0.00337105f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_X_c_502_n 0.00114174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VNB N_X_c_503_n 0.00114174f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_30 VNB X 0.00151968f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_637_n 0.00214417f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_638_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_639_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0.305 $Y2=1.16
cc_34 VNB N_VGND_c_640_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.212
cc_35 VNB N_VGND_c_641_n 3.19622e-19 $X=-0.19 $Y=-0.24 $X2=1.035 $Y2=1.16
cc_36 VNB N_VGND_c_642_n 0.0132714f $X=-0.19 $Y=-0.24 $X2=1.46 $Y2=1.212
cc_37 VNB N_VGND_c_643_n 0.0321553f $X=-0.19 $Y=-0.24 $X2=0.685 $Y2=1.175
cc_38 VNB N_VGND_c_644_n 0.0152765f $X=-0.19 $Y=-0.24 $X2=1.15 $Y2=1.175
cc_39 VNB N_VGND_c_645_n 0.013707f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_40 VNB N_VGND_c_646_n 0.0134547f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_41 VNB N_VGND_c_647_n 0.0126449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_42 VNB N_VGND_c_648_n 0.0126449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_43 VNB N_VGND_c_649_n 0.0143948f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_44 VNB N_VGND_c_650_n 0.308638f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_45 VNB N_VGND_c_651_n 0.00574292f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_46 VNB N_VGND_c_652_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_47 VNB N_VGND_c_653_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_48 VNB N_VGND_c_654_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_49 VNB N_VGND_c_655_n 0.00503278f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_50 VNB N_VGND_c_656_n 0.00577057f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_51 VPB N_A_c_103_n 0.0200897f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_52 VPB N_A_c_104_n 0.0158856f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_53 VPB N_A_c_105_n 0.0159691f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_54 VPB N_A_c_102_n 0.0283499f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_55 VPB N_A_27_47#_c_183_n 0.0164045f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.985
cc_56 VPB N_A_27_47#_c_184_n 0.0154215f $X=-0.19 $Y=1.305 $X2=1.065 $Y2=1.105
cc_57 VPB N_A_27_47#_c_185_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_58 VPB N_A_27_47#_c_186_n 0.0154404f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.212
cc_59 VPB N_A_27_47#_c_187_n 0.0157197f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_60 VPB N_A_27_47#_c_188_n 0.0154187f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_61 VPB N_A_27_47#_c_189_n 0.0155598f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_62 VPB N_A_27_47#_c_190_n 0.0198847f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_63 VPB N_A_27_47#_c_191_n 0.0331497f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_A_27_47#_c_192_n 0.00172363f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_A_27_47#_c_193_n 0.0107029f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_A_27_47#_c_194_n 8.69551e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_A_27_47#_c_178_n 0.00256049f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_A_27_47#_c_196_n 0.00177041f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_A_27_47#_c_182_n 0.0543892f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_396_n 0.00469739f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_397_n 0.0206409f $X=-0.19 $Y=1.305 $X2=0.6 $Y2=1.105
cc_72 VPB N_VPWR_c_398_n 0.00418552f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_399_n 3.32195e-19 $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.212
cc_74 VPB N_VPWR_c_400_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.212
cc_75 VPB N_VPWR_c_401_n 3.19622e-19 $X=-0.19 $Y=1.305 $X2=1.46 $Y2=1.212
cc_76 VPB N_VPWR_c_402_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 VPB N_VPWR_c_403_n 0.0461502f $X=-0.19 $Y=1.305 $X2=0.695 $Y2=1.19
cc_78 VPB N_VPWR_c_404_n 0.0176752f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_79 VPB N_VPWR_c_405_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_80 VPB N_VPWR_c_406_n 0.0140826f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_81 VPB N_VPWR_c_407_n 0.0143948f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_82 VPB N_VPWR_c_395_n 0.0559956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_83 VPB N_VPWR_c_409_n 0.0194569f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_84 VPB N_VPWR_c_410_n 0.00324069f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_85 VPB N_VPWR_c_411_n 0.00324402f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_86 VPB N_VPWR_c_412_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_87 VPB N_VPWR_c_413_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_88 VPB N_VPWR_c_414_n 0.00503453f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_89 VPB N_VPWR_c_415_n 0.00580385f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_90 VPB N_X_c_505_n 0.00254663f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.212
cc_91 VPB N_X_c_506_n 0.00144538f $X=-0.19 $Y=1.305 $X2=1.035 $Y2=1.16
cc_92 VPB N_X_c_507_n 0.00254663f $X=-0.19 $Y=1.305 $X2=1.05 $Y2=1.19
cc_93 VPB N_X_c_508_n 0.00241328f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_94 VPB N_X_c_509_n 0.00108853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_95 VPB N_X_c_510_n 0.00108853f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_96 VPB X 0.00138097f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_97 VPB X 4.42593e-19 $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_98 N_A_M1021_g N_A_27_47#_M1004_g 0.0204987f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_99 N_A_c_105_n N_A_27_47#_c_183_n 0.0219169f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_100 N_A_c_103_n N_A_27_47#_c_191_n 0.0115459f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_101 N_A_c_104_n N_A_27_47#_c_191_n 7.69893e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_102 N_A_M1002_g N_A_27_47#_c_202_n 0.00595153f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_103 N_A_M1002_g N_A_27_47#_c_174_n 0.01243f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_104 N_A_M1015_g N_A_27_47#_c_174_n 0.012417f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_105 A N_A_27_47#_c_174_n 0.0545384f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_106 N_A_c_102_n N_A_27_47#_c_174_n 0.00574557f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_107 A N_A_27_47#_c_175_n 0.0138086f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_108 N_A_c_102_n N_A_27_47#_c_175_n 0.00413894f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_109 N_A_c_103_n N_A_27_47#_c_192_n 0.0137916f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_110 N_A_c_104_n N_A_27_47#_c_192_n 0.0101048f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_111 A N_A_27_47#_c_192_n 0.0394547f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_112 N_A_c_102_n N_A_27_47#_c_192_n 0.00720931f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_113 N_A_c_103_n N_A_27_47#_c_193_n 0.00138874f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_114 A N_A_27_47#_c_193_n 0.0231493f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_115 N_A_c_102_n N_A_27_47#_c_193_n 0.00628911f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_116 N_A_c_103_n N_A_27_47#_c_216_n 8.07084e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_117 N_A_c_104_n N_A_27_47#_c_216_n 0.0141618f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_c_105_n N_A_27_47#_c_216_n 0.0116562f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_M1021_g N_A_27_47#_c_219_n 0.00438651f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_120 N_A_M1021_g N_A_27_47#_c_176_n 0.0123787f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_121 A N_A_27_47#_c_176_n 0.00394409f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_122 N_A_c_102_n N_A_27_47#_c_176_n 2.2583e-19 $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_123 N_A_c_105_n N_A_27_47#_c_194_n 0.0150852f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_124 N_A_c_102_n N_A_27_47#_c_194_n 3.58038e-19 $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_125 N_A_M1021_g N_A_27_47#_c_177_n 0.00420813f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_126 N_A_c_105_n N_A_27_47#_c_178_n 8.37329e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_127 A N_A_27_47#_c_178_n 0.00181689f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_128 N_A_c_102_n N_A_27_47#_c_178_n 0.00368389f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_129 N_A_c_104_n N_A_27_47#_c_196_n 0.00259297f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_c_105_n N_A_27_47#_c_196_n 0.00128924f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_131 A N_A_27_47#_c_196_n 0.0286323f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_132 N_A_c_102_n N_A_27_47#_c_196_n 0.00751302f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_133 A N_A_27_47#_c_180_n 0.0138008f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_134 N_A_c_102_n N_A_27_47#_c_180_n 0.00308219f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_135 A N_A_27_47#_c_181_n 0.01199f $X=1.065 $Y=1.105 $X2=0 $Y2=0
cc_136 N_A_c_102_n N_A_27_47#_c_181_n 0.00195556f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_137 N_A_c_102_n N_A_27_47#_c_182_n 0.0204987f $X=1.435 $Y=1.212 $X2=0 $Y2=0
cc_138 N_A_c_103_n N_VPWR_c_396_n 0.0052072f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_139 N_A_c_104_n N_VPWR_c_396_n 0.004751f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_c_104_n N_VPWR_c_397_n 0.00597712f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_c_105_n N_VPWR_c_397_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_142 N_A_c_105_n N_VPWR_c_398_n 0.0052072f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_143 N_A_c_103_n N_VPWR_c_395_n 0.0127552f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_144 N_A_c_104_n N_VPWR_c_395_n 0.00999457f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_c_105_n N_VPWR_c_395_n 0.011869f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_146 N_A_c_103_n N_VPWR_c_409_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_M1002_g N_VGND_c_637_n 0.0126564f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_148 N_A_M1015_g N_VGND_c_637_n 0.00162962f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_149 N_A_M1015_g N_VGND_c_638_n 6.55283e-19 $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_150 N_A_M1021_g N_VGND_c_638_n 0.011037f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_151 N_A_M1002_g N_VGND_c_644_n 0.0020416f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_152 N_A_M1015_g N_VGND_c_645_n 0.00439206f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_153 N_A_M1021_g N_VGND_c_645_n 0.0020416f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_154 N_A_M1002_g N_VGND_c_650_n 0.00378724f $X=0.52 $Y=0.56 $X2=0 $Y2=0
cc_155 N_A_M1015_g N_VGND_c_650_n 0.00613946f $X=0.99 $Y=0.56 $X2=0 $Y2=0
cc_156 N_A_M1021_g N_VGND_c_650_n 0.00288181f $X=1.46 $Y=0.56 $X2=0 $Y2=0
cc_157 N_A_27_47#_c_192_n N_VPWR_M1001_s 0.00199888f $X=0.985 $Y=1.53 $X2=-0.19
+ $Y2=-0.24
cc_158 N_A_27_47#_c_194_n N_VPWR_M1019_s 0.00365803f $X=1.57 $Y=1.53 $X2=0 $Y2=0
cc_159 N_A_27_47#_c_191_n N_VPWR_c_396_n 0.0381414f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_160 N_A_27_47#_c_192_n N_VPWR_c_396_n 0.0112848f $X=0.985 $Y=1.53 $X2=0 $Y2=0
cc_161 N_A_27_47#_c_216_n N_VPWR_c_396_n 0.0470327f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_162 N_A_27_47#_c_216_n N_VPWR_c_397_n 0.0223557f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_163 N_A_27_47#_c_183_n N_VPWR_c_398_n 0.00446011f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_164 N_A_27_47#_c_216_n N_VPWR_c_398_n 0.0385613f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_165 N_A_27_47#_c_194_n N_VPWR_c_398_n 0.0118234f $X=1.57 $Y=1.53 $X2=0 $Y2=0
cc_166 N_A_27_47#_c_179_n N_VPWR_c_398_n 2.86056e-19 $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_167 N_A_27_47#_c_183_n N_VPWR_c_399_n 7.31091e-19 $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_168 N_A_27_47#_c_184_n N_VPWR_c_399_n 0.0156322f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_169 N_A_27_47#_c_185_n N_VPWR_c_399_n 0.0117392f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_170 N_A_27_47#_c_186_n N_VPWR_c_399_n 6.61031e-19 $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_171 N_A_27_47#_c_185_n N_VPWR_c_400_n 6.99539e-19 $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_172 N_A_27_47#_c_186_n N_VPWR_c_400_n 0.0154534f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_173 N_A_27_47#_c_187_n N_VPWR_c_400_n 0.0117392f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_174 N_A_27_47#_c_188_n N_VPWR_c_400_n 6.61031e-19 $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_175 N_A_27_47#_c_187_n N_VPWR_c_401_n 6.99539e-19 $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_176 N_A_27_47#_c_188_n N_VPWR_c_401_n 0.0154534f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_177 N_A_27_47#_c_189_n N_VPWR_c_401_n 0.0117392f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_178 N_A_27_47#_c_190_n N_VPWR_c_401_n 6.61031e-19 $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_179 N_A_27_47#_c_189_n N_VPWR_c_402_n 0.00622633f $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_180 N_A_27_47#_c_190_n N_VPWR_c_402_n 0.00427505f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_181 N_A_27_47#_c_189_n N_VPWR_c_403_n 8.34825e-19 $X=4.725 $Y=1.41 $X2=0
+ $Y2=0
cc_182 N_A_27_47#_c_190_n N_VPWR_c_403_n 0.022204f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_183 N_A_27_47#_c_183_n N_VPWR_c_404_n 0.00702461f $X=1.905 $Y=1.41 $X2=0
+ $Y2=0
cc_184 N_A_27_47#_c_184_n N_VPWR_c_404_n 0.00427505f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_185 N_A_27_47#_c_185_n N_VPWR_c_405_n 0.00622633f $X=2.845 $Y=1.41 $X2=0
+ $Y2=0
cc_186 N_A_27_47#_c_186_n N_VPWR_c_405_n 0.00427505f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_187 N_A_27_47#_c_187_n N_VPWR_c_406_n 0.00622633f $X=3.785 $Y=1.41 $X2=0
+ $Y2=0
cc_188 N_A_27_47#_c_188_n N_VPWR_c_406_n 0.00427505f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_189 N_A_27_47#_M1001_d N_VPWR_c_395_n 0.00217517f $X=0.135 $Y=1.485 $X2=0
+ $Y2=0
cc_190 N_A_27_47#_M1008_d N_VPWR_c_395_n 0.00231261f $X=1.055 $Y=1.485 $X2=0
+ $Y2=0
cc_191 N_A_27_47#_c_183_n N_VPWR_c_395_n 0.0126126f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_27_47#_c_184_n N_VPWR_c_395_n 0.00740765f $X=2.375 $Y=1.41 $X2=0
+ $Y2=0
cc_193 N_A_27_47#_c_185_n N_VPWR_c_395_n 0.010479f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_27_47#_c_186_n N_VPWR_c_395_n 0.00740765f $X=3.315 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A_27_47#_c_187_n N_VPWR_c_395_n 0.010479f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_27_47#_c_188_n N_VPWR_c_395_n 0.00740765f $X=4.255 $Y=1.41 $X2=0
+ $Y2=0
cc_197 N_A_27_47#_c_189_n N_VPWR_c_395_n 0.010479f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_27_47#_c_190_n N_VPWR_c_395_n 0.00740765f $X=5.195 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A_27_47#_c_191_n N_VPWR_c_395_n 0.0124725f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_200 N_A_27_47#_c_216_n N_VPWR_c_395_n 0.0140101f $X=1.2 $Y=1.63 $X2=0 $Y2=0
cc_201 N_A_27_47#_c_191_n N_VPWR_c_409_n 0.0210596f $X=0.26 $Y=1.63 $X2=0 $Y2=0
cc_202 N_A_27_47#_M1004_g N_X_c_513_n 0.00462807f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_203 N_A_27_47#_c_183_n N_X_c_514_n 0.00771865f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_27_47#_c_184_n N_X_c_514_n 0.00657309f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_27_47#_M1005_g N_X_c_498_n 0.0115761f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_206 N_A_27_47#_M1009_g N_X_c_498_n 0.0120362f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_207 N_A_27_47#_c_179_n N_X_c_498_n 0.0538798f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_208 N_A_27_47#_c_182_n N_X_c_498_n 0.00342143f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_209 N_A_27_47#_M1004_g N_X_c_499_n 0.00167159f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_210 N_A_27_47#_c_176_n N_X_c_499_n 0.00988205f $X=1.57 $Y=0.82 $X2=0 $Y2=0
cc_211 N_A_27_47#_c_179_n N_X_c_499_n 0.0136633f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_212 N_A_27_47#_c_182_n N_X_c_499_n 0.00308294f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_213 N_A_27_47#_c_184_n N_X_c_505_n 0.0146085f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_214 N_A_27_47#_c_185_n N_X_c_505_n 0.0163255f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_215 N_A_27_47#_c_179_n N_X_c_505_n 0.0473195f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_216 N_A_27_47#_c_182_n N_X_c_505_n 0.0106248f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_217 N_A_27_47#_c_183_n N_X_c_506_n 0.00162552f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_27_47#_c_194_n N_X_c_506_n 0.00995523f $X=1.57 $Y=1.53 $X2=0 $Y2=0
cc_219 N_A_27_47#_c_179_n N_X_c_506_n 0.012145f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_220 N_A_27_47#_c_182_n N_X_c_506_n 0.00418485f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_221 N_A_27_47#_M1009_g N_X_c_532_n 0.00462807f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_222 N_A_27_47#_c_185_n N_X_c_533_n 0.00702928f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_27_47#_c_186_n N_X_c_533_n 0.00657309f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_27_47#_M1011_g N_X_c_500_n 0.0120914f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_225 N_A_27_47#_M1014_g N_X_c_500_n 0.0120914f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_226 N_A_27_47#_c_179_n N_X_c_500_n 0.0538798f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_27_47#_c_182_n N_X_c_500_n 0.00342143f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_228 N_A_27_47#_c_186_n N_X_c_507_n 0.0149392f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_27_47#_c_187_n N_X_c_507_n 0.0163685f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_27_47#_c_179_n N_X_c_507_n 0.0473195f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_231 N_A_27_47#_c_182_n N_X_c_507_n 0.0106248f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_232 N_A_27_47#_M1014_g N_X_c_543_n 0.00462807f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_233 N_A_27_47#_c_187_n N_X_c_544_n 0.00702928f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_234 N_A_27_47#_c_188_n N_X_c_544_n 0.00657309f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_27_47#_M1017_g N_X_c_501_n 0.0120914f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_236 N_A_27_47#_M1018_g N_X_c_501_n 0.00610685f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_237 N_A_27_47#_c_179_n N_X_c_501_n 0.027297f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_238 N_A_27_47#_c_182_n N_X_c_501_n 0.00336301f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_239 N_A_27_47#_c_188_n N_X_c_508_n 0.0148961f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_27_47#_c_189_n N_X_c_508_n 0.00612216f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_241 N_A_27_47#_c_179_n N_X_c_508_n 0.0239764f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_242 N_A_27_47#_c_182_n N_X_c_508_n 0.00950791f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_243 N_A_27_47#_M1018_g N_X_c_554_n 0.00469135f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_244 N_A_27_47#_M1020_g N_X_c_554_n 0.00174937f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_245 N_A_27_47#_c_179_n N_X_c_502_n 0.0136633f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_246 N_A_27_47#_c_182_n N_X_c_502_n 0.00308294f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_247 N_A_27_47#_c_179_n N_X_c_509_n 0.012145f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_27_47#_c_182_n N_X_c_509_n 0.00418485f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_249 N_A_27_47#_c_179_n N_X_c_503_n 0.0136633f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_250 N_A_27_47#_c_182_n N_X_c_503_n 0.00308294f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_251 N_A_27_47#_c_179_n N_X_c_510_n 0.012145f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_252 N_A_27_47#_c_182_n N_X_c_510_n 0.00418485f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_253 N_A_27_47#_M1017_g X 6.33396e-19 $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_254 N_A_27_47#_M1018_g X 0.00944399f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_255 N_A_27_47#_c_189_n X 0.0011912f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_256 N_A_27_47#_c_190_n X 9.39603e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_257 N_A_27_47#_M1020_g X 0.00500374f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_258 N_A_27_47#_c_179_n X 0.0120714f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_259 N_A_27_47#_c_182_n X 0.045751f $X=5.195 $Y=1.217 $X2=0 $Y2=0
cc_260 N_A_27_47#_c_189_n X 0.00945355f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_261 N_A_27_47#_c_190_n X 0.00210361f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_262 N_A_27_47#_c_189_n N_X_c_573_n 0.00702928f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_263 N_A_27_47#_c_190_n N_X_c_573_n 0.00289399f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_264 N_A_27_47#_c_174_n N_VGND_M1002_s 0.00213931f $X=1.115 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_265 N_A_27_47#_c_176_n N_VGND_M1021_s 0.00349935f $X=1.57 $Y=0.82 $X2=0 $Y2=0
cc_266 N_A_27_47#_c_202_n N_VGND_c_637_n 0.0231432f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_267 N_A_27_47#_c_174_n N_VGND_c_637_n 0.0219272f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_268 N_A_27_47#_M1004_g N_VGND_c_638_n 0.00850423f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_269 N_A_27_47#_M1005_g N_VGND_c_638_n 5.8773e-19 $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_270 N_A_27_47#_c_219_n N_VGND_c_638_n 0.0227699f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_271 N_A_27_47#_c_176_n N_VGND_c_638_n 0.0190274f $X=1.57 $Y=0.82 $X2=0 $Y2=0
cc_272 N_A_27_47#_c_179_n N_VGND_c_638_n 0.00197677f $X=4.28 $Y=1.16 $X2=0 $Y2=0
cc_273 N_A_27_47#_M1004_g N_VGND_c_639_n 5.66132e-19 $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_274 N_A_27_47#_M1005_g N_VGND_c_639_n 0.00806522f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_275 N_A_27_47#_M1009_g N_VGND_c_639_n 0.00842615f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_276 N_A_27_47#_M1011_g N_VGND_c_639_n 5.8773e-19 $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_277 N_A_27_47#_M1009_g N_VGND_c_640_n 5.66132e-19 $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_278 N_A_27_47#_M1011_g N_VGND_c_640_n 0.00806522f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_279 N_A_27_47#_M1014_g N_VGND_c_640_n 0.00842615f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_280 N_A_27_47#_M1017_g N_VGND_c_640_n 5.8773e-19 $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_281 N_A_27_47#_M1014_g N_VGND_c_641_n 5.66132e-19 $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_282 N_A_27_47#_M1017_g N_VGND_c_641_n 0.00806522f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_283 N_A_27_47#_M1018_g N_VGND_c_641_n 0.00845883f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_284 N_A_27_47#_M1020_g N_VGND_c_641_n 5.50819e-19 $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_285 N_A_27_47#_M1018_g N_VGND_c_642_n 0.00350486f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_286 N_A_27_47#_M1020_g N_VGND_c_642_n 0.00271402f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_287 N_A_27_47#_M1018_g N_VGND_c_643_n 7.50515e-19 $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_288 N_A_27_47#_M1020_g N_VGND_c_643_n 0.0177043f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_289 N_A_27_47#_c_202_n N_VGND_c_644_n 0.0117748f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_290 N_A_27_47#_c_174_n N_VGND_c_644_n 0.00193889f $X=1.115 $Y=0.82 $X2=0
+ $Y2=0
cc_291 N_A_27_47#_c_174_n N_VGND_c_645_n 0.00248202f $X=1.115 $Y=0.82 $X2=0
+ $Y2=0
cc_292 N_A_27_47#_c_219_n N_VGND_c_645_n 0.0112022f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_293 N_A_27_47#_c_176_n N_VGND_c_645_n 0.00193889f $X=1.57 $Y=0.82 $X2=0 $Y2=0
cc_294 N_A_27_47#_M1004_g N_VGND_c_646_n 0.0046653f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_295 N_A_27_47#_M1005_g N_VGND_c_646_n 0.00350562f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_296 N_A_27_47#_M1009_g N_VGND_c_647_n 0.00350562f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_297 N_A_27_47#_M1011_g N_VGND_c_647_n 0.00350562f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_298 N_A_27_47#_M1014_g N_VGND_c_648_n 0.00350562f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_299 N_A_27_47#_M1017_g N_VGND_c_648_n 0.00350562f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_300 N_A_27_47#_M1002_d N_VGND_c_650_n 0.00446387f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_301 N_A_27_47#_M1015_d N_VGND_c_650_n 0.00334116f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_302 N_A_27_47#_M1004_g N_VGND_c_650_n 0.00809951f $X=1.88 $Y=0.56 $X2=0 $Y2=0
cc_303 N_A_27_47#_M1005_g N_VGND_c_650_n 0.00431759f $X=2.35 $Y=0.56 $X2=0 $Y2=0
cc_304 N_A_27_47#_M1009_g N_VGND_c_650_n 0.00431759f $X=2.82 $Y=0.56 $X2=0 $Y2=0
cc_305 N_A_27_47#_M1011_g N_VGND_c_650_n 0.00431759f $X=3.29 $Y=0.56 $X2=0 $Y2=0
cc_306 N_A_27_47#_M1014_g N_VGND_c_650_n 0.00431759f $X=3.76 $Y=0.56 $X2=0 $Y2=0
cc_307 N_A_27_47#_M1017_g N_VGND_c_650_n 0.00431759f $X=4.23 $Y=0.56 $X2=0 $Y2=0
cc_308 N_A_27_47#_M1018_g N_VGND_c_650_n 0.00443596f $X=4.7 $Y=0.56 $X2=0 $Y2=0
cc_309 N_A_27_47#_M1020_g N_VGND_c_650_n 0.00522073f $X=5.22 $Y=0.56 $X2=0 $Y2=0
cc_310 N_A_27_47#_c_202_n N_VGND_c_650_n 0.0064623f $X=0.26 $Y=0.56 $X2=0 $Y2=0
cc_311 N_A_27_47#_c_174_n N_VGND_c_650_n 0.0104775f $X=1.115 $Y=0.82 $X2=0 $Y2=0
cc_312 N_A_27_47#_c_219_n N_VGND_c_650_n 0.00644569f $X=1.2 $Y=0.56 $X2=0 $Y2=0
cc_313 N_A_27_47#_c_176_n N_VGND_c_650_n 0.00526647f $X=1.57 $Y=0.82 $X2=0 $Y2=0
cc_314 N_VPWR_c_395_n N_X_M1000_d 0.00656398f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_315 N_VPWR_c_395_n N_X_M1006_d 0.00656398f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_316 N_VPWR_c_395_n N_X_M1010_d 0.00656398f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_317 N_VPWR_c_395_n N_X_M1013_d 0.00656398f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_318 N_VPWR_c_398_n N_X_c_514_n 0.0301172f $X=1.67 $Y=2 $X2=0 $Y2=0
cc_319 N_VPWR_c_399_n N_X_c_514_n 0.0470327f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_320 N_VPWR_c_404_n N_X_c_514_n 0.0118139f $X=2.395 $Y=2.72 $X2=0 $Y2=0
cc_321 N_VPWR_c_395_n N_X_c_514_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_322 N_VPWR_M1003_s N_X_c_505_n 0.00209407f $X=2.465 $Y=1.485 $X2=0 $Y2=0
cc_323 N_VPWR_c_399_n N_X_c_505_n 0.0172025f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_324 N_VPWR_c_399_n N_X_c_533_n 0.0385613f $X=2.61 $Y=2 $X2=0 $Y2=0
cc_325 N_VPWR_c_400_n N_X_c_533_n 0.0470327f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_326 N_VPWR_c_405_n N_X_c_533_n 0.0118139f $X=3.335 $Y=2.72 $X2=0 $Y2=0
cc_327 N_VPWR_c_395_n N_X_c_533_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_328 N_VPWR_M1007_s N_X_c_507_n 0.00209407f $X=3.405 $Y=1.485 $X2=0 $Y2=0
cc_329 N_VPWR_c_400_n N_X_c_507_n 0.0172025f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_330 N_VPWR_c_400_n N_X_c_544_n 0.0385613f $X=3.55 $Y=2 $X2=0 $Y2=0
cc_331 N_VPWR_c_401_n N_X_c_544_n 0.0470327f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_332 N_VPWR_c_406_n N_X_c_544_n 0.0118139f $X=4.275 $Y=2.72 $X2=0 $Y2=0
cc_333 N_VPWR_c_395_n N_X_c_544_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_334 N_VPWR_M1012_s N_X_c_508_n 0.00209407f $X=4.345 $Y=1.485 $X2=0 $Y2=0
cc_335 N_VPWR_c_401_n N_X_c_508_n 0.0172025f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_336 N_VPWR_c_403_n X 0.0108422f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_337 N_VPWR_c_401_n N_X_c_573_n 0.0385613f $X=4.49 $Y=2 $X2=0 $Y2=0
cc_338 N_VPWR_c_402_n N_X_c_573_n 0.0118139f $X=5.215 $Y=2.72 $X2=0 $Y2=0
cc_339 N_VPWR_c_403_n N_X_c_573_n 0.0634205f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_340 N_VPWR_c_395_n N_X_c_573_n 0.00646998f $X=5.75 $Y=2.72 $X2=0 $Y2=0
cc_341 N_VPWR_c_403_n N_VGND_c_643_n 0.0109366f $X=5.43 $Y=1.66 $X2=0 $Y2=0
cc_342 N_X_c_498_n N_VGND_M1005_s 0.00213931f $X=2.995 $Y=0.82 $X2=0 $Y2=0
cc_343 N_X_c_500_n N_VGND_M1011_s 0.00213931f $X=3.935 $Y=0.82 $X2=0 $Y2=0
cc_344 N_X_c_501_n N_VGND_M1017_s 0.00213931f $X=4.69 $Y=0.82 $X2=0 $Y2=0
cc_345 N_X_c_513_n N_VGND_c_638_n 0.0189749f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_346 N_X_c_498_n N_VGND_c_639_n 0.0203425f $X=2.995 $Y=0.82 $X2=0 $Y2=0
cc_347 N_X_c_532_n N_VGND_c_639_n 0.0189749f $X=3.08 $Y=0.56 $X2=0 $Y2=0
cc_348 N_X_c_500_n N_VGND_c_640_n 0.0203425f $X=3.935 $Y=0.82 $X2=0 $Y2=0
cc_349 N_X_c_543_n N_VGND_c_640_n 0.0189749f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_350 N_X_c_501_n N_VGND_c_641_n 0.0203425f $X=4.69 $Y=0.82 $X2=0 $Y2=0
cc_351 N_X_c_554_n N_VGND_c_641_n 0.0189749f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_352 N_X_c_501_n N_VGND_c_642_n 4.45603e-19 $X=4.69 $Y=0.82 $X2=0 $Y2=0
cc_353 N_X_c_554_n N_VGND_c_642_n 0.0118139f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_354 X N_VGND_c_642_n 0.00233077f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_355 N_X_c_554_n N_VGND_c_643_n 0.0357983f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_356 X N_VGND_c_643_n 0.0125104f $X=4.745 $Y=0.765 $X2=0 $Y2=0
cc_357 N_X_c_513_n N_VGND_c_646_n 0.0115672f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_358 N_X_c_498_n N_VGND_c_646_n 0.00193763f $X=2.995 $Y=0.82 $X2=0 $Y2=0
cc_359 N_X_c_498_n N_VGND_c_647_n 0.00259419f $X=2.995 $Y=0.82 $X2=0 $Y2=0
cc_360 N_X_c_532_n N_VGND_c_647_n 0.0115672f $X=3.08 $Y=0.56 $X2=0 $Y2=0
cc_361 N_X_c_500_n N_VGND_c_647_n 0.00193763f $X=3.935 $Y=0.82 $X2=0 $Y2=0
cc_362 N_X_c_500_n N_VGND_c_648_n 0.00259419f $X=3.935 $Y=0.82 $X2=0 $Y2=0
cc_363 N_X_c_543_n N_VGND_c_648_n 0.0115672f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_364 N_X_c_501_n N_VGND_c_648_n 0.00193763f $X=4.69 $Y=0.82 $X2=0 $Y2=0
cc_365 N_X_M1004_d N_VGND_c_650_n 0.00632385f $X=1.955 $Y=0.235 $X2=0 $Y2=0
cc_366 N_X_M1009_d N_VGND_c_650_n 0.00332158f $X=2.895 $Y=0.235 $X2=0 $Y2=0
cc_367 N_X_M1014_d N_VGND_c_650_n 0.00332158f $X=3.835 $Y=0.235 $X2=0 $Y2=0
cc_368 N_X_M1018_d N_VGND_c_650_n 0.00700694f $X=4.775 $Y=0.235 $X2=0 $Y2=0
cc_369 N_X_c_513_n N_VGND_c_650_n 0.0064623f $X=2.14 $Y=0.56 $X2=0 $Y2=0
cc_370 N_X_c_498_n N_VGND_c_650_n 0.0104569f $X=2.995 $Y=0.82 $X2=0 $Y2=0
cc_371 N_X_c_532_n N_VGND_c_650_n 0.0064623f $X=3.08 $Y=0.56 $X2=0 $Y2=0
cc_372 N_X_c_500_n N_VGND_c_650_n 0.0104569f $X=3.935 $Y=0.82 $X2=0 $Y2=0
cc_373 N_X_c_543_n N_VGND_c_650_n 0.0064623f $X=4.02 $Y=0.56 $X2=0 $Y2=0
cc_374 N_X_c_501_n N_VGND_c_650_n 0.00604001f $X=4.69 $Y=0.82 $X2=0 $Y2=0
cc_375 N_X_c_554_n N_VGND_c_650_n 0.00646998f $X=4.96 $Y=0.56 $X2=0 $Y2=0
cc_376 X N_VGND_c_650_n 0.00472011f $X=4.745 $Y=0.765 $X2=0 $Y2=0
