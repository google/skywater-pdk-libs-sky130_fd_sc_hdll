* File: sky130_fd_sc_hdll__nand2_6.pxi.spice
* Created: Thu Aug 27 19:13:02 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_6%B N_B_c_77_n N_B_M1002_g N_B_c_85_n N_B_M1001_g
+ N_B_c_86_n N_B_M1008_g N_B_c_78_n N_B_M1007_g N_B_c_79_n N_B_M1015_g
+ N_B_c_87_n N_B_M1010_g N_B_c_88_n N_B_M1012_g N_B_c_80_n N_B_M1017_g
+ N_B_c_81_n N_B_M1019_g N_B_c_89_n N_B_M1016_g N_B_c_90_n N_B_M1020_g
+ N_B_c_82_n N_B_M1021_g B N_B_c_83_n N_B_c_84_n PM_SKY130_FD_SC_HDLL__NAND2_6%B
x_PM_SKY130_FD_SC_HDLL__NAND2_6%A N_A_c_203_n N_A_M1005_g N_A_c_210_n
+ N_A_M1000_g N_A_c_204_n N_A_M1009_g N_A_c_211_n N_A_M1003_g N_A_c_205_n
+ N_A_M1011_g N_A_c_212_n N_A_M1004_g N_A_c_213_n N_A_M1006_g N_A_c_206_n
+ N_A_M1013_g N_A_c_207_n N_A_M1022_g N_A_c_214_n N_A_M1014_g N_A_c_215_n
+ N_A_M1018_g N_A_c_208_n N_A_M1023_g A N_A_c_248_p N_A_c_209_n
+ PM_SKY130_FD_SC_HDLL__NAND2_6%A
x_PM_SKY130_FD_SC_HDLL__NAND2_6%VPWR N_VPWR_M1001_d N_VPWR_M1008_d
+ N_VPWR_M1012_d N_VPWR_M1020_d N_VPWR_M1003_d N_VPWR_M1006_d N_VPWR_M1018_d
+ N_VPWR_c_309_n N_VPWR_c_310_n N_VPWR_c_311_n N_VPWR_c_312_n N_VPWR_c_313_n
+ N_VPWR_c_314_n N_VPWR_c_315_n N_VPWR_c_316_n N_VPWR_c_317_n N_VPWR_c_318_n
+ N_VPWR_c_319_n N_VPWR_c_320_n N_VPWR_c_321_n N_VPWR_c_322_n VPWR
+ N_VPWR_c_323_n N_VPWR_c_324_n N_VPWR_c_308_n N_VPWR_c_326_n N_VPWR_c_327_n
+ N_VPWR_c_328_n N_VPWR_c_329_n N_VPWR_c_330_n
+ PM_SKY130_FD_SC_HDLL__NAND2_6%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_6%Y N_Y_M1005_d N_Y_M1011_d N_Y_M1022_d
+ N_Y_M1001_s N_Y_M1010_s N_Y_M1016_s N_Y_M1000_s N_Y_M1004_s N_Y_M1014_s
+ N_Y_c_404_n N_Y_c_408_n N_Y_c_411_n N_Y_c_415_n N_Y_c_419_n N_Y_c_423_n
+ N_Y_c_426_n N_Y_c_427_n N_Y_c_444_n N_Y_c_450_n N_Y_c_454_n N_Y_c_458_n
+ N_Y_c_462_n N_Y_c_526_p N_Y_c_398_n N_Y_c_401_n N_Y_c_428_n N_Y_c_432_n
+ N_Y_c_471_n N_Y_c_472_n N_Y_c_475_n N_Y_c_479_n N_Y_c_399_n Y
+ PM_SKY130_FD_SC_HDLL__NAND2_6%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_6%A_27_47# N_A_27_47#_M1002_d N_A_27_47#_M1007_d
+ N_A_27_47#_M1017_d N_A_27_47#_M1021_d N_A_27_47#_M1009_s N_A_27_47#_M1013_s
+ N_A_27_47#_M1023_s N_A_27_47#_c_533_n N_A_27_47#_c_541_n N_A_27_47#_c_534_n
+ N_A_27_47#_c_547_n N_A_27_47#_c_551_n N_A_27_47#_c_555_n N_A_27_47#_c_559_n
+ N_A_27_47#_c_563_n N_A_27_47#_c_535_n N_A_27_47#_c_574_n N_A_27_47#_c_536_n
+ N_A_27_47#_c_537_n N_A_27_47#_c_538_n PM_SKY130_FD_SC_HDLL__NAND2_6%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_6%VGND N_VGND_M1002_s N_VGND_M1015_s
+ N_VGND_M1019_s N_VGND_c_629_n N_VGND_c_630_n N_VGND_c_631_n N_VGND_c_632_n
+ N_VGND_c_633_n VGND N_VGND_c_634_n N_VGND_c_635_n N_VGND_c_636_n
+ N_VGND_c_637_n N_VGND_c_638_n N_VGND_c_639_n
+ PM_SKY130_FD_SC_HDLL__NAND2_6%VGND
cc_1 VNB N_B_c_77_n 0.0228251f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_78_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B_c_79_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_B_c_80_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B_c_81_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_6 VNB N_B_c_82_n 0.0171127f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_7 VNB N_B_c_83_n 0.0101411f $X=-0.19 $Y=-0.24 $X2=2.6 $Y2=1.16
cc_8 VNB N_B_c_84_n 0.118032f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.202
cc_9 VNB N_A_c_203_n 0.0162568f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_10 VNB N_A_c_204_n 0.0168735f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_11 VNB N_A_c_205_n 0.0173555f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_12 VNB N_A_c_206_n 0.0168753f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_13 VNB N_A_c_207_n 0.0168204f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_14 VNB N_A_c_208_n 0.0227991f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_15 VNB N_A_c_209_n 0.119737f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.202
cc_16 VNB N_VPWR_c_308_n 0.269736f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_Y_c_398_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_Y_c_399_n 0.0113445f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB Y 0.00106016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB N_A_27_47#_c_533_n 0.0182048f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_21 VNB N_A_27_47#_c_534_n 0.0121122f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_22 VNB N_A_27_47#_c_535_n 0.00257277f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.202
cc_23 VNB N_A_27_47#_c_536_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=1.202
cc_24 VNB N_A_27_47#_c_537_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.202
cc_25 VNB N_A_27_47#_c_538_n 0.0292293f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.19
cc_26 VNB N_VGND_c_629_n 0.00466649f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.56
cc_27 VNB N_VGND_c_630_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.56
cc_28 VNB N_VGND_c_631_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=1.435 $Y2=1.985
cc_29 VNB N_VGND_c_632_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.985
cc_30 VNB N_VGND_c_633_n 0.00466098f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.56
cc_31 VNB N_VGND_c_634_n 0.0171658f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.41
cc_32 VNB N_VGND_c_635_n 0.0885447f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_636_n 0.325825f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_34 VNB N_VGND_c_637_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_35 VNB N_VGND_c_638_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_36 VNB N_VGND_c_639_n 0.00515836f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_37 VPB N_B_c_85_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_38 VPB N_B_c_86_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_39 VPB N_B_c_87_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_40 VPB N_B_c_88_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_41 VPB N_B_c_89_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_42 VPB N_B_c_90_n 0.0164383f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_43 VPB N_B_c_83_n 7.73822e-19 $X=-0.19 $Y=1.305 $X2=2.6 $Y2=1.16
cc_44 VPB N_B_c_84_n 0.074424f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.202
cc_45 VPB N_A_c_210_n 0.0161146f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_46 VPB N_A_c_211_n 0.0162386f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_47 VPB N_A_c_212_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_48 VPB N_A_c_213_n 0.0162606f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_49 VPB N_A_c_214_n 0.016238f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_50 VPB N_A_c_215_n 0.0207627f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_51 VPB N_A_c_209_n 0.0754428f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.202
cc_52 VPB N_VPWR_c_309_n 0.0113525f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.995
cc_53 VPB N_VPWR_c_310_n 0.0410822f $X=-0.19 $Y=1.305 $X2=1.93 $Y2=0.56
cc_54 VPB N_VPWR_c_311_n 0.0041373f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.985
cc_55 VPB N_VPWR_c_312_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.985
cc_56 VPB N_VPWR_c_313_n 0.0041373f $X=-0.19 $Y=1.305 $X2=2.87 $Y2=0.56
cc_57 VPB N_VPWR_c_314_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_58 VPB N_VPWR_c_315_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.16
cc_59 VPB N_VPWR_c_316_n 0.017949f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_60 VPB N_VPWR_c_317_n 0.0041373f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_61 VPB N_VPWR_c_318_n 0.017949f $X=-0.19 $Y=1.305 $X2=2.35 $Y2=1.202
cc_62 VPB N_VPWR_c_319_n 0.0041373f $X=-0.19 $Y=1.305 $X2=2.6 $Y2=1.16
cc_63 VPB N_VPWR_c_320_n 0.0410822f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_64 VPB N_VPWR_c_321_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_65 VPB N_VPWR_c_322_n 0.00516416f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_66 VPB N_VPWR_c_323_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_67 VPB N_VPWR_c_324_n 0.0150312f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_68 VPB N_VPWR_c_308_n 0.0575384f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_69 VPB N_VPWR_c_326_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_VPWR_c_327_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_71 VPB N_VPWR_c_328_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_72 VPB N_VPWR_c_329_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_73 VPB N_VPWR_c_330_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_74 VPB N_Y_c_401_n 0.0015125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_75 VPB N_Y_c_399_n 0.00213764f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_76 VPB Y 0.00155805f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_77 N_B_c_82_n N_A_c_203_n 0.0171779f $X=2.87 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_78 N_B_c_90_n N_A_c_210_n 0.0231397f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_79 N_B_c_83_n N_A_c_209_n 9.36964e-19 $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_80 N_B_c_84_n N_A_c_209_n 0.0171779f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_81 N_B_c_85_n N_VPWR_c_310_n 0.00354866f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_82 N_B_c_86_n N_VPWR_c_311_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_83 N_B_c_87_n N_VPWR_c_311_n 0.00173895f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_84 N_B_c_87_n N_VPWR_c_312_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_85 N_B_c_88_n N_VPWR_c_312_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_86 N_B_c_88_n N_VPWR_c_313_n 0.00173895f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_87 N_B_c_89_n N_VPWR_c_313_n 0.00173895f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_88 N_B_c_89_n N_VPWR_c_314_n 0.00673617f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_89 N_B_c_90_n N_VPWR_c_314_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_90 N_B_c_90_n N_VPWR_c_315_n 0.00173895f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_91 N_B_c_85_n N_VPWR_c_323_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_92 N_B_c_86_n N_VPWR_c_323_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_93 N_B_c_85_n N_VPWR_c_308_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_94 N_B_c_86_n N_VPWR_c_308_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_95 N_B_c_87_n N_VPWR_c_308_n 0.0117184f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_96 N_B_c_88_n N_VPWR_c_308_n 0.0117184f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_97 N_B_c_89_n N_VPWR_c_308_n 0.0117184f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_98 N_B_c_90_n N_VPWR_c_308_n 0.0117436f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_99 N_B_c_85_n N_Y_c_404_n 0.00215964f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_100 N_B_c_86_n N_Y_c_404_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_101 N_B_c_83_n N_Y_c_404_n 0.0215641f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_102 N_B_c_84_n N_Y_c_404_n 0.00631893f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_103 N_B_c_85_n N_Y_c_408_n 0.00897418f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_104 N_B_c_86_n N_Y_c_408_n 0.0100233f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_105 N_B_c_87_n N_Y_c_408_n 5.91934e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_106 N_B_c_86_n N_Y_c_411_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_107 N_B_c_87_n N_Y_c_411_n 0.0137916f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_108 N_B_c_83_n N_Y_c_411_n 0.0393642f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_109 N_B_c_84_n N_Y_c_411_n 0.00655651f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_110 N_B_c_86_n N_Y_c_415_n 5.91934e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_111 N_B_c_87_n N_Y_c_415_n 0.0100233f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_112 N_B_c_88_n N_Y_c_415_n 0.0100233f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_113 N_B_c_89_n N_Y_c_415_n 5.91934e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_114 N_B_c_88_n N_Y_c_419_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_115 N_B_c_89_n N_Y_c_419_n 0.0137916f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_116 N_B_c_83_n N_Y_c_419_n 0.0393642f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_117 N_B_c_84_n N_Y_c_419_n 0.00655651f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_118 N_B_c_88_n N_Y_c_423_n 5.91934e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_119 N_B_c_89_n N_Y_c_423_n 0.0100233f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_120 N_B_c_90_n N_Y_c_423_n 0.0100233f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_121 N_B_c_90_n N_Y_c_426_n 0.0159487f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_122 N_B_c_90_n N_Y_c_427_n 5.91934e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_123 N_B_c_87_n N_Y_c_428_n 5.79575e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_124 N_B_c_88_n N_Y_c_428_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_125 N_B_c_83_n N_Y_c_428_n 0.0215641f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_126 N_B_c_84_n N_Y_c_428_n 0.00631893f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_127 N_B_c_89_n N_Y_c_432_n 5.79575e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_128 N_B_c_90_n N_Y_c_432_n 7.27961e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_129 N_B_c_83_n N_Y_c_432_n 0.0207773f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_130 N_B_c_84_n N_Y_c_432_n 0.00631893f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_131 N_B_c_90_n Y 4.25242e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_132 N_B_c_82_n Y 0.00238668f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_133 N_B_c_83_n Y 0.00781726f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_134 N_B_c_77_n N_A_27_47#_c_533_n 0.00661134f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_135 N_B_c_78_n N_A_27_47#_c_533_n 5.22294e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_136 N_B_c_77_n N_A_27_47#_c_541_n 0.00899636f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_137 N_B_c_78_n N_A_27_47#_c_541_n 0.00899636f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_138 N_B_c_83_n N_A_27_47#_c_541_n 0.0395582f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_139 N_B_c_84_n N_A_27_47#_c_541_n 0.00457246f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_140 N_B_c_77_n N_A_27_47#_c_534_n 8.68782e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_141 N_B_c_83_n N_A_27_47#_c_534_n 0.00230475f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_142 N_B_c_77_n N_A_27_47#_c_547_n 5.22365e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_143 N_B_c_78_n N_A_27_47#_c_547_n 0.00661134f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_144 N_B_c_79_n N_A_27_47#_c_547_n 0.00661134f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_145 N_B_c_80_n N_A_27_47#_c_547_n 5.22365e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_146 N_B_c_79_n N_A_27_47#_c_551_n 0.00899636f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_147 N_B_c_80_n N_A_27_47#_c_551_n 0.00899636f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_148 N_B_c_83_n N_A_27_47#_c_551_n 0.0395582f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_149 N_B_c_84_n N_A_27_47#_c_551_n 0.00457246f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_150 N_B_c_79_n N_A_27_47#_c_555_n 5.22365e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_151 N_B_c_80_n N_A_27_47#_c_555_n 0.00661134f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_152 N_B_c_81_n N_A_27_47#_c_555_n 0.00661134f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_153 N_B_c_82_n N_A_27_47#_c_555_n 5.22365e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_154 N_B_c_81_n N_A_27_47#_c_559_n 0.00899636f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_155 N_B_c_82_n N_A_27_47#_c_559_n 0.0106433f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_156 N_B_c_83_n N_A_27_47#_c_559_n 0.0300673f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_157 N_B_c_84_n N_A_27_47#_c_559_n 0.00457246f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_158 N_B_c_82_n N_A_27_47#_c_563_n 0.00248145f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_159 N_B_c_81_n N_A_27_47#_c_535_n 4.7541e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_160 N_B_c_82_n N_A_27_47#_c_535_n 0.00541116f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_161 N_B_c_78_n N_A_27_47#_c_536_n 8.68782e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_162 N_B_c_79_n N_A_27_47#_c_536_n 8.68782e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_163 N_B_c_83_n N_A_27_47#_c_536_n 0.0214029f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_164 N_B_c_84_n N_A_27_47#_c_536_n 0.00224547f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_165 N_B_c_80_n N_A_27_47#_c_537_n 8.68782e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_166 N_B_c_81_n N_A_27_47#_c_537_n 8.68782e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_167 N_B_c_83_n N_A_27_47#_c_537_n 0.0214029f $X=2.6 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B_c_84_n N_A_27_47#_c_537_n 0.00224547f $X=2.845 $Y=1.202 $X2=0 $Y2=0
cc_169 N_B_c_77_n N_VGND_c_629_n 0.00296353f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_170 N_B_c_78_n N_VGND_c_629_n 0.00166854f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B_c_78_n N_VGND_c_630_n 0.00422241f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_172 N_B_c_79_n N_VGND_c_630_n 0.00422241f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_173 N_B_c_79_n N_VGND_c_631_n 0.00166854f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B_c_80_n N_VGND_c_631_n 0.00166854f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_175 N_B_c_80_n N_VGND_c_632_n 0.00422241f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_176 N_B_c_81_n N_VGND_c_632_n 0.00422241f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_177 N_B_c_81_n N_VGND_c_633_n 0.00166854f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_178 N_B_c_82_n N_VGND_c_633_n 0.00296353f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_179 N_B_c_77_n N_VGND_c_634_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_180 N_B_c_82_n N_VGND_c_635_n 0.00420723f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_181 N_B_c_77_n N_VGND_c_636_n 0.00689308f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_182 N_B_c_78_n N_VGND_c_636_n 0.00593887f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_183 N_B_c_79_n N_VGND_c_636_n 0.00593887f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_184 N_B_c_80_n N_VGND_c_636_n 0.00593887f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_185 N_B_c_81_n N_VGND_c_636_n 0.00593887f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_186 N_B_c_82_n N_VGND_c_636_n 0.00597515f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_187 N_A_c_210_n N_VPWR_c_315_n 0.00173895f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_188 N_A_c_210_n N_VPWR_c_316_n 0.00673617f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_189 N_A_c_211_n N_VPWR_c_316_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_190 N_A_c_211_n N_VPWR_c_317_n 0.00173895f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_191 N_A_c_212_n N_VPWR_c_317_n 0.00173895f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_192 N_A_c_212_n N_VPWR_c_318_n 0.00673617f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_193 N_A_c_213_n N_VPWR_c_318_n 0.00673617f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_194 N_A_c_213_n N_VPWR_c_319_n 0.00173895f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_195 N_A_c_214_n N_VPWR_c_319_n 0.00173895f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_196 N_A_c_215_n N_VPWR_c_320_n 0.00354866f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_197 N_A_c_214_n N_VPWR_c_321_n 0.00673617f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_198 N_A_c_215_n N_VPWR_c_321_n 0.00673617f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_199 N_A_c_210_n N_VPWR_c_308_n 0.0117436f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_200 N_A_c_211_n N_VPWR_c_308_n 0.0117184f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_201 N_A_c_212_n N_VPWR_c_308_n 0.0117184f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_202 N_A_c_213_n N_VPWR_c_308_n 0.0117184f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_203 N_A_c_214_n N_VPWR_c_308_n 0.0117184f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A_c_215_n N_VPWR_c_308_n 0.0128058f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_205 N_A_c_210_n N_Y_c_423_n 5.91934e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_206 N_A_c_210_n N_Y_c_426_n 0.0133907f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_207 N_A_c_210_n N_Y_c_427_n 0.0100233f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_208 N_A_c_211_n N_Y_c_427_n 0.0100233f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_209 N_A_c_212_n N_Y_c_427_n 5.91934e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_210 N_A_c_204_n N_Y_c_444_n 0.0124451f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_211 N_A_c_205_n N_Y_c_444_n 0.0109111f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_212 N_A_c_206_n N_Y_c_444_n 0.0104739f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_213 N_A_c_207_n N_Y_c_444_n 0.0116346f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_214 N_A_c_248_p N_Y_c_444_n 0.0868511f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_215 N_A_c_209_n N_Y_c_444_n 0.0102042f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_216 N_A_c_211_n N_Y_c_450_n 0.014973f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_217 N_A_c_212_n N_Y_c_450_n 0.0137916f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_218 N_A_c_248_p N_Y_c_450_n 0.0330732f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_219 N_A_c_209_n N_Y_c_450_n 0.00635951f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_220 N_A_c_211_n N_Y_c_454_n 5.91934e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_221 N_A_c_212_n N_Y_c_454_n 0.0100233f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_222 N_A_c_213_n N_Y_c_454_n 0.0100233f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_223 N_A_c_214_n N_Y_c_454_n 5.91934e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_224 N_A_c_213_n N_Y_c_458_n 0.0137916f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_225 N_A_c_214_n N_Y_c_458_n 0.0152385f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_226 N_A_c_248_p N_Y_c_458_n 0.0316677f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_227 N_A_c_209_n N_Y_c_458_n 0.00655651f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_228 N_A_c_213_n N_Y_c_462_n 5.91934e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_229 N_A_c_214_n N_Y_c_462_n 0.0100233f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_230 N_A_c_215_n N_Y_c_462_n 0.00897418f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_231 N_A_c_207_n N_Y_c_398_n 0.00286869f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_232 N_A_c_208_n N_Y_c_398_n 0.0031043f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_233 N_A_c_209_n N_Y_c_398_n 0.0106358f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_234 N_A_c_214_n N_Y_c_401_n 0.0019905f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_235 N_A_c_215_n N_Y_c_401_n 0.00423504f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_236 N_A_c_209_n N_Y_c_401_n 0.00694896f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_237 N_A_c_203_n N_Y_c_471_n 0.00303037f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_238 N_A_c_210_n N_Y_c_472_n 0.0036484f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_239 N_A_c_211_n N_Y_c_472_n 8.15944e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_240 N_A_c_209_n N_Y_c_472_n 0.00123735f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_241 N_A_c_212_n N_Y_c_475_n 5.79575e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_242 N_A_c_213_n N_Y_c_475_n 5.79575e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_243 N_A_c_248_p N_Y_c_475_n 0.0215641f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_244 N_A_c_209_n N_Y_c_475_n 0.00631893f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_245 N_A_c_214_n N_Y_c_479_n 8.15944e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_246 N_A_c_215_n N_Y_c_479_n 0.00188422f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_247 N_A_c_248_p N_Y_c_399_n 0.022444f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_248 N_A_c_209_n N_Y_c_399_n 0.0380526f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_249 N_A_c_203_n Y 0.00315482f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_250 N_A_c_210_n Y 0.00253311f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_251 N_A_c_204_n Y 0.00297134f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_252 N_A_c_211_n Y 0.00220286f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_253 N_A_c_248_p Y 0.0212466f $X=4.99 $Y=1.16 $X2=0 $Y2=0
cc_254 N_A_c_209_n Y 0.0346925f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_255 N_A_c_203_n N_A_27_47#_c_574_n 0.0127822f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_256 N_A_c_204_n N_A_27_47#_c_574_n 0.00903374f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_257 N_A_c_205_n N_A_27_47#_c_574_n 0.00935436f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_258 N_A_c_206_n N_A_27_47#_c_574_n 0.00935436f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_259 N_A_c_207_n N_A_27_47#_c_574_n 0.00935436f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_260 N_A_c_208_n N_A_27_47#_c_574_n 0.0113668f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_261 N_A_c_209_n N_A_27_47#_c_574_n 0.00110461f $X=5.665 $Y=1.202 $X2=0 $Y2=0
cc_262 N_A_c_203_n N_VGND_c_635_n 0.00357877f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_263 N_A_c_204_n N_VGND_c_635_n 0.00357877f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_264 N_A_c_205_n N_VGND_c_635_n 0.00357877f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_265 N_A_c_206_n N_VGND_c_635_n 0.00357877f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_266 N_A_c_207_n N_VGND_c_635_n 0.00357877f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_267 N_A_c_208_n N_VGND_c_635_n 0.00357877f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_268 N_A_c_203_n N_VGND_c_636_n 0.00538422f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_269 N_A_c_204_n N_VGND_c_636_n 0.00548399f $X=3.76 $Y=0.995 $X2=0 $Y2=0
cc_270 N_A_c_205_n N_VGND_c_636_n 0.00560377f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_271 N_A_c_206_n N_VGND_c_636_n 0.0054768f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_272 N_A_c_207_n N_VGND_c_636_n 0.0054768f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_273 N_A_c_208_n N_VGND_c_636_n 0.00661249f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_274 N_VPWR_c_308_n N_Y_M1001_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_275 N_VPWR_c_308_n N_Y_M1010_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_276 N_VPWR_c_308_n N_Y_M1016_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_277 N_VPWR_c_308_n N_Y_M1000_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_278 N_VPWR_c_308_n N_Y_M1004_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_279 N_VPWR_c_308_n N_Y_M1014_s 0.00231261f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_280 N_VPWR_c_323_n N_Y_c_408_n 0.0189467f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_281 N_VPWR_c_308_n N_Y_c_408_n 0.0123132f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_282 N_VPWR_M1008_d N_Y_c_411_n 0.00334388f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_283 N_VPWR_c_311_n N_Y_c_411_n 0.0143191f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_284 N_VPWR_c_312_n N_Y_c_415_n 0.0189467f $X=2.005 $Y=2.72 $X2=0 $Y2=0
cc_285 N_VPWR_c_308_n N_Y_c_415_n 0.0123132f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_286 N_VPWR_M1012_d N_Y_c_419_n 0.00334388f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_287 N_VPWR_c_313_n N_Y_c_419_n 0.0143191f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_288 N_VPWR_c_314_n N_Y_c_423_n 0.0189467f $X=2.945 $Y=2.72 $X2=0 $Y2=0
cc_289 N_VPWR_c_308_n N_Y_c_423_n 0.0123132f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_290 N_VPWR_M1020_d N_Y_c_426_n 0.00534233f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_291 N_VPWR_c_315_n N_Y_c_426_n 0.0143191f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_292 N_VPWR_c_316_n N_Y_c_427_n 0.0189467f $X=3.885 $Y=2.72 $X2=0 $Y2=0
cc_293 N_VPWR_c_308_n N_Y_c_427_n 0.0123132f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_294 N_VPWR_M1003_d N_Y_c_450_n 0.00334388f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_295 N_VPWR_c_317_n N_Y_c_450_n 0.0143191f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_296 N_VPWR_c_318_n N_Y_c_454_n 0.0189467f $X=4.825 $Y=2.72 $X2=0 $Y2=0
cc_297 N_VPWR_c_308_n N_Y_c_454_n 0.0123132f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_298 N_VPWR_M1006_d N_Y_c_458_n 0.00334388f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_299 N_VPWR_c_319_n N_Y_c_458_n 0.0143191f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_300 N_VPWR_c_321_n N_Y_c_462_n 0.0189467f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_301 N_VPWR_c_308_n N_Y_c_462_n 0.0123027f $X=6.21 $Y=2.72 $X2=0 $Y2=0
cc_302 N_VPWR_c_320_n N_Y_c_399_n 0.010666f $X=5.9 $Y=1.66 $X2=0 $Y2=0
cc_303 N_VPWR_c_310_n N_A_27_47#_c_534_n 0.00746809f $X=0.26 $Y=1.66 $X2=0 $Y2=0
cc_304 N_VPWR_c_320_n N_A_27_47#_c_538_n 0.00411041f $X=5.9 $Y=1.66 $X2=0 $Y2=0
cc_305 N_Y_c_444_n N_A_27_47#_M1009_s 0.00401355f $X=5.325 $Y=0.76 $X2=0 $Y2=0
cc_306 N_Y_c_444_n N_A_27_47#_M1013_s 0.00307883f $X=5.325 $Y=0.76 $X2=0 $Y2=0
cc_307 N_Y_c_426_n N_A_27_47#_c_559_n 0.00303452f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_308 N_Y_c_426_n N_A_27_47#_c_535_n 0.00572467f $X=3.335 $Y=1.58 $X2=0 $Y2=0
cc_309 N_Y_M1005_d N_A_27_47#_c_574_n 0.00399738f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_310 N_Y_M1011_d N_A_27_47#_c_574_n 0.00507102f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_311 N_Y_M1022_d N_A_27_47#_c_574_n 0.00506571f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_312 N_Y_c_444_n N_A_27_47#_c_574_n 0.0862528f $X=5.325 $Y=0.76 $X2=0 $Y2=0
cc_313 N_Y_c_526_p N_A_27_47#_c_574_n 0.018174f $X=5.46 $Y=0.885 $X2=0 $Y2=0
cc_314 N_Y_c_471_n N_A_27_47#_c_574_n 0.0182216f $X=3.485 $Y=0.885 $X2=0 $Y2=0
cc_315 N_Y_c_399_n N_A_27_47#_c_574_n 0.00406744f $X=5.46 $Y=1.19 $X2=0 $Y2=0
cc_316 N_Y_c_399_n N_A_27_47#_c_538_n 0.0101702f $X=5.46 $Y=1.19 $X2=0 $Y2=0
cc_317 N_Y_M1005_d N_VGND_c_636_n 0.00256987f $X=3.365 $Y=0.235 $X2=0 $Y2=0
cc_318 N_Y_M1011_d N_VGND_c_636_n 0.00297142f $X=4.305 $Y=0.235 $X2=0 $Y2=0
cc_319 N_Y_M1022_d N_VGND_c_636_n 0.00297142f $X=5.245 $Y=0.235 $X2=0 $Y2=0
cc_320 N_A_27_47#_c_541_n N_VGND_M1002_s 0.00500594f $X=1.035 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_321 N_A_27_47#_c_551_n N_VGND_M1015_s 0.00500594f $X=1.975 $Y=0.8 $X2=0 $Y2=0
cc_322 N_A_27_47#_c_559_n N_VGND_M1019_s 0.00500594f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_323 N_A_27_47#_c_541_n N_VGND_c_629_n 0.0199861f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_324 N_A_27_47#_c_541_n N_VGND_c_630_n 0.0020257f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_325 N_A_27_47#_c_547_n N_VGND_c_630_n 0.0188215f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_326 N_A_27_47#_c_551_n N_VGND_c_630_n 0.0020257f $X=1.975 $Y=0.8 $X2=0 $Y2=0
cc_327 N_A_27_47#_c_551_n N_VGND_c_631_n 0.0199861f $X=1.975 $Y=0.8 $X2=0 $Y2=0
cc_328 N_A_27_47#_c_551_n N_VGND_c_632_n 0.0020257f $X=1.975 $Y=0.8 $X2=0 $Y2=0
cc_329 N_A_27_47#_c_555_n N_VGND_c_632_n 0.0188215f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_330 N_A_27_47#_c_559_n N_VGND_c_632_n 0.0020257f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_331 N_A_27_47#_c_559_n N_VGND_c_633_n 0.0199861f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_332 N_A_27_47#_c_533_n N_VGND_c_634_n 0.0212882f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_333 N_A_27_47#_c_541_n N_VGND_c_634_n 0.0020257f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_334 N_A_27_47#_c_559_n N_VGND_c_635_n 0.0020257f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_335 N_A_27_47#_c_563_n N_VGND_c_635_n 0.0151813f $X=3.04 $Y=0.465 $X2=0 $Y2=0
cc_336 N_A_27_47#_c_574_n N_VGND_c_635_n 0.14729f $X=5.765 $Y=0.36 $X2=0 $Y2=0
cc_337 N_A_27_47#_c_538_n N_VGND_c_635_n 0.0190695f $X=5.9 $Y=0.38 $X2=0 $Y2=0
cc_338 N_A_27_47#_M1002_d N_VGND_c_636_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_339 N_A_27_47#_M1007_d N_VGND_c_636_n 0.00215201f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_340 N_A_27_47#_M1017_d N_VGND_c_636_n 0.00215201f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_341 N_A_27_47#_M1021_d N_VGND_c_636_n 0.00215206f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_342 N_A_27_47#_M1009_s N_VGND_c_636_n 0.00255381f $X=3.835 $Y=0.235 $X2=0
+ $Y2=0
cc_343 N_A_27_47#_M1013_s N_VGND_c_636_n 0.00215227f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_344 N_A_27_47#_M1023_s N_VGND_c_636_n 0.00209319f $X=5.765 $Y=0.235 $X2=0
+ $Y2=0
cc_345 N_A_27_47#_c_533_n N_VGND_c_636_n 0.0125939f $X=0.26 $Y=0.38 $X2=0 $Y2=0
cc_346 N_A_27_47#_c_541_n N_VGND_c_636_n 0.00880092f $X=1.035 $Y=0.8 $X2=0 $Y2=0
cc_347 N_A_27_47#_c_547_n N_VGND_c_636_n 0.0121968f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_348 N_A_27_47#_c_551_n N_VGND_c_636_n 0.00880092f $X=1.975 $Y=0.8 $X2=0 $Y2=0
cc_349 N_A_27_47#_c_555_n N_VGND_c_636_n 0.0121968f $X=2.14 $Y=0.38 $X2=0 $Y2=0
cc_350 N_A_27_47#_c_559_n N_VGND_c_636_n 0.00880092f $X=2.915 $Y=0.8 $X2=0 $Y2=0
cc_351 N_A_27_47#_c_563_n N_VGND_c_636_n 0.0093992f $X=3.04 $Y=0.465 $X2=0 $Y2=0
cc_352 N_A_27_47#_c_574_n N_VGND_c_636_n 0.092792f $X=5.765 $Y=0.36 $X2=0 $Y2=0
cc_353 N_A_27_47#_c_538_n N_VGND_c_636_n 0.0114921f $X=5.9 $Y=0.38 $X2=0 $Y2=0
