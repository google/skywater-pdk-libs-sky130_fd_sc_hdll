# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__probec_p_8
  CLASS CORE ;
  FOREIGN sky130_fd_sc_hdll__probec_p_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.832500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.140000 1.075000 1.240000 1.275000 ;
    END
  END A
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met5 ;
        RECT -1.260000 0.560000 1.060000 2.160000 ;
    END
  END X
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.930000 -0.895000 6.110000 0.285000 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360000 -1.170000 6.675000 -0.455000 ;
        RECT 4.360000 -0.155000 6.675000  0.560000 ;
        RECT 4.560000 -0.455000 6.675000 -0.155000 ;
    END
  END VGND
  PIN VNB
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER pwell ;
        RECT 0.150000 -0.085000 0.320000 0.085000 ;
    END
  END VNB
  PIN VPB
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT -0.190000 1.305000 6.170000 2.910000 ;
    END
  END VPB
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.930000 2.435000 6.110000 3.615000 ;
    END
    PORT
      LAYER met5 ;
        RECT 4.360000 2.160000 6.675000 2.875000 ;
        RECT 4.360000 3.175000 6.675000 3.890000 ;
        RECT 4.560000 2.875000 6.675000 3.175000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 5.980000 0.085000 ;
      RECT 0.000000  2.635000 5.980000 2.805000 ;
      RECT 0.095000  1.445000 1.595000 1.615000 ;
      RECT 0.095000  1.615000 0.425000 2.465000 ;
      RECT 0.145000  0.255000 0.445000 0.735000 ;
      RECT 0.145000  0.735000 1.595000 0.905000 ;
      RECT 0.595000  1.835000 0.865000 2.635000 ;
      RECT 0.615000  0.085000 0.895000 0.565000 ;
      RECT 1.035000  1.615000 1.365000 2.465000 ;
      RECT 1.065000  0.255000 1.335000 0.735000 ;
      RECT 1.420000  0.905000 1.595000 1.075000 ;
      RECT 1.420000  1.075000 4.045000 1.245000 ;
      RECT 1.420000  1.245000 1.595000 1.445000 ;
      RECT 1.505000  0.085000 1.805000 0.565000 ;
      RECT 1.535000  1.835000 1.805000 2.635000 ;
      RECT 1.975000  0.255000 2.305000 0.735000 ;
      RECT 1.975000  0.735000 5.125000 0.905000 ;
      RECT 1.975000  1.445000 5.125000 1.615000 ;
      RECT 1.975000  1.615000 2.305000 2.465000 ;
      RECT 2.475000  0.085000 2.745000 0.565000 ;
      RECT 2.475000  1.835000 2.745000 2.635000 ;
      RECT 2.915000  0.255000 3.245000 0.735000 ;
      RECT 2.915000  1.615000 3.245000 2.465000 ;
      RECT 3.415000  0.085000 3.685000 0.565000 ;
      RECT 3.415000  1.835000 3.685000 2.635000 ;
      RECT 3.855000  0.255000 4.185000 0.735000 ;
      RECT 3.855000  1.615000 4.185000 2.465000 ;
      RECT 4.290000  0.905000 5.125000 1.445000 ;
      RECT 4.355000  0.085000 4.625000 0.565000 ;
      RECT 4.355000  1.835000 4.625000 2.635000 ;
      RECT 4.795000  0.255000 5.125000 0.735000 ;
      RECT 4.795000  1.615000 5.125000 2.465000 ;
      RECT 5.295000  0.085000 5.545000 0.885000 ;
      RECT 5.295000  1.485000 5.595000 2.635000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
      RECT 4.285000 -0.085000 4.455000 0.085000 ;
      RECT 4.285000  2.635000 4.455000 2.805000 ;
      RECT 4.305000  1.105000 4.475000 1.275000 ;
      RECT 4.665000  1.105000 4.835000 1.275000 ;
      RECT 4.745000 -0.085000 4.915000 0.085000 ;
      RECT 4.745000  2.635000 4.915000 2.805000 ;
      RECT 5.205000 -0.085000 5.375000 0.085000 ;
      RECT 5.205000  2.635000 5.375000 2.805000 ;
      RECT 5.665000 -0.085000 5.835000 0.085000 ;
      RECT 5.665000  2.635000 5.835000 2.805000 ;
    LAYER met1 ;
      RECT 0.000000 -0.240000 5.980000 0.240000 ;
      RECT 0.000000  2.480000 5.980000 2.960000 ;
      RECT 2.020000  1.060000 2.660000 1.120000 ;
      RECT 2.020000  1.120000 4.895000 1.260000 ;
      RECT 2.020000  1.260000 2.660000 1.320000 ;
      RECT 4.245000  1.075000 4.895000 1.120000 ;
      RECT 4.245000  1.260000 4.895000 1.305000 ;
    LAYER met2 ;
      RECT 1.890000  1.050000 2.660000 1.330000 ;
      RECT 5.135000 -0.140000 5.905000 0.140000 ;
      RECT 5.135000  2.580000 5.905000 2.860000 ;
    LAYER met3 ;
      RECT -0.715000  1.030000 0.065000 1.350000 ;
      RECT  1.885000  1.025000 2.665000 1.355000 ;
      RECT  5.130000 -0.165000 5.910000 0.165000 ;
      RECT  5.130000  2.555000 5.910000 2.885000 ;
    LAYER met4 ;
      RECT -1.140000 0.770000 0.040000 1.950000 ;
      RECT  1.460000 0.770000 2.640000 1.950000 ;
    LAYER met5 ;
      RECT 1.160000 -1.105000 2.760000  3.825000 ;
      RECT 4.360000 -0.355000 4.460000 -0.255000 ;
      RECT 4.360000  2.975000 4.460000  3.075000 ;
    LAYER via ;
      RECT 2.050000  1.060000 2.310000 1.320000 ;
      RECT 2.370000  1.060000 2.630000 1.320000 ;
      RECT 5.230000 -0.130000 5.490000 0.130000 ;
      RECT 5.230000  2.590000 5.490000 2.850000 ;
      RECT 5.550000 -0.130000 5.810000 0.130000 ;
      RECT 5.550000  2.590000 5.810000 2.850000 ;
    LAYER via2 ;
      RECT 1.935000  1.050000 2.215000 1.330000 ;
      RECT 2.335000  1.050000 2.615000 1.330000 ;
      RECT 5.180000 -0.140000 5.460000 0.140000 ;
      RECT 5.180000  2.580000 5.460000 2.860000 ;
      RECT 5.580000 -0.140000 5.860000 0.140000 ;
      RECT 5.580000  2.580000 5.860000 2.860000 ;
    LAYER via3 ;
      RECT -0.685000  1.030000 -0.365000 1.350000 ;
      RECT -0.285000  1.030000  0.035000 1.350000 ;
      RECT  1.915000  1.030000  2.235000 1.350000 ;
      RECT  2.315000  1.030000  2.635000 1.350000 ;
      RECT  5.160000 -0.160000  5.480000 0.160000 ;
      RECT  5.160000  2.560000  5.480000 2.880000 ;
      RECT  5.560000 -0.160000  5.880000 0.160000 ;
      RECT  5.560000  2.560000  5.880000 2.880000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__probec_p_8
END LIBRARY
