* File: sky130_fd_sc_hdll__or4_1.spice
* Created: Wed Sep  2 08:49:12 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or4_1.pex.spice"
.subckt sky130_fd_sc_hdll__or4_1  VNB VPB D C B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* C	C
* D	D
* VPB	VPB
* VNB	VNB
MM1000 N_A_27_297#_M1000_d N_D_M1000_g N_VGND_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0798 AS=0.1302 PD=0.8 PS=1.46 NRD=7.14 NRS=12.852 M=1 R=2.8 SA=75000.2
+ SB=75002.4 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1005_d N_C_M1005_g N_A_27_297#_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0567 AS=0.0798 PD=0.69 PS=0.8 NRD=0 NRS=21.42 M=1 R=2.8 SA=75000.8
+ SB=75001.8 A=0.063 P=1.14 MULT=1
MM1007 N_A_27_297#_M1007_d N_B_M1007_g N_VGND_M1005_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0777 AS=0.0567 PD=0.79 PS=0.69 NRD=12.852 NRS=0 M=1 R=2.8 SA=75001.2
+ SB=75001.4 A=0.063 P=1.14 MULT=1
MM1002 N_VGND_M1002_d N_A_M1002_g N_A_27_297#_M1007_d VNB NSHORT L=0.15 W=0.42
+ AD=0.0927336 AS=0.0777 PD=0.816449 PS=0.79 NRD=12.852 NRS=12.852 M=1 R=2.8
+ SA=75001.7 SB=75000.9 A=0.063 P=1.14 MULT=1
MM1001 N_X_M1001_d N_A_27_297#_M1001_g N_VGND_M1002_d VNB NSHORT L=0.15 W=0.65
+ AD=0.273 AS=0.143516 PD=2.14 PS=1.26355 NRD=26.76 NRS=11.988 M=1 R=4.33333
+ SA=75001.5 SB=75000.3 A=0.0975 P=1.6 MULT=1
MM1003 A_117_297# N_D_M1003_g N_A_27_297#_M1003_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0735 AS=0.1134 PD=0.77 PS=1.38 NRD=56.2829 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90002.3 A=0.0756 P=1.2 MULT=1
MM1009 A_223_297# N_C_M1009_g A_117_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0504
+ AS=0.0735 PD=0.66 PS=0.77 NRD=30.4759 NRS=56.2829 M=1 R=2.33333 SA=90000.7
+ SB=90001.8 A=0.0756 P=1.2 MULT=1
MM1006 A_307_297# N_B_M1006_g A_223_297# VPB PHIGHVT L=0.18 W=0.42 AD=0.0714
+ AS=0.0504 PD=0.76 PS=0.66 NRD=53.9386 NRS=30.4759 M=1 R=2.33333 SA=90001.1
+ SB=90001.4 A=0.0756 P=1.2 MULT=1
MM1004 N_VPWR_M1004_d N_A_M1004_g A_307_297# VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0918972 AS=0.0714 PD=0.804507 PS=0.76 NRD=76.83 NRS=53.9386 M=1 R=2.33333
+ SA=90001.6 SB=90000.9 A=0.0756 P=1.2 MULT=1
MM1008 N_X_M1008_d N_A_27_297#_M1008_g N_VPWR_M1004_d VPB PHIGHVT L=0.18 W=1
+ AD=0.43 AS=0.218803 PD=2.86 PS=1.91549 NRD=30.535 NRS=1.9503 M=1 R=5.55556
+ SA=90001 SB=90000.3 A=0.18 P=2.36 MULT=1
DX10_noxref VNB VPB NWDIODE A=5.778 P=10.41
pX11_noxref noxref_14 C C PROBETYPE=1
pX12_noxref noxref_15 C C PROBETYPE=1
pX13_noxref noxref_16 B B PROBETYPE=1
pX14_noxref noxref_17 A A PROBETYPE=1
c_57 VPB 0 2.01548e-19 $X=0.15 $Y=2.635
*
.include "sky130_fd_sc_hdll__or4_1.pxi.spice"
*
.ends
*
*
