* File: sky130_fd_sc_hdll__and4bb_4.spice
* Created: Thu Aug 27 18:59:36 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__and4bb_4.pex.spice"
.subckt sky130_fd_sc_hdll__and4bb_4  VNB VPB B_N D C A_N VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A_N	A_N
* C	C
* D	D
* B_N	B_N
* VPB	VPB
* VNB	VNB
MM1014 N_VGND_M1014_d N_B_N_M1014_g N_A_27_47#_M1014_s VNB NSHORT L=0.15 W=0.42
+ AD=0.0761495 AS=0.1302 PD=0.765421 PS=1.46 NRD=14.28 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75004.3 A=0.063 P=1.14 MULT=1
MM1005 N_VGND_M1014_d N_A_184_21#_M1005_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.11785 AS=0.104 PD=1.18458 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.5 SB=75003.9 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1007_d N_A_184_21#_M1007_g N_X_M1005_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001
+ SB=75003.4 A=0.0975 P=1.6 MULT=1
MM1015 N_VGND_M1007_d N_A_184_21#_M1015_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75001.5
+ SB=75002.9 A=0.0975 P=1.6 MULT=1
MM1016 N_VGND_M1016_d N_A_184_21#_M1016_g N_X_M1015_s VNB NSHORT L=0.15 W=0.65
+ AD=0.13 AS=0.104 PD=1.05 PS=0.97 NRD=2.76 NRS=0 M=1 R=4.33333 SA=75001.9
+ SB=75002.5 A=0.0975 P=1.6 MULT=1
MM1000 A_606_47# N_D_M1000_g N_VGND_M1016_d VNB NSHORT L=0.15 W=0.65 AD=0.134875
+ AS=0.13 PD=1.065 PS=1.05 NRD=28.152 NRS=19.38 M=1 R=4.33333 SA=75002.5
+ SB=75001.9 A=0.0975 P=1.6 MULT=1
MM1017 A_719_47# N_C_M1017_g A_606_47# VNB NSHORT L=0.15 W=0.65 AD=0.141375
+ AS=0.134875 PD=1.085 PS=1.065 NRD=30 NRS=28.152 M=1 R=4.33333 SA=75003
+ SB=75001.3 A=0.0975 P=1.6 MULT=1
MM1009 A_836_47# N_A_27_47#_M1009_g A_719_47# VNB NSHORT L=0.15 W=0.65 AD=0.1235
+ AS=0.141375 PD=1.03 PS=1.085 NRD=24.912 NRS=30 M=1 R=4.33333 SA=75003.6
+ SB=75000.8 A=0.0975 P=1.6 MULT=1
MM1003 N_A_184_21#_M1003_d N_A_912_21#_M1003_g A_836_47# VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.1235 PD=1.92 PS=1.03 NRD=8.304 NRS=24.912 M=1 R=4.33333
+ SA=75004.2 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1012 N_A_912_21#_M1012_d N_A_N_M1012_g N_VGND_M1012_s VNB NSHORT L=0.15 W=0.42
+ AD=0.1302 AS=0.1932 PD=1.46 PS=1.76 NRD=12.852 NRS=44.28 M=1 R=2.8 SA=75000.4
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1002 N_VPWR_M1002_d N_B_N_M1002_g N_A_27_47#_M1002_s VPB PHIGHVT L=0.18 W=0.42
+ AD=0.0874606 AS=0.1134 PD=0.795634 PS=1.38 NRD=2.3443 NRS=2.3443 M=1 R=2.33333
+ SA=90000.2 SB=90005.6 A=0.0756 P=1.2 MULT=1
MM1008 N_VPWR_M1002_d N_A_184_21#_M1008_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.208239 AS=0.145 PD=1.89437 PS=1.29 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.4 SB=90004.4 A=0.18 P=2.36 MULT=1
MM1010 N_VPWR_M1010_d N_A_184_21#_M1010_g N_X_M1008_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.9 SB=90003.9 A=0.18 P=2.36 MULT=1
MM1013 N_VPWR_M1010_d N_A_184_21#_M1013_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.3 SB=90003.4 A=0.18 P=2.36 MULT=1
MM1019 N_VPWR_M1019_d N_A_184_21#_M1019_g N_X_M1013_s VPB PHIGHVT L=0.18 W=1
+ AD=0.185 AS=0.145 PD=1.37 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.8 SB=90002.9 A=0.18 P=2.36 MULT=1
MM1011 N_A_184_21#_M1011_d N_D_M1011_g N_VPWR_M1019_d VPB PHIGHVT L=0.18 W=1
+ AD=0.1925 AS=0.185 PD=1.385 PS=1.37 NRD=12.7853 NRS=16.7253 M=1 R=5.55556
+ SA=90002.4 SB=90002.4 A=0.18 P=2.36 MULT=1
MM1006 N_VPWR_M1006_d N_C_M1006_g N_A_184_21#_M1011_d VPB PHIGHVT L=0.18 W=1
+ AD=0.2025 AS=0.1925 PD=1.405 PS=1.385 NRD=13.7703 NRS=7.8603 M=1 R=5.55556
+ SA=90002.9 SB=90001.8 A=0.18 P=2.36 MULT=1
MM1004 N_A_184_21#_M1004_d N_A_27_47#_M1004_g N_VPWR_M1006_d VPB PHIGHVT L=0.18
+ W=1 AD=0.175 AS=0.2025 PD=1.35 PS=1.405 NRD=4.9053 NRS=10.8153 M=1 R=5.55556
+ SA=90003.5 SB=90001.2 A=0.18 P=2.36 MULT=1
MM1018 N_VPWR_M1018_d N_A_912_21#_M1018_g N_A_184_21#_M1004_d VPB PHIGHVT L=0.18
+ W=1 AD=0.437113 AS=0.175 PD=2.96479 PS=1.35 NRD=16.7253 NRS=8.8453 M=1
+ R=5.55556 SA=90004 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1001 N_A_912_21#_M1001_d N_A_N_M1001_g N_VPWR_M1018_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.183587 PD=1.38 PS=1.24521 NRD=2.3443 NRS=28.1316 M=1
+ R=2.33333 SA=90005.6 SB=90000.2 A=0.0756 P=1.2 MULT=1
DX20_noxref VNB VPB NWDIODE A=10.9461 P=16.85
pX21_noxref noxref_16 A_N A_N PROBETYPE=1
pX22_noxref noxref_17 A_N A_N PROBETYPE=1
*
.include "sky130_fd_sc_hdll__and4bb_4.pxi.spice"
*
.ends
*
*
