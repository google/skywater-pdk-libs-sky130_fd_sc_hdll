* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__sdlclkp_4 CLK GATE SCE VGND VNB VPB VPWR GCLK
X0 VPWR SCE a_117_369# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X1 a_1217_47# CLK VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X2 a_421_413# a_505_315# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X3 GCLK a_1125_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X4 GCLK a_1125_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 VGND a_1125_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X6 VPWR a_1125_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X7 VGND GATE a_27_47# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X8 VGND a_1125_47# GCLK VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X9 a_1125_47# a_505_315# a_1217_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X10 VGND CLK a_280_21# VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X11 VPWR a_310_47# a_505_315# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X12 a_27_47# SCE VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X13 VPWR CLK a_280_21# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X14 a_117_369# GATE a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X15 GCLK a_1125_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X16 GCLK a_1125_47# VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X17 a_310_47# a_280_21# a_421_413# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
X18 a_425_47# a_505_315# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X19 a_277_243# a_280_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=640000u l=180000u
X20 a_277_243# a_280_21# VGND VNB sky130_fd_pr__nfet_01v8 w=420000u l=150000u
X21 a_1125_47# CLK VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X22 a_27_47# a_280_21# a_310_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X23 VPWR a_1125_47# GCLK VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 a_310_47# a_277_243# a_425_47# VNB sky130_fd_pr__nfet_01v8 w=360000u l=150000u
X25 VGND a_310_47# a_505_315# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X26 VPWR a_505_315# a_1125_47# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X27 a_27_47# a_277_243# a_310_47# VPB sky130_fd_pr__pfet_01v8_hvt w=420000u l=180000u
.ends
