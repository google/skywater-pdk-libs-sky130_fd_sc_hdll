* Copyright 2020 The SkyWater PDK Authors
*
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0


.subckt sky130_fd_sc_hdll__xnor2_4 A B VGND VNB VPB VPWR Y
X0 Y B a_898_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X1 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X2 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X3 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X4 a_898_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X5 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X6 VGND A a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X7 VGND A a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X8 Y a_38_297# VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X9 a_898_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X10 VGND A a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X11 VGND B a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X12 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X13 VPWR A a_898_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X14 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X15 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X16 VPWR B a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X17 a_980_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X18 VGND B a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X19 Y B a_898_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X20 a_980_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X21 Y a_38_297# a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X22 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X23 a_898_297# B Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X24 Y a_38_297# a_980_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X25 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X26 a_980_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X27 a_980_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X28 a_38_297# B VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X29 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X30 a_38_47# A VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X31 VPWR A a_898_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X32 a_38_297# B a_38_47# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X33 a_980_47# B VGND VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X34 a_38_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X35 a_898_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X36 a_38_47# B a_38_297# VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
X37 VPWR a_38_297# Y VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X38 VPWR A a_38_297# VPB sky130_fd_pr__pfet_01v8_hvt w=1e+06u l=180000u
X39 a_980_47# a_38_297# Y VNB sky130_fd_pr__nfet_01v8 w=650000u l=150000u
.ends
