* File: sky130_fd_sc_hdll__mux2i_2.pex.spice
* Created: Thu Aug 27 19:11:08 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%S 1 3 4 6 7 9 10 12 13 15 16 18 19 20 30
r67 30 31 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=1.435 $Y=1.202
+ $X2=1.46 $Y2=1.202
r68 29 30 57.3503 $w=3.74e-07 $l=4.45e-07 $layer=POLY_cond $X=0.99 $Y=1.202
+ $X2=1.435 $Y2=1.202
r69 28 29 3.22193 $w=3.74e-07 $l=2.5e-08 $layer=POLY_cond $X=0.965 $Y=1.202
+ $X2=0.99 $Y2=1.202
r70 27 28 57.3503 $w=3.74e-07 $l=4.45e-07 $layer=POLY_cond $X=0.52 $Y=1.202
+ $X2=0.965 $Y2=1.202
r71 25 27 0.644385 $w=3.74e-07 $l=5e-09 $layer=POLY_cond $X=0.515 $Y=1.202
+ $X2=0.52 $Y2=1.202
r72 25 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.515
+ $Y=1.16 $X2=0.515 $Y2=1.16
r73 23 25 2.57754 $w=3.74e-07 $l=2e-08 $layer=POLY_cond $X=0.495 $Y=1.202
+ $X2=0.515 $Y2=1.202
r74 20 26 1.18065 $w=3.1e-07 $l=3e-08 $layer=LI1_cond $X=0.63 $Y=1.19 $X2=0.63
+ $Y2=1.16
r75 19 26 12.2 $w=3.1e-07 $l=3.1e-07 $layer=LI1_cond $X=0.63 $Y=0.85 $X2=0.63
+ $Y2=1.16
r76 16 31 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=1.202
r77 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.46 $Y=0.995
+ $X2=1.46 $Y2=0.56
r78 13 30 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.202
r79 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.435 $Y=1.41
+ $X2=1.435 $Y2=1.985
r80 10 29 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=1.202
r81 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.99 $Y=0.995
+ $X2=0.99 $Y2=0.56
r82 7 28 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.202
r83 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r84 4 27 24.2268 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.52 $Y2=1.202
r85 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r86 1 23 19.8678 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.202
r87 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A_27_47# 1 2 7 9 12 14 16 19 22 25 28 30
+ 32 35 37 38 41 43 48
c96 30 0 1.34758e-19 $X=1.545 $Y=1.24
c97 14 0 1.40621e-19 $X=2.375 $Y=1.41
r98 48 49 3.45272 $w=3.49e-07 $l=2.5e-08 $layer=POLY_cond $X=2.375 $Y=1.217
+ $X2=2.4 $Y2=1.217
r99 45 46 3.45272 $w=3.49e-07 $l=2.5e-08 $layer=POLY_cond $X=1.905 $Y=1.217
+ $X2=1.93 $Y2=1.217
r100 42 48 55.9341 $w=3.49e-07 $l=4.05e-07 $layer=POLY_cond $X=1.97 $Y=1.217
+ $X2=2.375 $Y2=1.217
r101 42 46 5.52436 $w=3.49e-07 $l=4e-08 $layer=POLY_cond $X=1.97 $Y=1.217
+ $X2=1.93 $Y2=1.217
r102 41 43 8.79328 $w=2.48e-07 $l=1.65e-07 $layer=LI1_cond $X=1.97 $Y=1.2
+ $X2=1.805 $Y2=1.2
r103 41 42 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r104 37 38 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=2.3
+ $X2=0.215 $Y2=2.135
r105 32 34 8.55024 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=0.215 $Y=0.51
+ $X2=0.215 $Y2=0.675
r106 30 43 16.9626 $w=1.68e-07 $l=2.6e-07 $layer=LI1_cond $X=1.545 $Y=1.24
+ $X2=1.805 $Y2=1.24
r107 27 30 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.435 $Y=1.325
+ $X2=1.545 $Y2=1.24
r108 27 28 8.90524 $w=2.18e-07 $l=1.7e-07 $layer=LI1_cond $X=1.435 $Y=1.325
+ $X2=1.435 $Y2=1.495
r109 26 35 1.44715 $w=1.7e-07 $l=8.8e-08 $layer=LI1_cond $X=0.26 $Y=1.58
+ $X2=0.172 $Y2=1.58
r110 25 28 6.96323 $w=1.7e-07 $l=1.46458e-07 $layer=LI1_cond $X=1.325 $Y=1.58
+ $X2=1.435 $Y2=1.495
r111 25 26 69.4813 $w=1.68e-07 $l=1.065e-06 $layer=LI1_cond $X=1.325 $Y=1.58
+ $X2=0.26 $Y2=1.58
r112 23 35 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.172 $Y=1.665
+ $X2=0.172 $Y2=1.58
r113 23 38 29.787 $w=1.73e-07 $l=4.7e-07 $layer=LI1_cond $X=0.172 $Y=1.665
+ $X2=0.172 $Y2=2.135
r114 22 35 5.04255 $w=1.75e-07 $l=8.5e-08 $layer=LI1_cond $X=0.172 $Y=1.495
+ $X2=0.172 $Y2=1.58
r115 22 34 51.9688 $w=1.73e-07 $l=8.2e-07 $layer=LI1_cond $X=0.172 $Y=1.495
+ $X2=0.172 $Y2=0.675
r116 17 49 22.56 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=2.4 $Y=1.025 $X2=2.4
+ $Y2=1.217
r117 17 19 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=2.4 $Y=1.025
+ $X2=2.4 $Y2=0.56
r118 14 48 18.24 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.217
r119 14 16 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.375 $Y=1.41
+ $X2=2.375 $Y2=1.985
r120 10 46 22.56 $w=1.5e-07 $l=1.92e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=1.217
r121 10 12 238.436 $w=1.5e-07 $l=4.65e-07 $layer=POLY_cond $X=1.93 $Y=1.025
+ $X2=1.93 $Y2=0.56
r122 7 45 18.24 $w=1.8e-07 $l=1.93e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.217
r123 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.905 $Y=1.41
+ $X2=1.905 $Y2=1.985
r124 2 37 600 $w=1.7e-07 $l=8.75271e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.3
r125 1 32 182 $w=1.7e-07 $l=3.31662e-07 $layer=licon1_NDIFF $count=1 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.51
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A0 1 3 4 6 7 9 10 12 13 14 15 19 29 34 36
+ 40
r54 34 36 22.7364 $w=1.98e-07 $l=4.1e-07 $layer=LI1_cond $X=3.015 $Y=1.175
+ $X2=3.425 $Y2=1.175
r55 29 30 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=3.835 $Y=1.202
+ $X2=3.86 $Y2=1.202
r56 28 40 15.8045 $w=1.98e-07 $l=2.85e-07 $layer=LI1_cond $X=3.615 $Y=1.175
+ $X2=3.9 $Y2=1.175
r57 27 29 28.0529 $w=3.78e-07 $l=2.2e-07 $layer=POLY_cond $X=3.615 $Y=1.202
+ $X2=3.835 $Y2=1.202
r58 27 28 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=3.615
+ $Y=1.16 $X2=3.615 $Y2=1.16
r59 25 27 28.6905 $w=3.78e-07 $l=2.25e-07 $layer=POLY_cond $X=3.39 $Y=1.202
+ $X2=3.615 $Y2=1.202
r60 24 25 3.18783 $w=3.78e-07 $l=2.5e-08 $layer=POLY_cond $X=3.365 $Y=1.202
+ $X2=3.39 $Y2=1.202
r61 19 24 14.9401 $w=3.78e-07 $l=1.253e-07 $layer=POLY_cond $X=3.265 $Y=1.145
+ $X2=3.365 $Y2=1.202
r62 19 21 75.9834 $w=3e-07 $l=3.8e-07 $layer=POLY_cond $X=3.265 $Y=1.145
+ $X2=2.885 $Y2=1.145
r63 15 40 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.905 $Y=1.175
+ $X2=3.9 $Y2=1.175
r64 14 28 10.2591 $w=1.98e-07 $l=1.85e-07 $layer=LI1_cond $X=3.43 $Y=1.175
+ $X2=3.615 $Y2=1.175
r65 14 36 0.277273 $w=1.98e-07 $l=5e-09 $layer=LI1_cond $X=3.43 $Y=1.175
+ $X2=3.425 $Y2=1.175
r66 13 34 7.20909 $w=1.98e-07 $l=1.3e-07 $layer=LI1_cond $X=2.885 $Y=1.175
+ $X2=3.015 $Y2=1.175
r67 13 21 96.8533 $w=1.7e-07 $l=2.55e-07 $layer=licon1_POLY $count=1 $X=2.885
+ $Y=1.16 $X2=2.885 $Y2=1.16
r68 10 30 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=1.202
r69 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.86 $Y=0.995
+ $X2=3.86 $Y2=0.56
r70 7 29 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.202
r71 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.835 $Y=1.41
+ $X2=3.835 $Y2=1.985
r72 4 25 24.4846 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.39 $Y=0.995
+ $X2=3.39 $Y2=1.202
r73 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.39 $Y=0.995 $X2=3.39
+ $Y2=0.56
r74 1 24 20.1192 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.202
r75 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.365 $Y=1.41
+ $X2=3.365 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A1 1 3 4 6 7 9 10 12 13 14 20 23
r43 22 23 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.95
+ $Y=1.16 $X2=4.95 $Y2=1.16
r44 20 22 17.0736 $w=3.67e-07 $l=1.3e-07 $layer=POLY_cond $X=4.82 $Y=1.202
+ $X2=4.95 $Y2=1.202
r45 19 20 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.795 $Y=1.202
+ $X2=4.82 $Y2=1.202
r46 18 19 59.1008 $w=3.67e-07 $l=4.5e-07 $layer=POLY_cond $X=4.345 $Y=1.202
+ $X2=4.795 $Y2=1.202
r47 17 18 3.28338 $w=3.67e-07 $l=2.5e-08 $layer=POLY_cond $X=4.32 $Y=1.202
+ $X2=4.345 $Y2=1.202
r48 13 14 10.4488 $w=3.73e-07 $l=3.4e-07 $layer=LI1_cond $X=4.897 $Y=1.19
+ $X2=4.897 $Y2=1.53
r49 13 23 0.921954 $w=3.73e-07 $l=3e-08 $layer=LI1_cond $X=4.897 $Y=1.19
+ $X2=4.897 $Y2=1.16
r50 10 20 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.202
r51 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.82 $Y=1.41
+ $X2=4.82 $Y2=1.985
r52 7 19 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.795 $Y=0.995
+ $X2=4.795 $Y2=1.202
r53 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.795 $Y=0.995
+ $X2=4.795 $Y2=0.56
r54 4 18 19.4219 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.345 $Y=1.41
+ $X2=4.345 $Y2=1.202
r55 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.345 $Y=1.41
+ $X2=4.345 $Y2=1.985
r56 1 17 23.77 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.32 $Y=0.995 $X2=4.32
+ $Y2=1.202
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.32 $Y=0.995 $X2=4.32
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%VPWR 1 2 3 10 14 16 18 23 33 34 37 44 51
r71 51 52 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r72 48 52 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=2.72
+ $X2=2.53 $Y2=2.72
r73 47 48 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r74 44 47 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=1.645 $Y=2.34
+ $X2=1.645 $Y2=2.72
r75 40 41 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=2.72
+ $X2=0.69 $Y2=2.72
r76 37 40 11.5244 $w=3.78e-07 $l=3.8e-07 $layer=LI1_cond $X=0.705 $Y=2.34
+ $X2=0.705 $Y2=2.72
r77 33 34 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r78 31 34 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r79 31 52 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=2.72
+ $X2=2.53 $Y2=2.72
r80 30 33 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=2.72
+ $X2=5.29 $Y2=2.72
r81 30 31 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=2.72
+ $X2=2.99 $Y2=2.72
r82 28 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.65 $Y2=2.72
r83 28 30 14.0267 $w=1.68e-07 $l=2.15e-07 $layer=LI1_cond $X=2.775 $Y=2.72
+ $X2=2.99 $Y2=2.72
r84 27 48 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=1.61 $Y2=2.72
r85 27 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=0.69 $Y2=2.72
r86 26 27 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 24 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=0.705 $Y2=2.72
r88 24 26 16.6364 $w=1.68e-07 $l=2.55e-07 $layer=LI1_cond $X=0.895 $Y=2.72
+ $X2=1.15 $Y2=2.72
r89 23 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.645 $Y2=2.72
r90 23 26 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=1.455 $Y=2.72
+ $X2=1.15 $Y2=2.72
r91 18 40 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.705 $Y2=2.72
r92 18 20 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=2.72
+ $X2=0.23 $Y2=2.72
r93 16 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=0.69 $Y2=2.72
r94 16 20 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r95 12 51 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=2.65 $Y=2.635
+ $X2=2.65 $Y2=2.72
r96 12 14 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=2.65 $Y=2.635
+ $X2=2.65 $Y2=2.34
r97 11 47 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.835 $Y=2.72
+ $X2=1.645 $Y2=2.72
r98 10 51 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=2.65 $Y2=2.72
r99 10 11 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.525 $Y=2.72
+ $X2=1.835 $Y2=2.72
r100 3 14 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=2.465
+ $Y=1.485 $X2=2.61 $Y2=2.34
r101 2 44 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=1.525
+ $Y=1.485 $X2=1.67 $Y2=2.34
r102 1 37 600 $w=1.7e-07 $l=9.24662e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A_211_297# 1 2 7 12 14 16 17
c47 7 0 1.40621e-19 $X=1.715 $Y=1.92
r48 16 17 11.8878 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=3.6 $Y=1.605
+ $X2=3.385 $Y2=1.605
r49 14 17 97.861 $w=1.68e-07 $l=1.5e-06 $layer=LI1_cond $X=1.885 $Y=1.58
+ $X2=3.385 $Y2=1.58
r50 11 14 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.8 $Y=1.665
+ $X2=1.885 $Y2=1.58
r51 11 12 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=1.8 $Y=1.665 $X2=1.8
+ $Y2=1.835
r52 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=1.715 $Y=1.92
+ $X2=1.8 $Y2=1.835
r53 7 9 33.5989 $w=1.68e-07 $l=5.15e-07 $layer=LI1_cond $X=1.715 $Y=1.92 $X2=1.2
+ $Y2=1.92
r54 2 16 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=3.455
+ $Y=1.485 $X2=3.6 $Y2=1.63
r55 1 9 600 $w=1.7e-07 $l=5.02295e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.92
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A_399_297# 1 2 11 13 16 17
r36 16 17 7.83661 $w=2.48e-07 $l=1.7e-07 $layer=LI1_cond $X=2.965 $Y=1.96
+ $X2=3.135 $Y2=1.96
r37 13 15 23.4141 $w=1.98e-07 $l=3.8e-07 $layer=LI1_cond $X=2.167 $Y=1.92
+ $X2=2.167 $Y2=2.3
r38 11 17 94.5989 $w=1.68e-07 $l=1.45e-06 $layer=LI1_cond $X=4.585 $Y=2
+ $X2=3.135 $Y2=2
r39 8 13 1.63057 $w=1.7e-07 $l=1.13e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=2.167 $Y2=1.92
r40 8 16 44.6898 $w=1.68e-07 $l=6.85e-07 $layer=LI1_cond $X=2.28 $Y=1.92
+ $X2=2.965 $Y2=1.92
r41 2 11 600 $w=1.7e-07 $l=5.85214e-07 $layer=licon1_PDIFF $count=1 $X=4.435
+ $Y=1.485 $X2=4.585 $Y2=2
r42 1 15 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.995
+ $Y=1.485 $X2=2.14 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%Y 1 2 3 4 5 6 19 28 29 37 41 56
r55 47 49 63.2834 $w=1.68e-07 $l=9.7e-07 $layer=LI1_cond $X=4.09 $Y=2.34
+ $X2=5.06 $Y2=2.34
r56 44 47 62.631 $w=1.68e-07 $l=9.6e-07 $layer=LI1_cond $X=3.13 $Y=2.34 $X2=4.09
+ $Y2=2.34
r57 37 41 2.30489 $w=2.23e-07 $l=4.5e-08 $layer=LI1_cond $X=5.312 $Y=2.255
+ $X2=5.312 $Y2=2.21
r58 36 56 1.38293 $w=2.23e-07 $l=2.7e-08 $layer=LI1_cond $X=5.312 $Y=1.897
+ $X2=5.312 $Y2=1.87
r59 29 37 3.0159 $w=2.25e-07 $l=8.5e-08 $layer=LI1_cond $X=5.312 $Y=2.34
+ $X2=5.312 $Y2=2.255
r60 29 49 7.82882 $w=2.08e-07 $l=1.4e-07 $layer=LI1_cond $X=5.2 $Y=2.34 $X2=5.06
+ $Y2=2.34
r61 29 41 1.02439 $w=2.23e-07 $l=2e-08 $layer=LI1_cond $X=5.312 $Y=2.19
+ $X2=5.312 $Y2=2.21
r62 28 56 1.48537 $w=2.23e-07 $l=2.9e-08 $layer=LI1_cond $X=5.312 $Y=1.841
+ $X2=5.312 $Y2=1.87
r63 28 29 13.522 $w=2.23e-07 $l=2.64e-07 $layer=LI1_cond $X=5.312 $Y=1.926
+ $X2=5.312 $Y2=2.19
r64 28 36 1.48537 $w=2.23e-07 $l=2.9e-08 $layer=LI1_cond $X=5.312 $Y=1.926
+ $X2=5.312 $Y2=1.897
r65 27 28 54.6137 $w=2.83e-07 $l=1.32e-06 $layer=LI1_cond $X=5.34 $Y=0.465
+ $X2=5.34 $Y2=1.785
r66 24 26 76.984 $w=1.68e-07 $l=1.18e-06 $layer=LI1_cond $X=4.07 $Y=0.38
+ $X2=5.25 $Y2=0.38
r67 21 24 61.3262 $w=1.68e-07 $l=9.4e-07 $layer=LI1_cond $X=3.13 $Y=0.38
+ $X2=4.07 $Y2=0.38
r68 19 27 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=5.255 $Y=0.38
+ $X2=5.34 $Y2=0.465
r69 19 26 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=5.255 $Y=0.38
+ $X2=5.25 $Y2=0.38
r70 6 49 600 $w=1.7e-07 $l=9.26971e-07 $layer=licon1_PDIFF $count=1 $X=4.91
+ $Y=1.485 $X2=5.06 $Y2=2.34
r71 5 47 600 $w=1.7e-07 $l=9.33863e-07 $layer=licon1_PDIFF $count=1 $X=3.925
+ $Y=1.485 $X2=4.09 $Y2=2.34
r72 4 44 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=3.005
+ $Y=1.485 $X2=3.13 $Y2=2.34
r73 3 26 182 $w=1.7e-07 $l=4.46654e-07 $layer=licon1_NDIFF $count=1 $X=4.87
+ $Y=0.235 $X2=5.25 $Y2=0.38
r74 2 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=3.935
+ $Y=0.235 $X2=4.07 $Y2=0.38
r75 1 21 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=3.005
+ $Y=0.235 $X2=3.13 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%VGND 1 2 3 12 14 18 20 24 26 28 38 39 42
+ 45 48
r74 48 49 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r75 46 49 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.61 $Y=0 $X2=2.53
+ $Y2=0
r76 45 46 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=0 $X2=1.61
+ $Y2=0
r77 43 46 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.69 $Y=0 $X2=1.61
+ $Y2=0
r78 42 43 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r79 38 39 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=5.29 $Y=0 $X2=5.29
+ $Y2=0
r80 36 39 0.654446 $w=4.8e-07 $l=2.3e-06 $layer=MET1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r81 36 49 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.99 $Y=0 $X2=2.53
+ $Y2=0
r82 35 38 150.053 $w=1.68e-07 $l=2.3e-06 $layer=LI1_cond $X=2.99 $Y=0 $X2=5.29
+ $Y2=0
r83 35 36 3.1 $w=1.7e-07 $l=5.1e-07 $layer=mcon $count=3 $X=2.99 $Y=0 $X2=2.99
+ $Y2=0
r84 33 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.61
+ $Y2=0
r85 33 35 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.695 $Y=0 $X2=2.99
+ $Y2=0
r86 28 42 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.7
+ $Y2=0
r87 28 30 18.5936 $w=1.68e-07 $l=2.85e-07 $layer=LI1_cond $X=0.515 $Y=0 $X2=0.23
+ $Y2=0
r88 26 43 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r89 26 30 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r90 22 48 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0
r91 22 24 19.246 $w=1.68e-07 $l=2.95e-07 $layer=LI1_cond $X=2.61 $Y=0.085
+ $X2=2.61 $Y2=0.38
r92 21 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.835 $Y=0 $X2=1.71
+ $Y2=0
r93 20 48 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.525 $Y=0 $X2=2.61
+ $Y2=0
r94 20 21 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=2.525 $Y=0 $X2=1.835
+ $Y2=0
r95 16 45 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0
r96 16 18 13.5988 $w=2.48e-07 $l=2.95e-07 $layer=LI1_cond $X=1.71 $Y=0.085
+ $X2=1.71 $Y2=0.38
r97 15 42 9.31531 $w=1.7e-07 $l=1.85e-07 $layer=LI1_cond $X=0.885 $Y=0 $X2=0.7
+ $Y2=0
r98 14 45 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=1.71
+ $Y2=0
r99 14 15 45.6684 $w=1.68e-07 $l=7e-07 $layer=LI1_cond $X=1.585 $Y=0 $X2=0.885
+ $Y2=0
r100 10 42 1.24149 $w=3.7e-07 $l=8.5e-08 $layer=LI1_cond $X=0.7 $Y=0.085 $X2=0.7
+ $Y2=0
r101 10 12 9.1884 $w=3.68e-07 $l=2.95e-07 $layer=LI1_cond $X=0.7 $Y=0.085
+ $X2=0.7 $Y2=0.38
r102 3 24 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=2.475
+ $Y=0.235 $X2=2.61 $Y2=0.38
r103 2 18 91 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=2 $X=1.535
+ $Y=0.235 $X2=1.67 $Y2=0.38
r104 1 12 182 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_NDIFF $count=1 $X=0.595
+ $Y=0.235 $X2=0.73 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A_213_47# 1 2 7 8 14 15 18
c64 7 0 1.45015e-19 $X=4.14 $Y=0.85
r65 15 23 15.5801 $w=2.31e-07 $l=2.95e-07 $layer=LI1_cond $X=4.285 $Y=0.795
+ $X2=4.58 $Y2=0.795
r66 14 15 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=4.285 $Y=0.85
+ $X2=4.285 $Y2=0.85
r67 10 18 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=1.255 $Y=0.85
+ $X2=1.255 $Y2=0.85
r68 8 10 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=1.4 $Y=0.85
+ $X2=1.255 $Y2=0.85
r69 7 14 0.115467 $w=2.3e-07 $l=1.45e-07 $layer=MET1_cond $X=4.14 $Y=0.85
+ $X2=4.285 $Y2=0.85
r70 7 8 3.39108 $w=1.4e-07 $l=2.74e-06 $layer=MET1_cond $X=4.14 $Y=0.85 $X2=1.4
+ $Y2=0.85
r71 2 23 182 $w=1.7e-07 $l=5.90297e-07 $layer=licon1_NDIFF $count=1 $X=4.395
+ $Y=0.235 $X2=4.58 $Y2=0.74
r72 1 18 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=1.065
+ $Y=0.235 $X2=1.2 $Y2=0.74
.ends

.subckt PM_SKY130_FD_SC_HDLL__MUX2I_2%A_401_47# 1 2 9 12 14 15
c37 2 0 1.45015e-19 $X=3.465 $Y=0.235
r38 14 15 11.0982 $w=2.48e-07 $l=2.15e-07 $layer=LI1_cond $X=3.6 $Y=0.78
+ $X2=3.385 $Y2=0.78
r39 12 15 75.6791 $w=1.68e-07 $l=1.16e-06 $layer=LI1_cond $X=2.225 $Y=0.82
+ $X2=3.385 $Y2=0.82
r40 7 12 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.225 $Y2=0.82
r41 7 9 17.9412 $w=1.68e-07 $l=2.75e-07 $layer=LI1_cond $X=2.14 $Y=0.735
+ $X2=2.14 $Y2=0.46
r42 2 14 182 $w=1.7e-07 $l=5.68507e-07 $layer=licon1_NDIFF $count=1 $X=3.465
+ $Y=0.235 $X2=3.6 $Y2=0.74
r43 1 9 182 $w=1.7e-07 $l=2.84605e-07 $layer=licon1_NDIFF $count=1 $X=2.005
+ $Y=0.235 $X2=2.14 $Y2=0.46
.ends

