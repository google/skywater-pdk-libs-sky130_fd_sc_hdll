* File: sky130_fd_sc_hdll__o2bb2ai_2.pex.spice
* Created: Thu Aug 27 19:22:11 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A1_N 1 3 4 6 7 9 10 12 13 16 21 30 32
c70 32 0 1.43188e-19 $X=0.675 $Y=1.345
c71 4 0 1.20797e-19 $X=0.54 $Y=0.995
r72 30 32 12.3152 $w=5.38e-07 $l=2.8e-07 $layer=LI1_cond $X=0.395 $Y=1.345
+ $X2=0.675 $Y2=1.345
r73 24 30 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.48
+ $Y=1.16 $X2=0.48 $Y2=1.16
r74 21 30 3.54394 $w=5.38e-07 $l=1.6e-07 $layer=LI1_cond $X=0.235 $Y=1.345
+ $X2=0.395 $Y2=1.345
r75 16 19 11.2212 $w=3.78e-07 $l=3.7e-07 $layer=LI1_cond $X=1.955 $Y=1.16
+ $X2=1.955 $Y2=1.53
r76 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.97
+ $Y=1.16 $X2=1.97 $Y2=1.16
r77 13 19 5.46774 $w=1.7e-07 $l=1.9e-07 $layer=LI1_cond $X=1.765 $Y=1.53
+ $X2=1.955 $Y2=1.53
r78 13 32 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=1.765 $Y=1.53
+ $X2=0.675 $Y2=1.53
r79 10 17 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.97 $Y2=1.16
r80 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.935 $Y=1.41
+ $X2=1.935 $Y2=1.985
r81 7 17 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.91 $Y=0.995
+ $X2=1.97 $Y2=1.16
r82 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.91 $Y=0.995 $X2=1.91
+ $Y2=0.56
r83 4 24 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.54 $Y=0.995
+ $X2=0.48 $Y2=1.16
r84 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.54 $Y=0.995 $X2=0.54
+ $Y2=0.56
r85 1 24 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.48 $Y2=1.16
r86 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.515 $Y=1.41
+ $X2=0.515 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A2_N 1 3 4 6 7 9 10 12 13 20
c44 1 0 6.98311e-20 $X=0.96 $Y=0.995
r45 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=1.455 $Y=1.202
+ $X2=1.48 $Y2=1.202
r46 18 20 30.4421 $w=3.8e-07 $l=2.4e-07 $layer=POLY_cond $X=1.215 $Y=1.202
+ $X2=1.455 $Y2=1.202
r47 16 18 29.1737 $w=3.8e-07 $l=2.3e-07 $layer=POLY_cond $X=0.985 $Y=1.202
+ $X2=1.215 $Y2=1.202
r48 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=0.96 $Y=1.202
+ $X2=0.985 $Y2=1.202
r49 13 18 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.215
+ $Y=1.16 $X2=1.215 $Y2=1.16
r50 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=1.202
r51 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.48 $Y=0.995
+ $X2=1.48 $Y2=0.56
r52 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.202
r53 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.455 $Y=1.41
+ $X2=1.455 $Y2=1.985
r54 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.202
r55 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.985 $Y=1.41
+ $X2=0.985 $Y2=1.985
r56 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=0.96 $Y=0.995
+ $X2=0.96 $Y2=1.202
r57 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.96 $Y=0.995 $X2=0.96
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_121_297# 1 2 3 10 12 13 15 16 18 19 21
+ 24 28 30 31 33 37 45
c95 37 0 1.20797e-19 $X=1.385 $Y=0.775
c96 19 0 1.98409e-19 $X=3.37 $Y=0.995
c97 2 0 1.43188e-19 $X=0.605 $Y=1.485
r98 45 46 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=3.345 $Y=1.202
+ $X2=3.37 $Y2=1.202
r99 44 45 58.7644 $w=3.65e-07 $l=4.45e-07 $layer=POLY_cond $X=2.9 $Y=1.202
+ $X2=3.345 $Y2=1.202
r100 43 44 3.30137 $w=3.65e-07 $l=2.5e-08 $layer=POLY_cond $X=2.875 $Y=1.202
+ $X2=2.9 $Y2=1.202
r101 41 43 31.0329 $w=3.65e-07 $l=2.35e-07 $layer=POLY_cond $X=2.64 $Y=1.202
+ $X2=2.875 $Y2=1.202
r102 40 41 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.64
+ $Y=1.16 $X2=2.64 $Y2=1.16
r103 35 37 8.41541 $w=2.58e-07 $l=1.65e-07 $layer=LI1_cond $X=1.22 $Y=0.775
+ $X2=1.385 $Y2=0.775
r104 30 40 8.97739 $w=3.02e-07 $l=2.16852e-07 $layer=LI1_cond $X=2.4 $Y=1.325
+ $X2=2.52 $Y2=1.16
r105 30 31 30.0107 $w=1.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.4 $Y=1.325
+ $X2=2.4 $Y2=1.785
r106 28 40 13.9371 $w=3.02e-07 $l=4.35603e-07 $layer=LI1_cond $X=2.315 $Y=0.815
+ $X2=2.52 $Y2=1.16
r107 28 37 57.303 $w=1.78e-07 $l=9.3e-07 $layer=LI1_cond $X=2.315 $Y=0.815
+ $X2=1.385 $Y2=0.815
r108 25 33 4.10122 $w=1.8e-07 $l=1.25e-07 $layer=LI1_cond $X=0.875 $Y=1.875
+ $X2=0.75 $Y2=1.875
r109 25 27 50.2172 $w=1.78e-07 $l=8.15e-07 $layer=LI1_cond $X=0.875 $Y=1.875
+ $X2=1.69 $Y2=1.875
r110 24 31 6.82373 $w=1.8e-07 $l=1.25499e-07 $layer=LI1_cond $X=2.315 $Y=1.875
+ $X2=2.4 $Y2=1.785
r111 24 27 38.5101 $w=1.78e-07 $l=6.25e-07 $layer=LI1_cond $X=2.315 $Y=1.875
+ $X2=1.69 $Y2=1.875
r112 19 46 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=1.202
r113 19 21 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.37 $Y=0.995
+ $X2=3.37 $Y2=0.56
r114 16 45 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=3.345 $Y=1.41
+ $X2=3.345 $Y2=1.202
r115 16 18 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.345 $Y=1.41
+ $X2=3.345 $Y2=1.985
r116 13 44 23.6381 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=2.9 $Y=0.995
+ $X2=2.9 $Y2=1.202
r117 13 15 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=2.9 $Y=0.995
+ $X2=2.9 $Y2=0.56
r118 10 43 19.2931 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=2.875 $Y=1.41
+ $X2=2.875 $Y2=1.202
r119 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.875 $Y=1.41
+ $X2=2.875 $Y2=1.985
r120 3 27 600 $w=1.7e-07 $l=4.51719e-07 $layer=licon1_PDIFF $count=1 $X=1.545
+ $Y=1.485 $X2=1.69 $Y2=1.87
r121 2 33 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.605
+ $Y=1.485 $X2=0.75 $Y2=1.96
r122 1 35 182 $w=1.7e-07 $l=5.80172e-07 $layer=licon1_NDIFF $count=1 $X=1.035
+ $Y=0.235 $X2=1.22 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B1 1 3 4 6 7 9 10 12 13 16 22
c74 4 0 2.98731e-20 $X=3.875 $Y=0.995
r75 22 26 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=5.295
+ $Y=1.16 $X2=5.295 $Y2=1.16
r76 21 22 9.95292 $w=3.28e-07 $l=2.85e-07 $layer=LI1_cond $X=5.295 $Y=1.445
+ $X2=5.295 $Y2=1.16
r77 16 19 10.9334 $w=3.88e-07 $l=3.7e-07 $layer=LI1_cond $X=3.845 $Y=1.16
+ $X2=3.845 $Y2=1.53
r78 16 17 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=3.815
+ $Y=1.16 $X2=3.815 $Y2=1.16
r79 14 19 5.6248 $w=1.7e-07 $l=1.95e-07 $layer=LI1_cond $X=4.04 $Y=1.53
+ $X2=3.845 $Y2=1.53
r80 13 21 7.76618 $w=1.7e-07 $l=2.03101e-07 $layer=LI1_cond $X=5.13 $Y=1.53
+ $X2=5.295 $Y2=1.445
r81 13 14 71.1123 $w=1.68e-07 $l=1.09e-06 $layer=LI1_cond $X=5.13 $Y=1.53
+ $X2=4.04 $Y2=1.53
r82 10 26 48.1208 $w=2.95e-07 $l=2.78388e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.32 $Y2=1.16
r83 10 12 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=5.26 $Y=1.41
+ $X2=5.26 $Y2=1.985
r84 7 26 38.578 $w=2.95e-07 $l=2.03101e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.32 $Y2=1.16
r85 7 9 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=5.235 $Y=0.995
+ $X2=5.235 $Y2=0.56
r86 4 17 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.815 $Y2=1.16
r87 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.875 $Y=0.995
+ $X2=3.875 $Y2=0.56
r88 1 17 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=3.85 $Y=1.41
+ $X2=3.815 $Y2=1.16
r89 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=3.85 $Y=1.41 $X2=3.85
+ $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%B2 1 3 4 6 7 9 10 12 13 20 24
r47 20 21 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.79 $Y=1.202
+ $X2=4.815 $Y2=1.202
r48 18 20 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.555 $Y=1.202
+ $X2=4.79 $Y2=1.202
r49 18 24 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=4.555
+ $Y=1.16 $X2=4.555 $Y2=1.16
r50 16 18 29.8079 $w=3.8e-07 $l=2.35e-07 $layer=POLY_cond $X=4.32 $Y=1.202
+ $X2=4.555 $Y2=1.202
r51 15 16 3.17105 $w=3.8e-07 $l=2.5e-08 $layer=POLY_cond $X=4.295 $Y=1.202
+ $X2=4.32 $Y2=1.202
r52 13 24 10.5364 $w=1.98e-07 $l=1.9e-07 $layer=LI1_cond $X=4.745 $Y=1.175
+ $X2=4.555 $Y2=1.175
r53 10 21 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=1.202
r54 10 12 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.815 $Y=0.995
+ $X2=4.815 $Y2=0.56
r55 7 20 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.79 $Y=1.41
+ $X2=4.79 $Y2=1.202
r56 7 9 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.79 $Y=1.41 $X2=4.79
+ $Y2=1.985
r57 4 16 20.2441 $w=1.8e-07 $l=2.08e-07 $layer=POLY_cond $X=4.32 $Y=1.41
+ $X2=4.32 $Y2=1.202
r58 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=4.32 $Y=1.41 $X2=4.32
+ $Y2=1.985
r59 1 15 24.6126 $w=1.5e-07 $l=2.07e-07 $layer=POLY_cond $X=4.295 $Y=0.995
+ $X2=4.295 $Y2=1.202
r60 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=4.295 $Y=0.995
+ $X2=4.295 $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VPWR 1 2 3 4 5 16 18 20 24 30 34 37 38
+ 40 41 42 55 56 62 67 73
r78 72 73 9.18355 $w=6.68e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=2.47
+ $X2=2.725 $Y2=2.47
r79 69 72 1.96371 $w=6.68e-07 $l=1.1e-07 $layer=LI1_cond $X=2.53 $Y=2.47
+ $X2=2.64 $Y2=2.47
r80 69 70 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r81 66 70 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.07 $Y=2.72
+ $X2=2.53 $Y2=2.72
r82 65 69 8.21188 $w=6.68e-07 $l=4.6e-07 $layer=LI1_cond $X=2.07 $Y=2.47
+ $X2=2.53 $Y2=2.47
r83 65 67 8.29096 $w=6.68e-07 $l=3.5e-08 $layer=LI1_cond $X=2.07 $Y=2.47
+ $X2=2.035 $Y2=2.47
r84 65 66 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=2.72
+ $X2=2.07 $Y2=2.72
r85 63 66 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=1.15 $Y=2.72
+ $X2=2.07 $Y2=2.72
r86 62 63 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.15 $Y=2.72
+ $X2=1.15 $Y2=2.72
r87 55 56 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=5.75 $Y=2.72
+ $X2=5.75 $Y2=2.72
r88 53 56 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=5.29 $Y=2.72
+ $X2=5.75 $Y2=2.72
r89 52 53 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.29 $Y=2.72
+ $X2=5.29 $Y2=2.72
r90 50 53 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r91 49 52 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=3.91 $Y=2.72
+ $X2=5.29 $Y2=2.72
r92 49 50 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=2.72
+ $X2=3.91 $Y2=2.72
r93 47 50 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=3.91 $Y2=2.72
r94 47 70 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.45 $Y=2.72
+ $X2=2.53 $Y2=2.72
r95 46 73 47.2995 $w=1.68e-07 $l=7.25e-07 $layer=LI1_cond $X=3.45 $Y=2.72
+ $X2=2.725 $Y2=2.72
r96 46 47 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r97 42 63 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.15 $Y2=2.72
r98 42 59 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r99 40 52 8.15508 $w=1.68e-07 $l=1.25e-07 $layer=LI1_cond $X=5.415 $Y=2.72
+ $X2=5.29 $Y2=2.72
r100 40 41 6.01921 $w=1.7e-07 $l=1.02e-07 $layer=LI1_cond $X=5.415 $Y=2.72
+ $X2=5.517 $Y2=2.72
r101 39 55 8.48128 $w=1.68e-07 $l=1.3e-07 $layer=LI1_cond $X=5.62 $Y=2.72
+ $X2=5.75 $Y2=2.72
r102 39 41 6.01921 $w=1.7e-07 $l=1.03e-07 $layer=LI1_cond $X=5.62 $Y=2.72
+ $X2=5.517 $Y2=2.72
r103 37 46 0.326203 $w=1.68e-07 $l=5e-09 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.45 $Y2=2.72
r104 37 38 7.75133 $w=1.7e-07 $l=1.42e-07 $layer=LI1_cond $X=3.455 $Y=2.72
+ $X2=3.597 $Y2=2.72
r105 36 49 11.0909 $w=1.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.74 $Y=2.72
+ $X2=3.91 $Y2=2.72
r106 36 38 7.75133 $w=1.7e-07 $l=1.43e-07 $layer=LI1_cond $X=3.74 $Y=2.72
+ $X2=3.597 $Y2=2.72
r107 32 41 0.677923 $w=2.05e-07 $l=8.5e-08 $layer=LI1_cond $X=5.517 $Y=2.635
+ $X2=5.517 $Y2=2.72
r108 32 34 36.5188 $w=2.03e-07 $l=6.75e-07 $layer=LI1_cond $X=5.517 $Y=2.635
+ $X2=5.517 $Y2=1.96
r109 28 38 0.432977 $w=2.85e-07 $l=8.5e-08 $layer=LI1_cond $X=3.597 $Y=2.635
+ $X2=3.597 $Y2=2.72
r110 28 30 13.5463 $w=2.83e-07 $l=3.35e-07 $layer=LI1_cond $X=3.597 $Y=2.635
+ $X2=3.597 $Y2=2.3
r111 27 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=1.22 $Y2=2.72
r112 27 67 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=1.345 $Y=2.72
+ $X2=2.035 $Y2=2.72
r113 22 62 0.00168595 $w=2.5e-07 $l=8.5e-08 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.72
r114 22 24 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=1.22 $Y=2.635
+ $X2=1.22 $Y2=2.3
r115 21 59 3.96842 $w=1.7e-07 $l=2e-07 $layer=LI1_cond $X=0.4 $Y=2.72 $X2=0.2
+ $Y2=2.72
r116 20 62 7.02821 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=1.22 $Y2=2.72
r117 20 21 45.3422 $w=1.68e-07 $l=6.95e-07 $layer=LI1_cond $X=1.095 $Y=2.72
+ $X2=0.4 $Y2=2.72
r118 16 59 3.17474 $w=2.5e-07 $l=1.16619e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.2 $Y2=2.72
r119 16 18 31.116 $w=2.48e-07 $l=6.75e-07 $layer=LI1_cond $X=0.275 $Y=2.635
+ $X2=0.275 $Y2=1.96
r120 5 34 300 $w=1.7e-07 $l=5.44862e-07 $layer=licon1_PDIFF $count=2 $X=5.35
+ $Y=1.485 $X2=5.5 $Y2=1.96
r121 4 30 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.435
+ $Y=1.485 $X2=3.58 $Y2=2.3
r122 3 72 300 $w=1.7e-07 $l=1.07956e-06 $layer=licon1_PDIFF $count=2 $X=2.025
+ $Y=1.485 $X2=2.64 $Y2=2.3
r123 2 24 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=1.075
+ $Y=1.485 $X2=1.22 $Y2=2.3
r124 1 18 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.28 $Y2=1.96
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%Y 1 2 3 12 16 18 20 23 24 29
r47 29 34 1.88854 $w=5.68e-07 $l=9e-08 $layer=LI1_cond $X=3.18 $Y=1.53 $X2=3.18
+ $Y2=1.62
r48 24 27 4.14879 $w=2.48e-07 $l=9e-08 $layer=LI1_cond $X=4.555 $Y=1.87
+ $X2=4.555 $Y2=1.96
r49 22 34 3.46233 $w=5.68e-07 $l=1.65e-07 $layer=LI1_cond $X=3.18 $Y=1.785
+ $X2=3.18 $Y2=1.62
r50 22 23 2.14437 $w=4.55e-07 $l=8.5e-08 $layer=LI1_cond $X=3.18 $Y=1.785
+ $X2=3.18 $Y2=1.87
r51 20 29 3.56725 $w=5.68e-07 $l=1.7e-07 $layer=LI1_cond $X=3.18 $Y=1.36
+ $X2=3.18 $Y2=1.53
r52 20 21 7.31248 $w=5.68e-07 $l=2.85e-07 $layer=LI1_cond $X=3.18 $Y=1.36
+ $X2=3.18 $Y2=1.075
r53 19 23 5.03717 $w=1.7e-07 $l=2.85e-07 $layer=LI1_cond $X=3.465 $Y=1.87
+ $X2=3.18 $Y2=1.87
r54 18 24 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.43 $Y=1.87
+ $X2=4.555 $Y2=1.87
r55 18 19 62.9572 $w=1.68e-07 $l=9.65e-07 $layer=LI1_cond $X=4.43 $Y=1.87
+ $X2=3.465 $Y2=1.87
r56 14 23 2.14437 $w=4.55e-07 $l=1.51658e-07 $layer=LI1_cond $X=3.065 $Y=1.955
+ $X2=3.18 $Y2=1.87
r57 14 16 0.169477 $w=3.38e-07 $l=5e-09 $layer=LI1_cond $X=3.065 $Y=1.955
+ $X2=3.065 $Y2=1.96
r58 12 21 10.463 $w=3.78e-07 $l=3.45e-07 $layer=LI1_cond $X=3.085 $Y=0.73
+ $X2=3.085 $Y2=1.075
r59 3 27 600 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=1 $X=4.41
+ $Y=1.485 $X2=4.555 $Y2=1.96
r60 2 34 600 $w=1.7e-07 $l=2.01494e-07 $layer=licon1_PDIFF $count=1 $X=2.965
+ $Y=1.485 $X2=3.11 $Y2=1.62
r61 2 16 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=2.965
+ $Y=1.485 $X2=3.11 $Y2=1.96
r62 1 12 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=2.975
+ $Y=0.235 $X2=3.11 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_788_297# 1 2 7 11 14
r17 14 16 3.68782 $w=2.48e-07 $l=8e-08 $layer=LI1_cond $X=4.085 $Y=2.3 $X2=4.085
+ $Y2=2.38
r18 9 11 15.4427 $w=2.48e-07 $l=3.35e-07 $layer=LI1_cond $X=5.025 $Y=2.295
+ $X2=5.025 $Y2=1.96
r19 8 16 2.99516 $w=1.7e-07 $l=1.25e-07 $layer=LI1_cond $X=4.21 $Y=2.38
+ $X2=4.085 $Y2=2.38
r20 7 9 7.14316 $w=1.7e-07 $l=1.62019e-07 $layer=LI1_cond $X=4.9 $Y=2.38
+ $X2=5.025 $Y2=2.295
r21 7 8 45.016 $w=1.68e-07 $l=6.9e-07 $layer=LI1_cond $X=4.9 $Y=2.38 $X2=4.21
+ $Y2=2.38
r22 2 11 300 $w=1.7e-07 $l=5.42679e-07 $layer=licon1_PDIFF $count=2 $X=4.88
+ $Y=1.485 $X2=5.025 $Y2=1.96
r23 1 14 600 $w=1.7e-07 $l=8.84534e-07 $layer=licon1_PDIFF $count=1 $X=3.94
+ $Y=1.485 $X2=4.085 $Y2=2.3
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%VGND 1 2 3 4 13 15 19 23 27 30 31 33 34
+ 35 37 53 54 60
r82 60 61 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.07 $Y=0 $X2=2.07
+ $Y2=0
r83 53 54 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=5.75 $Y=0 $X2=5.75
+ $Y2=0
r84 51 54 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=4.83 $Y=0 $X2=5.75
+ $Y2=0
r85 50 51 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=4.83 $Y=0 $X2=4.83
+ $Y2=0
r86 48 51 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=3.91 $Y=0 $X2=4.83
+ $Y2=0
r87 47 48 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.91 $Y=0 $X2=3.91
+ $Y2=0
r88 45 48 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r89 45 61 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=2.07
+ $Y2=0
r90 44 47 90.0321 $w=1.68e-07 $l=1.38e-06 $layer=LI1_cond $X=2.53 $Y=0 $X2=3.91
+ $Y2=0
r91 44 45 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r92 42 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.12
+ $Y2=0
r93 42 44 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=2.205 $Y=0 $X2=2.53
+ $Y2=0
r94 41 61 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.07
+ $Y2=0
r95 40 41 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r96 38 57 3.40825 $w=1.7e-07 $l=1.83e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.182
+ $Y2=0
r97 38 40 21.2032 $w=1.68e-07 $l=3.25e-07 $layer=LI1_cond $X=0.365 $Y=0 $X2=0.69
+ $Y2=0
r98 37 60 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.035 $Y=0 $X2=2.12
+ $Y2=0
r99 37 40 87.7487 $w=1.68e-07 $l=1.345e-06 $layer=LI1_cond $X=2.035 $Y=0
+ $X2=0.69 $Y2=0
r100 35 41 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r101 35 57 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r102 33 50 7.17647 $w=1.68e-07 $l=1.1e-07 $layer=LI1_cond $X=4.94 $Y=0 $X2=4.83
+ $Y2=0
r103 33 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.94 $Y=0 $X2=5.025
+ $Y2=0
r104 32 53 41.754 $w=1.68e-07 $l=6.4e-07 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.75
+ $Y2=0
r105 32 34 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.11 $Y=0 $X2=5.025
+ $Y2=0
r106 30 47 5.87166 $w=1.68e-07 $l=9e-08 $layer=LI1_cond $X=4 $Y=0 $X2=3.91 $Y2=0
r107 30 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4 $Y=0 $X2=4.085
+ $Y2=0
r108 29 50 43.0588 $w=1.68e-07 $l=6.6e-07 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.83
+ $Y2=0
r109 29 31 5.16603 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.17 $Y=0 $X2=4.085
+ $Y2=0
r110 25 34 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=5.025 $Y=0.085
+ $X2=5.025 $Y2=0
r111 25 27 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=5.025 $Y=0.085
+ $X2=5.025 $Y2=0.39
r112 21 31 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0
r113 21 23 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=4.085 $Y=0.085
+ $X2=4.085 $Y2=0.39
r114 17 60 1.34256 $w=1.7e-07 $l=8.5e-08 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0
r115 17 19 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=2.12 $Y=0.085
+ $X2=2.12 $Y2=0.39
r116 13 57 3.40825 $w=1.7e-07 $l=1.33918e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.182 $Y2=0
r117 13 15 19.8984 $w=1.68e-07 $l=3.05e-07 $layer=LI1_cond $X=0.28 $Y=0.085
+ $X2=0.28 $Y2=0.39
r118 4 27 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=4.89
+ $Y=0.235 $X2=5.025 $Y2=0.39
r119 3 23 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.95
+ $Y=0.235 $X2=4.085 $Y2=0.39
r120 2 19 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.985
+ $Y=0.235 $X2=2.12 $Y2=0.39
r121 1 15 91 $w=1.7e-07 $l=2.15639e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.28 $Y2=0.39
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_123_47# 1 2 7 9 13
c22 9 0 6.98311e-20 $X=0.75 $Y=0.73
r23 11 16 4.79851 $w=1.7e-07 $l=1.5e-07 $layer=LI1_cond $X=0.835 $Y=0.39
+ $X2=0.685 $Y2=0.39
r24 11 13 55.7807 $w=1.68e-07 $l=8.55e-07 $layer=LI1_cond $X=0.835 $Y=0.39
+ $X2=1.69 $Y2=0.39
r25 7 16 2.71916 $w=3e-07 $l=8.5e-08 $layer=LI1_cond $X=0.685 $Y=0.475 $X2=0.685
+ $Y2=0.39
r26 7 9 9.79577 $w=2.98e-07 $l=2.55e-07 $layer=LI1_cond $X=0.685 $Y=0.475
+ $X2=0.685 $Y2=0.73
r27 2 13 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=1.555
+ $Y=0.235 $X2=1.69 $Y2=0.39
r28 1 16 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.39
r29 1 9 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=0.615
+ $Y=0.235 $X2=0.75 $Y2=0.73
.ends

.subckt PM_SKY130_FD_SC_HDLL__O2BB2AI_2%A_503_47# 1 2 3 4 13 15 19 20 23 25 29
+ 34 37
c59 37 0 2.98731e-20 $X=4.53 $Y=0.815
c60 20 0 1.98409e-19 $X=3.78 $Y=0.82
r61 32 34 4.10683 $w=2.98e-07 $l=8.5e-08 $layer=LI1_cond $X=2.64 $Y=0.405
+ $X2=2.725 $Y2=0.405
r62 27 29 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=5.47 $Y=0.725
+ $X2=5.47 $Y2=0.39
r63 26 37 9.30075 $w=1.75e-07 $l=1.9e-07 $layer=LI1_cond $X=4.72 $Y=0.815
+ $X2=4.53 $Y2=0.815
r64 25 27 8.0135 $w=1.8e-07 $l=2.30651e-07 $layer=LI1_cond $X=5.28 $Y=0.815
+ $X2=5.47 $Y2=0.725
r65 25 26 34.5051 $w=1.78e-07 $l=5.6e-07 $layer=LI1_cond $X=5.28 $Y=0.815
+ $X2=4.72 $Y2=0.815
r66 21 37 1.23463 $w=3.8e-07 $l=9e-08 $layer=LI1_cond $X=4.53 $Y=0.725 $X2=4.53
+ $Y2=0.815
r67 21 23 10.1597 $w=3.78e-07 $l=3.35e-07 $layer=LI1_cond $X=4.53 $Y=0.725
+ $X2=4.53 $Y2=0.39
r68 19 37 9.30075 $w=1.75e-07 $l=1.92484e-07 $layer=LI1_cond $X=4.34 $Y=0.82
+ $X2=4.53 $Y2=0.815
r69 19 20 36.5348 $w=1.68e-07 $l=5.6e-07 $layer=LI1_cond $X=4.34 $Y=0.82
+ $X2=3.78 $Y2=0.82
r70 16 20 7.39867 $w=1.7e-07 $l=1.80566e-07 $layer=LI1_cond $X=3.637 $Y=0.735
+ $X2=3.78 $Y2=0.82
r71 16 18 0.202183 $w=2.83e-07 $l=5e-09 $layer=LI1_cond $X=3.637 $Y=0.735
+ $X2=3.637 $Y2=0.73
r72 15 36 3.04002 $w=2.85e-07 $l=1.1e-07 $layer=LI1_cond $X=3.637 $Y=0.475
+ $X2=3.637 $Y2=0.365
r73 15 18 10.3113 $w=2.83e-07 $l=2.55e-07 $layer=LI1_cond $X=3.637 $Y=0.475
+ $X2=3.637 $Y2=0.73
r74 13 36 3.92439 $w=2.2e-07 $l=1.42e-07 $layer=LI1_cond $X=3.495 $Y=0.365
+ $X2=3.637 $Y2=0.365
r75 13 34 40.3355 $w=2.18e-07 $l=7.7e-07 $layer=LI1_cond $X=3.495 $Y=0.365
+ $X2=2.725 $Y2=0.365
r76 4 29 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=5.31
+ $Y=0.235 $X2=5.495 $Y2=0.39
r77 3 23 91 $w=1.7e-07 $l=2.50799e-07 $layer=licon1_NDIFF $count=2 $X=4.37
+ $Y=0.235 $X2=4.555 $Y2=0.39
r78 2 36 182 $w=1.7e-07 $l=2.12014e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.235 $X2=3.58 $Y2=0.39
r79 2 18 182 $w=1.7e-07 $l=5.58435e-07 $layer=licon1_NDIFF $count=1 $X=3.445
+ $Y=0.235 $X2=3.58 $Y2=0.73
r80 1 32 182 $w=1.7e-07 $l=2.08327e-07 $layer=licon1_NDIFF $count=1 $X=2.515
+ $Y=0.235 $X2=2.64 $Y2=0.39
.ends

