* File: sky130_fd_sc_hdll__a2bb2oi_1.pxi.spice
* Created: Thu Aug 27 18:55:03 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A1_N N_A1_N_c_53_n N_A1_N_M1002_g
+ N_A1_N_c_54_n N_A1_N_M1007_g A1_N A1_N N_A1_N_c_55_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A2_N N_A2_N_c_77_n N_A2_N_M1001_g
+ N_A2_N_c_78_n N_A2_N_M1003_g A2_N A2_N PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_119_47# N_A_119_47#_M1007_d
+ N_A_119_47#_M1001_d N_A_119_47#_c_107_n N_A_119_47#_M1006_g
+ N_A_119_47#_c_108_n N_A_119_47#_M1004_g N_A_119_47#_c_120_n
+ N_A_119_47#_c_121_n N_A_119_47#_c_124_n N_A_119_47#_c_111_n
+ N_A_119_47#_c_112_n N_A_119_47#_c_113_n N_A_119_47#_c_109_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_119_47#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B2 N_B2_c_173_n N_B2_M1009_g N_B2_c_174_n
+ N_B2_M1000_g B2 B2 B2 B2 B2 PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B1 N_B1_c_213_n N_B1_M1008_g N_B1_c_214_n
+ N_B1_M1005_g B1 B1 PM_SKY130_FD_SC_HDLL__A2BB2OI_1%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VPWR N_VPWR_M1002_s N_VPWR_M1009_d
+ N_VPWR_c_240_n N_VPWR_c_241_n N_VPWR_c_242_n VPWR VPWR N_VPWR_c_244_n
+ N_VPWR_c_239_n N_VPWR_c_246_n PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%Y N_Y_M1004_d N_Y_M1006_s N_Y_c_285_n
+ N_Y_c_294_n Y Y Y N_Y_c_287_n Y N_Y_c_288_n PM_SKY130_FD_SC_HDLL__A2BB2OI_1%Y
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_409_297# N_A_409_297#_M1006_d
+ N_A_409_297#_M1005_d N_A_409_297#_c_324_n N_A_409_297#_c_327_n
+ N_A_409_297#_c_325_n N_A_409_297#_c_322_n N_A_409_297#_c_323_n
+ N_A_409_297#_c_331_n PM_SKY130_FD_SC_HDLL__A2BB2OI_1%A_409_297#
x_PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VGND N_VGND_M1007_s N_VGND_M1003_d
+ N_VGND_M1008_d N_VGND_c_355_n N_VGND_c_356_n N_VGND_c_357_n VGND VGND
+ N_VGND_c_359_n N_VGND_c_360_n N_VGND_c_361_n N_VGND_c_362_n N_VGND_c_363_n
+ PM_SKY130_FD_SC_HDLL__A2BB2OI_1%VGND
cc_1 VNB N_A1_N_c_53_n 0.0293922f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_2 VNB N_A1_N_c_54_n 0.0227688f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_3 VNB N_A1_N_c_55_n 0.0151164f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_4 VNB N_A2_N_c_77_n 0.0221726f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_A2_N_c_78_n 0.019998f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB A2_N 0.0110473f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_7 VNB N_A_119_47#_c_107_n 0.0385723f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_119_47#_c_108_n 0.0198871f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_9 VNB N_A_119_47#_c_109_n 0.00214269f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB N_B2_c_173_n 0.0234988f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_11 VNB N_B2_c_174_n 0.0163852f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_12 VNB B2 0.00199701f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_13 VNB B2 0.00321955f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB B2 0.00143542f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_B1_c_213_n 0.0214066f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_16 VNB N_B1_c_214_n 0.0248266f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_17 VNB B1 0.0145378f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_18 VNB N_VPWR_c_239_n 0.155873f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_Y_c_285_n 0.00290563f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.445
cc_20 VNB N_VGND_c_355_n 0.0277822f $X=-0.19 $Y=-0.24 $X2=0.41 $Y2=1.16
cc_21 VNB N_VGND_c_356_n 0.0355357f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB N_VGND_c_357_n 0.00606646f $X=-0.19 $Y=-0.24 $X2=0.335 $Y2=1.19
cc_23 VNB VGND 0.0115788f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_24 VNB N_VGND_c_359_n 0.0115308f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_25 VNB N_VGND_c_360_n 0.207304f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_26 VNB N_VGND_c_361_n 0.016052f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_27 VNB N_VGND_c_362_n 0.0162801f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_28 VNB N_VGND_c_363_n 0.0293343f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_29 VPB N_A1_N_c_53_n 0.0299451f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_30 VPB N_A1_N_c_55_n 0.00680297f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_31 VPB N_A2_N_c_77_n 0.0293154f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_32 VPB N_A_119_47#_c_107_n 0.0340465f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_33 VPB N_A_119_47#_c_111_n 0.00951556f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB N_A_119_47#_c_112_n 0.0141706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_A_119_47#_c_113_n 0.00299815f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 VPB N_A_119_47#_c_109_n 0.00241287f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_37 VPB N_B2_c_173_n 0.0245263f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_38 VPB B2 0.00248295f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_39 VPB N_B1_c_214_n 0.0285618f $X=-0.19 $Y=1.305 $X2=0.52 $Y2=0.995
cc_40 VPB B1 0.00808203f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_41 VPB N_VPWR_c_240_n 0.0023782f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_42 VPB N_VPWR_c_241_n 0.0586701f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_43 VPB N_VPWR_c_242_n 0.00359552f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_44 VPB VPWR 0.0103693f $X=-0.19 $Y=1.305 $X2=0.335 $Y2=1.16
cc_45 VPB N_VPWR_c_244_n 0.0230602f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_46 VPB N_VPWR_c_239_n 0.061956f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_47 VPB N_VPWR_c_246_n 0.0306634f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_48 VPB N_Y_c_285_n 0.00123769f $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.445
cc_49 VPB N_Y_c_287_n 0.00618859f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_50 VPB N_Y_c_288_n 0.00269924f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_51 VPB N_A_409_297#_c_322_n 0.00899863f $X=-0.19 $Y=1.305 $X2=0.435 $Y2=1.16
cc_52 VPB N_A_409_297#_c_323_n 0.0195283f $X=-0.19 $Y=1.305 $X2=0.41 $Y2=1.16
cc_53 N_A1_N_c_53_n N_A2_N_c_77_n 0.0919242f $X=0.495 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_54 N_A1_N_c_55_n N_A2_N_c_77_n 0.00188742f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_55 N_A1_N_c_54_n N_A2_N_c_78_n 0.0187856f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_56 N_A1_N_c_53_n A2_N 0.00186759f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_57 N_A1_N_c_55_n A2_N 0.0162612f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_58 N_A1_N_c_53_n N_A_119_47#_c_111_n 0.00296559f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_59 N_A1_N_c_53_n N_A_119_47#_c_113_n 4.83935e-19 $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_60 N_A1_N_c_55_n N_A_119_47#_c_113_n 0.00677707f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_61 N_A1_N_c_55_n N_VPWR_M1002_s 0.0081321f $X=0.41 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_62 N_A1_N_c_53_n N_VPWR_c_241_n 0.00622633f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_63 N_A1_N_c_53_n N_VPWR_c_239_n 0.0103479f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_64 N_A1_N_c_53_n N_VPWR_c_246_n 0.0181473f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_65 N_A1_N_c_55_n N_VPWR_c_246_n 0.017648f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_66 N_A1_N_c_54_n N_VGND_c_360_n 0.0117108f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_67 N_A1_N_c_54_n N_VGND_c_361_n 0.00585385f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_68 N_A1_N_c_54_n N_VGND_c_362_n 5.93551e-19 $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_69 N_A1_N_c_53_n N_VGND_c_363_n 0.00106812f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_70 N_A1_N_c_54_n N_VGND_c_363_n 0.00338835f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_71 N_A1_N_c_55_n N_VGND_c_363_n 0.0226315f $X=0.41 $Y=1.16 $X2=0 $Y2=0
cc_72 N_A2_N_c_77_n N_A_119_47#_c_107_n 0.00651131f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_73 A2_N N_A_119_47#_c_107_n 0.00274628f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_74 N_A2_N_c_78_n N_A_119_47#_c_120_n 0.00438427f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_75 N_A2_N_c_77_n N_A_119_47#_c_121_n 0.00279419f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_76 N_A2_N_c_78_n N_A_119_47#_c_121_n 0.0125248f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_77 A2_N N_A_119_47#_c_121_n 0.0331674f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_78 N_A2_N_c_77_n N_A_119_47#_c_124_n 2.455e-19 $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_79 A2_N N_A_119_47#_c_124_n 0.00319213f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_80 N_A2_N_c_77_n N_A_119_47#_c_111_n 0.0182521f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_81 A2_N N_A_119_47#_c_112_n 0.00268974f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_82 N_A2_N_c_77_n N_A_119_47#_c_113_n 0.00751953f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_83 A2_N N_A_119_47#_c_113_n 0.032179f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_84 N_A2_N_c_77_n N_A_119_47#_c_109_n 0.00315181f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A2_N_c_78_n N_A_119_47#_c_109_n 0.00370217f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_86 A2_N N_A_119_47#_c_109_n 0.0135327f $X=1.17 $Y=1.105 $X2=0 $Y2=0
cc_87 N_A2_N_c_77_n N_VPWR_c_241_n 0.00597712f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_88 N_A2_N_c_77_n N_VPWR_c_239_n 0.0113213f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_89 N_A2_N_c_77_n N_VPWR_c_246_n 0.00289871f $X=0.905 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A2_N_c_78_n N_VGND_c_360_n 0.00419427f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_91 N_A2_N_c_78_n N_VGND_c_361_n 0.00342263f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_92 N_A2_N_c_78_n N_VGND_c_362_n 0.00909388f $X=1 $Y=0.995 $X2=0 $Y2=0
cc_93 N_A_119_47#_c_107_n N_B2_c_173_n 0.047584f $X=1.955 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_94 N_A_119_47#_c_108_n N_B2_c_174_n 0.0195918f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_119_47#_c_108_n B2 4.13383e-19 $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_96 N_A_119_47#_c_107_n B2 3.33602e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_97 N_A_119_47#_c_107_n B2 5.60488e-19 $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_98 N_A_119_47#_c_107_n N_VPWR_c_241_n 0.00673617f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_99 N_A_119_47#_c_111_n N_VPWR_c_241_n 0.0244686f $X=1.14 $Y=1.64 $X2=0 $Y2=0
cc_100 N_A_119_47#_M1001_d N_VPWR_c_239_n 0.00217517f $X=0.995 $Y=1.485 $X2=0
+ $Y2=0
cc_101 N_A_119_47#_c_107_n N_VPWR_c_239_n 0.00856101f $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_102 N_A_119_47#_c_111_n N_VPWR_c_239_n 0.0141694f $X=1.14 $Y=1.64 $X2=0 $Y2=0
cc_103 N_A_119_47#_c_111_n N_VPWR_c_246_n 0.0207672f $X=1.14 $Y=1.64 $X2=0 $Y2=0
cc_104 N_A_119_47#_c_112_n N_Y_M1006_s 0.00354649f $X=1.645 $Y=1.53 $X2=0 $Y2=0
cc_105 N_A_119_47#_c_107_n N_Y_c_285_n 0.024332f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_106 N_A_119_47#_c_108_n N_Y_c_285_n 0.00372198f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_107 N_A_119_47#_c_112_n N_Y_c_285_n 0.00760687f $X=1.645 $Y=1.53 $X2=0 $Y2=0
cc_108 N_A_119_47#_c_109_n N_Y_c_285_n 0.0425355f $X=1.73 $Y=1.16 $X2=0 $Y2=0
cc_109 N_A_119_47#_c_108_n N_Y_c_294_n 0.00278677f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_110 N_A_119_47#_c_108_n Y 0.0138525f $X=1.98 $Y=0.995 $X2=0 $Y2=0
cc_111 N_A_119_47#_c_121_n Y 0.0138273f $X=1.645 $Y=0.745 $X2=0 $Y2=0
cc_112 N_A_119_47#_c_107_n N_Y_c_287_n 0.00729502f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_113 N_A_119_47#_c_111_n N_Y_c_287_n 0.0366936f $X=1.14 $Y=1.64 $X2=0 $Y2=0
cc_114 N_A_119_47#_c_107_n N_Y_c_288_n 0.0140497f $X=1.955 $Y=1.41 $X2=0 $Y2=0
cc_115 N_A_119_47#_c_111_n N_Y_c_288_n 0.0126567f $X=1.14 $Y=1.64 $X2=0 $Y2=0
cc_116 N_A_119_47#_c_112_n N_Y_c_288_n 0.0225044f $X=1.645 $Y=1.53 $X2=0 $Y2=0
cc_117 N_A_119_47#_c_107_n N_A_409_297#_c_324_n 0.00217158f $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_118 N_A_119_47#_c_107_n N_A_409_297#_c_325_n 5.51893e-19 $X=1.955 $Y=1.41
+ $X2=0 $Y2=0
cc_119 N_A_119_47#_c_121_n N_VGND_M1003_d 0.0219865f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_120 N_A_119_47#_c_109_n N_VGND_M1003_d 0.00132526f $X=1.73 $Y=1.16 $X2=0
+ $Y2=0
cc_121 N_A_119_47#_c_108_n N_VGND_c_356_n 0.00480635f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_122 N_A_119_47#_c_121_n N_VGND_c_356_n 0.00182296f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_123 N_A_119_47#_M1007_d N_VGND_c_360_n 0.00485355f $X=0.595 $Y=0.235 $X2=0
+ $Y2=0
cc_124 N_A_119_47#_c_108_n N_VGND_c_360_n 0.00996238f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_125 N_A_119_47#_c_120_n N_VGND_c_360_n 0.0064418f $X=0.73 $Y=0.66 $X2=0 $Y2=0
cc_126 N_A_119_47#_c_121_n N_VGND_c_360_n 0.0116102f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_127 N_A_119_47#_c_120_n N_VGND_c_361_n 0.0114662f $X=0.73 $Y=0.66 $X2=0 $Y2=0
cc_128 N_A_119_47#_c_121_n N_VGND_c_361_n 0.00323219f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_129 N_A_119_47#_c_107_n N_VGND_c_362_n 3.57259e-19 $X=1.955 $Y=1.41 $X2=0
+ $Y2=0
cc_130 N_A_119_47#_c_108_n N_VGND_c_362_n 0.00936866f $X=1.98 $Y=0.995 $X2=0
+ $Y2=0
cc_131 N_A_119_47#_c_120_n N_VGND_c_362_n 0.014533f $X=0.73 $Y=0.66 $X2=0 $Y2=0
cc_132 N_A_119_47#_c_121_n N_VGND_c_362_n 0.0472181f $X=1.645 $Y=0.745 $X2=0
+ $Y2=0
cc_133 N_B2_c_174_n N_B1_c_213_n 0.0284971f $X=2.53 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_134 B2 N_B1_c_213_n 0.00163618f $X=2.445 $Y=0.425 $X2=-0.19 $Y2=-0.24
cc_135 N_B2_c_173_n N_B1_c_214_n 0.0661818f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_136 B2 N_B1_c_214_n 0.00312973f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_137 B2 N_B1_c_214_n 3.54802e-19 $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_138 N_B2_c_173_n B1 8.9659e-19 $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_139 B2 B1 0.0270187f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_140 N_B2_c_173_n N_VPWR_c_240_n 0.00425183f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_141 N_B2_c_173_n N_VPWR_c_241_n 0.00581124f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_142 N_B2_c_173_n N_VPWR_c_239_n 0.0068111f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_143 N_B2_c_173_n N_Y_c_285_n 0.00645155f $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_144 N_B2_c_174_n N_Y_c_285_n 6.12594e-19 $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_145 B2 N_Y_c_285_n 0.0071097f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_146 B2 N_Y_c_285_n 0.0329494f $X=2.445 $Y=1.105 $X2=0 $Y2=0
cc_147 N_B2_c_174_n Y 0.00554269f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_148 N_B2_c_173_n N_Y_c_287_n 2.1132e-19 $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_149 N_B2_c_173_n N_Y_c_288_n 5.6527e-19 $X=2.505 $Y=1.41 $X2=0 $Y2=0
cc_150 N_B2_c_173_n N_A_409_297#_c_324_n 0.00750319f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_151 N_B2_c_173_n N_A_409_297#_c_327_n 0.00716825f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_152 B2 N_A_409_297#_c_327_n 0.00758348f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_153 N_B2_c_173_n N_A_409_297#_c_325_n 0.00483043f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_154 B2 N_A_409_297#_c_325_n 0.00655074f $X=2.525 $Y=1.19 $X2=0 $Y2=0
cc_155 N_B2_c_173_n N_A_409_297#_c_331_n 0.00427883f $X=2.505 $Y=1.41 $X2=0
+ $Y2=0
cc_156 N_B2_c_174_n N_VGND_c_355_n 0.00239844f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_157 N_B2_c_174_n N_VGND_c_356_n 0.00390689f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_158 B2 N_VGND_c_356_n 0.00505943f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_159 N_B2_c_174_n N_VGND_c_360_n 0.00580795f $X=2.53 $Y=0.995 $X2=0 $Y2=0
cc_160 B2 N_VGND_c_360_n 0.00512042f $X=2.445 $Y=0.425 $X2=0 $Y2=0
cc_161 N_B1_c_214_n N_VPWR_c_240_n 0.0097842f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_162 N_B1_c_214_n N_VPWR_c_244_n 0.00622633f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_163 N_B1_c_214_n N_VPWR_c_239_n 0.00653159f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_164 B1 N_A_409_297#_M1005_d 0.00635119f $X=2.99 $Y=1.105 $X2=0 $Y2=0
cc_165 N_B1_c_214_n N_A_409_297#_c_324_n 6.47949e-19 $X=2.985 $Y=1.41 $X2=0
+ $Y2=0
cc_166 N_B1_c_214_n N_A_409_297#_c_327_n 0.0111355f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_167 B1 N_A_409_297#_c_327_n 0.013636f $X=2.99 $Y=1.105 $X2=0 $Y2=0
cc_168 B1 N_A_409_297#_c_322_n 0.00802187f $X=2.99 $Y=1.105 $X2=0 $Y2=0
cc_169 N_B1_c_214_n N_A_409_297#_c_323_n 0.0037127f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B1_c_213_n N_VGND_c_355_n 0.0161804f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_171 N_B1_c_214_n N_VGND_c_355_n 0.00279043f $X=2.985 $Y=1.41 $X2=0 $Y2=0
cc_172 B1 N_VGND_c_355_n 0.0165536f $X=2.99 $Y=1.105 $X2=0 $Y2=0
cc_173 N_B1_c_213_n N_VGND_c_356_n 0.0046653f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_174 N_B1_c_213_n N_VGND_c_360_n 0.00802136f $X=2.96 $Y=0.995 $X2=0 $Y2=0
cc_175 N_VPWR_c_239_n A_117_297# 0.00983149f $X=3.45 $Y=2.72 $X2=-0.19 $Y2=-0.24
cc_176 N_VPWR_c_239_n N_Y_M1006_s 0.00217517f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_177 N_VPWR_c_241_n N_Y_c_287_n 0.0231203f $X=2.665 $Y=2.72 $X2=0 $Y2=0
cc_178 N_VPWR_c_239_n N_Y_c_287_n 0.0137178f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_179 N_VPWR_c_239_n N_Y_c_288_n 0.00538887f $X=3.45 $Y=2.72 $X2=0 $Y2=0
cc_180 N_VPWR_c_239_n N_A_409_297#_M1006_d 0.00301907f $X=3.45 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_181 N_VPWR_c_239_n N_A_409_297#_M1005_d 0.00249571f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_182 N_VPWR_c_240_n N_A_409_297#_c_324_n 0.00723635f $X=2.75 $Y=2.36 $X2=0
+ $Y2=0
cc_183 N_VPWR_M1009_d N_A_409_297#_c_327_n 0.00919602f $X=2.595 $Y=1.485 $X2=0
+ $Y2=0
cc_184 N_VPWR_c_240_n N_A_409_297#_c_327_n 0.0142813f $X=2.75 $Y=2.36 $X2=0
+ $Y2=0
cc_185 N_VPWR_c_239_n N_A_409_297#_c_327_n 0.0132153f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_186 N_VPWR_c_240_n N_A_409_297#_c_323_n 0.0201792f $X=2.75 $Y=2.36 $X2=0
+ $Y2=0
cc_187 N_VPWR_c_244_n N_A_409_297#_c_323_n 0.0178516f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_188 N_VPWR_c_239_n N_A_409_297#_c_323_n 0.00974347f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_189 N_VPWR_c_240_n N_A_409_297#_c_331_n 0.0177993f $X=2.75 $Y=2.36 $X2=0
+ $Y2=0
cc_190 N_VPWR_c_241_n N_A_409_297#_c_331_n 0.0252239f $X=2.665 $Y=2.72 $X2=0
+ $Y2=0
cc_191 N_VPWR_c_239_n N_A_409_297#_c_331_n 0.0160606f $X=3.45 $Y=2.72 $X2=0
+ $Y2=0
cc_192 N_Y_c_285_n N_A_409_297#_M1006_d 0.0035342f $X=2.07 $Y=1.785 $X2=-0.19
+ $Y2=-0.24
cc_193 N_Y_c_288_n N_A_409_297#_M1006_d 0.00233708f $X=2.07 $Y=1.87 $X2=-0.19
+ $Y2=-0.24
cc_194 N_Y_c_287_n N_A_409_297#_c_324_n 0.00996177f $X=1.72 $Y=1.98 $X2=0 $Y2=0
cc_195 N_Y_c_288_n N_A_409_297#_c_325_n 0.0150704f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_196 N_Y_c_288_n N_A_409_297#_c_331_n 0.00245726f $X=2.07 $Y=1.87 $X2=0 $Y2=0
cc_197 Y N_VGND_c_356_n 0.0180117f $X=2.105 $Y=0.425 $X2=0 $Y2=0
cc_198 N_Y_M1004_d N_VGND_c_360_n 0.00919186f $X=2.055 $Y=0.235 $X2=0 $Y2=0
cc_199 Y N_VGND_c_360_n 0.0107549f $X=2.105 $Y=0.425 $X2=0 $Y2=0
cc_200 Y N_VGND_c_362_n 0.0134065f $X=2.105 $Y=0.425 $X2=0 $Y2=0
cc_201 N_VGND_c_360_n A_521_47# 0.0116651f $X=3.45 $Y=0 $X2=-0.19 $Y2=-0.24
