* File: sky130_fd_sc_hdll__a22o_1.pex.spice
* Created: Wed Sep  2 08:18:30 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* Nominal Temperature: 27C
* Circuit Temperature: 27C
* 
.subckt PM_SKY130_FD_SC_HDLL__A22O_1%B2 1 3 4 6 7 11
r23 10 11 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=0.46
+ $Y=1.16 $X2=0.46 $Y2=1.16
r24 7 11 12.4773 $w=1.98e-07 $l=2.25e-07 $layer=LI1_cond $X=0.235 $Y=1.175
+ $X2=0.46 $Y2=1.175
r25 4 10 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.52 $Y=0.995
+ $X2=0.46 $Y2=1.16
r26 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.52 $Y=0.995 $X2=0.52
+ $Y2=0.56
r27 1 10 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.46 $Y2=1.16
r28 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.495 $Y=1.41
+ $X2=0.495 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%B1 1 3 4 6 7 8 21
c33 7 0 1.50529e-19 $X=1.155 $Y=0.85
r34 21 22 1.05628 $w=2.08e-07 $l=2e-08 $layer=LI1_cond $X=1.155 $Y=1.18
+ $X2=1.175 $Y2=1.18
r35 14 22 0.430812 $w=2.2e-07 $l=1.05e-07 $layer=LI1_cond $X=1.175 $Y=1.075
+ $X2=1.175 $Y2=1.18
r36 13 21 8.18615 $w=2.08e-07 $l=1.55e-07 $layer=LI1_cond $X=1 $Y=1.18 $X2=1.155
+ $Y2=1.18
r37 12 13 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1 $Y=1.16
+ $X2=1 $Y2=1.16
r38 8 22 1.32035 $w=2.08e-07 $l=2.5e-08 $layer=LI1_cond $X=1.2 $Y=1.18 $X2=1.175
+ $Y2=1.18
r39 7 14 11.7863 $w=2.18e-07 $l=2.25e-07 $layer=LI1_cond $X=1.175 $Y=0.85
+ $X2=1.175 $Y2=1.075
r40 4 12 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=1 $Y2=1.16
r41 4 6 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=0.965 $Y=1.41
+ $X2=0.965 $Y2=1.985
r42 1 12 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=0.94 $Y=0.995
+ $X2=1 $Y2=1.16
r43 1 3 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=0.94 $Y=0.995 $X2=0.94
+ $Y2=0.56
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%A1 1 3 4 6 7 8 14 15
c35 1 0 1.50529e-19 $X=1.955 $Y=1.41
r36 13 14 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=1.92
+ $Y=1.16 $X2=1.92 $Y2=1.16
r37 8 15 3.40825 $w=2.2e-07 $l=1.1e-07 $layer=LI1_cond $X=1.635 $Y=1.175
+ $X2=1.635 $Y2=1.065
r38 8 14 7.34307 $w=3.88e-07 $l=1.75e-07 $layer=LI1_cond $X=1.745 $Y=1.175
+ $X2=1.92 $Y2=1.175
r39 7 15 11.2625 $w=2.18e-07 $l=2.15e-07 $layer=LI1_cond $X=1.635 $Y=0.85
+ $X2=1.635 $Y2=1.065
r40 4 13 39.1435 $w=2.6e-07 $l=1.92678e-07 $layer=POLY_cond $X=1.98 $Y=0.995
+ $X2=1.92 $Y2=1.16
r41 4 6 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=1.98 $Y=0.995 $X2=1.98
+ $Y2=0.56
r42 1 13 50.9545 $w=2.6e-07 $l=2.66927e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.92 $Y2=1.16
r43 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=1.955 $Y=1.41
+ $X2=1.955 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%A2 1 3 4 6 7
c35 7 0 4.77488e-20 $X=2.4 $Y=1.19
r36 7 10 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.44
+ $Y=1.16 $X2=2.44 $Y2=1.16
r37 4 10 45.8513 $w=2.56e-07 $l=2.28035e-07 $layer=POLY_cond $X=2.5 $Y=0.96
+ $X2=2.44 $Y2=1.16
r38 4 6 128.533 $w=1.5e-07 $l=4e-07 $layer=POLY_cond $X=2.5 $Y=0.96 $X2=2.5
+ $Y2=0.56
r39 1 10 51.3767 $w=2.56e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.475 $Y=1.41
+ $X2=2.44 $Y2=1.16
r40 1 3 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.475 $Y=1.41
+ $X2=2.475 $Y2=1.985
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%A_27_297# 1 2 3 4 13 15 16 18 19 21 25 32
+ 33 34 38 43 44
c87 16 0 4.77488e-20 $X=3.01 $Y=0.995
r88 43 44 3.9534 $w=3.33e-07 $l=9.5e-08 $layer=LI1_cond $X=0.257 $Y=2.34
+ $X2=0.257 $Y2=2.245
r89 38 39 145.28 $w=1.7e-07 $l=1.7e-07 $layer=licon1_POLY $count=1 $X=2.95
+ $Y=1.16 $X2=2.95 $Y2=1.16
r90 36 38 21.8556 $w=1.68e-07 $l=3.35e-07 $layer=LI1_cond $X=2.95 $Y=1.495
+ $X2=2.95 $Y2=1.16
r91 35 38 24.4652 $w=1.68e-07 $l=3.75e-07 $layer=LI1_cond $X=2.95 $Y=0.785
+ $X2=2.95 $Y2=1.16
r92 33 35 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.865 $Y=0.7
+ $X2=2.95 $Y2=0.785
r93 33 34 38.1658 $w=1.68e-07 $l=5.85e-07 $layer=LI1_cond $X=2.865 $Y=0.7
+ $X2=2.28 $Y2=0.7
r94 32 34 6.81649 $w=1.7e-07 $l=1.20208e-07 $layer=LI1_cond $X=2.195 $Y=0.615
+ $X2=2.28 $Y2=0.7
r95 31 32 9.7861 $w=1.68e-07 $l=1.5e-07 $layer=LI1_cond $X=2.195 $Y=0.465
+ $X2=2.195 $Y2=0.615
r96 27 30 27.9913 $w=2.08e-07 $l=5.3e-07 $layer=LI1_cond $X=1.16 $Y=0.36
+ $X2=1.69 $Y2=0.36
r97 25 31 6.91519 $w=2.1e-07 $l=1.41244e-07 $layer=LI1_cond $X=2.11 $Y=0.36
+ $X2=2.195 $Y2=0.465
r98 25 30 22.1818 $w=2.08e-07 $l=4.2e-07 $layer=LI1_cond $X=2.11 $Y=0.36
+ $X2=1.69 $Y2=0.36
r99 22 41 3.69196 $w=2.2e-07 $l=1.28e-07 $layer=LI1_cond $X=0.345 $Y=1.605
+ $X2=0.217 $Y2=1.605
r100 22 24 44.7881 $w=2.18e-07 $l=8.55e-07 $layer=LI1_cond $X=0.345 $Y=1.605
+ $X2=1.2 $Y2=1.605
r101 21 36 6.96323 $w=2.2e-07 $l=1.46458e-07 $layer=LI1_cond $X=2.865 $Y=1.605
+ $X2=2.95 $Y2=1.495
r102 21 24 87.219 $w=2.18e-07 $l=1.665e-06 $layer=LI1_cond $X=2.865 $Y=1.605
+ $X2=1.2 $Y2=1.605
r103 19 41 3.17278 $w=2.55e-07 $l=1.1e-07 $layer=LI1_cond $X=0.217 $Y=1.715
+ $X2=0.217 $Y2=1.605
r104 19 44 23.9527 $w=2.53e-07 $l=5.3e-07 $layer=LI1_cond $X=0.217 $Y=1.715
+ $X2=0.217 $Y2=2.245
r105 16 39 39.2931 $w=2.55e-07 $l=1.92678e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=2.95 $Y2=1.16
r106 16 18 139.78 $w=1.5e-07 $l=4.35e-07 $layer=POLY_cond $X=3.01 $Y=0.995
+ $X2=3.01 $Y2=0.56
r107 13 39 51.486 $w=2.55e-07 $l=2.66927e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.95 $Y2=1.16
r108 13 15 153.972 $w=1.8e-07 $l=5.75e-07 $layer=POLY_cond $X=2.985 $Y=1.41
+ $X2=2.985 $Y2=1.985
r109 4 24 600 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_PDIFF $count=1 $X=1.055
+ $Y=1.485 $X2=1.2 $Y2=1.63
r110 3 43 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=2.34
r111 3 41 300 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_PDIFF $count=2 $X=0.135
+ $Y=1.485 $X2=0.26 $Y2=1.66
r112 2 30 182 $w=1.7e-07 $l=1.97864e-07 $layer=licon1_NDIFF $count=1 $X=1.565
+ $Y=0.235 $X2=1.69 $Y2=0.38
r113 1 27 182 $w=1.7e-07 $l=2.05061e-07 $layer=licon1_NDIFF $count=1 $X=1.015
+ $Y=0.235 $X2=1.16 $Y2=0.38
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%A_117_297# 1 2 7 11 13
r21 11 16 2.77883 $w=3.3e-07 $l=1e-07 $layer=LI1_cond $X=2.23 $Y=2.085 $X2=2.23
+ $Y2=1.985
r22 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.23 $Y=2.085
+ $X2=2.23 $Y2=2.36
r23 7 16 4.58506 $w=2e-07 $l=1.65e-07 $layer=LI1_cond $X=2.065 $Y=1.985 $X2=2.23
+ $Y2=1.985
r24 7 9 74.0318 $w=1.98e-07 $l=1.335e-06 $layer=LI1_cond $X=2.065 $Y=1.985
+ $X2=0.73 $Y2=1.985
r25 2 16 600 $w=1.7e-07 $l=5.8741e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.2 $Y2=2
r26 2 13 600 $w=1.7e-07 $l=9.63068e-07 $layer=licon1_PDIFF $count=1 $X=2.045
+ $Y=1.485 $X2=2.23 $Y2=2.36
r27 1 9 600 $w=1.7e-07 $l=5.83009e-07 $layer=licon1_PDIFF $count=1 $X=0.585
+ $Y=1.485 $X2=0.73 $Y2=2
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%VPWR 1 2 9 13 16 17 18 20 30 31 34
r44 34 35 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=1.61 $Y=2.72
+ $X2=1.61 $Y2=2.72
r45 30 31 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=2.72
+ $X2=3.45 $Y2=2.72
r46 28 31 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=3.45 $Y2=2.72
r47 28 35 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=2.72
+ $X2=1.61 $Y2=2.72
r48 27 28 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=2.53 $Y=2.72
+ $X2=2.53 $Y2=2.72
r49 25 34 9.05715 $w=1.7e-07 $l=1.78e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=1.717 $Y2=2.72
r50 25 27 41.4278 $w=1.68e-07 $l=6.35e-07 $layer=LI1_cond $X=1.895 $Y=2.72
+ $X2=2.53 $Y2=2.72
r51 20 34 9.05715 $w=1.7e-07 $l=1.77e-07 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=1.717 $Y2=2.72
r52 20 22 85.4652 $w=1.68e-07 $l=1.31e-06 $layer=LI1_cond $X=1.54 $Y=2.72
+ $X2=0.23 $Y2=2.72
r53 18 35 0.392668 $w=4.8e-07 $l=1.38e-06 $layer=MET1_cond $X=0.23 $Y=2.72
+ $X2=1.61 $Y2=2.72
r54 18 22 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=0.23 $Y=2.72
+ $X2=0.23 $Y2=2.72
r55 16 27 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=2.72
+ $X2=2.53 $Y2=2.72
r56 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=2.72
+ $X2=2.75 $Y2=2.72
r57 15 30 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=3.45 $Y2=2.72
r58 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=2.72
+ $X2=2.75 $Y2=2.72
r59 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.72
r60 11 13 21.4773 $w=3.28e-07 $l=6.15e-07 $layer=LI1_cond $X=2.75 $Y=2.635
+ $X2=2.75 $Y2=2.02
r61 7 34 1.11826 $w=3.55e-07 $l=8.5e-08 $layer=LI1_cond $X=1.717 $Y=2.635
+ $X2=1.717 $Y2=2.72
r62 7 9 9.57664 $w=3.53e-07 $l=2.95e-07 $layer=LI1_cond $X=1.717 $Y=2.635
+ $X2=1.717 $Y2=2.34
r63 2 13 300 $w=1.7e-07 $l=6.20645e-07 $layer=licon1_PDIFF $count=2 $X=2.565
+ $Y=1.485 $X2=2.75 $Y2=2.02
r64 1 9 600 $w=1.7e-07 $l=9.15369e-07 $layer=licon1_PDIFF $count=1 $X=1.595
+ $Y=1.485 $X2=1.72 $Y2=2.34
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%X 1 2 10 13 14 30
r16 19 30 1.99461 $w=2.58e-07 $l=4.5e-08 $layer=LI1_cond $X=3.405 $Y=1.915
+ $X2=3.405 $Y2=1.87
r17 13 30 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.405 $Y=1.85
+ $X2=3.405 $Y2=1.87
r18 13 14 12.1893 $w=2.58e-07 $l=2.75e-07 $layer=LI1_cond $X=3.405 $Y=1.935
+ $X2=3.405 $Y2=2.21
r19 13 19 0.886495 $w=2.58e-07 $l=2e-08 $layer=LI1_cond $X=3.405 $Y=1.935
+ $X2=3.405 $Y2=1.915
r20 11 13 50.6043 $w=2.78e-07 $l=1.2e-06 $layer=LI1_cond $X=3.45 $Y=0.585
+ $X2=3.45 $Y2=1.785
r21 10 11 4.62375 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=3.45 $Y=0.42
+ $X2=3.45 $Y2=0.585
r22 8 10 3.14303 $w=3.28e-07 $l=9e-08 $layer=LI1_cond $X=3.36 $Y=0.42 $X2=3.45
+ $Y2=0.42
r23 2 13 300 $w=1.7e-07 $l=6.00833e-07 $layer=licon1_PDIFF $count=2 $X=3.075
+ $Y=1.485 $X2=3.36 $Y2=1.96
r24 1 8 182 $w=1.7e-07 $l=3.55668e-07 $layer=licon1_NDIFF $count=1 $X=3.085
+ $Y=0.235 $X2=3.36 $Y2=0.42
.ends

.subckt PM_SKY130_FD_SC_HDLL__A22O_1%VGND 1 2 7 9 13 16 17 18 28 29
r39 28 29 4.65 $w=1.7e-07 $l=3.4e-07 $layer=mcon $count=2 $X=3.45 $Y=0 $X2=3.45
+ $Y2=0
r40 26 29 0.261778 $w=4.8e-07 $l=9.2e-07 $layer=MET1_cond $X=2.53 $Y=0 $X2=3.45
+ $Y2=0
r41 25 26 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=2.53 $Y=0 $X2=2.53
+ $Y2=0
r42 23 26 0.523557 $w=4.8e-07 $l=1.84e-06 $layer=MET1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r43 22 25 120.043 $w=1.68e-07 $l=1.84e-06 $layer=LI1_cond $X=0.69 $Y=0 $X2=2.53
+ $Y2=0
r44 22 23 3.72 $w=1.7e-07 $l=4.25e-07 $layer=mcon $count=2 $X=0.69 $Y=0 $X2=0.69
+ $Y2=0
r45 20 32 6.45619 $w=1.7e-07 $l=2.98e-07 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.297
+ $Y2=0
r46 20 22 6.19786 $w=1.68e-07 $l=9.5e-08 $layer=LI1_cond $X=0.595 $Y=0 $X2=0.69
+ $Y2=0
r47 18 23 0.130889 $w=4.8e-07 $l=4.6e-07 $layer=MET1_cond $X=0.23 $Y=0 $X2=0.69
+ $Y2=0
r48 18 32 9.3 $w=1.7e-07 $l=1.7e-07 $layer=mcon $count=1 $X=0.23 $Y=0 $X2=0.23
+ $Y2=0
r49 16 25 3.58824 $w=1.68e-07 $l=5.5e-08 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.53
+ $Y2=0
r50 16 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.585 $Y=0 $X2=2.75
+ $Y2=0
r51 15 28 34.9037 $w=1.68e-07 $l=5.35e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=3.45
+ $Y2=0
r52 15 17 8.61065 $w=1.7e-07 $l=1.65e-07 $layer=LI1_cond $X=2.915 $Y=0 $X2=2.75
+ $Y2=0
r53 11 17 0.89609 $w=3.3e-07 $l=8.5e-08 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0
r54 11 13 9.60369 $w=3.28e-07 $l=2.75e-07 $layer=LI1_cond $X=2.75 $Y=0.085
+ $X2=2.75 $Y2=0.36
r55 7 32 2.81646 $w=5.05e-07 $l=1.05119e-07 $layer=LI1_cond $X=0.342 $Y=0.085
+ $X2=0.297 $Y2=0
r56 7 9 7.46069 $w=5.03e-07 $l=3.15e-07 $layer=LI1_cond $X=0.342 $Y=0.085
+ $X2=0.342 $Y2=0.4
r57 2 13 182 $w=1.7e-07 $l=2.29129e-07 $layer=licon1_NDIFF $count=1 $X=2.575
+ $Y=0.235 $X2=2.75 $Y2=0.36
r58 1 9 91 $w=1.7e-07 $l=2.18746e-07 $layer=licon1_NDIFF $count=2 $X=0.135
+ $Y=0.235 $X2=0.26 $Y2=0.4
.ends

