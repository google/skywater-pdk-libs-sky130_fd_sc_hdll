# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
PROPERTYDEFINITIONS
  MACRO maskLayoutSubType STRING ;
  MACRO prCellType STRING ;
  MACRO originalViewName STRING ;
END PROPERTYDEFINITIONS
MACRO sky130_fd_sc_hdll__a21bo_1
  ORIGIN  0.000000  0.000000 ;
  CLASS CORE ;
  SYMMETRY X Y R90 ;
  SIZE  4.140000 BY  2.720000 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.900000 0.995000 2.275000 1.615000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.277500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.445000 0.995000 2.705000 1.615000 ;
    END
  END A2
  PIN B1_N
    ANTENNAGATEAREA  0.138600 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.105000 0.325000 0.335000 1.665000 ;
    END
  END B1_N
  PIN X
    ANTENNADIFFAREA  0.628800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.715000 0.265000 3.995000 2.455000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.140000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met1 ;
        RECT 0.000000 2.480000 4.140000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.000000 -0.085000 4.140000 0.085000 ;
      RECT 0.000000  2.635000 4.140000 2.805000 ;
      RECT 0.105000  1.845000 0.965000 2.045000 ;
      RECT 0.105000  2.045000 0.345000 2.435000 ;
      RECT 0.515000  0.265000 0.795000 1.165000 ;
      RECT 0.515000  1.165000 0.965000 1.845000 ;
      RECT 0.515000  2.225000 0.915000 2.635000 ;
      RECT 1.045000  0.085000 1.290000 0.865000 ;
      RECT 1.135000  1.045000 1.730000 1.345000 ;
      RECT 1.135000  1.345000 1.465000 2.455000 ;
      RECT 1.460000  0.265000 1.940000 0.625000 ;
      RECT 1.460000  0.625000 3.545000 0.815000 ;
      RECT 1.460000  0.815000 1.730000 1.045000 ;
      RECT 1.685000  1.785000 2.810000 1.985000 ;
      RECT 1.685000  1.985000 1.865000 2.455000 ;
      RECT 2.035000  2.155000 2.415000 2.635000 ;
      RECT 2.620000  0.085000 3.350000 0.455000 ;
      RECT 2.640000  1.985000 2.810000 2.455000 ;
      RECT 3.075000  1.495000 3.360000 2.635000 ;
      RECT 3.285000  0.815000 3.545000 1.325000 ;
    LAYER mcon ;
      RECT 0.145000 -0.085000 0.315000 0.085000 ;
      RECT 0.145000  2.635000 0.315000 2.805000 ;
      RECT 0.605000 -0.085000 0.775000 0.085000 ;
      RECT 0.605000  2.635000 0.775000 2.805000 ;
      RECT 1.065000 -0.085000 1.235000 0.085000 ;
      RECT 1.065000  2.635000 1.235000 2.805000 ;
      RECT 1.525000 -0.085000 1.695000 0.085000 ;
      RECT 1.525000  2.635000 1.695000 2.805000 ;
      RECT 1.985000 -0.085000 2.155000 0.085000 ;
      RECT 1.985000  2.635000 2.155000 2.805000 ;
      RECT 2.445000 -0.085000 2.615000 0.085000 ;
      RECT 2.445000  2.635000 2.615000 2.805000 ;
      RECT 2.905000 -0.085000 3.075000 0.085000 ;
      RECT 2.905000  2.635000 3.075000 2.805000 ;
      RECT 3.365000 -0.085000 3.535000 0.085000 ;
      RECT 3.365000  2.635000 3.535000 2.805000 ;
      RECT 3.825000 -0.085000 3.995000 0.085000 ;
      RECT 3.825000  2.635000 3.995000 2.805000 ;
  END
  PROPERTY maskLayoutSubType "abstract" ;
  PROPERTY prCellType "standard" ;
  PROPERTY originalViewName "layout" ;
END sky130_fd_sc_hdll__a21bo_1
END LIBRARY
