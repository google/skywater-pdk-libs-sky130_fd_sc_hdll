* File: sky130_fd_sc_hdll__nand2b_1.pxi.spice
* Created: Thu Aug 27 19:13:16 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%A_N N_A_N_c_39_n N_A_N_M1000_g N_A_N_c_36_n
+ N_A_N_M1002_g A_N N_A_N_c_38_n PM_SKY130_FD_SC_HDLL__NAND2B_1%A_N
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%B N_B_c_62_n N_B_M1003_g N_B_c_63_n N_B_M1005_g
+ B N_B_c_64_n B PM_SKY130_FD_SC_HDLL__NAND2B_1%B
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%A_27_93# N_A_27_93#_M1002_s N_A_27_93#_M1000_s
+ N_A_27_93#_c_90_n N_A_27_93#_M1004_g N_A_27_93#_c_91_n N_A_27_93#_M1001_g
+ N_A_27_93#_c_92_n N_A_27_93#_c_101_n N_A_27_93#_c_93_n N_A_27_93#_c_94_n
+ N_A_27_93#_c_97_n PM_SKY130_FD_SC_HDLL__NAND2B_1%A_27_93#
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%VPWR N_VPWR_M1000_d N_VPWR_M1001_d
+ N_VPWR_c_147_n N_VPWR_c_148_n N_VPWR_c_149_n N_VPWR_c_150_n VPWR
+ N_VPWR_c_151_n N_VPWR_c_146_n N_VPWR_c_153_n VPWR
+ PM_SKY130_FD_SC_HDLL__NAND2B_1%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%Y N_Y_M1004_d N_Y_M1003_d N_Y_c_186_n
+ N_Y_c_189_n N_Y_c_183_n Y Y Y Y Y N_Y_c_180_n N_Y_c_182_n
+ PM_SKY130_FD_SC_HDLL__NAND2B_1%Y
x_PM_SKY130_FD_SC_HDLL__NAND2B_1%VGND N_VGND_M1002_d N_VGND_c_216_n VGND
+ N_VGND_c_217_n N_VGND_c_218_n N_VGND_c_219_n VGND
+ PM_SKY130_FD_SC_HDLL__NAND2B_1%VGND
cc_1 VNB N_A_N_c_36_n 0.0240622f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_2 VNB A_N 0.0087467f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_3 VNB N_A_N_c_38_n 0.0390945f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.202
cc_4 VNB N_B_c_62_n 0.0206983f $X=-0.19 $Y=-0.24 $X2=0.495 $Y2=1.41
cc_5 VNB N_B_c_63_n 0.0192949f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=0.995
cc_6 VNB N_B_c_64_n 0.00461842f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_7 VNB N_A_27_93#_c_90_n 0.0200176f $X=-0.19 $Y=-0.24 $X2=0.15 $Y2=1.105
cc_8 VNB N_A_27_93#_c_91_n 0.0254925f $X=-0.19 $Y=-0.24 $X2=0.255 $Y2=1.16
cc_9 VNB N_A_27_93#_c_92_n 0.00746583f $X=-0.19 $Y=-0.24 $X2=0.52 $Y2=1.202
cc_10 VNB N_A_27_93#_c_93_n 8.65037e-19 $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_11 VNB N_A_27_93#_c_94_n 0.0166438f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_12 VNB N_VPWR_c_146_n 0.0989421f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB Y 0.04123f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_14 VNB N_Y_c_180_n 0.0177534f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_15 VNB N_VGND_c_216_n 0.0108309f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_16 VNB N_VGND_c_217_n 0.0353821f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_17 VNB N_VGND_c_218_n 0.151575f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_18 VNB N_VGND_c_219_n 0.0260346f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VPB N_A_N_c_39_n 0.0244803f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_20 VPB A_N 5.51043e-19 $X=-0.19 $Y=1.305 $X2=0.15 $Y2=1.105
cc_21 VPB N_A_N_c_38_n 0.0172642f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_22 VPB N_B_c_62_n 0.0279612f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_23 VPB N_B_c_64_n 0.00308028f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_24 VPB N_A_27_93#_c_91_n 0.0297152f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_25 VPB N_A_27_93#_c_93_n 0.0015454f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_26 VPB N_A_27_93#_c_97_n 0.0145649f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_27 VPB N_VPWR_c_147_n 0.0233057f $X=-0.19 $Y=1.305 $X2=0.255 $Y2=1.16
cc_28 VPB N_VPWR_c_148_n 0.0158916f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_29 VPB N_VPWR_c_149_n 0.0197985f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_30 VPB N_VPWR_c_150_n 0.00410791f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_31 VPB N_VPWR_c_151_n 0.0147471f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_32 VPB N_VPWR_c_146_n 0.0656045f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_33 VPB N_VPWR_c_153_n 0.0269706f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_34 VPB Y 0.0278693f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_35 VPB N_Y_c_182_n 0.0137276f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_36 N_A_N_c_39_n N_B_c_62_n 0.0175647f $X=0.495 $Y=1.41 $X2=-0.19 $Y2=-0.24
cc_37 N_A_N_c_38_n N_B_c_62_n 0.0210399f $X=0.495 $Y=1.202 $X2=-0.19 $Y2=-0.24
cc_38 N_A_N_c_36_n N_B_c_63_n 0.0166248f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_39 A_N N_B_c_64_n 0.0187966f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_40 N_A_N_c_38_n N_B_c_64_n 0.00634897f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_41 N_A_N_c_36_n N_A_27_93#_c_92_n 0.012567f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_42 A_N N_A_27_93#_c_92_n 0.00435033f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_43 N_A_N_c_38_n N_A_27_93#_c_92_n 0.00240586f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_44 N_A_N_c_39_n N_A_27_93#_c_101_n 0.0170092f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_45 A_N N_A_27_93#_c_101_n 0.0021049f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_46 A_N N_A_27_93#_c_94_n 0.0212525f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_47 N_A_N_c_38_n N_A_27_93#_c_94_n 0.00626797f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_48 A_N N_A_27_93#_c_97_n 0.0196991f $X=0.15 $Y=1.105 $X2=0 $Y2=0
cc_49 N_A_N_c_38_n N_A_27_93#_c_97_n 0.00588109f $X=0.495 $Y=1.202 $X2=0 $Y2=0
cc_50 N_A_N_c_39_n N_VPWR_c_147_n 0.00390207f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_51 N_A_N_c_39_n N_VPWR_c_146_n 0.00500987f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_52 N_A_N_c_39_n N_VPWR_c_153_n 0.00393512f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_53 N_A_N_c_36_n N_VGND_c_216_n 0.0042306f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_54 N_A_N_c_36_n N_VGND_c_218_n 0.00512902f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_55 N_A_N_c_36_n N_VGND_c_219_n 0.00399957f $X=0.52 $Y=0.995 $X2=0 $Y2=0
cc_56 N_B_c_63_n N_A_27_93#_c_90_n 0.0307109f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_57 N_B_c_62_n N_A_27_93#_c_91_n 0.0551998f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_58 N_B_c_64_n N_A_27_93#_c_91_n 0.00176242f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_59 N_B_c_62_n N_A_27_93#_c_92_n 0.00314143f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_60 N_B_c_63_n N_A_27_93#_c_92_n 0.0126703f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_61 N_B_c_64_n N_A_27_93#_c_92_n 0.0443393f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_62 N_B_c_62_n N_A_27_93#_c_101_n 0.0170695f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_63 N_B_c_64_n N_A_27_93#_c_101_n 0.036075f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_64 N_B_c_62_n N_A_27_93#_c_93_n 0.00132101f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_65 N_B_c_63_n N_A_27_93#_c_93_n 9.99298e-19 $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_66 N_B_c_64_n N_A_27_93#_c_93_n 0.0136458f $X=0.995 $Y=1.16 $X2=0 $Y2=0
cc_67 N_B_c_62_n N_VPWR_c_147_n 0.00672788f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_68 N_B_c_62_n N_VPWR_c_149_n 0.00597712f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_69 N_B_c_62_n N_VPWR_c_146_n 0.0113021f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_70 N_B_c_62_n N_Y_c_183_n 0.0106076f $X=1.03 $Y=1.41 $X2=0 $Y2=0
cc_71 N_B_c_63_n N_VGND_c_216_n 0.00482545f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_72 N_B_c_63_n N_VGND_c_217_n 0.00439206f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_73 N_B_c_63_n N_VGND_c_218_n 0.00723496f $X=1.055 $Y=0.995 $X2=0 $Y2=0
cc_74 N_A_27_93#_c_101_n N_VPWR_M1000_d 0.00509529f $X=1.45 $Y=1.58 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_27_93#_c_101_n N_VPWR_c_147_n 0.019282f $X=1.45 $Y=1.58 $X2=0 $Y2=0
cc_76 N_A_27_93#_c_91_n N_VPWR_c_148_n 0.00584657f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_77 N_A_27_93#_c_91_n N_VPWR_c_149_n 0.00514793f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_78 N_A_27_93#_c_91_n N_VPWR_c_146_n 0.00789758f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_79 N_A_27_93#_c_92_n N_Y_M1004_d 0.00193245f $X=1.45 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_27_93#_c_101_n N_Y_M1003_d 0.00506813f $X=1.45 $Y=1.58 $X2=0 $Y2=0
cc_81 N_A_27_93#_c_90_n N_Y_c_186_n 0.00868471f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_82 N_A_27_93#_c_91_n N_Y_c_186_n 0.001689f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_83 N_A_27_93#_c_92_n N_Y_c_186_n 0.010852f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_84 N_A_27_93#_c_91_n N_Y_c_189_n 0.0135727f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_85 N_A_27_93#_c_101_n N_Y_c_189_n 0.0119102f $X=1.45 $Y=1.58 $X2=0 $Y2=0
cc_86 N_A_27_93#_c_91_n N_Y_c_183_n 0.011734f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_87 N_A_27_93#_c_101_n N_Y_c_183_n 0.0209598f $X=1.45 $Y=1.58 $X2=0 $Y2=0
cc_88 N_A_27_93#_c_90_n Y 0.00757532f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_89 N_A_27_93#_c_91_n Y 0.0159933f $X=1.5 $Y=1.41 $X2=0 $Y2=0
cc_90 N_A_27_93#_c_92_n Y 0.0129994f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_91 N_A_27_93#_c_93_n Y 0.04042f $X=1.535 $Y=1.16 $X2=0 $Y2=0
cc_92 N_A_27_93#_c_92_n N_VGND_M1002_d 0.00315224f $X=1.45 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_93 N_A_27_93#_c_92_n N_VGND_c_216_n 0.0193134f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_94 N_A_27_93#_c_90_n N_VGND_c_217_n 0.00357877f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_95 N_A_27_93#_c_92_n N_VGND_c_217_n 0.004883f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_96 N_A_27_93#_c_90_n N_VGND_c_218_n 0.00657948f $X=1.475 $Y=0.995 $X2=0 $Y2=0
cc_97 N_A_27_93#_c_92_n N_VGND_c_218_n 0.0180715f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_98 N_A_27_93#_c_94_n N_VGND_c_218_n 0.00852335f $X=0.26 $Y=0.69 $X2=0 $Y2=0
cc_99 N_A_27_93#_c_92_n N_VGND_c_219_n 0.00304573f $X=1.45 $Y=0.82 $X2=0 $Y2=0
cc_100 N_A_27_93#_c_94_n N_VGND_c_219_n 0.00647838f $X=0.26 $Y=0.69 $X2=0 $Y2=0
cc_101 N_A_27_93#_c_92_n A_226_47# 0.00302426f $X=1.45 $Y=0.82 $X2=-0.19
+ $Y2=-0.24
cc_102 N_VPWR_c_146_n N_Y_M1003_d 0.00231261f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_103 N_VPWR_M1001_d N_Y_c_189_n 0.00823846f $X=1.59 $Y=1.485 $X2=0 $Y2=0
cc_104 N_VPWR_c_148_n N_Y_c_189_n 0.0131603f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_105 N_VPWR_c_149_n N_Y_c_189_n 0.00267292f $X=1.65 $Y=2.72 $X2=0 $Y2=0
cc_106 N_VPWR_c_146_n N_Y_c_189_n 0.00570853f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_107 N_VPWR_c_147_n N_Y_c_183_n 0.0490267f $X=0.795 $Y=2 $X2=0 $Y2=0
cc_108 N_VPWR_c_148_n N_Y_c_183_n 0.0180622f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_109 N_VPWR_c_149_n N_Y_c_183_n 0.0222542f $X=1.65 $Y=2.72 $X2=0 $Y2=0
cc_110 N_VPWR_c_146_n N_Y_c_183_n 0.0139813f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_111 N_VPWR_M1001_d Y 0.00468004f $X=1.59 $Y=1.485 $X2=0 $Y2=0
cc_112 N_VPWR_M1001_d N_Y_c_182_n 7.9691e-19 $X=1.59 $Y=1.485 $X2=0 $Y2=0
cc_113 N_VPWR_c_148_n N_Y_c_182_n 0.00376703f $X=1.735 $Y=2.34 $X2=0 $Y2=0
cc_114 N_VPWR_c_151_n N_Y_c_182_n 0.00561964f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_115 N_VPWR_c_146_n N_Y_c_182_n 0.00944587f $X=2.07 $Y=2.72 $X2=0 $Y2=0
cc_116 N_Y_c_186_n N_VGND_c_217_n 0.0269271f $X=1.82 $Y=0.4 $X2=0 $Y2=0
cc_117 N_Y_c_180_n N_VGND_c_217_n 0.0264722f $X=2.005 $Y=0.545 $X2=0 $Y2=0
cc_118 N_Y_M1004_d N_VGND_c_218_n 0.00250335f $X=1.55 $Y=0.235 $X2=0 $Y2=0
cc_119 N_Y_c_186_n N_VGND_c_218_n 0.0165764f $X=1.82 $Y=0.4 $X2=0 $Y2=0
cc_120 N_Y_c_180_n N_VGND_c_218_n 0.0142494f $X=2.005 $Y=0.545 $X2=0 $Y2=0
cc_121 N_VGND_c_218_n A_226_47# 0.00334583f $X=2.07 $Y=0 $X2=-0.19 $Y2=-0.24
