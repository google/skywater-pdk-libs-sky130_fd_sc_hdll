* File: sky130_fd_sc_hdll__muxb4to1_4.spice
* Created: Thu Aug 27 19:11:59 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__muxb4to1_4.pex.spice"
.subckt sky130_fd_sc_hdll__muxb4to1_4  VNB VPB D[0] S[0] S[1] D[1] D[2] S[2]
+ S[3] D[3] VPWR Z VGND
* 
* VGND	VGND
* Z	Z
* VPWR	VPWR
* D[3]	D[3]
* S[3]	S[3]
* S[2]	S[2]
* D[2]	D[2]
* D[1]	D[1]
* S[1]	S[1]
* S[0]	S[0]
* D[0]	D[0]
* VPB	VPB
* VNB	VNB
MM1024 N_VGND_M1024_d N_D[0]_M1024_g N_A_119_47#_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1057 N_VGND_M1057_d N_D[0]_M1057_g N_A_119_47#_M1024_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1073 N_VGND_M1057_d N_D[0]_M1073_g N_A_119_47#_M1073_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1078 N_VGND_M1078_d N_D[0]_M1078_g N_A_119_47#_M1073_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1015 N_A_119_47#_M1015_d N_S[0]_M1015_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1023 N_A_119_47#_M1023_d N_S[0]_M1023_g N_Z_M1015_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1028 N_A_119_47#_M1023_d N_S[0]_M1028_g N_Z_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1037 N_A_119_47#_M1037_d N_S[0]_M1037_g N_Z_M1028_s VNB NSHORT L=0.15 W=0.52
+ AD=0.1352 AS=0.0702 PD=1.56 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1046 N_A_559_265#_M1046_d N_S[0]_M1046_g N_VGND_M1046_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1053 N_A_559_265#_M1046_d N_S[0]_M1053_g N_VGND_M1053_s VNB NSHORT L=0.15
+ W=0.42 AD=0.0567 AS=0.1092 PD=0.69 PS=1.36 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1061 N_VGND_M1061_d N_S[1]_M1061_g N_A_1430_325#_M1061_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1069 N_VGND_M1069_d N_S[1]_M1069_g N_A_1430_325#_M1061_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1007 N_Z_M1007_d N_S[1]_M1007_g N_A_1693_66#_M1007_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1016 N_Z_M1007_d N_S[1]_M1016_g N_A_1693_66#_M1016_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1026 N_Z_M1026_d N_S[1]_M1026_g N_A_1693_66#_M1016_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1033 N_Z_M1026_d N_S[1]_M1033_g N_A_1693_66#_M1033_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1017 N_VGND_M1017_d N_D[1]_M1017_g N_A_1693_66#_M1017_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1029 N_VGND_M1029_d N_D[1]_M1029_g N_A_1693_66#_M1017_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1049 N_VGND_M1029_d N_D[1]_M1049_g N_A_1693_66#_M1049_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1079 N_VGND_M1079_d N_D[1]_M1079_g N_A_1693_66#_M1049_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1002 N_A_2695_47#_M1002_d N_D[2]_M1002_g N_VGND_M1002_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.5 A=0.0975 P=1.6 MULT=1
MM1021 N_A_2695_47#_M1002_d N_D[2]_M1021_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75000.7 SB=75001.1 A=0.0975 P=1.6 MULT=1
MM1034 N_A_2695_47#_M1034_d N_D[2]_M1034_g N_VGND_M1021_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75000.6 A=0.0975 P=1.6 MULT=1
MM1052 N_A_2695_47#_M1034_d N_D[2]_M1052_g N_VGND_M1052_s VNB NSHORT L=0.15
+ W=0.65 AD=0.08775 AS=0.169 PD=0.92 PS=1.82 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.6 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1008 N_Z_M1008_d N_S[2]_M1008_g N_A_2695_47#_M1008_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1009 N_Z_M1008_d N_S[2]_M1009_g N_A_2695_47#_M1009_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1030 N_Z_M1030_d N_S[2]_M1030_g N_A_2695_47#_M1009_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1077 N_Z_M1030_d N_S[2]_M1077_g N_A_2695_47#_M1077_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1058 N_VGND_M1058_d N_S[2]_M1058_g N_A_3135_265#_M1058_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1062 N_VGND_M1062_d N_S[2]_M1062_g N_A_3135_265#_M1058_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1059 N_VGND_M1059_d N_S[3]_M1059_g N_A_4006_325#_M1059_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.2
+ SB=75000.6 A=0.063 P=1.14 MULT=1
MM1075 N_VGND_M1075_d N_S[3]_M1075_g N_A_4006_325#_M1059_s VNB NSHORT L=0.15
+ W=0.42 AD=0.1092 AS=0.0567 PD=1.36 PS=0.69 NRD=0 NRS=0 M=1 R=2.8 SA=75000.6
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1011 N_Z_M1011_d N_S[3]_M1011_g N_A_4269_66#_M1011_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.2
+ SB=75001.4 A=0.078 P=1.34 MULT=1
MM1012 N_Z_M1011_d N_S[3]_M1012_g N_A_4269_66#_M1012_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75000.6
+ SB=75001 A=0.078 P=1.34 MULT=1
MM1022 N_Z_M1022_d N_S[3]_M1022_g N_A_4269_66#_M1012_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.0702 PD=0.79 PS=0.79 NRD=0 NRS=0 M=1 R=3.46667 SA=75001
+ SB=75000.6 A=0.078 P=1.34 MULT=1
MM1031 N_Z_M1022_d N_S[3]_M1031_g N_A_4269_66#_M1031_s VNB NSHORT L=0.15 W=0.52
+ AD=0.0702 AS=0.1352 PD=0.79 PS=1.56 NRD=0 NRS=0 M=1 R=3.46667 SA=75001.4
+ SB=75000.2 A=0.078 P=1.34 MULT=1
MM1013 N_VGND_M1013_d N_D[3]_M1013_g N_A_4269_66#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.169 AS=0.08775 PD=1.82 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75000.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1032 N_VGND_M1032_d N_D[3]_M1032_g N_A_4269_66#_M1013_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75000.6 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1040 N_VGND_M1032_d N_D[3]_M1040_g N_A_4269_66#_M1040_s VNB NSHORT L=0.15
+ W=0.65 AD=0.12025 AS=0.08775 PD=1.02 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333
+ SA=75001.1 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1054 N_VGND_M1054_d N_D[3]_M1054_g N_A_4269_66#_M1040_s VNB NSHORT L=0.15
+ W=0.65 AD=0.2015 AS=0.08775 PD=1.92 PS=0.92 NRD=0 NRS=0 M=1 R=4.33333
+ SA=75001.5 SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_D[0]_M1003_g N_A_117_297#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1041 N_VPWR_M1041_d N_D[0]_M1041_g N_A_117_297#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1055 N_VPWR_M1041_d N_D[0]_M1055_g N_A_117_297#_M1055_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1071 N_VPWR_M1071_d N_D[0]_M1071_g N_A_117_297#_M1055_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1042 N_A_117_297#_M1042_d N_A_559_265#_M1042_g N_Z_M1042_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1056 N_A_117_297#_M1056_d N_A_559_265#_M1056_g N_Z_M1042_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1063 N_A_117_297#_M1056_d N_A_559_265#_M1063_g N_Z_M1063_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1072 N_A_117_297#_M1072_d N_A_559_265#_M1072_g N_Z_M1063_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1004 N_VPWR_M1004_d N_S[0]_M1004_g N_A_559_265#_M1004_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1018 N_VPWR_M1018_d N_S[0]_M1018_g N_A_559_265#_M1004_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1036 N_VPWR_M1036_d N_S[1]_M1036_g N_A_1430_325#_M1036_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1050 N_VPWR_M1050_d N_S[1]_M1050_g N_A_1430_325#_M1036_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1000 N_Z_M1000_d N_A_1430_325#_M1000_g N_A_1643_311#_M1000_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1014 N_Z_M1000_d N_A_1430_325#_M1014_g N_A_1643_311#_M1014_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1043 N_Z_M1043_d N_A_1430_325#_M1043_g N_A_1643_311#_M1014_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1066 N_Z_M1043_d N_A_1430_325#_M1066_g N_A_1643_311#_M1066_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1001 N_A_1643_311#_M1001_d N_D[1]_M1001_g N_VPWR_M1001_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_A_1643_311#_M1001_d N_D[1]_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1038 N_A_1643_311#_M1038_d N_D[1]_M1038_g N_VPWR_M1006_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1065 N_A_1643_311#_M1038_d N_D[1]_M1065_g N_VPWR_M1065_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_2693_297#_M1005_d N_D[2]_M1005_g N_VPWR_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1019 N_A_2693_297#_M1005_d N_D[2]_M1019_g N_VPWR_M1019_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1047 N_A_2693_297#_M1047_d N_D[2]_M1047_g N_VPWR_M1019_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1074 N_A_2693_297#_M1047_d N_D[2]_M1074_g N_VPWR_M1074_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.27 PD=1.29 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
MM1025 N_A_2693_297#_M1025_d N_A_3135_265#_M1025_g N_Z_M1025_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1044 N_A_2693_297#_M1044_d N_A_3135_265#_M1044_g N_Z_M1025_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1051 N_A_2693_297#_M1044_d N_A_3135_265#_M1051_g N_Z_M1051_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1064 N_A_2693_297#_M1064_d N_A_3135_265#_M1064_g N_Z_M1051_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1020 N_A_3135_265#_M1020_d N_S[2]_M1020_g N_VPWR_M1020_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1076 N_A_3135_265#_M1020_d N_S[2]_M1076_g N_VPWR_M1076_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1045 N_A_4006_325#_M1045_d N_S[3]_M1045_g N_VPWR_M1045_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.2 SB=90000.6 A=0.1476 P=2 MULT=1
MM1067 N_A_4006_325#_M1045_d N_S[3]_M1067_g N_VPWR_M1067_s VPB PHIGHVT L=0.18
+ W=0.82 AD=0.1189 AS=0.2214 PD=1.11 PS=2.18 NRD=1.182 NRS=1.182 M=1 R=4.55556
+ SA=90000.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1039 N_A_4219_311#_M1039_d N_A_4006_325#_M1039_g N_Z_M1039_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.2 SB=90001.6 A=0.1476 P=2 MULT=1
MM1048 N_A_4219_311#_M1048_d N_A_4006_325#_M1048_g N_Z_M1039_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90000.6 SB=90001.1 A=0.1476 P=2 MULT=1
MM1060 N_A_4219_311#_M1048_d N_A_4006_325#_M1060_g N_Z_M1060_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.1189 AS=0.1189 PD=1.11 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.1 SB=90000.6 A=0.1476 P=2 MULT=1
MM1068 N_A_4219_311#_M1068_d N_A_4006_325#_M1068_g N_Z_M1060_s VPB PHIGHVT
+ L=0.18 W=0.82 AD=0.2214 AS=0.1189 PD=2.18 PS=1.11 NRD=1.182 NRS=1.182 M=1
+ R=4.55556 SA=90001.6 SB=90000.2 A=0.1476 P=2 MULT=1
MM1010 N_VPWR_M1010_d N_D[3]_M1010_g N_A_4219_311#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1027 N_VPWR_M1027_d N_D[3]_M1027_g N_A_4219_311#_M1010_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1035 N_VPWR_M1027_d N_D[3]_M1035_g N_A_4219_311#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.1 SB=90000.6 A=0.18 P=2.36 MULT=1
MM1070 N_VPWR_M1070_d N_D[3]_M1070_g N_A_4219_311#_M1035_s VPB PHIGHVT L=0.18
+ W=1 AD=0.27 AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX80_noxref VNB VPB NWDIODE A=41.9547 P=55.49
c_485 VPB 0 4.83259e-19 $X=25.445 $Y=2.635
*
.include "sky130_fd_sc_hdll__muxb4to1_4.pxi.spice"
*
.ends
*
*
