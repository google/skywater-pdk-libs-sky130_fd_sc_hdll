* File: sky130_fd_sc_hdll__or2_4.spice
* Created: Wed Sep  2 08:47:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__or2_4.pex.spice"
.subckt sky130_fd_sc_hdll__or2_4  VNB VPB B A VPWR X VGND
* 
* VGND	VGND
* X	X
* VPWR	VPWR
* A	A
* B	B
* VPB	VPB
* VNB	VNB
MM1009 N_A_35_297#_M1009_d N_B_M1009_g N_VGND_M1009_s VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.2015 PD=0.92 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75002.6 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_A_35_297#_M1009_d VNB NSHORT L=0.15 W=0.65
+ AD=0.131625 AS=0.08775 PD=1.055 PS=0.92 NRD=16.608 NRS=0 M=1 R=4.33333
+ SA=75000.7 SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1000 N_VGND_M1004_d N_A_35_297#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.131625 AS=0.104 PD=1.055 PS=0.97 NRD=6.456 NRS=8.304 M=1 R=4.33333
+ SA=75001.2 SB=75001.6 A=0.0975 P=1.6 MULT=1
MM1005 N_VGND_M1005_d N_A_35_297#_M1005_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.104 PD=0.97 PS=0.97 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7
+ SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 N_VGND_M1005_d N_A_35_297#_M1007_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.104 AS=0.12025 PD=0.97 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.1
+ SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1008 N_VGND_M1008_d N_A_35_297#_M1008_g N_X_M1007_s VNB NSHORT L=0.15 W=0.65
+ AD=0.169 AS=0.12025 PD=1.82 PS=1.02 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75002.7
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 A_129_297# N_B_M1003_g N_A_35_297#_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.115 AS=0.29 PD=1.23 PS=2.58 NRD=11.8003 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90002.6 A=0.18 P=2.36 MULT=1
MM1001 N_VPWR_M1001_d N_A_M1001_g A_129_297# VPB PHIGHVT L=0.18 W=1 AD=0.1875
+ AS=0.115 PD=1.375 PS=1.23 NRD=9.8303 NRS=11.8003 M=1 R=5.55556 SA=90000.6
+ SB=90002.2 A=0.18 P=2.36 MULT=1
MM1002 N_X_M1002_d N_A_35_297#_M1002_g N_VPWR_M1001_d VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.1875 PD=1.29 PS=1.375 NRD=0.9653 NRS=8.8453 M=1 R=5.55556
+ SA=90001.2 SB=90001.6 A=0.18 P=2.36 MULT=1
MM1006 N_X_M1002_d N_A_35_297#_M1006_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90001.6 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1010 N_X_M1010_d N_A_35_297#_M1010_g N_VPWR_M1006_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.145 PD=1.29 PS=1.29 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.1 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1011 N_X_M1010_d N_A_35_297#_M1011_g N_VPWR_M1011_s VPB PHIGHVT L=0.18 W=1
+ AD=0.145 AS=0.29 PD=1.29 PS=2.58 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90002.6 SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=6.5163 P=11.33
c_234 A_129_297# 0 1.05688e-19 $X=0.645 $Y=1.485
*
.include "sky130_fd_sc_hdll__or2_4.pxi.spice"
*
.ends
*
*
