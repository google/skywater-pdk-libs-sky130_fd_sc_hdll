* File: sky130_fd_sc_hdll__nand2_16.pxi.spice
* Created: Thu Aug 27 19:12:35 2020
* 
x_PM_SKY130_FD_SC_HDLL__NAND2_16%B N_B_c_165_n N_B_M1004_g N_B_c_183_n
+ N_B_M1000_g N_B_c_184_n N_B_M1002_g N_B_c_166_n N_B_M1005_g N_B_c_167_n
+ N_B_M1014_g N_B_c_185_n N_B_M1007_g N_B_c_186_n N_B_M1009_g N_B_c_168_n
+ N_B_M1016_g N_B_c_169_n N_B_M1020_g N_B_c_187_n N_B_M1010_g N_B_c_188_n
+ N_B_M1015_g N_B_c_170_n N_B_M1025_g N_B_c_171_n N_B_M1034_g N_B_c_189_n
+ N_B_M1019_g N_B_c_190_n N_B_M1028_g N_B_c_172_n N_B_M1035_g N_B_c_173_n
+ N_B_M1039_g N_B_c_191_n N_B_M1033_g N_B_c_192_n N_B_M1037_g N_B_c_174_n
+ N_B_M1040_g N_B_c_175_n N_B_M1046_g N_B_c_193_n N_B_M1042_g N_B_c_194_n
+ N_B_M1045_g N_B_c_176_n N_B_M1053_g N_B_c_177_n N_B_M1055_g N_B_c_195_n
+ N_B_M1050_g N_B_c_196_n N_B_M1051_g N_B_c_178_n N_B_M1056_g N_B_c_179_n
+ N_B_M1057_g N_B_c_197_n N_B_M1054_g N_B_c_198_n N_B_M1060_g N_B_c_180_n
+ N_B_M1058_g B N_B_c_181_n N_B_c_182_n PM_SKY130_FD_SC_HDLL__NAND2_16%B
x_PM_SKY130_FD_SC_HDLL__NAND2_16%A N_A_c_493_n N_A_M1001_g N_A_c_510_n
+ N_A_M1003_g N_A_c_494_n N_A_M1006_g N_A_c_511_n N_A_M1008_g N_A_c_495_n
+ N_A_M1011_g N_A_c_512_n N_A_M1012_g N_A_c_513_n N_A_M1013_g N_A_c_496_n
+ N_A_M1017_g N_A_c_497_n N_A_M1018_g N_A_c_514_n N_A_M1021_g N_A_c_515_n
+ N_A_M1022_g N_A_c_498_n N_A_M1024_g N_A_c_499_n N_A_M1026_g N_A_c_516_n
+ N_A_M1023_g N_A_c_500_n N_A_M1027_g N_A_c_517_n N_A_M1029_g N_A_c_501_n
+ N_A_M1030_g N_A_c_518_n N_A_M1031_g N_A_c_519_n N_A_M1038_g N_A_c_502_n
+ N_A_M1032_g N_A_c_503_n N_A_M1036_g N_A_c_520_n N_A_M1041_g N_A_c_521_n
+ N_A_M1048_g N_A_c_504_n N_A_M1043_g N_A_c_505_n N_A_M1044_g N_A_c_522_n
+ N_A_M1049_g N_A_c_523_n N_A_M1052_g N_A_c_506_n N_A_M1047_g N_A_c_507_n
+ N_A_M1059_g N_A_c_524_n N_A_M1061_g N_A_c_525_n N_A_M1063_g N_A_c_508_n
+ N_A_M1062_g A N_A_c_598_p N_A_c_509_n PM_SKY130_FD_SC_HDLL__NAND2_16%A
x_PM_SKY130_FD_SC_HDLL__NAND2_16%VPWR N_VPWR_M1000_d N_VPWR_M1002_d
+ N_VPWR_M1009_d N_VPWR_M1015_d N_VPWR_M1028_d N_VPWR_M1037_d N_VPWR_M1045_d
+ N_VPWR_M1051_d N_VPWR_M1060_d N_VPWR_M1008_d N_VPWR_M1013_d N_VPWR_M1022_d
+ N_VPWR_M1029_d N_VPWR_M1038_d N_VPWR_M1048_d N_VPWR_M1052_d N_VPWR_M1063_d
+ N_VPWR_c_749_n N_VPWR_c_750_n N_VPWR_c_751_n N_VPWR_c_752_n N_VPWR_c_753_n
+ N_VPWR_c_754_n N_VPWR_c_755_n N_VPWR_c_756_n N_VPWR_c_757_n N_VPWR_c_758_n
+ N_VPWR_c_759_n N_VPWR_c_760_n N_VPWR_c_761_n N_VPWR_c_762_n N_VPWR_c_763_n
+ N_VPWR_c_764_n N_VPWR_c_765_n N_VPWR_c_766_n N_VPWR_c_767_n N_VPWR_c_768_n
+ N_VPWR_c_769_n N_VPWR_c_770_n N_VPWR_c_771_n N_VPWR_c_772_n N_VPWR_c_773_n
+ N_VPWR_c_774_n N_VPWR_c_775_n N_VPWR_c_776_n N_VPWR_c_777_n N_VPWR_c_778_n
+ N_VPWR_c_779_n N_VPWR_c_780_n N_VPWR_c_781_n N_VPWR_c_782_n N_VPWR_c_783_n
+ N_VPWR_c_784_n N_VPWR_c_785_n N_VPWR_c_786_n N_VPWR_c_787_n N_VPWR_c_788_n
+ N_VPWR_c_789_n N_VPWR_c_790_n N_VPWR_c_791_n VPWR N_VPWR_c_792_n
+ N_VPWR_c_793_n N_VPWR_c_794_n N_VPWR_c_795_n N_VPWR_c_796_n N_VPWR_c_797_n
+ N_VPWR_c_798_n N_VPWR_c_748_n PM_SKY130_FD_SC_HDLL__NAND2_16%VPWR
x_PM_SKY130_FD_SC_HDLL__NAND2_16%Y N_Y_M1001_d N_Y_M1011_d N_Y_M1018_d
+ N_Y_M1026_d N_Y_M1030_d N_Y_M1036_d N_Y_M1044_d N_Y_M1059_d N_Y_M1000_s
+ N_Y_M1007_s N_Y_M1010_s N_Y_M1019_s N_Y_M1033_s N_Y_M1042_s N_Y_M1050_s
+ N_Y_M1054_s N_Y_M1003_s N_Y_M1012_s N_Y_M1021_s N_Y_M1023_s N_Y_M1031_s
+ N_Y_M1041_s N_Y_M1049_s N_Y_M1061_s N_Y_c_980_n N_Y_c_984_n N_Y_c_987_n
+ N_Y_c_991_n N_Y_c_995_n N_Y_c_999_n N_Y_c_1003_n N_Y_c_1007_n N_Y_c_1011_n
+ N_Y_c_1015_n N_Y_c_1019_n N_Y_c_1023_n N_Y_c_1027_n N_Y_c_1031_n N_Y_c_1035_n
+ N_Y_c_1039_n N_Y_c_1042_n N_Y_c_1078_n N_Y_c_1044_n N_Y_c_1082_n N_Y_c_1098_n
+ N_Y_c_1102_n N_Y_c_1106_n N_Y_c_1110_n N_Y_c_1114_n N_Y_c_1118_n N_Y_c_1122_n
+ N_Y_c_1126_n N_Y_c_1130_n N_Y_c_1134_n N_Y_c_1138_n N_Y_c_1142_n N_Y_c_1146_n
+ N_Y_c_1150_n N_Y_c_1294_p N_Y_c_978_n N_Y_c_1045_n N_Y_c_1049_n N_Y_c_1053_n
+ N_Y_c_1057_n N_Y_c_1061_n N_Y_c_1065_n N_Y_c_1069_n N_Y_c_1156_n N_Y_c_1159_n
+ N_Y_c_1163_n N_Y_c_1167_n N_Y_c_1171_n N_Y_c_1175_n N_Y_c_1179_n N_Y_c_1183_n
+ N_Y_c_976_n N_Y_c_1188_n Y N_Y_c_977_n Y PM_SKY130_FD_SC_HDLL__NAND2_16%Y
x_PM_SKY130_FD_SC_HDLL__NAND2_16%A_27_47# N_A_27_47#_M1004_d N_A_27_47#_M1005_d
+ N_A_27_47#_M1016_d N_A_27_47#_M1025_d N_A_27_47#_M1035_d N_A_27_47#_M1040_d
+ N_A_27_47#_M1053_d N_A_27_47#_M1056_d N_A_27_47#_M1058_d N_A_27_47#_M1006_s
+ N_A_27_47#_M1017_s N_A_27_47#_M1024_s N_A_27_47#_M1027_s N_A_27_47#_M1032_s
+ N_A_27_47#_M1043_s N_A_27_47#_M1047_s N_A_27_47#_M1062_s N_A_27_47#_c_1305_n
+ N_A_27_47#_c_1319_n N_A_27_47#_c_1306_n N_A_27_47#_c_1325_n
+ N_A_27_47#_c_1329_n N_A_27_47#_c_1333_n N_A_27_47#_c_1337_n
+ N_A_27_47#_c_1341_n N_A_27_47#_c_1345_n N_A_27_47#_c_1349_n
+ N_A_27_47#_c_1353_n N_A_27_47#_c_1357_n N_A_27_47#_c_1361_n
+ N_A_27_47#_c_1365_n N_A_27_47#_c_1369_n N_A_27_47#_c_1373_n
+ N_A_27_47#_c_1377_n N_A_27_47#_c_1381_n N_A_27_47#_c_1307_n
+ N_A_27_47#_c_1412_n N_A_27_47#_c_1308_n N_A_27_47#_c_1309_n
+ N_A_27_47#_c_1310_n N_A_27_47#_c_1311_n N_A_27_47#_c_1312_n
+ N_A_27_47#_c_1313_n N_A_27_47#_c_1314_n N_A_27_47#_c_1315_n
+ N_A_27_47#_c_1316_n PM_SKY130_FD_SC_HDLL__NAND2_16%A_27_47#
x_PM_SKY130_FD_SC_HDLL__NAND2_16%VGND N_VGND_M1004_s N_VGND_M1014_s
+ N_VGND_M1020_s N_VGND_M1034_s N_VGND_M1039_s N_VGND_M1046_s N_VGND_M1055_s
+ N_VGND_M1057_s N_VGND_c_1532_n N_VGND_c_1533_n N_VGND_c_1534_n N_VGND_c_1535_n
+ N_VGND_c_1536_n N_VGND_c_1537_n N_VGND_c_1538_n N_VGND_c_1539_n
+ N_VGND_c_1540_n N_VGND_c_1541_n N_VGND_c_1542_n N_VGND_c_1543_n
+ N_VGND_c_1544_n N_VGND_c_1545_n N_VGND_c_1546_n N_VGND_c_1547_n
+ N_VGND_c_1548_n N_VGND_c_1549_n VGND N_VGND_c_1550_n N_VGND_c_1551_n
+ N_VGND_c_1552_n N_VGND_c_1553_n N_VGND_c_1554_n N_VGND_c_1555_n
+ N_VGND_c_1556_n N_VGND_c_1557_n PM_SKY130_FD_SC_HDLL__NAND2_16%VGND
cc_1 VNB N_B_c_165_n 0.0228251f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_2 VNB N_B_c_166_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=0.995
cc_3 VNB N_B_c_167_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_4 VNB N_B_c_168_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_5 VNB N_B_c_169_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_6 VNB N_B_c_170_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_7 VNB N_B_c_171_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.995
cc_8 VNB N_B_c_172_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.995
cc_9 VNB N_B_c_173_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.995
cc_10 VNB N_B_c_174_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.995
cc_11 VNB N_B_c_175_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.995
cc_12 VNB N_B_c_176_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_13 VNB N_B_c_177_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=0.995
cc_14 VNB N_B_c_178_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=6.63 $Y2=0.995
cc_15 VNB N_B_c_179_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=7.05 $Y2=0.995
cc_16 VNB N_B_c_180_n 0.0171127f $X=-0.19 $Y=-0.24 $X2=7.57 $Y2=0.995
cc_17 VNB N_B_c_181_n 0.0101411f $X=-0.19 $Y=-0.24 $X2=7.36 $Y2=1.16
cc_18 VNB N_B_c_182_n 0.305486f $X=-0.19 $Y=-0.24 $X2=7.545 $Y2=1.202
cc_19 VNB N_A_c_493_n 0.0162568f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=0.995
cc_20 VNB N_A_c_494_n 0.0168735f $X=-0.19 $Y=-0.24 $X2=0.965 $Y2=1.41
cc_21 VNB N_A_c_495_n 0.0173555f $X=-0.19 $Y=-0.24 $X2=1.41 $Y2=0.995
cc_22 VNB N_A_c_496_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=1.93 $Y2=0.995
cc_23 VNB N_A_c_497_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.995
cc_24 VNB N_A_c_498_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.995
cc_25 VNB N_A_c_499_n 0.0164369f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.995
cc_26 VNB N_A_c_500_n 0.0169186f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.41
cc_27 VNB N_A_c_501_n 0.0173608f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.995
cc_28 VNB N_A_c_502_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.995
cc_29 VNB N_A_c_503_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.995
cc_30 VNB N_A_c_504_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_31 VNB N_A_c_505_n 0.0168791f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=0.995
cc_32 VNB N_A_c_506_n 0.0168753f $X=-0.19 $Y=-0.24 $X2=6.63 $Y2=0.995
cc_33 VNB N_A_c_507_n 0.0168204f $X=-0.19 $Y=-0.24 $X2=7.05 $Y2=0.995
cc_34 VNB N_A_c_508_n 0.0228463f $X=-0.19 $Y=-0.24 $X2=7.57 $Y2=0.995
cc_35 VNB N_A_c_509_n 0.313864f $X=-0.19 $Y=-0.24 $X2=7.545 $Y2=1.202
cc_36 VNB N_VPWR_c_748_n 0.649277f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_37 VNB N_Y_c_976_n 0.00209731f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_38 VNB N_Y_c_977_n 0.00106016f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_39 VNB N_A_27_47#_c_1305_n 0.018052f $X=-0.19 $Y=-0.24 $X2=4.255 $Y2=1.985
cc_40 VNB N_A_27_47#_c_1306_n 0.011879f $X=-0.19 $Y=-0.24 $X2=4.725 $Y2=1.985
cc_41 VNB N_A_27_47#_c_1307_n 0.00257277f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.202
cc_42 VNB N_A_27_47#_c_1308_n 0.00914706f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=1.202
cc_43 VNB N_A_27_47#_c_1309_n 0.0204013f $X=-0.19 $Y=-0.24 $X2=4.725 $Y2=1.202
cc_44 VNB N_A_27_47#_c_1310_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=1.202
cc_45 VNB N_A_27_47#_c_1311_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=5.195 $Y2=1.202
cc_46 VNB N_A_27_47#_c_1312_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.202
cc_47 VNB N_A_27_47#_c_1313_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=1.202
cc_48 VNB N_A_27_47#_c_1314_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=1.202
cc_49 VNB N_A_27_47#_c_1315_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=6.135 $Y2=1.202
cc_50 VNB N_A_27_47#_c_1316_n 0.00115812f $X=-0.19 $Y=-0.24 $X2=6.605 $Y2=1.202
cc_51 VNB N_VGND_c_1532_n 0.00466649f $X=-0.19 $Y=-0.24 $X2=2.35 $Y2=0.56
cc_52 VNB N_VGND_c_1533_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.985
cc_53 VNB N_VGND_c_1534_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=2.845 $Y2=1.985
cc_54 VNB N_VGND_c_1535_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=0.56
cc_55 VNB N_VGND_c_1536_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=3.29 $Y2=0.56
cc_56 VNB N_VGND_c_1537_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.315 $Y2=1.985
cc_57 VNB N_VGND_c_1538_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=3.785 $Y2=1.985
cc_58 VNB N_VGND_c_1539_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=3.81 $Y2=0.56
cc_59 VNB N_VGND_c_1540_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=4.23 $Y2=0.56
cc_60 VNB N_VGND_c_1541_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=4.725 $Y2=1.41
cc_61 VNB N_VGND_c_1542_n 0.00414011f $X=-0.19 $Y=-0.24 $X2=4.75 $Y2=0.56
cc_62 VNB N_VGND_c_1543_n 0.00466098f $X=-0.19 $Y=-0.24 $X2=5.17 $Y2=0.56
cc_63 VNB N_VGND_c_1544_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=5.195 $Y2=1.985
cc_64 VNB N_VGND_c_1545_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.41
cc_65 VNB N_VGND_c_1546_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=5.665 $Y2=1.985
cc_66 VNB N_VGND_c_1547_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.995
cc_67 VNB N_VGND_c_1548_n 0.0166431f $X=-0.19 $Y=-0.24 $X2=5.69 $Y2=0.56
cc_68 VNB N_VGND_c_1549_n 0.00515836f $X=-0.19 $Y=-0.24 $X2=6.11 $Y2=0.995
cc_69 VNB N_VGND_c_1550_n 0.0172128f $X=-0.19 $Y=-0.24 $X2=6.135 $Y2=1.41
cc_70 VNB N_VGND_c_1551_n 0.186236f $X=-0.19 $Y=-0.24 $X2=7.57 $Y2=0.56
cc_71 VNB N_VGND_c_1552_n 0.698664f $X=-0.19 $Y=-0.24 $X2=7.57 $Y2=0.56
cc_72 VNB N_VGND_c_1553_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.47 $Y2=1.202
cc_73 VNB N_VGND_c_1554_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.56 $Y2=1.16
cc_74 VNB N_VGND_c_1555_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=0.99 $Y2=1.202
cc_75 VNB N_VGND_c_1556_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=1.905 $Y2=1.202
cc_76 VNB N_VGND_c_1557_n 0.00515873f $X=-0.19 $Y=-0.24 $X2=2.375 $Y2=1.202
cc_77 VPB N_B_c_183_n 0.0210879f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_78 VPB N_B_c_184_n 0.0162635f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.41
cc_79 VPB N_B_c_185_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_80 VPB N_B_c_186_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_81 VPB N_B_c_187_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_82 VPB N_B_c_188_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_83 VPB N_B_c_189_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_84 VPB N_B_c_190_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.41
cc_85 VPB N_B_c_191_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_86 VPB N_B_c_192_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.41
cc_87 VPB N_B_c_193_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.41
cc_88 VPB N_B_c_194_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.41
cc_89 VPB N_B_c_195_n 0.0162635f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.41
cc_90 VPB N_B_c_196_n 0.0162635f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.41
cc_91 VPB N_B_c_197_n 0.0162635f $X=-0.19 $Y=1.305 $X2=7.075 $Y2=1.41
cc_92 VPB N_B_c_198_n 0.0164324f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.41
cc_93 VPB N_B_c_181_n 7.73822e-19 $X=-0.19 $Y=1.305 $X2=7.36 $Y2=1.16
cc_94 VPB N_B_c_182_n 0.204034f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.202
cc_95 VPB N_A_c_510_n 0.0160834f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.41
cc_96 VPB N_A_c_511_n 0.0162386f $X=-0.19 $Y=1.305 $X2=0.99 $Y2=0.995
cc_97 VPB N_A_c_512_n 0.016261f $X=-0.19 $Y=1.305 $X2=1.435 $Y2=1.41
cc_98 VPB N_A_c_513_n 0.0162635f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.41
cc_99 VPB N_A_c_514_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.375 $Y2=1.41
cc_100 VPB N_A_c_515_n 0.0162635f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.41
cc_101 VPB N_A_c_516_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.315 $Y2=1.41
cc_102 VPB N_A_c_517_n 0.0162635f $X=-0.19 $Y=1.305 $X2=3.81 $Y2=0.995
cc_103 VPB N_A_c_518_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_104 VPB N_A_c_519_n 0.0162635f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.41
cc_105 VPB N_A_c_520_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.41
cc_106 VPB N_A_c_521_n 0.0162635f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.41
cc_107 VPB N_A_c_522_n 0.0162635f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.41
cc_108 VPB N_A_c_523_n 0.0162606f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.41
cc_109 VPB N_A_c_524_n 0.016238f $X=-0.19 $Y=1.305 $X2=7.075 $Y2=1.41
cc_110 VPB N_A_c_525_n 0.0207627f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.41
cc_111 VPB N_A_c_509_n 0.205595f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.202
cc_112 VPB N_VPWR_c_749_n 0.0113525f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.41
cc_113 VPB N_VPWR_c_750_n 0.0410822f $X=-0.19 $Y=1.305 $X2=4.255 $Y2=1.985
cc_114 VPB N_VPWR_c_751_n 0.0041373f $X=-0.19 $Y=1.305 $X2=4.75 $Y2=0.56
cc_115 VPB N_VPWR_c_752_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.17 $Y2=0.56
cc_116 VPB N_VPWR_c_753_n 0.0041373f $X=-0.19 $Y=1.305 $X2=5.195 $Y2=1.985
cc_117 VPB N_VPWR_c_754_n 0.017949f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.985
cc_118 VPB N_VPWR_c_755_n 0.0041373f $X=-0.19 $Y=1.305 $X2=5.69 $Y2=0.56
cc_119 VPB N_VPWR_c_756_n 0.017949f $X=-0.19 $Y=1.305 $X2=6.11 $Y2=0.56
cc_120 VPB N_VPWR_c_757_n 0.0041373f $X=-0.19 $Y=1.305 $X2=6.135 $Y2=1.985
cc_121 VPB N_VPWR_c_758_n 0.017949f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.985
cc_122 VPB N_VPWR_c_759_n 0.0041373f $X=-0.19 $Y=1.305 $X2=6.63 $Y2=0.56
cc_123 VPB N_VPWR_c_760_n 0.0041373f $X=-0.19 $Y=1.305 $X2=7.075 $Y2=1.41
cc_124 VPB N_VPWR_c_761_n 0.0041373f $X=-0.19 $Y=1.305 $X2=7.545 $Y2=1.985
cc_125 VPB N_VPWR_c_762_n 0.0041373f $X=-0.19 $Y=1.305 $X2=7.57 $Y2=0.56
cc_126 VPB N_VPWR_c_763_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.495 $Y2=1.202
cc_127 VPB N_VPWR_c_764_n 0.0041373f $X=-0.19 $Y=1.305 $X2=0.965 $Y2=1.202
cc_128 VPB N_VPWR_c_765_n 0.0041373f $X=-0.19 $Y=1.305 $X2=1.905 $Y2=1.202
cc_129 VPB N_VPWR_c_766_n 0.0041373f $X=-0.19 $Y=1.305 $X2=2.845 $Y2=1.202
cc_130 VPB N_VPWR_c_767_n 0.0041373f $X=-0.19 $Y=1.305 $X2=3.785 $Y2=1.202
cc_131 VPB N_VPWR_c_768_n 0.0041373f $X=-0.19 $Y=1.305 $X2=4.725 $Y2=1.202
cc_132 VPB N_VPWR_c_769_n 0.0041373f $X=-0.19 $Y=1.305 $X2=5.665 $Y2=1.202
cc_133 VPB N_VPWR_c_770_n 0.0139043f $X=-0.19 $Y=1.305 $X2=6.11 $Y2=1.202
cc_134 VPB N_VPWR_c_771_n 0.0410822f $X=-0.19 $Y=1.305 $X2=6.605 $Y2=1.202
cc_135 VPB N_VPWR_c_772_n 0.017949f $X=-0.19 $Y=1.305 $X2=7.36 $Y2=1.16
cc_136 VPB N_VPWR_c_773_n 0.00516083f $X=-0.19 $Y=1.305 $X2=7.36 $Y2=1.16
cc_137 VPB N_VPWR_c_774_n 0.017949f $X=-0.19 $Y=1.305 $X2=7.57 $Y2=1.202
cc_138 VPB N_VPWR_c_775_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0.56 $Y2=1.19
cc_139 VPB N_VPWR_c_776_n 0.017949f $X=-0.19 $Y=1.305 $X2=3.91 $Y2=1.19
cc_140 VPB N_VPWR_c_777_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_141 VPB N_VPWR_c_778_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_142 VPB N_VPWR_c_779_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_143 VPB N_VPWR_c_780_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_144 VPB N_VPWR_c_781_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_145 VPB N_VPWR_c_782_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_146 VPB N_VPWR_c_783_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_147 VPB N_VPWR_c_784_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_148 VPB N_VPWR_c_785_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_149 VPB N_VPWR_c_786_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_150 VPB N_VPWR_c_787_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_151 VPB N_VPWR_c_788_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_152 VPB N_VPWR_c_789_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_153 VPB N_VPWR_c_790_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_154 VPB N_VPWR_c_791_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_155 VPB N_VPWR_c_792_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_156 VPB N_VPWR_c_793_n 0.017949f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_157 VPB N_VPWR_c_794_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_158 VPB N_VPWR_c_795_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_159 VPB N_VPWR_c_796_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_160 VPB N_VPWR_c_797_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_161 VPB N_VPWR_c_798_n 0.00516083f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_162 VPB N_VPWR_c_748_n 0.050553f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_163 VPB N_Y_c_978_n 0.0015125f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_164 VPB Y 0.00161879f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_165 N_B_c_180_n N_A_c_493_n 0.0168484f $X=7.57 $Y=0.995 $X2=-0.19 $Y2=-0.24
cc_166 N_B_c_198_n N_A_c_510_n 0.0230419f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_167 N_B_c_181_n N_A_c_509_n 9.92551e-19 $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_168 N_B_c_182_n N_A_c_509_n 0.0168484f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_169 N_B_c_183_n N_VPWR_c_750_n 0.00354866f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_170 N_B_c_184_n N_VPWR_c_751_n 0.00173895f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_171 N_B_c_185_n N_VPWR_c_751_n 0.00173895f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_172 N_B_c_185_n N_VPWR_c_752_n 0.00673617f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_173 N_B_c_186_n N_VPWR_c_752_n 0.00673617f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_174 N_B_c_186_n N_VPWR_c_753_n 0.00173895f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_175 N_B_c_187_n N_VPWR_c_753_n 0.00173895f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_176 N_B_c_187_n N_VPWR_c_754_n 0.00673617f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_177 N_B_c_188_n N_VPWR_c_754_n 0.00673617f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_178 N_B_c_188_n N_VPWR_c_755_n 0.00173895f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_179 N_B_c_189_n N_VPWR_c_755_n 0.00173895f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_180 N_B_c_189_n N_VPWR_c_756_n 0.00673617f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_181 N_B_c_190_n N_VPWR_c_756_n 0.00673617f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_182 N_B_c_190_n N_VPWR_c_757_n 0.00173895f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_183 N_B_c_191_n N_VPWR_c_757_n 0.00173895f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_184 N_B_c_191_n N_VPWR_c_758_n 0.00673617f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_185 N_B_c_192_n N_VPWR_c_758_n 0.00673617f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_186 N_B_c_192_n N_VPWR_c_759_n 0.00173895f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_187 N_B_c_193_n N_VPWR_c_759_n 0.00173895f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_188 N_B_c_194_n N_VPWR_c_760_n 0.00173895f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_189 N_B_c_195_n N_VPWR_c_760_n 0.00173895f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_190 N_B_c_196_n N_VPWR_c_761_n 0.00173895f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_191 N_B_c_197_n N_VPWR_c_761_n 0.00173895f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_192 N_B_c_198_n N_VPWR_c_762_n 0.00173895f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_193 N_B_c_193_n N_VPWR_c_772_n 0.00673617f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_194 N_B_c_194_n N_VPWR_c_772_n 0.00673617f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_195 N_B_c_195_n N_VPWR_c_774_n 0.00673617f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_196 N_B_c_196_n N_VPWR_c_774_n 0.00673617f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_197 N_B_c_197_n N_VPWR_c_776_n 0.00673617f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_198 N_B_c_198_n N_VPWR_c_776_n 0.00673617f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_199 N_B_c_183_n N_VPWR_c_792_n 0.00673617f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_200 N_B_c_184_n N_VPWR_c_792_n 0.00673617f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_201 N_B_c_183_n N_VPWR_c_748_n 0.0126298f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_202 N_B_c_184_n N_VPWR_c_748_n 0.0117184f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_203 N_B_c_185_n N_VPWR_c_748_n 0.0117184f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_204 N_B_c_186_n N_VPWR_c_748_n 0.0117184f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_205 N_B_c_187_n N_VPWR_c_748_n 0.0117184f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_206 N_B_c_188_n N_VPWR_c_748_n 0.0117184f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_207 N_B_c_189_n N_VPWR_c_748_n 0.0117184f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_208 N_B_c_190_n N_VPWR_c_748_n 0.0117184f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_209 N_B_c_191_n N_VPWR_c_748_n 0.0117184f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_210 N_B_c_192_n N_VPWR_c_748_n 0.0117184f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_211 N_B_c_193_n N_VPWR_c_748_n 0.0117184f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_212 N_B_c_194_n N_VPWR_c_748_n 0.0117184f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_213 N_B_c_195_n N_VPWR_c_748_n 0.0117184f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_214 N_B_c_196_n N_VPWR_c_748_n 0.0117184f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_215 N_B_c_197_n N_VPWR_c_748_n 0.0117184f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_216 N_B_c_198_n N_VPWR_c_748_n 0.0117436f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_217 N_B_c_183_n N_Y_c_980_n 0.00215964f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_218 N_B_c_184_n N_Y_c_980_n 5.79575e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_219 N_B_c_181_n N_Y_c_980_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_220 N_B_c_182_n N_Y_c_980_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_221 N_B_c_183_n N_Y_c_984_n 0.00897418f $X=0.495 $Y=1.41 $X2=0 $Y2=0
cc_222 N_B_c_184_n N_Y_c_984_n 0.0100233f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_223 N_B_c_185_n N_Y_c_984_n 5.91934e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_224 N_B_c_184_n N_Y_c_987_n 0.0137916f $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_225 N_B_c_185_n N_Y_c_987_n 0.0137916f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_226 N_B_c_181_n N_Y_c_987_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_227 N_B_c_182_n N_Y_c_987_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_228 N_B_c_184_n N_Y_c_991_n 5.91934e-19 $X=0.965 $Y=1.41 $X2=0 $Y2=0
cc_229 N_B_c_185_n N_Y_c_991_n 0.0100233f $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_230 N_B_c_186_n N_Y_c_991_n 0.0100233f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_231 N_B_c_187_n N_Y_c_991_n 5.91934e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_232 N_B_c_186_n N_Y_c_995_n 0.0137916f $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_233 N_B_c_187_n N_Y_c_995_n 0.0137916f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_234 N_B_c_181_n N_Y_c_995_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_235 N_B_c_182_n N_Y_c_995_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_236 N_B_c_186_n N_Y_c_999_n 5.91934e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_237 N_B_c_187_n N_Y_c_999_n 0.0100233f $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_238 N_B_c_188_n N_Y_c_999_n 0.0100233f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_239 N_B_c_189_n N_Y_c_999_n 5.91934e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_240 N_B_c_188_n N_Y_c_1003_n 0.0137916f $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_241 N_B_c_189_n N_Y_c_1003_n 0.0137916f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_242 N_B_c_181_n N_Y_c_1003_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_243 N_B_c_182_n N_Y_c_1003_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_244 N_B_c_188_n N_Y_c_1007_n 5.91934e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_245 N_B_c_189_n N_Y_c_1007_n 0.0100233f $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_246 N_B_c_190_n N_Y_c_1007_n 0.0100233f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_247 N_B_c_191_n N_Y_c_1007_n 5.91934e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_248 N_B_c_190_n N_Y_c_1011_n 0.0137916f $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_249 N_B_c_191_n N_Y_c_1011_n 0.0137916f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_250 N_B_c_181_n N_Y_c_1011_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_251 N_B_c_182_n N_Y_c_1011_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_252 N_B_c_190_n N_Y_c_1015_n 5.91934e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_253 N_B_c_191_n N_Y_c_1015_n 0.0100233f $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_254 N_B_c_192_n N_Y_c_1015_n 0.0100233f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_255 N_B_c_193_n N_Y_c_1015_n 5.91934e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_256 N_B_c_192_n N_Y_c_1019_n 0.0137916f $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_257 N_B_c_193_n N_Y_c_1019_n 0.0137916f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_258 N_B_c_181_n N_Y_c_1019_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_259 N_B_c_182_n N_Y_c_1019_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_260 N_B_c_192_n N_Y_c_1023_n 5.91934e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_261 N_B_c_193_n N_Y_c_1023_n 0.0100233f $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_262 N_B_c_194_n N_Y_c_1023_n 0.0100233f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_263 N_B_c_195_n N_Y_c_1023_n 5.91934e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_264 N_B_c_194_n N_Y_c_1027_n 0.0137916f $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_265 N_B_c_195_n N_Y_c_1027_n 0.0137916f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_266 N_B_c_181_n N_Y_c_1027_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_267 N_B_c_182_n N_Y_c_1027_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_268 N_B_c_194_n N_Y_c_1031_n 5.91934e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_269 N_B_c_195_n N_Y_c_1031_n 0.0100233f $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_270 N_B_c_196_n N_Y_c_1031_n 0.0100233f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_271 N_B_c_197_n N_Y_c_1031_n 5.91934e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_272 N_B_c_196_n N_Y_c_1035_n 0.0137916f $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_273 N_B_c_197_n N_Y_c_1035_n 0.0137916f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_274 N_B_c_181_n N_Y_c_1035_n 0.0393642f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_275 N_B_c_182_n N_Y_c_1035_n 0.00655651f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_276 N_B_c_196_n N_Y_c_1039_n 5.91934e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_277 N_B_c_197_n N_Y_c_1039_n 0.0100233f $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_278 N_B_c_198_n N_Y_c_1039_n 0.0100233f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_279 N_B_c_198_n N_Y_c_1042_n 0.0152705f $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_280 N_B_c_181_n N_Y_c_1042_n 0.00347994f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_281 N_B_c_198_n N_Y_c_1044_n 5.91934e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_282 N_B_c_185_n N_Y_c_1045_n 5.79575e-19 $X=1.435 $Y=1.41 $X2=0 $Y2=0
cc_283 N_B_c_186_n N_Y_c_1045_n 5.79575e-19 $X=1.905 $Y=1.41 $X2=0 $Y2=0
cc_284 N_B_c_181_n N_Y_c_1045_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_285 N_B_c_182_n N_Y_c_1045_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_286 N_B_c_187_n N_Y_c_1049_n 5.79575e-19 $X=2.375 $Y=1.41 $X2=0 $Y2=0
cc_287 N_B_c_188_n N_Y_c_1049_n 5.79575e-19 $X=2.845 $Y=1.41 $X2=0 $Y2=0
cc_288 N_B_c_181_n N_Y_c_1049_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_289 N_B_c_182_n N_Y_c_1049_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_290 N_B_c_189_n N_Y_c_1053_n 5.79575e-19 $X=3.315 $Y=1.41 $X2=0 $Y2=0
cc_291 N_B_c_190_n N_Y_c_1053_n 5.79575e-19 $X=3.785 $Y=1.41 $X2=0 $Y2=0
cc_292 N_B_c_181_n N_Y_c_1053_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_293 N_B_c_182_n N_Y_c_1053_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_294 N_B_c_191_n N_Y_c_1057_n 5.79575e-19 $X=4.255 $Y=1.41 $X2=0 $Y2=0
cc_295 N_B_c_192_n N_Y_c_1057_n 5.79575e-19 $X=4.725 $Y=1.41 $X2=0 $Y2=0
cc_296 N_B_c_181_n N_Y_c_1057_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_297 N_B_c_182_n N_Y_c_1057_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_298 N_B_c_193_n N_Y_c_1061_n 5.79575e-19 $X=5.195 $Y=1.41 $X2=0 $Y2=0
cc_299 N_B_c_194_n N_Y_c_1061_n 5.79575e-19 $X=5.665 $Y=1.41 $X2=0 $Y2=0
cc_300 N_B_c_181_n N_Y_c_1061_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_301 N_B_c_182_n N_Y_c_1061_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_302 N_B_c_195_n N_Y_c_1065_n 5.79575e-19 $X=6.135 $Y=1.41 $X2=0 $Y2=0
cc_303 N_B_c_196_n N_Y_c_1065_n 5.79575e-19 $X=6.605 $Y=1.41 $X2=0 $Y2=0
cc_304 N_B_c_181_n N_Y_c_1065_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_305 N_B_c_182_n N_Y_c_1065_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_306 N_B_c_197_n N_Y_c_1069_n 5.79575e-19 $X=7.075 $Y=1.41 $X2=0 $Y2=0
cc_307 N_B_c_198_n N_Y_c_1069_n 5.79575e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_308 N_B_c_181_n N_Y_c_1069_n 0.0215641f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_309 N_B_c_182_n N_Y_c_1069_n 0.00631893f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_310 N_B_c_198_n Y 5.27102e-19 $X=7.545 $Y=1.41 $X2=0 $Y2=0
cc_311 N_B_c_181_n Y 0.0108577f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_312 N_B_c_182_n Y 0.00179199f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_313 N_B_c_180_n N_Y_c_977_n 8.84206e-19 $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_314 N_B_c_165_n N_A_27_47#_c_1305_n 0.00661134f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_315 N_B_c_166_n N_A_27_47#_c_1305_n 5.22365e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_316 N_B_c_165_n N_A_27_47#_c_1319_n 0.00899636f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_317 N_B_c_166_n N_A_27_47#_c_1319_n 0.00899636f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_318 N_B_c_181_n N_A_27_47#_c_1319_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_319 N_B_c_182_n N_A_27_47#_c_1319_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_320 N_B_c_165_n N_A_27_47#_c_1306_n 8.68782e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_321 N_B_c_181_n N_A_27_47#_c_1306_n 0.00230475f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_322 N_B_c_165_n N_A_27_47#_c_1325_n 5.22365e-19 $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_323 N_B_c_166_n N_A_27_47#_c_1325_n 0.00661134f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_324 N_B_c_167_n N_A_27_47#_c_1325_n 0.00661134f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_325 N_B_c_168_n N_A_27_47#_c_1325_n 5.22365e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_326 N_B_c_167_n N_A_27_47#_c_1329_n 0.00899636f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_327 N_B_c_168_n N_A_27_47#_c_1329_n 0.00899636f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_328 N_B_c_181_n N_A_27_47#_c_1329_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_329 N_B_c_182_n N_A_27_47#_c_1329_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_330 N_B_c_167_n N_A_27_47#_c_1333_n 5.22365e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_331 N_B_c_168_n N_A_27_47#_c_1333_n 0.00661134f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_332 N_B_c_169_n N_A_27_47#_c_1333_n 0.00661134f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_333 N_B_c_170_n N_A_27_47#_c_1333_n 5.22365e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_334 N_B_c_169_n N_A_27_47#_c_1337_n 0.00899636f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_335 N_B_c_170_n N_A_27_47#_c_1337_n 0.00899636f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_336 N_B_c_181_n N_A_27_47#_c_1337_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_337 N_B_c_182_n N_A_27_47#_c_1337_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_338 N_B_c_169_n N_A_27_47#_c_1341_n 5.22365e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_339 N_B_c_170_n N_A_27_47#_c_1341_n 0.00661134f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_340 N_B_c_171_n N_A_27_47#_c_1341_n 0.00661134f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_341 N_B_c_172_n N_A_27_47#_c_1341_n 5.22365e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_342 N_B_c_171_n N_A_27_47#_c_1345_n 0.00899636f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_343 N_B_c_172_n N_A_27_47#_c_1345_n 0.00899636f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_344 N_B_c_181_n N_A_27_47#_c_1345_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_345 N_B_c_182_n N_A_27_47#_c_1345_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_346 N_B_c_171_n N_A_27_47#_c_1349_n 5.22365e-19 $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_347 N_B_c_172_n N_A_27_47#_c_1349_n 0.00661134f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_348 N_B_c_173_n N_A_27_47#_c_1349_n 0.00661134f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_349 N_B_c_174_n N_A_27_47#_c_1349_n 5.22365e-19 $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_350 N_B_c_173_n N_A_27_47#_c_1353_n 0.00899636f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_351 N_B_c_174_n N_A_27_47#_c_1353_n 0.00899636f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_352 N_B_c_181_n N_A_27_47#_c_1353_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_353 N_B_c_182_n N_A_27_47#_c_1353_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_354 N_B_c_173_n N_A_27_47#_c_1357_n 5.22365e-19 $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_355 N_B_c_174_n N_A_27_47#_c_1357_n 0.00661134f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_356 N_B_c_175_n N_A_27_47#_c_1357_n 0.00661134f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_357 N_B_c_176_n N_A_27_47#_c_1357_n 5.22365e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_358 N_B_c_175_n N_A_27_47#_c_1361_n 0.00899636f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_359 N_B_c_176_n N_A_27_47#_c_1361_n 0.00899636f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_360 N_B_c_181_n N_A_27_47#_c_1361_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_361 N_B_c_182_n N_A_27_47#_c_1361_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_362 N_B_c_175_n N_A_27_47#_c_1365_n 5.22365e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_363 N_B_c_176_n N_A_27_47#_c_1365_n 0.00661134f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_364 N_B_c_177_n N_A_27_47#_c_1365_n 0.00661134f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_365 N_B_c_178_n N_A_27_47#_c_1365_n 5.22365e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_366 N_B_c_177_n N_A_27_47#_c_1369_n 0.00899636f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_367 N_B_c_178_n N_A_27_47#_c_1369_n 0.00899636f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_368 N_B_c_181_n N_A_27_47#_c_1369_n 0.0395582f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_369 N_B_c_182_n N_A_27_47#_c_1369_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_370 N_B_c_177_n N_A_27_47#_c_1373_n 5.22365e-19 $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_371 N_B_c_178_n N_A_27_47#_c_1373_n 0.00661134f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_372 N_B_c_179_n N_A_27_47#_c_1373_n 0.00661134f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_373 N_B_c_180_n N_A_27_47#_c_1373_n 5.22365e-19 $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_374 N_B_c_179_n N_A_27_47#_c_1377_n 0.00899636f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_375 N_B_c_180_n N_A_27_47#_c_1377_n 0.0102281f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_376 N_B_c_181_n N_A_27_47#_c_1377_n 0.0332672f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_377 N_B_c_182_n N_A_27_47#_c_1377_n 0.00457246f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_378 N_B_c_180_n N_A_27_47#_c_1381_n 0.00248145f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_379 N_B_c_179_n N_A_27_47#_c_1307_n 4.7541e-19 $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_380 N_B_c_180_n N_A_27_47#_c_1307_n 0.00541116f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_381 N_B_c_166_n N_A_27_47#_c_1310_n 8.68782e-19 $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_382 N_B_c_167_n N_A_27_47#_c_1310_n 8.68782e-19 $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_383 N_B_c_181_n N_A_27_47#_c_1310_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_384 N_B_c_182_n N_A_27_47#_c_1310_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_385 N_B_c_168_n N_A_27_47#_c_1311_n 8.68782e-19 $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_386 N_B_c_169_n N_A_27_47#_c_1311_n 8.68782e-19 $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_387 N_B_c_181_n N_A_27_47#_c_1311_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_388 N_B_c_182_n N_A_27_47#_c_1311_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_389 N_B_c_170_n N_A_27_47#_c_1312_n 8.68782e-19 $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_390 N_B_c_171_n N_A_27_47#_c_1312_n 8.68782e-19 $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_391 N_B_c_181_n N_A_27_47#_c_1312_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_392 N_B_c_182_n N_A_27_47#_c_1312_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_393 N_B_c_172_n N_A_27_47#_c_1313_n 8.68782e-19 $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_394 N_B_c_173_n N_A_27_47#_c_1313_n 8.68782e-19 $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_395 N_B_c_181_n N_A_27_47#_c_1313_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_396 N_B_c_182_n N_A_27_47#_c_1313_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_397 N_B_c_174_n N_A_27_47#_c_1314_n 8.68782e-19 $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_398 N_B_c_175_n N_A_27_47#_c_1314_n 8.68782e-19 $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_399 N_B_c_181_n N_A_27_47#_c_1314_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_400 N_B_c_182_n N_A_27_47#_c_1314_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_401 N_B_c_176_n N_A_27_47#_c_1315_n 8.68782e-19 $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_402 N_B_c_177_n N_A_27_47#_c_1315_n 8.68782e-19 $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_403 N_B_c_181_n N_A_27_47#_c_1315_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_404 N_B_c_182_n N_A_27_47#_c_1315_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_405 N_B_c_178_n N_A_27_47#_c_1316_n 8.68782e-19 $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_406 N_B_c_179_n N_A_27_47#_c_1316_n 8.68782e-19 $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_407 N_B_c_181_n N_A_27_47#_c_1316_n 0.0214029f $X=7.36 $Y=1.16 $X2=0 $Y2=0
cc_408 N_B_c_182_n N_A_27_47#_c_1316_n 0.00224547f $X=7.545 $Y=1.202 $X2=0 $Y2=0
cc_409 N_B_c_165_n N_VGND_c_1532_n 0.00296353f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_410 N_B_c_166_n N_VGND_c_1532_n 0.00166854f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_411 N_B_c_166_n N_VGND_c_1533_n 0.00422241f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_412 N_B_c_167_n N_VGND_c_1533_n 0.00422241f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_413 N_B_c_167_n N_VGND_c_1534_n 0.00166854f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_414 N_B_c_168_n N_VGND_c_1534_n 0.00166854f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_415 N_B_c_168_n N_VGND_c_1535_n 0.00422241f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_416 N_B_c_169_n N_VGND_c_1535_n 0.00422241f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_417 N_B_c_169_n N_VGND_c_1536_n 0.00166854f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_418 N_B_c_170_n N_VGND_c_1536_n 0.00166854f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_419 N_B_c_170_n N_VGND_c_1537_n 0.00422241f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_420 N_B_c_171_n N_VGND_c_1537_n 0.00422241f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_421 N_B_c_171_n N_VGND_c_1538_n 0.00166854f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_422 N_B_c_172_n N_VGND_c_1538_n 0.00166854f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_423 N_B_c_172_n N_VGND_c_1539_n 0.00422241f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_424 N_B_c_173_n N_VGND_c_1539_n 0.00422241f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_425 N_B_c_173_n N_VGND_c_1540_n 0.00166854f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_426 N_B_c_174_n N_VGND_c_1540_n 0.00166854f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_427 N_B_c_175_n N_VGND_c_1541_n 0.00166854f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_428 N_B_c_176_n N_VGND_c_1541_n 0.00166854f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_429 N_B_c_177_n N_VGND_c_1542_n 0.00166854f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_430 N_B_c_178_n N_VGND_c_1542_n 0.00166854f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_431 N_B_c_179_n N_VGND_c_1543_n 0.00166854f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_432 N_B_c_180_n N_VGND_c_1543_n 0.00296353f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_433 N_B_c_174_n N_VGND_c_1544_n 0.00422241f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_434 N_B_c_175_n N_VGND_c_1544_n 0.00422241f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_435 N_B_c_176_n N_VGND_c_1546_n 0.00422241f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_436 N_B_c_177_n N_VGND_c_1546_n 0.00422241f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_437 N_B_c_178_n N_VGND_c_1548_n 0.00422241f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_438 N_B_c_179_n N_VGND_c_1548_n 0.00422241f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_439 N_B_c_165_n N_VGND_c_1550_n 0.00422241f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_440 N_B_c_180_n N_VGND_c_1551_n 0.00420723f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_441 N_B_c_165_n N_VGND_c_1552_n 0.00689308f $X=0.47 $Y=0.995 $X2=0 $Y2=0
cc_442 N_B_c_166_n N_VGND_c_1552_n 0.00593887f $X=0.99 $Y=0.995 $X2=0 $Y2=0
cc_443 N_B_c_167_n N_VGND_c_1552_n 0.00593887f $X=1.41 $Y=0.995 $X2=0 $Y2=0
cc_444 N_B_c_168_n N_VGND_c_1552_n 0.00593887f $X=1.93 $Y=0.995 $X2=0 $Y2=0
cc_445 N_B_c_169_n N_VGND_c_1552_n 0.00593887f $X=2.35 $Y=0.995 $X2=0 $Y2=0
cc_446 N_B_c_170_n N_VGND_c_1552_n 0.00593887f $X=2.87 $Y=0.995 $X2=0 $Y2=0
cc_447 N_B_c_171_n N_VGND_c_1552_n 0.00593887f $X=3.29 $Y=0.995 $X2=0 $Y2=0
cc_448 N_B_c_172_n N_VGND_c_1552_n 0.00593887f $X=3.81 $Y=0.995 $X2=0 $Y2=0
cc_449 N_B_c_173_n N_VGND_c_1552_n 0.00593887f $X=4.23 $Y=0.995 $X2=0 $Y2=0
cc_450 N_B_c_174_n N_VGND_c_1552_n 0.00593887f $X=4.75 $Y=0.995 $X2=0 $Y2=0
cc_451 N_B_c_175_n N_VGND_c_1552_n 0.00593887f $X=5.17 $Y=0.995 $X2=0 $Y2=0
cc_452 N_B_c_176_n N_VGND_c_1552_n 0.00593887f $X=5.69 $Y=0.995 $X2=0 $Y2=0
cc_453 N_B_c_177_n N_VGND_c_1552_n 0.00593887f $X=6.11 $Y=0.995 $X2=0 $Y2=0
cc_454 N_B_c_178_n N_VGND_c_1552_n 0.00593887f $X=6.63 $Y=0.995 $X2=0 $Y2=0
cc_455 N_B_c_179_n N_VGND_c_1552_n 0.00593887f $X=7.05 $Y=0.995 $X2=0 $Y2=0
cc_456 N_B_c_180_n N_VGND_c_1552_n 0.00597515f $X=7.57 $Y=0.995 $X2=0 $Y2=0
cc_457 N_A_c_510_n N_VPWR_c_762_n 0.00173895f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_458 N_A_c_511_n N_VPWR_c_763_n 0.00173895f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_459 N_A_c_512_n N_VPWR_c_763_n 0.00173895f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_460 N_A_c_513_n N_VPWR_c_764_n 0.00173895f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_461 N_A_c_514_n N_VPWR_c_764_n 0.00173895f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_462 N_A_c_515_n N_VPWR_c_765_n 0.00173895f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_463 N_A_c_516_n N_VPWR_c_765_n 0.00173895f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_464 N_A_c_517_n N_VPWR_c_766_n 0.00173895f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_465 N_A_c_518_n N_VPWR_c_766_n 0.00173895f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_466 N_A_c_519_n N_VPWR_c_767_n 0.00173895f $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_467 N_A_c_520_n N_VPWR_c_767_n 0.00173895f $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_468 N_A_c_521_n N_VPWR_c_768_n 0.00173895f $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_469 N_A_c_522_n N_VPWR_c_768_n 0.00173895f $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_470 N_A_c_523_n N_VPWR_c_769_n 0.00173895f $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_471 N_A_c_524_n N_VPWR_c_769_n 0.00173895f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_472 N_A_c_525_n N_VPWR_c_771_n 0.00354866f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_473 N_A_c_510_n N_VPWR_c_778_n 0.00673617f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_474 N_A_c_511_n N_VPWR_c_778_n 0.00673617f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_475 N_A_c_512_n N_VPWR_c_780_n 0.00673617f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_476 N_A_c_513_n N_VPWR_c_780_n 0.00673617f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_477 N_A_c_514_n N_VPWR_c_782_n 0.00673617f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_478 N_A_c_515_n N_VPWR_c_782_n 0.00673617f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_479 N_A_c_516_n N_VPWR_c_784_n 0.00673617f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_480 N_A_c_517_n N_VPWR_c_784_n 0.00673617f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_481 N_A_c_518_n N_VPWR_c_786_n 0.00673617f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_482 N_A_c_519_n N_VPWR_c_786_n 0.00673617f $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_483 N_A_c_520_n N_VPWR_c_788_n 0.00673617f $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_484 N_A_c_521_n N_VPWR_c_788_n 0.00673617f $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_485 N_A_c_522_n N_VPWR_c_790_n 0.00673617f $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_486 N_A_c_523_n N_VPWR_c_790_n 0.00673617f $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_487 N_A_c_524_n N_VPWR_c_793_n 0.00673617f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_488 N_A_c_525_n N_VPWR_c_793_n 0.00673617f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_489 N_A_c_510_n N_VPWR_c_748_n 0.0117436f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_490 N_A_c_511_n N_VPWR_c_748_n 0.0117184f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_491 N_A_c_512_n N_VPWR_c_748_n 0.0117184f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_492 N_A_c_513_n N_VPWR_c_748_n 0.0117184f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_493 N_A_c_514_n N_VPWR_c_748_n 0.0117184f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_494 N_A_c_515_n N_VPWR_c_748_n 0.0117184f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_495 N_A_c_516_n N_VPWR_c_748_n 0.0117184f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_496 N_A_c_517_n N_VPWR_c_748_n 0.0117184f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_497 N_A_c_518_n N_VPWR_c_748_n 0.0117184f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_498 N_A_c_519_n N_VPWR_c_748_n 0.0117184f $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_499 N_A_c_520_n N_VPWR_c_748_n 0.0117184f $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_500 N_A_c_521_n N_VPWR_c_748_n 0.0117184f $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_501 N_A_c_522_n N_VPWR_c_748_n 0.0117184f $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_502 N_A_c_523_n N_VPWR_c_748_n 0.0117184f $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_503 N_A_c_524_n N_VPWR_c_748_n 0.0117184f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_504 N_A_c_525_n N_VPWR_c_748_n 0.0126961f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_505 N_A_c_510_n N_Y_c_1039_n 5.91934e-19 $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_506 N_A_c_493_n N_Y_c_1078_n 0.00303037f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_507 N_A_c_510_n N_Y_c_1044_n 0.0100233f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_508 N_A_c_511_n N_Y_c_1044_n 0.0100233f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_509 N_A_c_512_n N_Y_c_1044_n 5.91934e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_510 N_A_c_494_n N_Y_c_1082_n 0.0124451f $X=8.46 $Y=0.995 $X2=0 $Y2=0
cc_511 N_A_c_495_n N_Y_c_1082_n 0.0109111f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_512 N_A_c_496_n N_Y_c_1082_n 0.0104739f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_513 N_A_c_497_n N_Y_c_1082_n 0.0104739f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_514 N_A_c_498_n N_Y_c_1082_n 0.0104739f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_515 N_A_c_499_n N_Y_c_1082_n 0.0104739f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_516 N_A_c_500_n N_Y_c_1082_n 0.0109111f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_517 N_A_c_501_n N_Y_c_1082_n 0.0109111f $X=11.75 $Y=0.995 $X2=0 $Y2=0
cc_518 N_A_c_502_n N_Y_c_1082_n 0.0104739f $X=12.27 $Y=0.995 $X2=0 $Y2=0
cc_519 N_A_c_503_n N_Y_c_1082_n 0.0104739f $X=12.69 $Y=0.995 $X2=0 $Y2=0
cc_520 N_A_c_504_n N_Y_c_1082_n 0.0104739f $X=13.21 $Y=0.995 $X2=0 $Y2=0
cc_521 N_A_c_505_n N_Y_c_1082_n 0.0104739f $X=13.63 $Y=0.995 $X2=0 $Y2=0
cc_522 N_A_c_506_n N_Y_c_1082_n 0.0104739f $X=14.15 $Y=0.995 $X2=0 $Y2=0
cc_523 N_A_c_507_n N_Y_c_1082_n 0.0123979f $X=14.57 $Y=0.995 $X2=0 $Y2=0
cc_524 N_A_c_598_p N_Y_c_1082_n 0.372356f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_525 N_A_c_509_n N_Y_c_1082_n 0.0447032f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_526 N_A_c_511_n N_Y_c_1098_n 0.014973f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_527 N_A_c_512_n N_Y_c_1098_n 0.0137916f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_528 N_A_c_598_p N_Y_c_1098_n 0.0330732f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_529 N_A_c_509_n N_Y_c_1098_n 0.00635951f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_530 N_A_c_511_n N_Y_c_1102_n 5.91934e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_531 N_A_c_512_n N_Y_c_1102_n 0.0100233f $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_532 N_A_c_513_n N_Y_c_1102_n 0.0100233f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_533 N_A_c_514_n N_Y_c_1102_n 5.91934e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_534 N_A_c_513_n N_Y_c_1106_n 0.0137916f $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_535 N_A_c_514_n N_Y_c_1106_n 0.0137916f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_536 N_A_c_598_p N_Y_c_1106_n 0.0393642f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_537 N_A_c_509_n N_Y_c_1106_n 0.00655651f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_538 N_A_c_513_n N_Y_c_1110_n 5.91934e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_539 N_A_c_514_n N_Y_c_1110_n 0.0100233f $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_540 N_A_c_515_n N_Y_c_1110_n 0.0100233f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_541 N_A_c_516_n N_Y_c_1110_n 5.91934e-19 $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_542 N_A_c_515_n N_Y_c_1114_n 0.0137916f $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_543 N_A_c_516_n N_Y_c_1114_n 0.0137916f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_544 N_A_c_598_p N_Y_c_1114_n 0.0393642f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_545 N_A_c_509_n N_Y_c_1114_n 0.00655651f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_546 N_A_c_515_n N_Y_c_1118_n 5.91934e-19 $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_547 N_A_c_516_n N_Y_c_1118_n 0.0100233f $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_548 N_A_c_517_n N_Y_c_1118_n 0.0100233f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_549 N_A_c_518_n N_Y_c_1118_n 5.91934e-19 $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_550 N_A_c_517_n N_Y_c_1122_n 0.0137916f $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_551 N_A_c_518_n N_Y_c_1122_n 0.0137916f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_552 N_A_c_598_p N_Y_c_1122_n 0.0393642f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_553 N_A_c_509_n N_Y_c_1122_n 0.00635951f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_554 N_A_c_517_n N_Y_c_1126_n 5.91934e-19 $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_555 N_A_c_518_n N_Y_c_1126_n 0.0100233f $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_556 N_A_c_519_n N_Y_c_1126_n 0.0100233f $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_557 N_A_c_520_n N_Y_c_1126_n 5.91934e-19 $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_558 N_A_c_519_n N_Y_c_1130_n 0.0137916f $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_559 N_A_c_520_n N_Y_c_1130_n 0.0137916f $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_560 N_A_c_598_p N_Y_c_1130_n 0.0393642f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_561 N_A_c_509_n N_Y_c_1130_n 0.00655651f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_562 N_A_c_519_n N_Y_c_1134_n 5.91934e-19 $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_563 N_A_c_520_n N_Y_c_1134_n 0.0100233f $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_564 N_A_c_521_n N_Y_c_1134_n 0.0100233f $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_565 N_A_c_522_n N_Y_c_1134_n 5.91934e-19 $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_566 N_A_c_521_n N_Y_c_1138_n 0.0137916f $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_567 N_A_c_522_n N_Y_c_1138_n 0.0137916f $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_568 N_A_c_598_p N_Y_c_1138_n 0.0393642f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_569 N_A_c_509_n N_Y_c_1138_n 0.00655651f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_570 N_A_c_521_n N_Y_c_1142_n 5.91934e-19 $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_571 N_A_c_522_n N_Y_c_1142_n 0.0100233f $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_572 N_A_c_523_n N_Y_c_1142_n 0.0100233f $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_573 N_A_c_524_n N_Y_c_1142_n 5.91934e-19 $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_574 N_A_c_523_n N_Y_c_1146_n 0.0137916f $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_575 N_A_c_524_n N_Y_c_1146_n 0.0159022f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_576 N_A_c_598_p N_Y_c_1146_n 0.0135025f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_577 N_A_c_509_n N_Y_c_1146_n 0.00732298f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_578 N_A_c_523_n N_Y_c_1150_n 5.91934e-19 $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_579 N_A_c_524_n N_Y_c_1150_n 0.0100233f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_580 N_A_c_525_n N_Y_c_1150_n 0.00897418f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_581 N_A_c_524_n N_Y_c_978_n 0.0019905f $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_582 N_A_c_525_n N_Y_c_978_n 0.00423504f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_583 N_A_c_509_n N_Y_c_978_n 0.00694896f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_584 N_A_c_510_n N_Y_c_1156_n 0.0130984f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_585 N_A_c_511_n N_Y_c_1156_n 8.15944e-19 $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_586 N_A_c_509_n N_Y_c_1156_n 0.00123735f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_587 N_A_c_512_n N_Y_c_1159_n 5.79575e-19 $X=8.955 $Y=1.41 $X2=0 $Y2=0
cc_588 N_A_c_513_n N_Y_c_1159_n 5.79575e-19 $X=9.425 $Y=1.41 $X2=0 $Y2=0
cc_589 N_A_c_598_p N_Y_c_1159_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_590 N_A_c_509_n N_Y_c_1159_n 0.00631893f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_591 N_A_c_514_n N_Y_c_1163_n 5.79575e-19 $X=9.895 $Y=1.41 $X2=0 $Y2=0
cc_592 N_A_c_515_n N_Y_c_1163_n 5.79575e-19 $X=10.365 $Y=1.41 $X2=0 $Y2=0
cc_593 N_A_c_598_p N_Y_c_1163_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_594 N_A_c_509_n N_Y_c_1163_n 0.00631893f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_595 N_A_c_516_n N_Y_c_1167_n 5.79575e-19 $X=10.835 $Y=1.41 $X2=0 $Y2=0
cc_596 N_A_c_517_n N_Y_c_1167_n 5.79575e-19 $X=11.305 $Y=1.41 $X2=0 $Y2=0
cc_597 N_A_c_598_p N_Y_c_1167_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_598 N_A_c_509_n N_Y_c_1167_n 0.00651614f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_599 N_A_c_518_n N_Y_c_1171_n 5.79575e-19 $X=11.775 $Y=1.41 $X2=0 $Y2=0
cc_600 N_A_c_519_n N_Y_c_1171_n 5.79575e-19 $X=12.245 $Y=1.41 $X2=0 $Y2=0
cc_601 N_A_c_598_p N_Y_c_1171_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_602 N_A_c_509_n N_Y_c_1171_n 0.00631893f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_603 N_A_c_520_n N_Y_c_1175_n 5.79575e-19 $X=12.715 $Y=1.41 $X2=0 $Y2=0
cc_604 N_A_c_521_n N_Y_c_1175_n 5.79575e-19 $X=13.185 $Y=1.41 $X2=0 $Y2=0
cc_605 N_A_c_598_p N_Y_c_1175_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_606 N_A_c_509_n N_Y_c_1175_n 0.00631893f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_607 N_A_c_522_n N_Y_c_1179_n 5.79575e-19 $X=13.655 $Y=1.41 $X2=0 $Y2=0
cc_608 N_A_c_523_n N_Y_c_1179_n 5.79575e-19 $X=14.125 $Y=1.41 $X2=0 $Y2=0
cc_609 N_A_c_598_p N_Y_c_1179_n 0.0215641f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_610 N_A_c_509_n N_Y_c_1179_n 0.00631893f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_611 N_A_c_524_n N_Y_c_1183_n 8.15944e-19 $X=14.595 $Y=1.41 $X2=0 $Y2=0
cc_612 N_A_c_525_n N_Y_c_1183_n 0.00188422f $X=15.065 $Y=1.41 $X2=0 $Y2=0
cc_613 N_A_c_507_n N_Y_c_976_n 0.00286869f $X=14.57 $Y=0.995 $X2=0 $Y2=0
cc_614 N_A_c_508_n N_Y_c_976_n 0.0031043f $X=15.09 $Y=0.995 $X2=0 $Y2=0
cc_615 N_A_c_509_n N_Y_c_976_n 0.0106358f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_616 N_A_c_598_p N_Y_c_1188_n 0.00981282f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_617 N_A_c_509_n N_Y_c_1188_n 0.0421699f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_618 N_A_c_510_n Y 0.00326841f $X=8.015 $Y=1.41 $X2=0 $Y2=0
cc_619 N_A_c_511_n Y 0.00234191f $X=8.485 $Y=1.41 $X2=0 $Y2=0
cc_620 N_A_c_598_p Y 0.0216953f $X=14.11 $Y=1.16 $X2=0 $Y2=0
cc_621 N_A_c_509_n Y 0.0313911f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_622 N_A_c_493_n N_Y_c_977_n 0.00315482f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_623 N_A_c_494_n N_Y_c_977_n 0.00297134f $X=8.46 $Y=0.995 $X2=0 $Y2=0
cc_624 N_A_c_509_n N_Y_c_977_n 0.00830622f $X=15.065 $Y=1.202 $X2=0 $Y2=0
cc_625 N_A_c_493_n N_A_27_47#_c_1412_n 0.0108171f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_626 N_A_c_494_n N_A_27_47#_c_1412_n 0.00903374f $X=8.46 $Y=0.995 $X2=0 $Y2=0
cc_627 N_A_c_495_n N_A_27_47#_c_1412_n 0.00935436f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_628 N_A_c_496_n N_A_27_47#_c_1412_n 0.00935436f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_629 N_A_c_497_n N_A_27_47#_c_1412_n 0.00935436f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_630 N_A_c_498_n N_A_27_47#_c_1412_n 0.00935436f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_631 N_A_c_499_n N_A_27_47#_c_1412_n 0.00903374f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_632 N_A_c_500_n N_A_27_47#_c_1412_n 0.00903374f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_633 N_A_c_501_n N_A_27_47#_c_1412_n 0.00935436f $X=11.75 $Y=0.995 $X2=0 $Y2=0
cc_634 N_A_c_502_n N_A_27_47#_c_1412_n 0.00935436f $X=12.27 $Y=0.995 $X2=0 $Y2=0
cc_635 N_A_c_503_n N_A_27_47#_c_1412_n 0.00935436f $X=12.69 $Y=0.995 $X2=0 $Y2=0
cc_636 N_A_c_504_n N_A_27_47#_c_1412_n 0.00935436f $X=13.21 $Y=0.995 $X2=0 $Y2=0
cc_637 N_A_c_505_n N_A_27_47#_c_1412_n 0.00935436f $X=13.63 $Y=0.995 $X2=0 $Y2=0
cc_638 N_A_c_506_n N_A_27_47#_c_1412_n 0.00935436f $X=14.15 $Y=0.995 $X2=0 $Y2=0
cc_639 N_A_c_507_n N_A_27_47#_c_1412_n 0.00935436f $X=14.57 $Y=0.995 $X2=0 $Y2=0
cc_640 N_A_c_508_n N_A_27_47#_c_1412_n 0.0122646f $X=15.09 $Y=0.995 $X2=0 $Y2=0
cc_641 N_A_c_509_n N_A_27_47#_c_1412_n 0.00110461f $X=15.065 $Y=1.202 $X2=0
+ $Y2=0
cc_642 N_A_c_493_n N_VGND_c_1551_n 0.00357877f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_643 N_A_c_494_n N_VGND_c_1551_n 0.00357877f $X=8.46 $Y=0.995 $X2=0 $Y2=0
cc_644 N_A_c_495_n N_VGND_c_1551_n 0.00357877f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_645 N_A_c_496_n N_VGND_c_1551_n 0.00357877f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_646 N_A_c_497_n N_VGND_c_1551_n 0.00357877f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_647 N_A_c_498_n N_VGND_c_1551_n 0.00357877f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_648 N_A_c_499_n N_VGND_c_1551_n 0.00357877f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_649 N_A_c_500_n N_VGND_c_1551_n 0.00357877f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_650 N_A_c_501_n N_VGND_c_1551_n 0.00357877f $X=11.75 $Y=0.995 $X2=0 $Y2=0
cc_651 N_A_c_502_n N_VGND_c_1551_n 0.00357877f $X=12.27 $Y=0.995 $X2=0 $Y2=0
cc_652 N_A_c_503_n N_VGND_c_1551_n 0.00357877f $X=12.69 $Y=0.995 $X2=0 $Y2=0
cc_653 N_A_c_504_n N_VGND_c_1551_n 0.00357877f $X=13.21 $Y=0.995 $X2=0 $Y2=0
cc_654 N_A_c_505_n N_VGND_c_1551_n 0.00357877f $X=13.63 $Y=0.995 $X2=0 $Y2=0
cc_655 N_A_c_506_n N_VGND_c_1551_n 0.00357877f $X=14.15 $Y=0.995 $X2=0 $Y2=0
cc_656 N_A_c_507_n N_VGND_c_1551_n 0.00357877f $X=14.57 $Y=0.995 $X2=0 $Y2=0
cc_657 N_A_c_508_n N_VGND_c_1551_n 0.00357877f $X=15.09 $Y=0.995 $X2=0 $Y2=0
cc_658 N_A_c_493_n N_VGND_c_1552_n 0.00538422f $X=7.99 $Y=0.995 $X2=0 $Y2=0
cc_659 N_A_c_494_n N_VGND_c_1552_n 0.00548399f $X=8.46 $Y=0.995 $X2=0 $Y2=0
cc_660 N_A_c_495_n N_VGND_c_1552_n 0.00560377f $X=8.93 $Y=0.995 $X2=0 $Y2=0
cc_661 N_A_c_496_n N_VGND_c_1552_n 0.0054768f $X=9.45 $Y=0.995 $X2=0 $Y2=0
cc_662 N_A_c_497_n N_VGND_c_1552_n 0.0054768f $X=9.87 $Y=0.995 $X2=0 $Y2=0
cc_663 N_A_c_498_n N_VGND_c_1552_n 0.0054768f $X=10.39 $Y=0.995 $X2=0 $Y2=0
cc_664 N_A_c_499_n N_VGND_c_1552_n 0.00535702f $X=10.81 $Y=0.995 $X2=0 $Y2=0
cc_665 N_A_c_500_n N_VGND_c_1552_n 0.00548399f $X=11.28 $Y=0.995 $X2=0 $Y2=0
cc_666 N_A_c_501_n N_VGND_c_1552_n 0.00560377f $X=11.75 $Y=0.995 $X2=0 $Y2=0
cc_667 N_A_c_502_n N_VGND_c_1552_n 0.0054768f $X=12.27 $Y=0.995 $X2=0 $Y2=0
cc_668 N_A_c_503_n N_VGND_c_1552_n 0.0054768f $X=12.69 $Y=0.995 $X2=0 $Y2=0
cc_669 N_A_c_504_n N_VGND_c_1552_n 0.0054768f $X=13.21 $Y=0.995 $X2=0 $Y2=0
cc_670 N_A_c_505_n N_VGND_c_1552_n 0.0054768f $X=13.63 $Y=0.995 $X2=0 $Y2=0
cc_671 N_A_c_506_n N_VGND_c_1552_n 0.0054768f $X=14.15 $Y=0.995 $X2=0 $Y2=0
cc_672 N_A_c_507_n N_VGND_c_1552_n 0.0054768f $X=14.57 $Y=0.995 $X2=0 $Y2=0
cc_673 N_A_c_508_n N_VGND_c_1552_n 0.00649939f $X=15.09 $Y=0.995 $X2=0 $Y2=0
cc_674 N_VPWR_c_748_n N_Y_M1000_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_675 N_VPWR_c_748_n N_Y_M1007_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_676 N_VPWR_c_748_n N_Y_M1010_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_677 N_VPWR_c_748_n N_Y_M1019_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_678 N_VPWR_c_748_n N_Y_M1033_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_679 N_VPWR_c_748_n N_Y_M1042_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_680 N_VPWR_c_748_n N_Y_M1050_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_681 N_VPWR_c_748_n N_Y_M1054_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_682 N_VPWR_c_748_n N_Y_M1003_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_683 N_VPWR_c_748_n N_Y_M1012_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_684 N_VPWR_c_748_n N_Y_M1021_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_685 N_VPWR_c_748_n N_Y_M1023_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_686 N_VPWR_c_748_n N_Y_M1031_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_687 N_VPWR_c_748_n N_Y_M1041_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_688 N_VPWR_c_748_n N_Y_M1049_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_689 N_VPWR_c_748_n N_Y_M1061_s 0.00231261f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_690 N_VPWR_c_792_n N_Y_c_984_n 0.0189467f $X=1.065 $Y=2.72 $X2=0 $Y2=0
cc_691 N_VPWR_c_748_n N_Y_c_984_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_692 N_VPWR_M1002_d N_Y_c_987_n 0.00334388f $X=1.055 $Y=1.485 $X2=0 $Y2=0
cc_693 N_VPWR_c_751_n N_Y_c_987_n 0.0143191f $X=1.2 $Y=2 $X2=0 $Y2=0
cc_694 N_VPWR_c_752_n N_Y_c_991_n 0.0189467f $X=2.005 $Y=2.72 $X2=0 $Y2=0
cc_695 N_VPWR_c_748_n N_Y_c_991_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_696 N_VPWR_M1009_d N_Y_c_995_n 0.00334388f $X=1.995 $Y=1.485 $X2=0 $Y2=0
cc_697 N_VPWR_c_753_n N_Y_c_995_n 0.0143191f $X=2.14 $Y=2 $X2=0 $Y2=0
cc_698 N_VPWR_c_754_n N_Y_c_999_n 0.0189467f $X=2.945 $Y=2.72 $X2=0 $Y2=0
cc_699 N_VPWR_c_748_n N_Y_c_999_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_700 N_VPWR_M1015_d N_Y_c_1003_n 0.00334388f $X=2.935 $Y=1.485 $X2=0 $Y2=0
cc_701 N_VPWR_c_755_n N_Y_c_1003_n 0.0143191f $X=3.08 $Y=2 $X2=0 $Y2=0
cc_702 N_VPWR_c_756_n N_Y_c_1007_n 0.0189467f $X=3.885 $Y=2.72 $X2=0 $Y2=0
cc_703 N_VPWR_c_748_n N_Y_c_1007_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_704 N_VPWR_M1028_d N_Y_c_1011_n 0.00334388f $X=3.875 $Y=1.485 $X2=0 $Y2=0
cc_705 N_VPWR_c_757_n N_Y_c_1011_n 0.0143191f $X=4.02 $Y=2 $X2=0 $Y2=0
cc_706 N_VPWR_c_758_n N_Y_c_1015_n 0.0189467f $X=4.825 $Y=2.72 $X2=0 $Y2=0
cc_707 N_VPWR_c_748_n N_Y_c_1015_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_708 N_VPWR_M1037_d N_Y_c_1019_n 0.00334388f $X=4.815 $Y=1.485 $X2=0 $Y2=0
cc_709 N_VPWR_c_759_n N_Y_c_1019_n 0.0143191f $X=4.96 $Y=2 $X2=0 $Y2=0
cc_710 N_VPWR_c_772_n N_Y_c_1023_n 0.0189467f $X=5.765 $Y=2.72 $X2=0 $Y2=0
cc_711 N_VPWR_c_748_n N_Y_c_1023_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_712 N_VPWR_M1045_d N_Y_c_1027_n 0.00334388f $X=5.755 $Y=1.485 $X2=0 $Y2=0
cc_713 N_VPWR_c_760_n N_Y_c_1027_n 0.0143191f $X=5.9 $Y=2 $X2=0 $Y2=0
cc_714 N_VPWR_c_774_n N_Y_c_1031_n 0.0189467f $X=6.705 $Y=2.72 $X2=0 $Y2=0
cc_715 N_VPWR_c_748_n N_Y_c_1031_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_716 N_VPWR_M1051_d N_Y_c_1035_n 0.00334388f $X=6.695 $Y=1.485 $X2=0 $Y2=0
cc_717 N_VPWR_c_761_n N_Y_c_1035_n 0.0143191f $X=6.84 $Y=2 $X2=0 $Y2=0
cc_718 N_VPWR_c_776_n N_Y_c_1039_n 0.0189467f $X=7.645 $Y=2.72 $X2=0 $Y2=0
cc_719 N_VPWR_c_748_n N_Y_c_1039_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_720 N_VPWR_M1060_d N_Y_c_1042_n 0.00534233f $X=7.635 $Y=1.485 $X2=0 $Y2=0
cc_721 N_VPWR_c_762_n N_Y_c_1042_n 0.0143191f $X=7.78 $Y=2 $X2=0 $Y2=0
cc_722 N_VPWR_c_778_n N_Y_c_1044_n 0.0189467f $X=8.585 $Y=2.72 $X2=0 $Y2=0
cc_723 N_VPWR_c_748_n N_Y_c_1044_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_724 N_VPWR_M1008_d N_Y_c_1098_n 0.00334388f $X=8.575 $Y=1.485 $X2=0 $Y2=0
cc_725 N_VPWR_c_763_n N_Y_c_1098_n 0.0143191f $X=8.72 $Y=2 $X2=0 $Y2=0
cc_726 N_VPWR_c_780_n N_Y_c_1102_n 0.0189467f $X=9.525 $Y=2.72 $X2=0 $Y2=0
cc_727 N_VPWR_c_748_n N_Y_c_1102_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_728 N_VPWR_M1013_d N_Y_c_1106_n 0.00334388f $X=9.515 $Y=1.485 $X2=0 $Y2=0
cc_729 N_VPWR_c_764_n N_Y_c_1106_n 0.0143191f $X=9.66 $Y=2 $X2=0 $Y2=0
cc_730 N_VPWR_c_782_n N_Y_c_1110_n 0.0189467f $X=10.465 $Y=2.72 $X2=0 $Y2=0
cc_731 N_VPWR_c_748_n N_Y_c_1110_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_732 N_VPWR_M1022_d N_Y_c_1114_n 0.00334388f $X=10.455 $Y=1.485 $X2=0 $Y2=0
cc_733 N_VPWR_c_765_n N_Y_c_1114_n 0.0143191f $X=10.6 $Y=2 $X2=0 $Y2=0
cc_734 N_VPWR_c_784_n N_Y_c_1118_n 0.0189467f $X=11.405 $Y=2.72 $X2=0 $Y2=0
cc_735 N_VPWR_c_748_n N_Y_c_1118_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_736 N_VPWR_M1029_d N_Y_c_1122_n 0.00334388f $X=11.395 $Y=1.485 $X2=0 $Y2=0
cc_737 N_VPWR_c_766_n N_Y_c_1122_n 0.0143191f $X=11.54 $Y=2 $X2=0 $Y2=0
cc_738 N_VPWR_c_786_n N_Y_c_1126_n 0.0189467f $X=12.345 $Y=2.72 $X2=0 $Y2=0
cc_739 N_VPWR_c_748_n N_Y_c_1126_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_740 N_VPWR_M1038_d N_Y_c_1130_n 0.00334388f $X=12.335 $Y=1.485 $X2=0 $Y2=0
cc_741 N_VPWR_c_767_n N_Y_c_1130_n 0.0143191f $X=12.48 $Y=2 $X2=0 $Y2=0
cc_742 N_VPWR_c_788_n N_Y_c_1134_n 0.0189467f $X=13.285 $Y=2.72 $X2=0 $Y2=0
cc_743 N_VPWR_c_748_n N_Y_c_1134_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_744 N_VPWR_M1048_d N_Y_c_1138_n 0.00334388f $X=13.275 $Y=1.485 $X2=0 $Y2=0
cc_745 N_VPWR_c_768_n N_Y_c_1138_n 0.0143191f $X=13.42 $Y=2 $X2=0 $Y2=0
cc_746 N_VPWR_c_790_n N_Y_c_1142_n 0.0189467f $X=14.225 $Y=2.72 $X2=0 $Y2=0
cc_747 N_VPWR_c_748_n N_Y_c_1142_n 0.0123132f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_748 N_VPWR_M1052_d N_Y_c_1146_n 0.00419101f $X=14.215 $Y=1.485 $X2=0 $Y2=0
cc_749 N_VPWR_c_769_n N_Y_c_1146_n 0.0143191f $X=14.36 $Y=2 $X2=0 $Y2=0
cc_750 N_VPWR_c_793_n N_Y_c_1150_n 0.0189467f $X=15.165 $Y=2.72 $X2=0 $Y2=0
cc_751 N_VPWR_c_748_n N_Y_c_1150_n 0.0123027f $X=15.41 $Y=2.72 $X2=0 $Y2=0
cc_752 N_VPWR_c_750_n N_A_27_47#_c_1306_n 0.00746809f $X=0.26 $Y=1.66 $X2=0
+ $Y2=0
cc_753 N_VPWR_c_771_n N_A_27_47#_c_1309_n 0.00739919f $X=15.3 $Y=1.66 $X2=0
+ $Y2=0
cc_754 N_Y_c_1082_n N_A_27_47#_M1006_s 0.00401355f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_755 N_Y_c_1082_n N_A_27_47#_M1017_s 0.00307883f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_756 N_Y_c_1082_n N_A_27_47#_M1024_s 0.00307883f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_757 N_Y_c_1082_n N_A_27_47#_M1027_s 0.00401355f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_758 N_Y_c_1082_n N_A_27_47#_M1032_s 0.00307883f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_759 N_Y_c_1082_n N_A_27_47#_M1043_s 0.00307883f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_760 N_Y_c_1082_n N_A_27_47#_M1047_s 0.00404759f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_761 N_Y_c_1042_n N_A_27_47#_c_1377_n 0.00210535f $X=7.925 $Y=1.58 $X2=0 $Y2=0
cc_762 N_Y_c_1042_n N_A_27_47#_c_1307_n 0.00572467f $X=7.925 $Y=1.58 $X2=0 $Y2=0
cc_763 N_Y_M1001_d N_A_27_47#_c_1412_n 0.00399738f $X=8.065 $Y=0.235 $X2=0 $Y2=0
cc_764 N_Y_M1011_d N_A_27_47#_c_1412_n 0.00507102f $X=9.005 $Y=0.235 $X2=0 $Y2=0
cc_765 N_Y_M1018_d N_A_27_47#_c_1412_n 0.00507102f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_766 N_Y_M1026_d N_A_27_47#_c_1412_n 0.00400219f $X=10.885 $Y=0.235 $X2=0
+ $Y2=0
cc_767 N_Y_M1030_d N_A_27_47#_c_1412_n 0.00507102f $X=11.825 $Y=0.235 $X2=0
+ $Y2=0
cc_768 N_Y_M1036_d N_A_27_47#_c_1412_n 0.00507102f $X=12.765 $Y=0.235 $X2=0
+ $Y2=0
cc_769 N_Y_M1044_d N_A_27_47#_c_1412_n 0.00507102f $X=13.705 $Y=0.235 $X2=0
+ $Y2=0
cc_770 N_Y_M1059_d N_A_27_47#_c_1412_n 0.00506571f $X=14.645 $Y=0.235 $X2=0
+ $Y2=0
cc_771 N_Y_c_1078_n N_A_27_47#_c_1412_n 0.0182216f $X=8.185 $Y=0.885 $X2=0 $Y2=0
cc_772 N_Y_c_1082_n N_A_27_47#_c_1412_n 0.334928f $X=14.725 $Y=0.76 $X2=0 $Y2=0
cc_773 N_Y_c_1294_p N_A_27_47#_c_1412_n 0.018174f $X=14.86 $Y=0.885 $X2=0 $Y2=0
cc_774 N_Y_c_1188_n N_A_27_47#_c_1412_n 0.00279601f $X=14.92 $Y=1.325 $X2=0
+ $Y2=0
cc_775 Y N_A_27_47#_c_1412_n 0.00297886f $X=7.965 $Y=1.105 $X2=0 $Y2=0
cc_776 N_Y_M1001_d N_VGND_c_1552_n 0.00256987f $X=8.065 $Y=0.235 $X2=0 $Y2=0
cc_777 N_Y_M1011_d N_VGND_c_1552_n 0.00297142f $X=9.005 $Y=0.235 $X2=0 $Y2=0
cc_778 N_Y_M1018_d N_VGND_c_1552_n 0.00297142f $X=9.945 $Y=0.235 $X2=0 $Y2=0
cc_779 N_Y_M1026_d N_VGND_c_1552_n 0.00256987f $X=10.885 $Y=0.235 $X2=0 $Y2=0
cc_780 N_Y_M1030_d N_VGND_c_1552_n 0.00297142f $X=11.825 $Y=0.235 $X2=0 $Y2=0
cc_781 N_Y_M1036_d N_VGND_c_1552_n 0.00297142f $X=12.765 $Y=0.235 $X2=0 $Y2=0
cc_782 N_Y_M1044_d N_VGND_c_1552_n 0.00297142f $X=13.705 $Y=0.235 $X2=0 $Y2=0
cc_783 N_Y_M1059_d N_VGND_c_1552_n 0.00297142f $X=14.645 $Y=0.235 $X2=0 $Y2=0
cc_784 N_A_27_47#_c_1319_n N_VGND_M1004_s 0.00500594f $X=1.035 $Y=0.8 $X2=-0.19
+ $Y2=-0.24
cc_785 N_A_27_47#_c_1329_n N_VGND_M1014_s 0.00500594f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_786 N_A_27_47#_c_1337_n N_VGND_M1020_s 0.00500594f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_787 N_A_27_47#_c_1345_n N_VGND_M1034_s 0.00500594f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_788 N_A_27_47#_c_1353_n N_VGND_M1039_s 0.00500594f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_789 N_A_27_47#_c_1361_n N_VGND_M1046_s 0.00500594f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_790 N_A_27_47#_c_1369_n N_VGND_M1055_s 0.00500594f $X=6.675 $Y=0.8 $X2=0
+ $Y2=0
cc_791 N_A_27_47#_c_1377_n N_VGND_M1057_s 0.00500594f $X=7.615 $Y=0.8 $X2=0
+ $Y2=0
cc_792 N_A_27_47#_c_1319_n N_VGND_c_1532_n 0.0199861f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_793 N_A_27_47#_c_1319_n N_VGND_c_1533_n 0.0020257f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_794 N_A_27_47#_c_1325_n N_VGND_c_1533_n 0.0188215f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_795 N_A_27_47#_c_1329_n N_VGND_c_1533_n 0.0020257f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_796 N_A_27_47#_c_1329_n N_VGND_c_1534_n 0.0199861f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_797 N_A_27_47#_c_1329_n N_VGND_c_1535_n 0.0020257f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_798 N_A_27_47#_c_1333_n N_VGND_c_1535_n 0.0188215f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_799 N_A_27_47#_c_1337_n N_VGND_c_1535_n 0.0020257f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_800 N_A_27_47#_c_1337_n N_VGND_c_1536_n 0.0199861f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_801 N_A_27_47#_c_1337_n N_VGND_c_1537_n 0.0020257f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_802 N_A_27_47#_c_1341_n N_VGND_c_1537_n 0.0188215f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_803 N_A_27_47#_c_1345_n N_VGND_c_1537_n 0.0020257f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_804 N_A_27_47#_c_1345_n N_VGND_c_1538_n 0.0199861f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_805 N_A_27_47#_c_1345_n N_VGND_c_1539_n 0.0020257f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_806 N_A_27_47#_c_1349_n N_VGND_c_1539_n 0.0188215f $X=4.02 $Y=0.38 $X2=0
+ $Y2=0
cc_807 N_A_27_47#_c_1353_n N_VGND_c_1539_n 0.0020257f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_808 N_A_27_47#_c_1353_n N_VGND_c_1540_n 0.0199861f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_809 N_A_27_47#_c_1361_n N_VGND_c_1541_n 0.0199861f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_810 N_A_27_47#_c_1369_n N_VGND_c_1542_n 0.0199861f $X=6.675 $Y=0.8 $X2=0
+ $Y2=0
cc_811 N_A_27_47#_c_1377_n N_VGND_c_1543_n 0.0199861f $X=7.615 $Y=0.8 $X2=0
+ $Y2=0
cc_812 N_A_27_47#_c_1353_n N_VGND_c_1544_n 0.0020257f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_813 N_A_27_47#_c_1357_n N_VGND_c_1544_n 0.0188215f $X=4.96 $Y=0.38 $X2=0
+ $Y2=0
cc_814 N_A_27_47#_c_1361_n N_VGND_c_1544_n 0.0020257f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_815 N_A_27_47#_c_1361_n N_VGND_c_1546_n 0.0020257f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_816 N_A_27_47#_c_1365_n N_VGND_c_1546_n 0.0188215f $X=5.9 $Y=0.38 $X2=0 $Y2=0
cc_817 N_A_27_47#_c_1369_n N_VGND_c_1546_n 0.0020257f $X=6.675 $Y=0.8 $X2=0
+ $Y2=0
cc_818 N_A_27_47#_c_1369_n N_VGND_c_1548_n 0.0020257f $X=6.675 $Y=0.8 $X2=0
+ $Y2=0
cc_819 N_A_27_47#_c_1373_n N_VGND_c_1548_n 0.0188215f $X=6.84 $Y=0.38 $X2=0
+ $Y2=0
cc_820 N_A_27_47#_c_1377_n N_VGND_c_1548_n 0.0020257f $X=7.615 $Y=0.8 $X2=0
+ $Y2=0
cc_821 N_A_27_47#_c_1305_n N_VGND_c_1550_n 0.0209318f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_822 N_A_27_47#_c_1319_n N_VGND_c_1550_n 0.0020257f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_823 N_A_27_47#_c_1377_n N_VGND_c_1551_n 0.0020257f $X=7.615 $Y=0.8 $X2=0
+ $Y2=0
cc_824 N_A_27_47#_c_1381_n N_VGND_c_1551_n 0.0151813f $X=7.74 $Y=0.465 $X2=0
+ $Y2=0
cc_825 N_A_27_47#_c_1412_n N_VGND_c_1551_n 0.415017f $X=15.215 $Y=0.36 $X2=0
+ $Y2=0
cc_826 N_A_27_47#_c_1308_n N_VGND_c_1551_n 0.0172955f $X=15.34 $Y=0.465 $X2=0
+ $Y2=0
cc_827 N_A_27_47#_M1004_d N_VGND_c_1552_n 0.00209319f $X=0.135 $Y=0.235 $X2=0
+ $Y2=0
cc_828 N_A_27_47#_M1005_d N_VGND_c_1552_n 0.00215201f $X=1.065 $Y=0.235 $X2=0
+ $Y2=0
cc_829 N_A_27_47#_M1016_d N_VGND_c_1552_n 0.00215201f $X=2.005 $Y=0.235 $X2=0
+ $Y2=0
cc_830 N_A_27_47#_M1025_d N_VGND_c_1552_n 0.00215201f $X=2.945 $Y=0.235 $X2=0
+ $Y2=0
cc_831 N_A_27_47#_M1035_d N_VGND_c_1552_n 0.00215201f $X=3.885 $Y=0.235 $X2=0
+ $Y2=0
cc_832 N_A_27_47#_M1040_d N_VGND_c_1552_n 0.00215201f $X=4.825 $Y=0.235 $X2=0
+ $Y2=0
cc_833 N_A_27_47#_M1053_d N_VGND_c_1552_n 0.00215201f $X=5.765 $Y=0.235 $X2=0
+ $Y2=0
cc_834 N_A_27_47#_M1056_d N_VGND_c_1552_n 0.00215201f $X=6.705 $Y=0.235 $X2=0
+ $Y2=0
cc_835 N_A_27_47#_M1058_d N_VGND_c_1552_n 0.00215206f $X=7.645 $Y=0.235 $X2=0
+ $Y2=0
cc_836 N_A_27_47#_M1006_s N_VGND_c_1552_n 0.00255381f $X=8.535 $Y=0.235 $X2=0
+ $Y2=0
cc_837 N_A_27_47#_M1017_s N_VGND_c_1552_n 0.00215227f $X=9.525 $Y=0.235 $X2=0
+ $Y2=0
cc_838 N_A_27_47#_M1024_s N_VGND_c_1552_n 0.00215227f $X=10.465 $Y=0.235 $X2=0
+ $Y2=0
cc_839 N_A_27_47#_M1027_s N_VGND_c_1552_n 0.00255381f $X=11.355 $Y=0.235 $X2=0
+ $Y2=0
cc_840 N_A_27_47#_M1032_s N_VGND_c_1552_n 0.00215227f $X=12.345 $Y=0.235 $X2=0
+ $Y2=0
cc_841 N_A_27_47#_M1043_s N_VGND_c_1552_n 0.00215227f $X=13.285 $Y=0.235 $X2=0
+ $Y2=0
cc_842 N_A_27_47#_M1047_s N_VGND_c_1552_n 0.00215227f $X=14.225 $Y=0.235 $X2=0
+ $Y2=0
cc_843 N_A_27_47#_M1062_s N_VGND_c_1552_n 0.00209324f $X=15.165 $Y=0.235 $X2=0
+ $Y2=0
cc_844 N_A_27_47#_c_1305_n N_VGND_c_1552_n 0.0124017f $X=0.26 $Y=0.38 $X2=0
+ $Y2=0
cc_845 N_A_27_47#_c_1319_n N_VGND_c_1552_n 0.00880092f $X=1.035 $Y=0.8 $X2=0
+ $Y2=0
cc_846 N_A_27_47#_c_1325_n N_VGND_c_1552_n 0.0121968f $X=1.2 $Y=0.38 $X2=0 $Y2=0
cc_847 N_A_27_47#_c_1329_n N_VGND_c_1552_n 0.00880092f $X=1.975 $Y=0.8 $X2=0
+ $Y2=0
cc_848 N_A_27_47#_c_1333_n N_VGND_c_1552_n 0.0121968f $X=2.14 $Y=0.38 $X2=0
+ $Y2=0
cc_849 N_A_27_47#_c_1337_n N_VGND_c_1552_n 0.00880092f $X=2.915 $Y=0.8 $X2=0
+ $Y2=0
cc_850 N_A_27_47#_c_1341_n N_VGND_c_1552_n 0.0121968f $X=3.08 $Y=0.38 $X2=0
+ $Y2=0
cc_851 N_A_27_47#_c_1345_n N_VGND_c_1552_n 0.00880092f $X=3.855 $Y=0.8 $X2=0
+ $Y2=0
cc_852 N_A_27_47#_c_1349_n N_VGND_c_1552_n 0.0121968f $X=4.02 $Y=0.38 $X2=0
+ $Y2=0
cc_853 N_A_27_47#_c_1353_n N_VGND_c_1552_n 0.00880092f $X=4.795 $Y=0.8 $X2=0
+ $Y2=0
cc_854 N_A_27_47#_c_1357_n N_VGND_c_1552_n 0.0121968f $X=4.96 $Y=0.38 $X2=0
+ $Y2=0
cc_855 N_A_27_47#_c_1361_n N_VGND_c_1552_n 0.00880092f $X=5.735 $Y=0.8 $X2=0
+ $Y2=0
cc_856 N_A_27_47#_c_1365_n N_VGND_c_1552_n 0.0121968f $X=5.9 $Y=0.38 $X2=0 $Y2=0
cc_857 N_A_27_47#_c_1369_n N_VGND_c_1552_n 0.00880092f $X=6.675 $Y=0.8 $X2=0
+ $Y2=0
cc_858 N_A_27_47#_c_1373_n N_VGND_c_1552_n 0.0121968f $X=6.84 $Y=0.38 $X2=0
+ $Y2=0
cc_859 N_A_27_47#_c_1377_n N_VGND_c_1552_n 0.00880092f $X=7.615 $Y=0.8 $X2=0
+ $Y2=0
cc_860 N_A_27_47#_c_1381_n N_VGND_c_1552_n 0.0093992f $X=7.74 $Y=0.465 $X2=0
+ $Y2=0
cc_861 N_A_27_47#_c_1412_n N_VGND_c_1552_n 0.262938f $X=15.215 $Y=0.36 $X2=0
+ $Y2=0
cc_862 N_A_27_47#_c_1308_n N_VGND_c_1552_n 0.00960883f $X=15.34 $Y=0.465 $X2=0
+ $Y2=0
