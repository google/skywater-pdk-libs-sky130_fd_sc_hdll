* File: sky130_fd_sc_hdll__nor4bb_1.spice
* Created: Thu Aug 27 19:17:49 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__nor4bb_1.pex.spice"
.subckt sky130_fd_sc_hdll__nor4bb_1  VNB VPB C_N D_N B A VPWR Y VGND
* 
* VGND	VGND
* Y	Y
* VPWR	VPWR
* A	A
* B	B
* D_N	D_N
* C_N	C_N
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_C_N_M1000_g N_A_27_410#_M1000_s VNB NSHORT L=0.15 W=0.42
+ AD=0.06195 AS=0.1302 PD=0.715 PS=1.46 NRD=4.284 NRS=12.852 M=1 R=2.8
+ SA=75000.2 SB=75000.7 A=0.063 P=1.14 MULT=1
MM1002 N_A_216_93#_M1002_d N_D_N_M1002_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.42
+ AD=0.1281 AS=0.06195 PD=1.45 PS=0.715 NRD=11.424 NRS=0 M=1 R=2.8 SA=75000.7
+ SB=75000.2 A=0.063 P=1.14 MULT=1
MM1003 N_Y_M1003_d N_A_216_93#_M1003_g N_VGND_M1003_s VNB NSHORT L=0.15 W=0.65
+ AD=0.10725 AS=0.2015 PD=0.98 PS=1.92 NRD=0 NRS=8.304 M=1 R=4.33333 SA=75000.2
+ SB=75001.7 A=0.0975 P=1.6 MULT=1
MM1006 N_VGND_M1006_d N_A_27_410#_M1006_g N_Y_M1003_d VNB NSHORT L=0.15 W=0.65
+ AD=0.12025 AS=0.10725 PD=1.02 PS=0.98 NRD=2.76 NRS=10.152 M=1 R=4.33333
+ SA=75000.7 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1001 N_Y_M1001_d N_B_M1001_g N_VGND_M1006_d VNB NSHORT L=0.15 W=0.65
+ AD=0.08775 AS=0.12025 PD=0.92 PS=1.02 NRD=0 NRS=13.836 M=1 R=4.33333
+ SA=75001.2 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A_M1004_g N_Y_M1001_d VNB NSHORT L=0.15 W=0.65 AD=0.2015
+ AS=0.08775 PD=1.92 PS=0.92 NRD=8.304 NRS=0 M=1 R=4.33333 SA=75001.7 SB=75000.2
+ A=0.0975 P=1.6 MULT=1
MM1008 N_VPWR_M1008_d N_C_N_M1008_g N_A_27_410#_M1008_s VPB PHIGHVT L=0.18
+ W=0.42 AD=0.126812 AS=0.1134 PD=1.34 PS=1.38 NRD=2.3443 NRS=2.3443 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1009 N_A_216_93#_M1009_d N_D_N_M1009_g N_VPWR_M1008_d VPB PHIGHVT L=0.18
+ W=0.42 AD=0.1134 AS=0.126812 PD=1.38 PS=1.34 NRD=2.3443 NRS=115.816 M=1
+ R=2.33333 SA=90000.2 SB=90000.2 A=0.0756 P=1.2 MULT=1
MM1005 A_422_297# N_A_216_93#_M1005_g N_Y_M1005_s VPB PHIGHVT L=0.18 W=1 AD=0.15
+ AS=0.27 PD=1.3 PS=2.54 NRD=18.6953 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90001.6 A=0.18 P=2.36 MULT=1
MM1011 A_518_297# N_A_27_410#_M1011_g A_422_297# VPB PHIGHVT L=0.18 W=1 AD=0.17
+ AS=0.15 PD=1.34 PS=1.3 NRD=22.6353 NRS=18.6953 M=1 R=5.55556 SA=90000.7
+ SB=90001.2 A=0.18 P=2.36 MULT=1
MM1010 A_622_297# N_B_M1010_g A_518_297# VPB PHIGHVT L=0.18 W=1 AD=0.145 AS=0.17
+ PD=1.29 PS=1.34 NRD=17.7103 NRS=22.6353 M=1 R=5.55556 SA=90001.2 SB=90000.6
+ A=0.18 P=2.36 MULT=1
MM1007 N_VPWR_M1007_d N_A_M1007_g A_622_297# VPB PHIGHVT L=0.18 W=1 AD=0.27
+ AS=0.145 PD=2.54 PS=1.29 NRD=0.9653 NRS=17.7103 M=1 R=5.55556 SA=90001.6
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX12_noxref VNB VPB NWDIODE A=7.2546 P=12.25
pX13_noxref noxref_15 D_N D_N PROBETYPE=1
*
.include "sky130_fd_sc_hdll__nor4bb_1.pxi.spice"
*
.ends
*
*
