* File: sky130_fd_sc_hdll__a2bb2o_2.pxi.spice
* Created: Wed Sep  2 08:19:18 2020
* 
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_82_21# N_A_82_21#_M1013_d N_A_82_21#_M1007_s
+ N_A_82_21#_c_74_n N_A_82_21#_M1003_g N_A_82_21#_c_81_n N_A_82_21#_M1000_g
+ N_A_82_21#_c_75_n N_A_82_21#_M1011_g N_A_82_21#_c_82_n N_A_82_21#_M1010_g
+ N_A_82_21#_c_83_n N_A_82_21#_c_92_p N_A_82_21#_c_133_p N_A_82_21#_c_84_n
+ N_A_82_21#_c_85_n N_A_82_21#_c_86_n N_A_82_21#_c_76_n N_A_82_21#_c_77_n
+ N_A_82_21#_c_78_n N_A_82_21#_c_88_n N_A_82_21#_c_79_n N_A_82_21#_c_80_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_82_21#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%A1_N N_A1_N_c_189_n N_A1_N_M1008_g
+ N_A1_N_M1006_g A1_N A1_N PM_SKY130_FD_SC_HDLL__A2BB2O_2%A1_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%A2_N N_A2_N_c_224_n N_A2_N_M1002_g
+ N_A2_N_M1005_g A2_N PM_SKY130_FD_SC_HDLL__A2BB2O_2%A2_N
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_343_47# N_A_343_47#_M1006_d
+ N_A_343_47#_M1002_d N_A_343_47#_c_256_n N_A_343_47#_M1013_g
+ N_A_343_47#_c_257_n N_A_343_47#_c_261_n N_A_343_47#_c_262_n
+ N_A_343_47#_M1007_g N_A_343_47#_c_290_n N_A_343_47#_c_258_n
+ N_A_343_47#_c_259_n N_A_343_47#_c_263_n N_A_343_47#_c_264_n
+ N_A_343_47#_c_280_n PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_343_47#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%B2 N_B2_M1001_g N_B2_c_322_n N_B2_M1009_g B2
+ PM_SKY130_FD_SC_HDLL__A2BB2O_2%B2
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%B1 N_B1_M1012_g N_B1_c_360_n N_B1_c_361_n
+ N_B1_M1004_g B1 B1 B1 N_B1_c_359_n PM_SKY130_FD_SC_HDLL__A2BB2O_2%B1
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%VPWR N_VPWR_M1000_s N_VPWR_M1010_s
+ N_VPWR_M1009_d N_VPWR_c_389_n N_VPWR_c_390_n N_VPWR_c_391_n N_VPWR_c_392_n
+ VPWR VPWR N_VPWR_c_394_n N_VPWR_c_395_n N_VPWR_c_388_n N_VPWR_c_397_n
+ N_VPWR_c_398_n VPWR PM_SKY130_FD_SC_HDLL__A2BB2O_2%VPWR
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%X N_X_M1003_s N_X_M1000_d N_X_c_456_n
+ N_X_c_458_n N_X_c_454_n X X X N_X_c_470_n PM_SKY130_FD_SC_HDLL__A2BB2O_2%X
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_622_369# N_A_622_369#_M1007_d
+ N_A_622_369#_M1004_d N_A_622_369#_c_486_n N_A_622_369#_c_484_n
+ N_A_622_369#_c_485_n N_A_622_369#_c_501_n N_A_622_369#_c_496_n
+ PM_SKY130_FD_SC_HDLL__A2BB2O_2%A_622_369#
x_PM_SKY130_FD_SC_HDLL__A2BB2O_2%VGND N_VGND_M1003_d N_VGND_M1011_d
+ N_VGND_M1005_d N_VGND_M1012_d N_VGND_c_516_n N_VGND_c_517_n VGND VGND
+ N_VGND_c_519_n N_VGND_c_520_n N_VGND_c_521_n N_VGND_c_522_n N_VGND_c_523_n
+ N_VGND_c_524_n N_VGND_c_525_n VGND PM_SKY130_FD_SC_HDLL__A2BB2O_2%VGND
cc_1 VNB N_A_82_21#_c_74_n 0.0208267f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_2 VNB N_A_82_21#_c_75_n 0.0184072f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_3 VNB N_A_82_21#_c_76_n 0.0020092f $X=-0.19 $Y=-0.24 $X2=2.99 $Y2=1.895
cc_4 VNB N_A_82_21#_c_77_n 0.00127915f $X=-0.19 $Y=-0.24 $X2=3.195 $Y2=0.445
cc_5 VNB N_A_82_21#_c_78_n 0.00477711f $X=-0.19 $Y=-0.24 $X2=1 $Y2=1.16
cc_6 VNB N_A_82_21#_c_79_n 0.00975046f $X=-0.19 $Y=-0.24 $X2=3.195 $Y2=0.785
cc_7 VNB N_A_82_21#_c_80_n 0.0539915f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.202
cc_8 VNB N_A1_N_c_189_n 0.023739f $X=-0.19 $Y=-0.24 $X2=3.06 $Y2=0.235
cc_9 VNB N_A1_N_M1006_g 0.0336449f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_10 VNB A1_N 0.00825275f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.56
cc_11 VNB N_A2_N_c_224_n 0.0249656f $X=-0.19 $Y=-0.24 $X2=3.06 $Y2=0.235
cc_12 VNB N_A2_N_M1005_g 0.0314369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_13 VNB A2_N 0.00382657f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.56
cc_14 VNB N_A_343_47#_c_256_n 0.0195396f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.995
cc_15 VNB N_A_343_47#_c_257_n 0.0655469f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_16 VNB N_A_343_47#_c_258_n 0.0122742f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.325
cc_17 VNB N_A_343_47#_c_259_n 0.00732265f $X=-0.19 $Y=-0.24 $X2=1.11 $Y2=1.805
cc_18 VNB N_B2_M1001_g 0.0435654f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_19 VNB N_B2_c_322_n 0.00485315f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_20 VNB B2 0.0161759f $X=-0.19 $Y=-0.24 $X2=0.485 $Y2=0.56
cc_21 VNB N_B1_M1012_g 0.0351328f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_22 VNB B1 0.0274058f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.41
cc_23 VNB N_B1_c_359_n 0.0445339f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.985
cc_24 VNB N_VPWR_c_388_n 0.193827f $X=-0.19 $Y=-0.24 $X2=2.87 $Y2=2.285
cc_25 VNB N_X_c_454_n 0.00106626f $X=-0.19 $Y=-0.24 $X2=0.51 $Y2=1.985
cc_26 VNB N_VGND_c_516_n 0.0169736f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.995
cc_27 VNB N_VGND_c_517_n 0.0192442f $X=-0.19 $Y=-0.24 $X2=0.955 $Y2=0.56
cc_28 VNB VGND 0.0113688f $X=-0.19 $Y=-0.24 $X2=0.98 $Y2=1.985
cc_29 VNB N_VGND_c_519_n 0.0164623f $X=-0.19 $Y=-0.24 $X2=1.22 $Y2=1.89
cc_30 VNB N_VGND_c_520_n 0.0287369f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_31 VNB N_VGND_c_521_n 0.0110256f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_32 VNB N_VGND_c_522_n 0.017867f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_33 VNB N_VGND_c_523_n 0.0178809f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_34 VNB N_VGND_c_524_n 0.242525f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_35 VNB N_VGND_c_525_n 0.00874672f $X=-0.19 $Y=-0.24 $X2=0 $Y2=0
cc_36 VPB N_A_82_21#_c_81_n 0.0197071f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_37 VPB N_A_82_21#_c_82_n 0.0177824f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_38 VPB N_A_82_21#_c_83_n 0.00112304f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.805
cc_39 VPB N_A_82_21#_c_84_n 6.97853e-19 $X=-0.19 $Y=1.305 $X2=1.75 $Y2=2.2
cc_40 VPB N_A_82_21#_c_85_n 0.0194012f $X=-0.19 $Y=1.305 $X2=2.64 $Y2=2.285
cc_41 VPB N_A_82_21#_c_86_n 0.00289098f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=2.285
cc_42 VPB N_A_82_21#_c_76_n 0.00452542f $X=-0.19 $Y=1.305 $X2=2.99 $Y2=1.895
cc_43 VPB N_A_82_21#_c_88_n 0.00496563f $X=-0.19 $Y=1.305 $X2=2.785 $Y2=2.275
cc_44 VPB N_A_82_21#_c_80_n 0.0282372f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_45 VPB N_A1_N_c_189_n 0.0256674f $X=-0.19 $Y=1.305 $X2=3.06 $Y2=0.235
cc_46 VPB A1_N 0.00272922f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_47 VPB N_A2_N_c_224_n 0.0289618f $X=-0.19 $Y=1.305 $X2=3.06 $Y2=0.235
cc_48 VPB A2_N 0.00384954f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_49 VPB N_A_343_47#_c_257_n 0.0264053f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_50 VPB N_A_343_47#_c_261_n 0.0155514f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_51 VPB N_A_343_47#_c_262_n 0.027906f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_52 VPB N_A_343_47#_c_263_n 0.0103697f $X=-0.19 $Y=1.305 $X2=1.64 $Y2=1.89
cc_53 VPB N_A_343_47#_c_264_n 0.00197279f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=2.285
cc_54 VPB N_B2_c_322_n 0.0518635f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_55 VPB B2 0.00733785f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_56 VPB N_B1_c_360_n 0.023488f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_57 VPB N_B1_c_361_n 0.0301327f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.995
cc_58 VPB B1 0.0220074f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_59 VPB N_B1_c_359_n 0.00765335f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.985
cc_60 VPB N_VPWR_c_389_n 0.00921986f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_61 VPB N_VPWR_c_390_n 0.00242779f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.41
cc_62 VPB N_VPWR_c_391_n 0.0574928f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.325
cc_63 VPB N_VPWR_c_392_n 0.00359728f $X=-0.19 $Y=1.305 $X2=1.11 $Y2=1.805
cc_64 VPB VPWR 0.0113429f $X=-0.19 $Y=1.305 $X2=1.64 $Y2=1.89
cc_65 VPB N_VPWR_c_394_n 0.0164231f $X=-0.19 $Y=1.305 $X2=1.86 $Y2=2.285
cc_66 VPB N_VPWR_c_395_n 0.0201535f $X=-0.19 $Y=1.305 $X2=2.785 $Y2=2.275
cc_67 VPB N_VPWR_c_388_n 0.0640558f $X=-0.19 $Y=1.305 $X2=2.87 $Y2=2.285
cc_68 VPB N_VPWR_c_397_n 0.005797f $X=-0.19 $Y=1.305 $X2=0.98 $Y2=1.202
cc_69 VPB N_VPWR_c_398_n 0.00853175f $X=-0.19 $Y=1.305 $X2=0 $Y2=0
cc_70 VPB N_X_c_454_n 0.00108723f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.985
cc_71 VPB N_A_622_369#_c_484_n 0.00628852f $X=-0.19 $Y=1.305 $X2=0.485 $Y2=0.56
cc_72 VPB N_A_622_369#_c_485_n 0.00156978f $X=-0.19 $Y=1.305 $X2=0.51 $Y2=1.41
cc_73 N_A_82_21#_c_82_n N_A1_N_c_189_n 0.0176388f $X=0.98 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_74 N_A_82_21#_c_83_n N_A1_N_c_189_n 0.00473761f $X=1.11 $Y=1.805 $X2=-0.19
+ $Y2=-0.24
cc_75 N_A_82_21#_c_92_p N_A1_N_c_189_n 0.0134648f $X=1.64 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_76 N_A_82_21#_c_84_n N_A1_N_c_189_n 0.00668216f $X=1.75 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_77 N_A_82_21#_c_86_n N_A1_N_c_189_n 0.00286009f $X=1.86 $Y=2.285 $X2=-0.19
+ $Y2=-0.24
cc_78 N_A_82_21#_c_78_n N_A1_N_c_189_n 0.00205895f $X=1 $Y=1.16 $X2=-0.19
+ $Y2=-0.24
cc_79 N_A_82_21#_c_80_n N_A1_N_c_189_n 0.0227547f $X=0.98 $Y=1.202 $X2=-0.19
+ $Y2=-0.24
cc_80 N_A_82_21#_c_75_n N_A1_N_M1006_g 0.0161481f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_81 N_A_82_21#_c_82_n A1_N 6.26543e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_82 N_A_82_21#_c_92_p A1_N 0.0186991f $X=1.64 $Y=1.89 $X2=0 $Y2=0
cc_83 N_A_82_21#_c_78_n A1_N 0.040211f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_84 N_A_82_21#_c_80_n A1_N 6.22435e-19 $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_85 N_A_82_21#_c_92_p N_A2_N_c_224_n 0.00312323f $X=1.64 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_86 N_A_82_21#_c_84_n N_A2_N_c_224_n 0.00534531f $X=1.75 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_87 N_A_82_21#_c_85_n N_A2_N_c_224_n 0.0136956f $X=2.64 $Y=2.285 $X2=-0.19
+ $Y2=-0.24
cc_88 N_A_82_21#_c_88_n N_A2_N_c_224_n 0.00775922f $X=2.785 $Y=2.275 $X2=-0.19
+ $Y2=-0.24
cc_89 N_A_82_21#_c_79_n N_A2_N_M1005_g 2.0633e-19 $X=3.195 $Y=0.785 $X2=0 $Y2=0
cc_90 N_A_82_21#_c_77_n N_A_343_47#_c_256_n 5.08356e-19 $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_91 N_A_82_21#_c_79_n N_A_343_47#_c_256_n 0.00605921f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_92 N_A_82_21#_c_76_n N_A_343_47#_c_257_n 0.0235829f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_93 N_A_82_21#_c_88_n N_A_343_47#_c_257_n 0.00602719f $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_94 N_A_82_21#_c_79_n N_A_343_47#_c_257_n 0.00615575f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_95 N_A_82_21#_c_76_n N_A_343_47#_c_261_n 0.00877171f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_96 N_A_82_21#_c_76_n N_A_343_47#_c_262_n 0.00972423f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_97 N_A_82_21#_c_88_n N_A_343_47#_c_262_n 0.0142243f $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_98 N_A_82_21#_c_77_n N_A_343_47#_c_258_n 0.0020691f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_99 N_A_82_21#_c_79_n N_A_343_47#_c_258_n 0.0106477f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_100 N_A_82_21#_c_85_n N_A_343_47#_c_263_n 0.0110871f $X=2.64 $Y=2.285 $X2=0
+ $Y2=0
cc_101 N_A_82_21#_c_76_n N_A_343_47#_c_263_n 0.0139127f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_102 N_A_82_21#_c_88_n N_A_343_47#_c_263_n 0.00605907f $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_103 N_A_82_21#_c_76_n N_A_343_47#_c_264_n 0.0474799f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_104 N_A_82_21#_c_79_n N_A_343_47#_c_264_n 0.00317388f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_105 N_A_82_21#_c_92_p N_A_343_47#_c_280_n 0.0051555f $X=1.64 $Y=1.89 $X2=0
+ $Y2=0
cc_106 N_A_82_21#_c_85_n N_A_343_47#_c_280_n 0.00805606f $X=2.64 $Y=2.285 $X2=0
+ $Y2=0
cc_107 N_A_82_21#_c_76_n N_A_343_47#_c_280_n 0.00510251f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_108 N_A_82_21#_c_88_n N_A_343_47#_c_280_n 5.4232e-19 $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_109 N_A_82_21#_c_76_n N_B2_M1001_g 0.00431132f $X=2.99 $Y=1.895 $X2=0 $Y2=0
cc_110 N_A_82_21#_c_77_n N_B2_M1001_g 0.00111676f $X=3.195 $Y=0.445 $X2=0 $Y2=0
cc_111 N_A_82_21#_c_79_n N_B2_M1001_g 0.00474495f $X=3.195 $Y=0.785 $X2=0 $Y2=0
cc_112 N_A_82_21#_c_76_n N_B2_c_322_n 0.0011701f $X=2.99 $Y=1.895 $X2=0 $Y2=0
cc_113 N_A_82_21#_c_76_n B2 0.0423355f $X=2.99 $Y=1.895 $X2=0 $Y2=0
cc_114 N_A_82_21#_c_83_n N_VPWR_M1010_s 0.00380992f $X=1.11 $Y=1.805 $X2=0 $Y2=0
cc_115 N_A_82_21#_c_92_p N_VPWR_M1010_s 0.0122086f $X=1.64 $Y=1.89 $X2=0 $Y2=0
cc_116 N_A_82_21#_c_133_p N_VPWR_M1010_s 0.00120001f $X=1.22 $Y=1.89 $X2=0 $Y2=0
cc_117 N_A_82_21#_c_81_n N_VPWR_c_389_n 6.49455e-19 $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_118 N_A_82_21#_c_82_n N_VPWR_c_389_n 0.0111791f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_119 N_A_82_21#_c_92_p N_VPWR_c_389_n 0.00862919f $X=1.64 $Y=1.89 $X2=0 $Y2=0
cc_120 N_A_82_21#_c_133_p N_VPWR_c_389_n 0.00918694f $X=1.22 $Y=1.89 $X2=0 $Y2=0
cc_121 N_A_82_21#_c_86_n N_VPWR_c_389_n 0.00886738f $X=1.86 $Y=2.285 $X2=0 $Y2=0
cc_122 N_A_82_21#_c_92_p N_VPWR_c_391_n 0.00310724f $X=1.64 $Y=1.89 $X2=0 $Y2=0
cc_123 N_A_82_21#_c_85_n N_VPWR_c_391_n 0.0314683f $X=2.64 $Y=2.285 $X2=0 $Y2=0
cc_124 N_A_82_21#_c_86_n N_VPWR_c_391_n 0.00969682f $X=1.86 $Y=2.285 $X2=0 $Y2=0
cc_125 N_A_82_21#_c_88_n N_VPWR_c_391_n 0.0178604f $X=2.785 $Y=2.275 $X2=0 $Y2=0
cc_126 N_A_82_21#_c_81_n N_VPWR_c_394_n 0.00590121f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_127 N_A_82_21#_c_82_n N_VPWR_c_394_n 0.00427505f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_128 N_A_82_21#_M1007_s N_VPWR_c_388_n 0.00243299f $X=2.66 $Y=1.845 $X2=0
+ $Y2=0
cc_129 N_A_82_21#_c_81_n N_VPWR_c_388_n 0.0107882f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_130 N_A_82_21#_c_82_n N_VPWR_c_388_n 0.00740765f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_131 N_A_82_21#_c_92_p N_VPWR_c_388_n 0.00737713f $X=1.64 $Y=1.89 $X2=0 $Y2=0
cc_132 N_A_82_21#_c_133_p N_VPWR_c_388_n 0.00110043f $X=1.22 $Y=1.89 $X2=0 $Y2=0
cc_133 N_A_82_21#_c_85_n N_VPWR_c_388_n 0.0273188f $X=2.64 $Y=2.285 $X2=0 $Y2=0
cc_134 N_A_82_21#_c_86_n N_VPWR_c_388_n 0.00800038f $X=1.86 $Y=2.285 $X2=0 $Y2=0
cc_135 N_A_82_21#_c_88_n N_VPWR_c_388_n 0.0145966f $X=2.785 $Y=2.275 $X2=0 $Y2=0
cc_136 N_A_82_21#_c_81_n N_VPWR_c_398_n 0.00680281f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_137 N_A_82_21#_c_74_n N_X_c_456_n 0.00232185f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_138 N_A_82_21#_c_80_n N_X_c_456_n 0.00190599f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_139 N_A_82_21#_c_81_n N_X_c_458_n 0.00263447f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_140 N_A_82_21#_c_82_n N_X_c_458_n 0.00866396f $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_141 N_A_82_21#_c_83_n N_X_c_458_n 0.0208954f $X=1.11 $Y=1.805 $X2=0 $Y2=0
cc_142 N_A_82_21#_c_80_n N_X_c_458_n 0.0037632f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_143 N_A_82_21#_c_74_n N_X_c_454_n 0.00573813f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_144 N_A_82_21#_c_81_n N_X_c_454_n 0.00359097f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_145 N_A_82_21#_c_75_n N_X_c_454_n 0.00425752f $X=0.955 $Y=0.995 $X2=0 $Y2=0
cc_146 N_A_82_21#_c_82_n N_X_c_454_n 8.33442e-19 $X=0.98 $Y=1.41 $X2=0 $Y2=0
cc_147 N_A_82_21#_c_83_n N_X_c_454_n 0.0108589f $X=1.11 $Y=1.805 $X2=0 $Y2=0
cc_148 N_A_82_21#_c_78_n N_X_c_454_n 0.02387f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_149 N_A_82_21#_c_80_n N_X_c_454_n 0.0352171f $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_150 N_A_82_21#_c_74_n X 0.00604588f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_151 N_A_82_21#_c_81_n N_X_c_470_n 0.0134485f $X=0.51 $Y=1.41 $X2=0 $Y2=0
cc_152 N_A_82_21#_c_133_p N_X_c_470_n 0.0139285f $X=1.22 $Y=1.89 $X2=0 $Y2=0
cc_153 N_A_82_21#_c_92_p A_341_297# 0.00463816f $X=1.64 $Y=1.89 $X2=-0.19
+ $Y2=-0.24
cc_154 N_A_82_21#_c_84_n A_341_297# 0.00169863f $X=1.75 $Y=2.2 $X2=-0.19
+ $Y2=-0.24
cc_155 N_A_82_21#_c_88_n N_A_622_369#_c_486_n 0.0117549f $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_156 N_A_82_21#_c_76_n N_A_622_369#_c_485_n 0.00449826f $X=2.99 $Y=1.895 $X2=0
+ $Y2=0
cc_157 N_A_82_21#_c_88_n N_A_622_369#_c_485_n 0.0087494f $X=2.785 $Y=2.275 $X2=0
+ $Y2=0
cc_158 N_A_82_21#_c_74_n N_VGND_c_519_n 0.00533769f $X=0.485 $Y=0.995 $X2=0
+ $Y2=0
cc_159 N_A_82_21#_c_75_n N_VGND_c_519_n 0.00468308f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_160 N_A_82_21#_c_77_n N_VGND_c_520_n 0.0110645f $X=3.195 $Y=0.445 $X2=0 $Y2=0
cc_161 N_A_82_21#_c_79_n N_VGND_c_520_n 0.00326385f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_162 N_A_82_21#_c_74_n N_VGND_c_521_n 6.4445e-19 $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_163 N_A_82_21#_c_75_n N_VGND_c_521_n 0.00892418f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_164 N_A_82_21#_c_78_n N_VGND_c_521_n 0.00749638f $X=1 $Y=1.16 $X2=0 $Y2=0
cc_165 N_A_82_21#_c_80_n N_VGND_c_521_n 7.89286e-19 $X=0.98 $Y=1.202 $X2=0 $Y2=0
cc_166 N_A_82_21#_M1013_d N_VGND_c_524_n 0.00413042f $X=3.06 $Y=0.235 $X2=0
+ $Y2=0
cc_167 N_A_82_21#_c_74_n N_VGND_c_524_n 0.0104682f $X=0.485 $Y=0.995 $X2=0 $Y2=0
cc_168 N_A_82_21#_c_75_n N_VGND_c_524_n 0.00809956f $X=0.955 $Y=0.995 $X2=0
+ $Y2=0
cc_169 N_A_82_21#_c_77_n N_VGND_c_524_n 0.00640047f $X=3.195 $Y=0.445 $X2=0
+ $Y2=0
cc_170 N_A_82_21#_c_79_n N_VGND_c_524_n 0.00521813f $X=3.195 $Y=0.785 $X2=0
+ $Y2=0
cc_171 N_A_82_21#_c_74_n N_VGND_c_525_n 0.00408879f $X=0.485 $Y=0.995 $X2=0
+ $Y2=0
cc_172 N_A1_N_c_189_n N_A2_N_c_224_n 0.0713926f $X=1.615 $Y=1.41 $X2=-0.19
+ $Y2=-0.24
cc_173 A1_N N_A2_N_c_224_n 0.00732684f $X=1.535 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_174 N_A1_N_M1006_g N_A2_N_M1005_g 0.0199256f $X=1.64 $Y=0.445 $X2=0 $Y2=0
cc_175 N_A1_N_c_189_n A2_N 3.54483e-19 $X=1.615 $Y=1.41 $X2=0 $Y2=0
cc_176 A1_N A2_N 0.0304754f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_177 N_A1_N_M1006_g N_A_343_47#_c_259_n 0.00547454f $X=1.64 $Y=0.445 $X2=0
+ $Y2=0
cc_178 A1_N N_A_343_47#_c_259_n 0.00450064f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_179 A1_N N_A_343_47#_c_280_n 0.00310541f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_180 A1_N N_VPWR_M1010_s 0.00160587f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_181 N_A1_N_c_189_n N_VPWR_c_391_n 0.00288394f $X=1.615 $Y=1.41 $X2=0 $Y2=0
cc_182 N_A1_N_c_189_n N_VPWR_c_388_n 0.00364146f $X=1.615 $Y=1.41 $X2=0 $Y2=0
cc_183 A1_N A_341_297# 0.00213836f $X=1.535 $Y=1.105 $X2=-0.19 $Y2=-0.24
cc_184 N_A1_N_c_189_n N_VGND_c_521_n 0.0018495f $X=1.615 $Y=1.41 $X2=0 $Y2=0
cc_185 N_A1_N_M1006_g N_VGND_c_521_n 0.00543324f $X=1.64 $Y=0.445 $X2=0 $Y2=0
cc_186 A1_N N_VGND_c_521_n 0.00129799f $X=1.535 $Y=1.105 $X2=0 $Y2=0
cc_187 N_A1_N_M1006_g N_VGND_c_522_n 0.00585385f $X=1.64 $Y=0.445 $X2=0 $Y2=0
cc_188 N_A1_N_M1006_g N_VGND_c_523_n 6.07118e-19 $X=1.64 $Y=0.445 $X2=0 $Y2=0
cc_189 N_A1_N_M1006_g N_VGND_c_524_n 0.0114959f $X=1.64 $Y=0.445 $X2=0 $Y2=0
cc_190 N_A2_N_c_224_n N_A_343_47#_c_257_n 0.0233422f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_191 N_A2_N_M1005_g N_A_343_47#_c_257_n 0.0103075f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_192 A2_N N_A_343_47#_c_257_n 0.00279244f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_193 N_A2_N_M1005_g N_A_343_47#_c_290_n 0.00397472f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_194 N_A2_N_c_224_n N_A_343_47#_c_258_n 0.00300425f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_195 N_A2_N_M1005_g N_A_343_47#_c_258_n 0.0126745f $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_196 A2_N N_A_343_47#_c_258_n 0.0262975f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_197 N_A2_N_c_224_n N_A_343_47#_c_259_n 4.43981e-19 $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_198 N_A2_N_c_224_n N_A_343_47#_c_264_n 0.00323675f $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_199 N_A2_N_M1005_g N_A_343_47#_c_264_n 9.47693e-19 $X=2.11 $Y=0.445 $X2=0
+ $Y2=0
cc_200 A2_N N_A_343_47#_c_264_n 0.025075f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_201 N_A2_N_c_224_n N_A_343_47#_c_280_n 5.79699e-19 $X=2.025 $Y=1.41 $X2=0
+ $Y2=0
cc_202 A2_N N_A_343_47#_c_280_n 0.0132635f $X=1.995 $Y=1.105 $X2=0 $Y2=0
cc_203 N_A2_N_c_224_n N_VPWR_c_391_n 7.74976e-19 $X=2.025 $Y=1.41 $X2=0 $Y2=0
cc_204 N_A2_N_M1005_g N_VGND_c_522_n 0.00341689f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_205 N_A2_N_M1005_g N_VGND_c_523_n 0.00913044f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_206 N_A2_N_M1005_g N_VGND_c_524_n 0.00416126f $X=2.11 $Y=0.445 $X2=0 $Y2=0
cc_207 N_A_343_47#_c_256_n N_B2_M1001_g 0.0249681f $X=2.985 $Y=0.765 $X2=0 $Y2=0
cc_208 N_A_343_47#_c_257_n N_B2_M1001_g 0.0184608f $X=3.02 $Y=1.435 $X2=0 $Y2=0
cc_209 N_A_343_47#_c_261_n N_B2_c_322_n 0.0240785f $X=3.02 $Y=1.67 $X2=0 $Y2=0
cc_210 N_A_343_47#_c_262_n N_B2_c_322_n 0.018501f $X=3.02 $Y=1.77 $X2=0 $Y2=0
cc_211 N_A_343_47#_c_257_n B2 0.00384201f $X=3.02 $Y=1.435 $X2=0 $Y2=0
cc_212 N_A_343_47#_c_262_n N_VPWR_c_391_n 0.00523952f $X=3.02 $Y=1.77 $X2=0
+ $Y2=0
cc_213 N_A_343_47#_c_262_n N_VPWR_c_388_n 0.00858269f $X=3.02 $Y=1.77 $X2=0
+ $Y2=0
cc_214 N_A_343_47#_c_262_n N_A_622_369#_c_486_n 0.00159931f $X=3.02 $Y=1.77
+ $X2=0 $Y2=0
cc_215 N_A_343_47#_c_262_n N_A_622_369#_c_485_n 0.00122308f $X=3.02 $Y=1.77
+ $X2=0 $Y2=0
cc_216 N_A_343_47#_c_258_n N_VGND_M1005_d 0.00182057f $X=2.54 $Y=0.74 $X2=0
+ $Y2=0
cc_217 N_A_343_47#_c_256_n N_VGND_c_520_n 0.00434414f $X=2.985 $Y=0.765 $X2=0
+ $Y2=0
cc_218 N_A_343_47#_c_290_n N_VGND_c_522_n 0.011459f $X=1.85 $Y=0.445 $X2=0 $Y2=0
cc_219 N_A_343_47#_c_258_n N_VGND_c_522_n 0.00361022f $X=2.54 $Y=0.74 $X2=0
+ $Y2=0
cc_220 N_A_343_47#_c_256_n N_VGND_c_523_n 0.00509285f $X=2.985 $Y=0.765 $X2=0
+ $Y2=0
cc_221 N_A_343_47#_c_257_n N_VGND_c_523_n 0.00780208f $X=3.02 $Y=1.435 $X2=0
+ $Y2=0
cc_222 N_A_343_47#_c_290_n N_VGND_c_523_n 0.0147362f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_223 N_A_343_47#_c_258_n N_VGND_c_523_n 0.0414636f $X=2.54 $Y=0.74 $X2=0 $Y2=0
cc_224 N_A_343_47#_M1006_d N_VGND_c_524_n 0.00472584f $X=1.715 $Y=0.235 $X2=0
+ $Y2=0
cc_225 N_A_343_47#_c_256_n N_VGND_c_524_n 0.00714603f $X=2.985 $Y=0.765 $X2=0
+ $Y2=0
cc_226 N_A_343_47#_c_290_n N_VGND_c_524_n 0.00644035f $X=1.85 $Y=0.445 $X2=0
+ $Y2=0
cc_227 N_A_343_47#_c_258_n N_VGND_c_524_n 0.0080021f $X=2.54 $Y=0.74 $X2=0 $Y2=0
cc_228 N_B2_M1001_g N_B1_M1012_g 0.0401131f $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_229 N_B2_c_322_n N_B1_c_360_n 0.00714349f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_230 N_B2_c_322_n N_B1_c_361_n 0.0223311f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_231 N_B2_M1001_g B1 3.76865e-19 $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_232 N_B2_c_322_n B1 2.93445e-19 $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_233 B2 B1 0.0309756f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_234 N_B2_M1001_g N_B1_c_359_n 0.00392512f $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_235 N_B2_c_322_n N_B1_c_359_n 0.0162779f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_236 B2 N_B1_c_359_n 0.00608499f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_237 N_B2_c_322_n N_VPWR_c_390_n 0.00499199f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_238 N_B2_c_322_n N_VPWR_c_391_n 0.00514401f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_239 N_B2_c_322_n N_VPWR_c_388_n 0.00690865f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_240 N_B2_c_322_n N_A_622_369#_c_486_n 0.00515995f $X=3.525 $Y=1.77 $X2=0
+ $Y2=0
cc_241 N_B2_c_322_n N_A_622_369#_c_484_n 0.0112023f $X=3.525 $Y=1.77 $X2=0 $Y2=0
cc_242 B2 N_A_622_369#_c_484_n 0.023014f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_243 N_B2_c_322_n N_A_622_369#_c_485_n 0.00300185f $X=3.525 $Y=1.77 $X2=0
+ $Y2=0
cc_244 B2 N_A_622_369#_c_485_n 0.0130284f $X=3.365 $Y=1.445 $X2=0 $Y2=0
cc_245 N_B2_c_322_n N_A_622_369#_c_496_n 0.00222466f $X=3.525 $Y=1.77 $X2=0
+ $Y2=0
cc_246 N_B2_M1001_g N_VGND_c_517_n 0.00221199f $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_247 N_B2_M1001_g N_VGND_c_520_n 0.00585385f $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_248 N_B2_M1001_g N_VGND_c_524_n 0.0109909f $X=3.405 $Y=0.445 $X2=0 $Y2=0
cc_249 N_B1_c_361_n N_VPWR_c_390_n 0.00894644f $X=3.995 $Y=1.77 $X2=0 $Y2=0
cc_250 N_B1_c_361_n N_VPWR_c_395_n 0.00464801f $X=3.995 $Y=1.77 $X2=0 $Y2=0
cc_251 N_B1_c_361_n N_VPWR_c_388_n 0.00643063f $X=3.995 $Y=1.77 $X2=0 $Y2=0
cc_252 N_B1_c_361_n N_A_622_369#_c_486_n 7.29534e-19 $X=3.995 $Y=1.77 $X2=0
+ $Y2=0
cc_253 N_B1_c_361_n N_A_622_369#_c_484_n 0.0208762f $X=3.995 $Y=1.77 $X2=0 $Y2=0
cc_254 B1 N_A_622_369#_c_484_n 0.0202805f $X=4.245 $Y=0.765 $X2=0 $Y2=0
cc_255 N_B1_c_359_n N_A_622_369#_c_484_n 0.0030871f $X=3.995 $Y=1.16 $X2=0 $Y2=0
cc_256 N_B1_c_361_n N_A_622_369#_c_501_n 0.00580049f $X=3.995 $Y=1.77 $X2=0
+ $Y2=0
cc_257 B1 N_VGND_c_516_n 0.00157103f $X=4.245 $Y=0.765 $X2=0 $Y2=0
cc_258 N_B1_M1012_g N_VGND_c_517_n 0.0162078f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_259 B1 N_VGND_c_517_n 0.0244597f $X=4.245 $Y=0.765 $X2=0 $Y2=0
cc_260 N_B1_c_359_n N_VGND_c_517_n 0.00489451f $X=3.995 $Y=1.16 $X2=0 $Y2=0
cc_261 N_B1_M1012_g N_VGND_c_520_n 0.00407992f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_262 N_B1_M1012_g N_VGND_c_524_n 0.00719726f $X=3.875 $Y=0.445 $X2=0 $Y2=0
cc_263 B1 N_VGND_c_524_n 0.00385325f $X=4.245 $Y=0.765 $X2=0 $Y2=0
cc_264 N_VPWR_c_388_n N_X_M1000_d 0.00444633f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_265 N_VPWR_c_398_n N_X_c_454_n 0.0746891f $X=0.27 $Y=1.64 $X2=0 $Y2=0
cc_266 N_VPWR_c_389_n N_X_c_470_n 0.0179342f $X=1.215 $Y=2.32 $X2=0 $Y2=0
cc_267 N_VPWR_c_394_n N_X_c_470_n 0.0191629f $X=1 $Y=2.72 $X2=0 $Y2=0
cc_268 N_VPWR_c_388_n N_X_c_470_n 0.0113307f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_269 N_VPWR_c_388_n N_A_622_369#_M1007_d 0.00310751f $X=4.37 $Y=2.72 $X2=-0.19
+ $Y2=-0.24
cc_270 N_VPWR_c_388_n N_A_622_369#_M1004_d 0.00388786f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_271 N_VPWR_c_390_n N_A_622_369#_c_486_n 0.00474967f $X=3.76 $Y=2.34 $X2=0
+ $Y2=0
cc_272 N_VPWR_M1009_d N_A_622_369#_c_484_n 0.00178166f $X=3.615 $Y=1.845 $X2=0
+ $Y2=0
cc_273 N_VPWR_c_390_n N_A_622_369#_c_484_n 0.0147753f $X=3.76 $Y=2.34 $X2=0
+ $Y2=0
cc_274 N_VPWR_c_391_n N_A_622_369#_c_484_n 0.00267292f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_275 N_VPWR_c_395_n N_A_622_369#_c_484_n 0.00265818f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_276 N_VPWR_c_388_n N_A_622_369#_c_484_n 0.0110849f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_277 N_VPWR_c_390_n N_A_622_369#_c_501_n 0.0171884f $X=3.76 $Y=2.34 $X2=0
+ $Y2=0
cc_278 N_VPWR_c_395_n N_A_622_369#_c_501_n 0.0117479f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_279 N_VPWR_c_388_n N_A_622_369#_c_501_n 0.00645703f $X=4.37 $Y=2.72 $X2=0
+ $Y2=0
cc_280 N_VPWR_c_390_n N_A_622_369#_c_496_n 0.0105122f $X=3.76 $Y=2.34 $X2=0
+ $Y2=0
cc_281 N_VPWR_c_391_n N_A_622_369#_c_496_n 0.014461f $X=3.675 $Y=2.72 $X2=0
+ $Y2=0
cc_282 N_VPWR_c_388_n N_A_622_369#_c_496_n 0.011831f $X=4.37 $Y=2.72 $X2=0 $Y2=0
cc_283 N_VPWR_c_398_n N_VGND_c_525_n 0.00726759f $X=0.27 $Y=1.64 $X2=0 $Y2=0
cc_284 X N_VGND_c_519_n 0.0189588f $X=0.635 $Y=0.425 $X2=0 $Y2=0
cc_285 N_X_M1003_s N_VGND_c_524_n 0.00434007f $X=0.56 $Y=0.235 $X2=0 $Y2=0
cc_286 X N_VGND_c_524_n 0.0114966f $X=0.635 $Y=0.425 $X2=0 $Y2=0
cc_287 X N_VGND_c_525_n 0.0263896f $X=0.635 $Y=0.425 $X2=0 $Y2=0
cc_288 N_VGND_c_524_n A_696_47# 0.0136786f $X=4.37 $Y=0 $X2=-0.19 $Y2=-0.24
