* File: sky130_fd_sc_hdll__a21o_1.spice
* Created: Thu Aug 27 18:52:43 2020
* Program "Calibre xRC"
* Version "v2018.4_34.26"
* 
.include "sky130_fd_sc_hdll__a21o_1.pex.spice"
.subckt sky130_fd_sc_hdll__a21o_1  VNB VPB B1 A1 A2 X VPWR VGND
* 
* VGND	VGND
* VPWR	VPWR
* X	X
* A2	A2
* A1	A1
* B1	B1
* VPB	VPB
* VNB	VNB
MM1000 N_VGND_M1000_d N_A_81_21#_M1000_g N_X_M1000_s VNB NSHORT L=0.15 W=0.65
+ AD=0.28925 AS=0.169 PD=1.54 PS=1.82 NRD=24.912 NRS=0 M=1 R=4.33333 SA=75000.2
+ SB=75002.2 A=0.0975 P=1.6 MULT=1
MM1001 N_A_81_21#_M1001_d N_B1_M1001_g N_VGND_M1000_d VNB NSHORT L=0.15 W=0.65
+ AD=0.108875 AS=0.28925 PD=0.985 PS=1.54 NRD=0 NRS=24.912 M=1 R=4.33333
+ SA=75001.2 SB=75001.2 A=0.0975 P=1.6 MULT=1
MM1007 A_416_47# N_A1_M1007_g N_A_81_21#_M1001_d VNB NSHORT L=0.15 W=0.65
+ AD=0.091 AS=0.108875 PD=0.93 PS=0.985 NRD=15.684 NRS=11.076 M=1 R=4.33333
+ SA=75001.7 SB=75000.7 A=0.0975 P=1.6 MULT=1
MM1004 N_VGND_M1004_d N_A2_M1004_g A_416_47# VNB NSHORT L=0.15 W=0.65 AD=0.20475
+ AS=0.091 PD=1.93 PS=0.93 NRD=9.228 NRS=15.684 M=1 R=4.33333 SA=75002.1
+ SB=75000.2 A=0.0975 P=1.6 MULT=1
MM1003 N_VPWR_M1003_d N_A_81_21#_M1003_g N_X_M1003_s VPB PHIGHVT L=0.18 W=1
+ AD=0.27 AS=0.27 PD=2.54 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556 SA=90000.2
+ SB=90000.2 A=0.18 P=2.36 MULT=1
MM1005 N_A_317_297#_M1005_d N_B1_M1005_g N_A_81_21#_M1005_s VPB PHIGHVT L=0.18
+ W=1 AD=0.1525 AS=0.27 PD=1.305 PS=2.54 NRD=0.9653 NRS=0.9653 M=1 R=5.55556
+ SA=90000.2 SB=90001.1 A=0.18 P=2.36 MULT=1
MM1002 N_VPWR_M1002_d N_A1_M1002_g N_A_317_297#_M1005_d VPB PHIGHVT L=0.18 W=1
+ AD=0.15 AS=0.1525 PD=1.3 PS=1.305 NRD=1.9503 NRS=3.9203 M=1 R=5.55556
+ SA=90000.7 SB=90000.7 A=0.18 P=2.36 MULT=1
MM1006 N_A_317_297#_M1006_d N_A2_M1006_g N_VPWR_M1002_d VPB PHIGHVT L=0.18 W=1
+ AD=0.275 AS=0.15 PD=2.55 PS=1.3 NRD=1.9503 NRS=1.9503 M=1 R=5.55556 SA=90001.1
+ SB=90000.2 A=0.18 P=2.36 MULT=1
DX8_noxref VNB VPB NWDIODE A=5.778 P=10.41
*
.include "sky130_fd_sc_hdll__a21o_1.pxi.spice"
*
.ends
*
*
